# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_io__top_xres4v2
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 200 ;
  SYMMETRY R90 ;
  PIN AMUXBUS_A
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN DISABLE_PULLUP_H
    ANTENNAPARTIALCUTAREA  0.045000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 28.635000 28.540000 33.025000 28.580000 ;
        RECT 28.635000 28.580000 28.950000 28.650000 ;
        RECT 28.635000 28.650000 28.880000 28.720000 ;
        RECT 28.635000 28.720000 28.865000 28.735000 ;
        RECT 28.635000 28.735000 28.865000 32.435000 ;
        RECT 28.685000 28.490000 33.025000 28.540000 ;
        RECT 28.755000 28.420000 33.025000 28.490000 ;
        RECT 28.825000 28.350000 33.025000 28.420000 ;
        RECT 32.555000 28.340000 33.025000 28.350000 ;
        RECT 32.625000 28.270000 33.025000 28.340000 ;
        RECT 32.695000 28.200000 33.025000 28.270000 ;
        RECT 32.760000  0.000000 33.020000  8.720000 ;
        RECT 32.760000  8.720000 33.020000  8.725000 ;
        RECT 32.760000  8.725000 33.025000  8.830000 ;
        RECT 32.765000  8.830000 33.025000  8.835000 ;
        RECT 32.765000  8.835000 33.025000 28.130000 ;
        RECT 32.765000 28.130000 33.025000 28.200000 ;
    END
    PORT
      LAYER met2 ;
        RECT 32.760000 0.000000 33.020000 0.640000 ;
    END
  END DISABLE_PULLUP_H
  PIN ENABLE_H
    ANTENNAPARTIALCUTAREA  0.180000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 12.145000  6.635000 12.545000  6.665000 ;
        RECT 12.215000  6.565000 12.545000  6.635000 ;
        RECT 12.285000  0.000000 12.545000  6.495000 ;
        RECT 12.285000  6.495000 12.545000  6.565000 ;
        RECT 12.370000  6.665000 12.545000  6.775000 ;
        RECT 12.370000  6.775000 12.545000  6.845000 ;
        RECT 12.370000  6.845000 12.615000  6.915000 ;
        RECT 12.370000  6.915000 12.685000  6.925000 ;
        RECT 12.440000  6.925000 12.695000  6.995000 ;
        RECT 12.510000  6.995000 12.765000  7.065000 ;
        RECT 12.575000  7.065000 12.835000  7.130000 ;
        RECT 12.635000  7.130000 12.900000  7.190000 ;
        RECT 12.695000  7.190000 12.900000  7.250000 ;
        RECT 12.695000  7.250000 12.900000 10.230000 ;
        RECT 12.800000 10.230000 12.865000 10.265000 ;
        RECT 12.800000 10.265000 12.830000 10.300000 ;
        RECT 12.800000 10.300000 12.825000 10.305000 ;
    END
    PORT
      LAYER met2 ;
        RECT 12.285000 0.000000 12.545000 1.470000 ;
    END
  END ENABLE_H
  PIN ENABLE_VDDIO
    ANTENNAPARTIALCUTAREA  0.200000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.425000 0.000000 8.895000 1.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.775000 17.410000  7.400000 17.515000 ;
        RECT 6.775000 17.515000  7.295000 17.620000 ;
        RECT 6.775000 17.620000  7.295000 31.295000 ;
        RECT 6.775000 31.295000  7.295000 31.400000 ;
        RECT 6.775000 31.400000  7.400000 31.505000 ;
        RECT 6.840000 17.345000  7.505000 17.410000 ;
        RECT 6.925000 31.505000  7.505000 31.655000 ;
        RECT 6.990000 17.195000  7.570000 17.345000 ;
        RECT 7.075000 31.655000  7.655000 31.805000 ;
        RECT 7.140000 17.045000  7.720000 17.195000 ;
        RECT 7.225000 31.805000  7.805000 31.955000 ;
        RECT 7.290000 16.895000  7.870000 17.045000 ;
        RECT 7.375000 31.955000  7.955000 32.105000 ;
        RECT 7.440000 16.745000  8.020000 16.895000 ;
        RECT 7.525000 32.105000  8.105000 32.255000 ;
        RECT 7.590000 16.595000  8.170000 16.745000 ;
        RECT 7.675000 32.255000  8.255000 32.405000 ;
        RECT 7.740000 16.445000  8.320000 16.595000 ;
        RECT 7.825000 32.405000  8.405000 32.555000 ;
        RECT 7.890000 16.295000  8.470000 16.445000 ;
        RECT 7.975000 32.555000  8.555000 32.705000 ;
        RECT 8.040000 16.145000  8.620000 16.295000 ;
        RECT 8.125000 32.705000  8.705000 32.855000 ;
        RECT 8.190000 15.995000  8.770000 16.145000 ;
        RECT 8.275000 32.855000  8.855000 33.005000 ;
        RECT 8.295000 15.890000  8.920000 15.995000 ;
        RECT 8.400000  0.000000  8.920000 15.785000 ;
        RECT 8.400000 15.785000  8.920000 15.890000 ;
        RECT 8.425000 33.005000  9.005000 33.155000 ;
        RECT 8.575000 33.155000  9.155000 33.305000 ;
        RECT 8.665000 33.305000  9.305000 33.395000 ;
        RECT 8.815000 33.395000 22.275000 33.545000 ;
        RECT 8.965000 33.545000 22.275000 33.695000 ;
        RECT 9.115000 33.695000 22.275000 33.845000 ;
        RECT 9.265000 33.845000 22.275000 33.995000 ;
        RECT 9.395000 33.995000 22.275000 34.125000 ;
    END
  END ENABLE_VDDIO
  PIN EN_VDDIO_SIG_H
    ANTENNAPARTIALCUTAREA  0.157500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 22.360000 0.000000 22.660000 1.205000 ;
    END
    PORT
      LAYER met2 ;
        RECT  9.735000  4.520000 10.050000  4.575000 ;
        RECT  9.735000  4.575000  9.995000  4.630000 ;
        RECT  9.735000  4.630000  9.995000  8.860000 ;
        RECT  9.735000  8.860000  9.995000  8.915000 ;
        RECT  9.735000  8.915000 10.050000  8.970000 ;
        RECT  9.790000  4.465000 10.105000  4.520000 ;
        RECT  9.805000  8.970000 10.105000  9.040000 ;
        RECT  9.860000  4.395000 10.160000  4.465000 ;
        RECT  9.875000  9.040000 10.175000  9.110000 ;
        RECT  9.930000  4.325000 10.230000  4.395000 ;
        RECT  9.945000  9.110000 10.245000  9.180000 ;
        RECT 10.000000  4.255000 10.300000  4.325000 ;
        RECT 10.015000  9.180000 10.315000  9.250000 ;
        RECT 10.070000  4.185000 10.370000  4.255000 ;
        RECT 10.085000  9.250000 10.385000  9.320000 ;
        RECT 10.140000  4.115000 10.440000  4.185000 ;
        RECT 10.155000  9.320000 10.455000  9.390000 ;
        RECT 10.210000  4.045000 10.510000  4.115000 ;
        RECT 10.225000  9.390000 10.525000  9.460000 ;
        RECT 10.280000  3.975000 10.580000  4.045000 ;
        RECT 10.295000  9.460000 10.595000  9.530000 ;
        RECT 10.350000  3.905000 10.650000  3.975000 ;
        RECT 10.365000  9.530000 10.665000  9.600000 ;
        RECT 10.420000  3.835000 10.720000  3.905000 ;
        RECT 10.435000  9.600000 10.735000  9.670000 ;
        RECT 10.490000  3.765000 10.790000  3.835000 ;
        RECT 10.505000  9.670000 10.805000  9.740000 ;
        RECT 10.560000  3.695000 10.860000  3.765000 ;
        RECT 10.575000  9.740000 10.875000  9.810000 ;
        RECT 10.610000  3.645000 15.095000  3.695000 ;
        RECT 10.645000  9.810000 10.945000  9.880000 ;
        RECT 10.650000 26.825000 11.125000 27.085000 ;
        RECT 10.650000 27.085000 11.055000 27.155000 ;
        RECT 10.650000 27.155000 10.985000 27.225000 ;
        RECT 10.650000 27.225000 10.915000 27.295000 ;
        RECT 10.650000 27.295000 10.910000 27.300000 ;
        RECT 10.650000 27.300000 10.910000 27.935000 ;
        RECT 10.650000 27.935000 10.910000 28.005000 ;
        RECT 10.650000 28.005000 10.980000 28.075000 ;
        RECT 10.650000 28.075000 11.050000 28.145000 ;
        RECT 10.650000 28.145000 11.120000 28.150000 ;
        RECT 10.650000 28.150000 11.125000 28.410000 ;
        RECT 10.655000 26.820000 11.125000 26.825000 ;
        RECT 10.680000  3.575000 15.025000  3.645000 ;
        RECT 10.715000  9.880000 11.015000  9.950000 ;
        RECT 10.720000 28.410000 11.125000 28.480000 ;
        RECT 10.725000 26.750000 11.125000 26.820000 ;
        RECT 10.750000  3.505000 14.955000  3.575000 ;
        RECT 10.755000  9.950000 11.085000  9.990000 ;
        RECT 10.790000 28.480000 11.125000 28.550000 ;
        RECT 10.795000 26.680000 11.125000 26.750000 ;
        RECT 10.810000  9.990000 11.125000 10.045000 ;
        RECT 10.820000  3.435000 14.885000  3.505000 ;
        RECT 10.860000 28.550000 11.125000 28.620000 ;
        RECT 10.865000 10.045000 11.125000 10.100000 ;
        RECT 10.865000 10.100000 11.125000 26.610000 ;
        RECT 10.865000 26.610000 11.125000 26.680000 ;
        RECT 10.865000 28.620000 11.125000 28.625000 ;
        RECT 10.865000 28.625000 11.125000 31.085000 ;
        RECT 10.865000 31.085000 11.125000 31.140000 ;
        RECT 10.865000 31.140000 11.180000 31.195000 ;
        RECT 10.935000 31.195000 11.235000 31.265000 ;
        RECT 11.005000 31.265000 11.305000 31.335000 ;
        RECT 11.075000 31.335000 11.375000 31.405000 ;
        RECT 11.145000 31.405000 11.445000 31.475000 ;
        RECT 11.150000 31.475000 11.515000 31.480000 ;
        RECT 11.205000 31.480000 11.520000 31.535000 ;
        RECT 11.260000 31.535000 11.520000 31.590000 ;
        RECT 11.260000 31.590000 11.520000 36.020000 ;
        RECT 11.260000 36.020000 12.150000 36.280000 ;
        RECT 14.845000  3.695000 15.145000  3.765000 ;
        RECT 14.915000  3.765000 15.215000  3.835000 ;
        RECT 14.985000  3.835000 15.285000  3.905000 ;
        RECT 15.055000  3.905000 15.355000  3.975000 ;
        RECT 15.125000  3.975000 15.425000  4.045000 ;
        RECT 15.195000  4.045000 15.495000  4.115000 ;
        RECT 15.265000  4.115000 15.565000  4.185000 ;
        RECT 15.335000  4.185000 15.635000  4.255000 ;
        RECT 15.405000  4.255000 15.705000  4.325000 ;
        RECT 15.475000  4.325000 15.775000  4.395000 ;
        RECT 15.545000  4.395000 15.845000  4.465000 ;
        RECT 15.615000  4.465000 15.915000  4.535000 ;
        RECT 15.625000  4.535000 15.985000  4.545000 ;
        RECT 15.695000  4.545000 28.765000  4.615000 ;
        RECT 15.765000  4.615000 28.835000  4.685000 ;
        RECT 15.835000  4.685000 28.905000  4.755000 ;
        RECT 15.885000  4.755000 28.975000  4.805000 ;
        RECT 22.065000  4.540000 22.940000  4.545000 ;
        RECT 22.135000  4.470000 22.870000  4.540000 ;
        RECT 22.205000  4.400000 22.800000  4.470000 ;
        RECT 22.275000  4.330000 22.730000  4.400000 ;
        RECT 22.345000  4.260000 22.660000  4.330000 ;
        RECT 22.350000  4.255000 22.660000  4.260000 ;
        RECT 22.355000  4.250000 22.660000  4.255000 ;
        RECT 22.360000  0.000000 22.660000  4.245000 ;
        RECT 22.360000  4.245000 22.660000  4.250000 ;
        RECT 28.725000  4.805000 29.025000  4.875000 ;
        RECT 28.795000  4.875000 29.095000  4.945000 ;
        RECT 28.865000  4.945000 29.165000  5.015000 ;
        RECT 28.935000  5.015000 29.235000  5.085000 ;
        RECT 29.005000  5.085000 29.305000  5.155000 ;
        RECT 29.075000  5.155000 29.375000  5.225000 ;
        RECT 29.145000  5.225000 29.445000  5.295000 ;
        RECT 29.210000  5.295000 29.515000  5.360000 ;
        RECT 29.265000  5.360000 29.580000  5.415000 ;
        RECT 29.320000  5.415000 29.580000  5.470000 ;
        RECT 29.320000  5.470000 29.580000 10.975000 ;
        RECT 29.320000 10.975000 29.580000 11.030000 ;
        RECT 29.320000 11.030000 29.635000 11.085000 ;
        RECT 29.390000 11.085000 29.690000 11.155000 ;
        RECT 29.460000 11.155000 29.760000 11.225000 ;
        RECT 29.530000 11.225000 29.830000 11.295000 ;
        RECT 29.600000 11.295000 29.900000 11.365000 ;
        RECT 29.660000 11.365000 29.970000 11.425000 ;
        RECT 29.715000 11.425000 30.030000 11.480000 ;
        RECT 29.770000 11.480000 30.030000 11.535000 ;
        RECT 29.770000 11.535000 30.030000 15.645000 ;
        RECT 29.770000 15.645000 30.030000 15.700000 ;
        RECT 29.770000 15.700000 30.085000 15.755000 ;
        RECT 29.840000 15.755000 30.140000 15.825000 ;
        RECT 29.910000 15.825000 30.210000 15.895000 ;
        RECT 29.980000 15.895000 30.280000 15.965000 ;
        RECT 30.050000 15.965000 30.350000 16.035000 ;
        RECT 30.120000 16.035000 30.420000 16.105000 ;
        RECT 30.190000 16.105000 30.490000 16.175000 ;
        RECT 30.255000 16.175000 30.560000 16.240000 ;
        RECT 30.310000 16.240000 30.625000 16.295000 ;
        RECT 30.365000 16.295000 30.625000 16.350000 ;
        RECT 30.365000 16.350000 30.625000 20.495000 ;
    END
  END EN_VDDIO_SIG_H
  PIN FILT_IN_H
    ANTENNAPARTIALCUTAREA  0.960000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.075000 0.000000 21.225000 3.455000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.075000 0.000000 21.225000  6.670000 ;
        RECT 20.075000 6.670000 21.225000  6.820000 ;
        RECT 20.075000 6.820000 21.375000  6.970000 ;
        RECT 20.075000 6.970000 21.525000  7.120000 ;
        RECT 20.075000 7.120000 21.675000  7.150000 ;
        RECT 20.225000 7.150000 21.705000  7.300000 ;
        RECT 20.375000 7.300000 21.855000  7.450000 ;
        RECT 20.525000 7.450000 22.005000  7.600000 ;
        RECT 20.675000 7.600000 22.155000  7.750000 ;
        RECT 20.825000 7.750000 22.305000  7.900000 ;
        RECT 20.975000 7.900000 22.455000  8.050000 ;
        RECT 21.125000 8.050000 22.605000  8.200000 ;
        RECT 21.275000 8.200000 22.755000  8.350000 ;
        RECT 21.425000 8.350000 22.905000  8.500000 ;
        RECT 21.575000 8.500000 23.055000  8.650000 ;
        RECT 21.725000 8.650000 23.205000  8.800000 ;
        RECT 21.875000 8.800000 23.355000  8.950000 ;
        RECT 22.025000 8.950000 23.505000  9.100000 ;
        RECT 22.175000 9.100000 23.655000  9.250000 ;
        RECT 22.325000 9.250000 23.805000  9.400000 ;
        RECT 22.420000 9.400000 23.955000  9.495000 ;
        RECT 22.570000 9.495000 24.050000  9.645000 ;
        RECT 22.720000 9.645000 24.050000  9.795000 ;
        RECT 22.870000 9.795000 24.050000  9.945000 ;
        RECT 22.905000 9.945000 24.050000  9.980000 ;
        RECT 22.905000 9.980000 24.050000 12.265000 ;
    END
  END FILT_IN_H
  PIN INP_SEL_H
    ANTENNAGATEAREA  6.240000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.600000 11.420000 16.830000 12.310000 ;
        RECT 16.600000 12.310000 16.830000 12.360000 ;
        RECT 16.600000 12.360000 16.880000 12.410000 ;
        RECT 16.670000 12.410000 16.930000 12.480000 ;
        RECT 16.740000 12.480000 17.000000 12.550000 ;
        RECT 16.810000 12.550000 17.070000 12.620000 ;
        RECT 16.825000 12.620000 17.140000 12.635000 ;
        RECT 16.870000 12.635000 25.295000 12.680000 ;
        RECT 16.915000 12.680000 25.340000 12.725000 ;
        RECT 16.985000 12.725000 25.385000 12.795000 ;
        RECT 17.055000 12.795000 25.385000 12.865000 ;
        RECT 24.640000 12.615000 25.275000 12.635000 ;
        RECT 24.710000 12.545000 25.205000 12.615000 ;
        RECT 24.780000 12.475000 25.135000 12.545000 ;
        RECT 24.785000 12.470000 25.135000 12.475000 ;
        RECT 24.845000 12.410000 25.135000 12.470000 ;
        RECT 24.905000  0.000000 25.135000 12.350000 ;
        RECT 24.905000 12.350000 25.135000 12.410000 ;
        RECT 24.975000 12.865000 25.385000 12.935000 ;
        RECT 25.045000 12.935000 25.385000 13.005000 ;
        RECT 25.115000 13.005000 25.385000 13.075000 ;
        RECT 25.155000 13.075000 25.385000 13.115000 ;
        RECT 25.155000 13.115000 25.385000 15.035000 ;
        RECT 25.155000 15.035000 25.385000 15.085000 ;
        RECT 25.155000 15.085000 25.435000 15.135000 ;
        RECT 25.225000 15.135000 25.485000 15.205000 ;
        RECT 25.295000 15.205000 25.555000 15.275000 ;
        RECT 25.365000 15.275000 25.625000 15.345000 ;
        RECT 25.435000 15.345000 25.695000 15.415000 ;
        RECT 25.505000 15.415000 25.765000 15.485000 ;
        RECT 25.575000 15.485000 25.835000 15.555000 ;
        RECT 25.635000 15.555000 25.905000 15.615000 ;
        RECT 25.705000 15.615000 29.965000 15.685000 ;
        RECT 25.775000 15.685000 30.035000 15.755000 ;
        RECT 25.845000 15.755000 30.105000 15.825000 ;
        RECT 25.865000 15.825000 30.175000 15.845000 ;
        RECT 29.935000 15.845000 30.195000 15.915000 ;
        RECT 30.005000 15.915000 30.265000 15.985000 ;
        RECT 30.075000 15.985000 30.335000 16.055000 ;
        RECT 30.145000 16.055000 30.405000 16.125000 ;
        RECT 30.215000 16.125000 30.475000 16.195000 ;
        RECT 30.285000 16.195000 30.545000 16.265000 ;
        RECT 30.355000 16.265000 30.615000 16.335000 ;
        RECT 30.425000 16.335000 30.685000 16.405000 ;
        RECT 30.495000 16.405000 30.755000 16.475000 ;
        RECT 30.565000 16.475000 30.825000 16.545000 ;
        RECT 30.635000 16.545000 30.895000 16.615000 ;
        RECT 30.705000 16.615000 30.965000 16.685000 ;
        RECT 30.755000 16.685000 31.035000 16.735000 ;
        RECT 30.805000 16.735000 31.035000 16.785000 ;
        RECT 30.805000 16.785000 31.035000 19.345000 ;
    END
  END INP_SEL_H
  PIN PAD
    ANTENNAPARTIALMETALSIDEAREA  245.6270 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 29.695000 127.115000 41.990000 145.625000 ;
    END
  END PAD
  PIN PAD_A_ESD_H
    ANTENNAPARTIALCUTAREA  0.960000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.245000 0.000000 18.910000 3.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.245000 0.000000 18.910000 3.135000 ;
    END
  END PAD_A_ESD_H
  PIN PULLUP_H
    ANTENNAPARTIALCUTAREA  0.270000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  6.065000 43.285000 24.570000 43.355000 ;
        RECT  6.065000 43.355000 24.500000 43.425000 ;
        RECT  6.065000 43.425000 24.430000 43.495000 ;
        RECT  6.065000 43.495000 24.380000 43.545000 ;
        RECT 14.555000  0.000000 15.135000 12.210000 ;
        RECT 14.555000 12.210000 15.135000 12.275000 ;
        RECT 14.555000 12.275000 15.200000 12.340000 ;
        RECT 14.625000 12.340000 15.265000 12.410000 ;
        RECT 14.695000 12.410000 15.335000 12.480000 ;
        RECT 14.765000 12.480000 15.405000 12.550000 ;
        RECT 14.835000 12.550000 15.475000 12.620000 ;
        RECT 14.905000 12.620000 15.545000 12.690000 ;
        RECT 14.975000 12.690000 15.615000 12.760000 ;
        RECT 15.045000 12.760000 15.685000 12.830000 ;
        RECT 15.115000 12.830000 15.755000 12.900000 ;
        RECT 15.185000 12.900000 15.825000 12.970000 ;
        RECT 15.255000 12.970000 15.895000 13.040000 ;
        RECT 15.325000 13.040000 15.965000 13.110000 ;
        RECT 15.395000 13.110000 16.035000 13.180000 ;
        RECT 15.465000 13.180000 16.105000 13.250000 ;
        RECT 15.535000 13.250000 16.175000 13.320000 ;
        RECT 15.605000 13.320000 16.245000 13.390000 ;
        RECT 15.675000 13.390000 16.315000 13.460000 ;
        RECT 15.745000 13.460000 16.385000 13.530000 ;
        RECT 15.815000 13.530000 16.455000 13.600000 ;
        RECT 15.885000 13.600000 16.525000 13.670000 ;
        RECT 15.955000 13.670000 16.595000 13.740000 ;
        RECT 16.025000 13.740000 16.665000 13.810000 ;
        RECT 16.095000 13.810000 16.735000 13.880000 ;
        RECT 16.165000 13.880000 16.805000 13.950000 ;
        RECT 16.235000 13.950000 16.875000 14.020000 ;
        RECT 16.305000 14.020000 16.945000 14.090000 ;
        RECT 16.375000 14.090000 17.015000 14.160000 ;
        RECT 16.445000 14.160000 17.085000 14.230000 ;
        RECT 16.515000 14.230000 17.155000 14.300000 ;
        RECT 16.585000 14.300000 17.225000 14.370000 ;
        RECT 16.655000 14.370000 17.295000 14.440000 ;
        RECT 16.725000 14.440000 17.365000 14.510000 ;
        RECT 16.795000 14.510000 17.435000 14.580000 ;
        RECT 16.865000 14.580000 17.505000 14.650000 ;
        RECT 16.935000 14.650000 17.575000 14.720000 ;
        RECT 17.005000 14.720000 17.645000 14.790000 ;
        RECT 17.075000 14.790000 17.715000 14.860000 ;
        RECT 17.145000 14.860000 17.785000 14.930000 ;
        RECT 17.215000 14.930000 17.855000 15.000000 ;
        RECT 17.285000 15.000000 17.925000 15.070000 ;
        RECT 17.355000 15.070000 17.995000 15.140000 ;
        RECT 17.425000 15.140000 18.065000 15.210000 ;
        RECT 17.495000 15.210000 18.135000 15.280000 ;
        RECT 17.565000 15.280000 18.205000 15.350000 ;
        RECT 17.635000 15.350000 18.275000 15.420000 ;
        RECT 17.705000 15.420000 21.745000 15.490000 ;
        RECT 17.775000 15.490000 21.815000 15.560000 ;
        RECT 17.845000 15.560000 21.885000 15.630000 ;
        RECT 17.915000 15.630000 21.955000 15.700000 ;
        RECT 17.985000 15.700000 22.025000 15.770000 ;
        RECT 18.055000 15.770000 22.095000 15.840000 ;
        RECT 18.125000 15.840000 22.165000 15.910000 ;
        RECT 18.135000 15.910000 22.235000 15.920000 ;
        RECT 21.605000 15.920000 22.245000 15.990000 ;
        RECT 21.675000 15.990000 22.315000 16.060000 ;
        RECT 21.745000 16.060000 22.385000 16.130000 ;
        RECT 21.815000 16.130000 22.455000 16.200000 ;
        RECT 21.885000 16.200000 22.525000 16.270000 ;
        RECT 21.955000 16.270000 22.595000 16.340000 ;
        RECT 22.025000 16.340000 22.665000 16.410000 ;
        RECT 22.095000 16.410000 22.735000 16.480000 ;
        RECT 22.165000 16.480000 22.805000 16.550000 ;
        RECT 22.235000 16.550000 22.875000 16.620000 ;
        RECT 22.305000 16.620000 22.945000 16.690000 ;
        RECT 22.375000 16.690000 23.015000 16.760000 ;
        RECT 22.445000 16.760000 23.085000 16.830000 ;
        RECT 22.515000 16.830000 23.155000 16.900000 ;
        RECT 22.585000 16.900000 23.225000 16.970000 ;
        RECT 22.655000 16.970000 23.295000 17.040000 ;
        RECT 22.725000 17.040000 23.365000 17.110000 ;
        RECT 22.795000 17.110000 23.435000 17.180000 ;
        RECT 22.865000 17.180000 23.505000 17.250000 ;
        RECT 22.935000 17.250000 23.575000 17.320000 ;
        RECT 23.005000 17.320000 23.645000 17.390000 ;
        RECT 23.075000 17.390000 23.715000 17.460000 ;
        RECT 23.145000 17.460000 23.785000 17.530000 ;
        RECT 23.215000 17.530000 23.855000 17.600000 ;
        RECT 23.285000 17.600000 23.925000 17.670000 ;
        RECT 23.355000 17.670000 23.995000 17.740000 ;
        RECT 23.425000 17.740000 24.065000 17.810000 ;
        RECT 23.495000 17.810000 24.135000 17.880000 ;
        RECT 23.565000 17.880000 24.205000 17.950000 ;
        RECT 23.635000 17.950000 24.275000 18.020000 ;
        RECT 23.705000 18.020000 24.345000 18.090000 ;
        RECT 23.775000 18.090000 24.415000 18.160000 ;
        RECT 23.845000 18.160000 24.485000 18.230000 ;
        RECT 23.915000 18.230000 24.555000 18.300000 ;
        RECT 23.985000 18.300000 24.625000 18.370000 ;
        RECT 24.015000 18.370000 24.695000 18.400000 ;
        RECT 24.085000 18.400000 24.725000 18.470000 ;
        RECT 24.155000 18.470000 24.725000 18.540000 ;
        RECT 24.225000 18.540000 24.725000 18.610000 ;
        RECT 24.225000 18.610000 24.725000 25.145000 ;
        RECT 24.225000 25.145000 24.725000 25.215000 ;
        RECT 24.225000 25.215000 24.795000 25.285000 ;
        RECT 24.225000 25.285000 24.865000 25.355000 ;
        RECT 24.295000 25.355000 24.935000 25.425000 ;
        RECT 24.325000 43.230000 24.640000 43.285000 ;
        RECT 24.365000 25.425000 25.005000 25.495000 ;
        RECT 24.395000 43.160000 24.695000 43.230000 ;
        RECT 24.435000 25.495000 25.075000 25.565000 ;
        RECT 24.465000 43.090000 24.765000 43.160000 ;
        RECT 24.505000 25.565000 25.145000 25.635000 ;
        RECT 24.535000 43.020000 24.835000 43.090000 ;
        RECT 24.575000 25.635000 25.215000 25.705000 ;
        RECT 24.605000 25.705000 25.285000 25.735000 ;
        RECT 24.605000 42.950000 24.905000 43.020000 ;
        RECT 24.675000 25.735000 25.315000 25.805000 ;
        RECT 24.675000 42.880000 24.975000 42.950000 ;
        RECT 24.745000 25.805000 25.315000 25.875000 ;
        RECT 24.745000 42.810000 25.045000 42.880000 ;
        RECT 24.815000 25.875000 25.315000 25.945000 ;
        RECT 24.815000 25.945000 25.315000 42.610000 ;
        RECT 24.815000 42.610000 25.250000 42.675000 ;
        RECT 24.815000 42.675000 25.185000 42.740000 ;
        RECT 24.815000 42.740000 25.115000 42.810000 ;
    END
    PORT
      LAYER met2 ;
        RECT 14.555000 0.000000 15.135000 0.985000 ;
    END
  END PULLUP_H
  PIN TIE_HI_ESD
    ANTENNAPARTIALCUTAREA  0.045000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 28.185000 4.895000 30.220000 4.965000 ;
        RECT 28.185000 4.965000 30.150000 5.035000 ;
        RECT 28.185000 5.035000 30.080000 5.105000 ;
        RECT 28.185000 5.105000 30.010000 5.175000 ;
        RECT 28.185000 5.175000 29.940000 5.245000 ;
        RECT 28.185000 5.245000 29.870000 5.315000 ;
        RECT 28.185000 5.315000 29.800000 5.385000 ;
        RECT 28.185000 5.385000 29.730000 5.455000 ;
        RECT 28.185000 5.455000 29.660000 5.525000 ;
        RECT 28.185000 5.525000 29.640000 5.545000 ;
        RECT 29.395000 4.870000 30.290000 4.895000 ;
        RECT 29.465000 4.800000 30.315000 4.870000 ;
        RECT 29.535000 4.730000 30.385000 4.800000 ;
        RECT 29.605000 4.660000 30.455000 4.730000 ;
        RECT 29.675000 4.590000 30.525000 4.660000 ;
        RECT 29.745000 4.520000 30.595000 4.590000 ;
        RECT 29.815000 4.450000 30.665000 4.520000 ;
        RECT 29.885000 4.380000 30.735000 4.450000 ;
        RECT 29.955000 4.310000 30.805000 4.380000 ;
        RECT 30.025000 4.240000 30.875000 4.310000 ;
        RECT 30.095000 4.170000 30.945000 4.240000 ;
        RECT 30.165000 4.100000 31.015000 4.170000 ;
        RECT 30.235000 4.030000 31.085000 4.100000 ;
        RECT 30.295000 3.970000 31.155000 4.030000 ;
        RECT 30.365000 3.900000 31.155000 3.970000 ;
        RECT 30.435000 3.830000 31.155000 3.900000 ;
        RECT 30.505000 0.000000 31.155000 3.760000 ;
        RECT 30.505000 3.760000 31.155000 3.830000 ;
    END
    PORT
      LAYER met2 ;
        RECT 30.505000 0.000000 31.155000 0.330000 ;
    END
  END TIE_HI_ESD
  PIN TIE_LO_ESD
    ANTENNAPARTIALCUTAREA  0.045000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 27.580000 0.000000 28.230000 2.855000 ;
        RECT 27.580000 2.855000 28.230000 2.925000 ;
        RECT 27.580000 2.925000 28.300000 2.995000 ;
        RECT 27.580000 2.995000 28.370000 3.065000 ;
        RECT 27.580000 3.065000 28.440000 3.125000 ;
        RECT 27.650000 3.125000 28.500000 3.195000 ;
        RECT 27.720000 3.195000 28.570000 3.265000 ;
        RECT 27.790000 3.265000 28.640000 3.335000 ;
        RECT 27.860000 3.335000 28.710000 3.405000 ;
        RECT 27.915000 3.405000 28.780000 3.460000 ;
        RECT 27.985000 3.460000 28.835000 3.530000 ;
        RECT 28.055000 3.530000 28.835000 3.600000 ;
        RECT 28.125000 3.600000 28.835000 3.670000 ;
        RECT 28.185000 3.670000 28.835000 3.730000 ;
        RECT 28.185000 3.730000 28.835000 4.105000 ;
    END
    PORT
      LAYER met2 ;
        RECT 27.580000 0.000000 28.230000 0.330000 ;
    END
  END TIE_LO_ESD
  PIN TIE_WEAK_HI_H
    ANTENNAPARTIALCUTAREA  0.520000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.215000 0.000000 73.235000 0.770000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.860000 71.930000 66.310000 72.080000 ;
        RECT 64.860000 72.080000 66.160000 72.230000 ;
        RECT 64.860000 72.230000 66.010000 72.380000 ;
        RECT 64.860000 72.380000 65.990000 72.400000 ;
        RECT 64.860000 72.400000 65.990000 94.645000 ;
        RECT 64.990000 71.800000 66.460000 71.930000 ;
        RECT 65.140000 71.650000 66.590000 71.800000 ;
        RECT 65.290000 71.500000 66.740000 71.650000 ;
        RECT 65.440000 71.350000 66.890000 71.500000 ;
        RECT 65.590000 71.200000 67.040000 71.350000 ;
        RECT 65.740000 71.050000 67.190000 71.200000 ;
        RECT 65.890000 70.900000 67.340000 71.050000 ;
        RECT 66.040000 70.750000 67.490000 70.900000 ;
        RECT 66.190000 70.600000 67.640000 70.750000 ;
        RECT 66.340000 70.450000 67.790000 70.600000 ;
        RECT 66.490000 70.300000 67.940000 70.450000 ;
        RECT 66.640000 70.150000 68.090000 70.300000 ;
        RECT 66.790000 70.000000 68.240000 70.150000 ;
        RECT 66.940000 69.850000 68.390000 70.000000 ;
        RECT 67.090000 69.700000 68.540000 69.850000 ;
        RECT 67.240000 69.550000 68.690000 69.700000 ;
        RECT 67.390000 69.400000 68.840000 69.550000 ;
        RECT 67.540000 69.250000 68.990000 69.400000 ;
        RECT 67.690000 69.100000 69.140000 69.250000 ;
        RECT 67.840000 68.950000 69.290000 69.100000 ;
        RECT 67.990000 68.800000 69.440000 68.950000 ;
        RECT 68.140000 68.650000 69.590000 68.800000 ;
        RECT 68.290000 68.500000 69.740000 68.650000 ;
        RECT 68.440000 68.350000 69.890000 68.500000 ;
        RECT 68.590000 68.200000 70.040000 68.350000 ;
        RECT 68.740000 68.050000 70.190000 68.200000 ;
        RECT 68.890000 67.900000 70.340000 68.050000 ;
        RECT 69.040000 67.750000 70.490000 67.900000 ;
        RECT 69.190000 67.600000 70.640000 67.750000 ;
        RECT 69.340000 67.450000 70.790000 67.600000 ;
        RECT 69.490000 67.300000 70.940000 67.450000 ;
        RECT 69.640000 67.150000 71.090000 67.300000 ;
        RECT 69.790000 67.000000 71.240000 67.150000 ;
        RECT 69.940000 66.850000 71.390000 67.000000 ;
        RECT 70.090000 66.700000 71.540000 66.850000 ;
        RECT 70.240000 66.550000 71.690000 66.700000 ;
        RECT 70.390000 66.400000 71.840000 66.550000 ;
        RECT 70.540000 66.250000 71.990000 66.400000 ;
        RECT 70.690000 66.100000 72.140000 66.250000 ;
        RECT 70.840000 65.950000 72.290000 66.100000 ;
        RECT 70.990000 65.800000 72.440000 65.950000 ;
        RECT 71.140000 65.650000 72.590000 65.800000 ;
        RECT 71.290000 65.500000 72.740000 65.650000 ;
        RECT 71.440000 65.350000 72.890000 65.500000 ;
        RECT 71.590000 65.200000 73.040000 65.350000 ;
        RECT 71.740000 65.050000 73.190000 65.200000 ;
        RECT 71.890000 64.900000 73.340000 65.050000 ;
        RECT 72.040000 64.750000 73.490000 64.900000 ;
        RECT 72.190000  0.000000 73.260000 49.320000 ;
        RECT 72.190000 49.320000 73.260000 49.470000 ;
        RECT 72.190000 49.470000 73.410000 49.620000 ;
        RECT 72.190000 49.620000 73.560000 49.770000 ;
        RECT 72.190000 49.770000 73.710000 49.920000 ;
        RECT 72.190000 49.920000 73.860000 49.985000 ;
        RECT 72.190000 49.985000 73.925000 64.465000 ;
        RECT 72.190000 64.465000 73.860000 64.530000 ;
        RECT 72.190000 64.530000 73.795000 64.595000 ;
        RECT 72.190000 64.595000 73.790000 64.600000 ;
        RECT 72.190000 64.600000 73.640000 64.750000 ;
    END
  END TIE_WEAK_HI_H
  PIN XRES_H_N
    ANTENNAPARTIALCUTAREA  0.240000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.915000 0.000000 29.685000 0.335000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.170000 10.610000 29.050000 10.760000 ;
        RECT 28.170000 10.760000 28.900000 10.910000 ;
        RECT 28.170000 10.910000 28.900000 14.770000 ;
        RECT 28.185000 10.595000 29.200000 10.610000 ;
        RECT 28.335000 10.445000 29.215000 10.595000 ;
        RECT 28.485000 10.295000 29.365000 10.445000 ;
        RECT 28.635000 10.145000 29.515000 10.295000 ;
        RECT 28.785000  9.995000 29.665000 10.145000 ;
        RECT 28.935000  0.000000 29.665000  9.845000 ;
        RECT 28.935000  9.845000 29.665000  9.995000 ;
    END
  END XRES_H_N
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 1.270000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 8.885000 75.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 1.270000 13.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 2.035000 75.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 1.270000 7.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 14.935000 75.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 0.965000 18.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 1.270000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 19.785000 75.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 70.035000 75.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 1.270000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 1.270000 94.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 19.885000 75.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 1.270000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 64.085000 75.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 1.270000 68.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 1.270000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 1.270000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 36.735000 75.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 47.735000 75.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.645000 75.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.405000 75.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.840000 1.270000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 1.270000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 36.840000 75.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 1.270000 41.655000 ;
        RECT 0.000000 41.655000 3.720000 46.170000 ;
        RECT 0.000000 46.170000 1.270000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.655000 41.630000 75.000000 46.190000 ;
        RECT 73.730000 41.585000 75.000000 41.630000 ;
        RECT 73.730000 46.190000 75.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 1.270000 46.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 1.270000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 25.835000 75.000000 30.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 1.270000 30.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 1.270000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 58.235000 75.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 1.270000 62.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 31.885000 75.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 1.270000 35.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT -0.265000 125.265000 75.000000 129.185000 ;
      RECT -0.265000 129.185000 41.620000 130.225000 ;
      RECT -0.160000 140.815000 75.160000 144.435000 ;
      RECT  0.000000  96.860000 58.340000  96.865000 ;
      RECT  0.000000  96.865000 75.000000  97.865000 ;
      RECT  0.000000  97.865000 58.340000  99.360000 ;
      RECT  0.000000  99.360000 75.000000 101.740000 ;
      RECT  0.000000 101.740000 58.340000 101.780000 ;
      RECT  0.000000 101.780000  0.165000 102.385000 ;
      RECT  0.000000 102.385000  0.455000 102.395000 ;
      RECT  0.000000 102.395000  0.595000 125.265000 ;
      RECT  0.000000 130.995000 38.355000 131.325000 ;
      RECT  0.000000 131.325000 13.200000 134.390000 ;
      RECT  0.000000 134.390000 75.000000 134.950000 ;
      RECT  0.000000 134.950000 52.445000 136.970000 ;
      RECT  0.000000 136.970000  1.045000 138.600000 ;
      RECT  0.000000 138.600000 75.000000 140.050000 ;
      RECT  0.700000 130.425000 42.015000 130.795000 ;
      RECT  0.700000 130.795000 38.355000 130.995000 ;
      RECT  0.985000   0.185000 33.890000   0.645000 ;
      RECT  0.985000   0.645000  4.525000   3.740000 ;
      RECT  0.985000   3.740000  7.065000   4.105000 ;
      RECT  0.985000 101.780000  2.645000 102.395000 ;
      RECT  1.015000   4.105000  7.065000   8.600000 ;
      RECT  1.015000   8.600000  5.625000  12.860000 ;
      RECT  1.015000  12.860000  6.055000  13.870000 ;
      RECT  1.015000  13.870000  5.625000  17.770000 ;
      RECT  1.015000  17.770000 14.130000  18.870000 ;
      RECT  1.015000  18.870000  5.605000  37.435000 ;
      RECT  1.015000  37.435000 14.270000  38.625000 ;
      RECT  1.015000  38.625000  4.525000  71.780000 ;
      RECT  1.015000  71.780000 31.450000  84.665000 ;
      RECT  1.100000  85.320000  2.790000  96.860000 ;
      RECT  1.145000  84.665000 31.450000  85.320000 ;
      RECT 11.005000  17.765000 11.270000  17.770000 ;
      RECT 11.270000  18.870000 14.130000  25.580000 ;
      RECT 13.095000   3.770000 16.800000   6.465000 ;
      RECT 13.095000   6.465000 32.410000   6.520000 ;
      RECT 13.095000   6.520000 32.395000   8.665000 ;
      RECT 13.460000  25.580000 14.130000  27.375000 ;
      RECT 13.460000  27.375000 20.685000  27.545000 ;
      RECT 13.460000  27.545000 14.130000  34.045000 ;
      RECT 14.130000 136.970000 52.445000 137.930000 ;
      RECT 14.130000 137.930000 75.000000 138.600000 ;
      RECT 14.165000  13.360000 14.435000  13.735000 ;
      RECT 14.185000   8.665000 14.385000  12.750000 ;
      RECT 14.480000  13.050000 24.760000  15.670000 ;
      RECT 16.115000  10.105000 16.285000  10.160000 ;
      RECT 16.115000  10.160000 16.800000  10.330000 ;
      RECT 16.115000  10.330000 16.285000  10.635000 ;
      RECT 16.130000  11.590000 16.800000  11.760000 ;
      RECT 16.630000  11.480000 16.800000  11.590000 ;
      RECT 16.630000  11.760000 16.800000  12.010000 ;
      RECT 16.950000  15.670000 24.760000  15.930000 ;
      RECT 16.950000  15.930000 32.350000  16.600000 ;
      RECT 16.950000  16.600000 26.460000  18.815000 ;
      RECT 17.885000   0.645000 33.890000   3.235000 ;
      RECT 18.700000  18.815000 26.460000  20.255000 ;
      RECT 18.885000  24.405000 20.685000  27.375000 ;
      RECT 19.155000  39.220000 26.270000  41.890000 ;
      RECT 19.155000  41.890000 32.495000  42.120000 ;
      RECT 19.155000  42.120000 32.435000  43.020000 ;
      RECT 20.685000  20.255000 26.460000  20.490000 ;
      RECT 20.855000  20.490000 26.460000  21.035000 ;
      RECT 20.855000  24.480000 26.460000  25.800000 ;
      RECT 21.135000  37.530000 26.270000  39.220000 ;
      RECT 23.730000  21.035000 26.460000  24.480000 ;
      RECT 24.035000 131.325000 25.835000 134.390000 ;
      RECT 24.435000  11.465000 25.140000  11.995000 ;
      RECT 24.470000   9.975000 25.105000  10.160000 ;
      RECT 24.470000  10.160000 25.140000  10.330000 ;
      RECT 24.470000  10.330000 25.105000  10.505000 ;
      RECT 25.070000  25.800000 26.460000  26.780000 ;
      RECT 25.070000  26.780000 32.625000  27.950000 ;
      RECT 25.070000  27.950000 27.385000  33.830000 ;
      RECT 25.070000  33.830000 32.435000  33.940000 ;
      RECT 25.070000  33.940000 32.495000  34.170000 ;
      RECT 25.070000  34.170000 26.270000  37.530000 ;
      RECT 25.140000  47.770000 31.450000  71.780000 ;
      RECT 26.480000  14.880000 26.650000  15.410000 ;
      RECT 26.975000  34.730000 31.525000  34.960000 ;
      RECT 26.975000  34.960000 27.205000  40.965000 ;
      RECT 26.975000  40.965000 31.525000  41.195000 ;
      RECT 27.370000  17.445000 27.540000  25.820000 ;
      RECT 27.760000  14.880000 27.930000  15.410000 ;
      RECT 27.850000  35.215000 30.690000  35.385000 ;
      RECT 28.665000  30.760000 28.835000  31.290000 ;
      RECT 28.665000  31.845000 28.835000  32.375000 ;
      RECT 29.035000  28.960000 29.205000  29.490000 ;
      RECT 29.035000  30.070000 29.205000  30.600000 ;
      RECT 29.065000  31.460000 29.595000  31.630000 ;
      RECT 29.150000  18.365000 29.680000  18.535000 ;
      RECT 29.150000  20.125000 29.680000  20.295000 ;
      RECT 29.330000  24.890000 30.490000  25.220000 ;
      RECT 29.455000   3.235000 32.410000   6.465000 ;
      RECT 30.105000  25.405000 30.635000  25.575000 ;
      RECT 30.115000  29.700000 30.645000  29.870000 ;
      RECT 30.215000  14.720000 30.385000  15.250000 ;
      RECT 30.415000  19.390000 30.585000  19.920000 ;
      RECT 30.415000  20.510000 30.585000  21.040000 ;
      RECT 30.835000  17.635000 31.005000  18.165000 ;
      RECT 30.835000  18.755000 31.005000  19.285000 ;
      RECT 30.960000  46.750000 31.490000  46.920000 ;
      RECT 31.130000  46.485000 31.490000  46.750000 ;
      RECT 31.130000  46.920000 31.490000  47.155000 ;
      RECT 31.295000  34.960000 31.525000  40.965000 ;
      RECT 31.495000  14.720000 31.665000  15.250000 ;
      RECT 32.155000  28.780000 32.325000  32.550000 ;
      RECT 32.265000  34.170000 32.495000  41.890000 ;
      RECT 33.420000  73.960000 33.870000  81.465000 ;
      RECT 33.445000  82.260000 34.600000  83.340000 ;
      RECT 33.535000  81.905000 34.065000  82.075000 ;
      RECT 34.850000  83.100000 35.380000  83.270000 ;
      RECT 35.090000   0.900000 38.860000   1.070000 ;
      RECT 35.160000   1.070000 38.860000   1.080000 ;
      RECT 36.555000 131.325000 38.355000 134.390000 ;
      RECT 38.970000 133.145000 40.600000 133.825000 ;
      RECT 40.040000   0.195000 74.560000   5.755000 ;
      RECT 40.335000   5.755000 74.560000   5.960000 ;
      RECT 40.495000 130.795000 42.015000 130.995000 ;
      RECT 40.495000 130.995000 75.000000 132.595000 ;
      RECT 42.840000 129.770000 43.730000 130.440000 ;
      RECT 43.350000  60.495000 43.720000  78.760000 ;
      RECT 48.290000 129.770000 50.440000 130.440000 ;
      RECT 51.880000 133.145000 52.770000 133.815000 ;
      RECT 53.575000 135.430000 55.095000 137.450000 ;
      RECT 53.970000   5.960000 74.560000   6.580000 ;
      RECT 55.000000 129.770000 56.460000 130.440000 ;
      RECT 58.340000 102.310000 72.060000 102.395000 ;
      RECT 60.770000 133.145000 61.800000 133.815000 ;
      RECT 60.855000 129.760000 61.780000 130.430000 ;
      RECT 62.040000 129.185000 75.000000 130.225000 ;
      RECT 62.065000 132.595000 75.000000 134.390000 ;
      RECT 62.730000   6.580000 63.170000  59.670000 ;
      RECT 63.130000  60.940000 63.180000  85.005000 ;
      RECT 67.105000 134.950000 75.000000 137.930000 ;
      RECT 68.960000  85.895000 71.490000  86.125000 ;
      RECT 68.960000  86.125000 74.315000  94.410000 ;
      RECT 69.260000  94.410000 74.315000  96.865000 ;
      RECT 72.060000  97.865000 75.000000  99.360000 ;
      RECT 72.060000 101.740000 75.000000 101.780000 ;
      RECT 73.265000   6.580000 74.560000  84.995000 ;
      RECT 73.265000  84.995000 73.855000  85.020000 ;
      RECT 74.355000 101.780000 75.000000 125.265000 ;
    LAYER met1 ;
      RECT -0.145000  95.895000  2.680000  95.965000 ;
      RECT -0.145000  95.965000  2.750000  96.035000 ;
      RECT -0.145000  96.035000  2.820000  96.105000 ;
      RECT -0.145000  96.105000  2.890000  96.175000 ;
      RECT -0.145000  96.175000  2.960000  96.245000 ;
      RECT -0.145000  96.245000  3.030000  96.315000 ;
      RECT -0.145000  96.315000  3.100000  96.385000 ;
      RECT -0.145000  96.385000  3.170000  96.455000 ;
      RECT -0.145000  96.455000  3.240000  96.525000 ;
      RECT -0.145000  96.525000  3.310000  96.595000 ;
      RECT -0.145000  96.543000  3.328000  96.610000 ;
      RECT -0.145000  96.543000  3.328000  96.610000 ;
      RECT -0.145000  96.595000  3.380000  96.665000 ;
      RECT -0.145000  96.610000  3.395000  96.680000 ;
      RECT -0.145000  96.610000  3.395000  96.680000 ;
      RECT -0.145000  96.665000  3.450000  96.735000 ;
      RECT -0.145000  96.680000  3.465000  96.750000 ;
      RECT -0.145000  96.680000  3.465000  96.750000 ;
      RECT -0.145000  96.735000  3.520000  96.805000 ;
      RECT -0.145000  96.750000  3.535000  96.820000 ;
      RECT -0.145000  96.750000  3.535000  96.820000 ;
      RECT -0.145000  96.805000  3.590000  96.875000 ;
      RECT -0.145000  96.820000  3.605000  96.890000 ;
      RECT -0.145000  96.820000  3.605000  96.890000 ;
      RECT -0.145000  96.875000  3.660000  96.945000 ;
      RECT -0.145000  96.890000  3.675000  96.960000 ;
      RECT -0.145000  96.890000  3.675000  96.960000 ;
      RECT -0.145000  96.945000  3.730000  97.015000 ;
      RECT -0.145000  96.960000  3.745000  97.030000 ;
      RECT -0.145000  96.960000  3.745000  97.030000 ;
      RECT -0.145000  97.015000  3.800000  97.085000 ;
      RECT -0.145000  97.030000  3.815000  97.100000 ;
      RECT -0.145000  97.030000  3.815000  97.100000 ;
      RECT -0.145000  97.085000  3.870000  97.155000 ;
      RECT -0.145000  97.100000  3.885000  97.170000 ;
      RECT -0.145000  97.100000  3.885000  97.170000 ;
      RECT -0.145000  97.155000  3.940000  97.225000 ;
      RECT -0.145000  97.170000  3.955000  97.240000 ;
      RECT -0.145000  97.170000  3.955000  97.240000 ;
      RECT -0.145000  97.225000  4.010000  97.295000 ;
      RECT -0.145000  97.240000  4.025000  97.310000 ;
      RECT -0.145000  97.240000  4.025000  97.310000 ;
      RECT -0.145000  97.295000  4.080000  97.365000 ;
      RECT -0.145000  97.310000  4.095000  97.380000 ;
      RECT -0.145000  97.310000  4.095000  97.380000 ;
      RECT -0.145000  97.365000  4.150000  97.435000 ;
      RECT -0.145000  97.380000  4.165000  97.450000 ;
      RECT -0.145000  97.380000  4.165000  97.450000 ;
      RECT -0.145000  97.435000  4.220000  97.505000 ;
      RECT -0.145000  97.450000  4.235000  97.520000 ;
      RECT -0.145000  97.450000  4.235000  97.520000 ;
      RECT -0.145000  97.505000  4.290000  97.530000 ;
      RECT -0.145000  97.520000  4.305000  97.530000 ;
      RECT -0.145000  97.520000  4.305000  97.530000 ;
      RECT -0.145000  97.530000 56.545000 100.330000 ;
      RECT -0.145000 100.330000 56.545000 101.420000 ;
      RECT -0.145000 125.440000 14.680000 125.510000 ;
      RECT -0.145000 125.440000 14.680000 125.510000 ;
      RECT -0.145000 125.510000 14.610000 125.580000 ;
      RECT -0.145000 125.510000 14.610000 125.580000 ;
      RECT -0.145000 125.580000 14.540000 125.650000 ;
      RECT -0.145000 125.580000 14.540000 125.650000 ;
      RECT -0.145000 125.650000 14.470000 125.720000 ;
      RECT -0.145000 125.650000 14.470000 125.720000 ;
      RECT -0.145000 125.720000 14.400000 125.790000 ;
      RECT -0.145000 125.720000 14.400000 125.790000 ;
      RECT -0.145000 125.790000 14.330000 125.860000 ;
      RECT -0.145000 125.790000 14.330000 125.860000 ;
      RECT -0.145000 125.860000 14.260000 125.930000 ;
      RECT -0.145000 125.860000 14.260000 125.930000 ;
      RECT -0.145000 125.930000 14.190000 126.000000 ;
      RECT -0.145000 125.930000 14.190000 126.000000 ;
      RECT -0.145000 126.000000 14.120000 126.070000 ;
      RECT -0.145000 126.000000 14.120000 126.070000 ;
      RECT -0.145000 126.070000 14.050000 126.140000 ;
      RECT -0.145000 126.070000 14.050000 126.140000 ;
      RECT -0.145000 126.140000 13.980000 126.210000 ;
      RECT -0.145000 126.140000 13.980000 126.210000 ;
      RECT -0.145000 126.210000 13.910000 126.280000 ;
      RECT -0.145000 126.210000 13.910000 126.280000 ;
      RECT -0.145000 126.280000 13.840000 126.350000 ;
      RECT -0.145000 126.280000 13.840000 126.350000 ;
      RECT -0.145000 126.350000 13.770000 126.420000 ;
      RECT -0.145000 126.350000 13.770000 126.420000 ;
      RECT -0.145000 126.420000 13.700000 126.490000 ;
      RECT -0.145000 126.420000 13.700000 126.490000 ;
      RECT -0.145000 126.490000 13.630000 126.560000 ;
      RECT -0.145000 126.490000 13.630000 126.560000 ;
      RECT -0.145000 126.560000 13.560000 126.630000 ;
      RECT -0.145000 126.560000 13.560000 126.630000 ;
      RECT -0.145000 126.630000 13.490000 126.700000 ;
      RECT -0.145000 126.630000 13.490000 126.700000 ;
      RECT -0.145000 126.700000 13.420000 126.770000 ;
      RECT -0.145000 126.700000 13.420000 126.770000 ;
      RECT -0.145000 126.770000 13.350000 126.840000 ;
      RECT -0.145000 126.770000 13.350000 126.840000 ;
      RECT -0.145000 126.840000 13.280000 126.910000 ;
      RECT -0.145000 126.840000 13.280000 126.910000 ;
      RECT -0.145000 126.910000 13.210000 126.980000 ;
      RECT -0.145000 126.910000 13.210000 126.980000 ;
      RECT -0.145000 126.980000 13.140000 127.050000 ;
      RECT -0.145000 126.980000 13.140000 127.050000 ;
      RECT -0.145000 127.050000 13.070000 127.120000 ;
      RECT -0.145000 127.050000 13.070000 127.120000 ;
      RECT -0.145000 127.120000 13.000000 127.190000 ;
      RECT -0.145000 127.120000 13.000000 127.190000 ;
      RECT -0.145000 127.190000 12.930000 127.260000 ;
      RECT -0.145000 127.190000 12.930000 127.260000 ;
      RECT -0.145000 127.260000 12.860000 127.330000 ;
      RECT -0.145000 127.260000 12.860000 127.330000 ;
      RECT -0.145000 127.330000 12.790000 127.400000 ;
      RECT -0.145000 127.330000 12.790000 127.400000 ;
      RECT -0.145000 127.400000 12.720000 127.470000 ;
      RECT -0.145000 127.400000 12.720000 127.470000 ;
      RECT -0.145000 127.470000 12.650000 127.540000 ;
      RECT -0.145000 127.470000 12.650000 127.540000 ;
      RECT -0.145000 127.540000 12.580000 127.610000 ;
      RECT -0.145000 127.540000 12.580000 127.610000 ;
      RECT -0.145000 127.610000 12.510000 127.680000 ;
      RECT -0.145000 127.610000 12.510000 127.680000 ;
      RECT -0.145000 127.680000 12.440000 127.750000 ;
      RECT -0.145000 127.680000 12.440000 127.750000 ;
      RECT -0.145000 127.750000 12.370000 127.820000 ;
      RECT -0.145000 127.750000 12.370000 127.820000 ;
      RECT -0.145000 127.820000 12.300000 127.890000 ;
      RECT -0.145000 127.820000 12.300000 127.890000 ;
      RECT -0.145000 127.890000 12.230000 127.960000 ;
      RECT -0.145000 127.890000 12.230000 127.960000 ;
      RECT -0.145000 127.960000 12.160000 128.030000 ;
      RECT -0.145000 127.960000 12.160000 128.030000 ;
      RECT -0.145000 128.030000 12.090000 128.100000 ;
      RECT -0.145000 128.030000 12.090000 128.100000 ;
      RECT -0.145000 128.100000 12.020000 128.170000 ;
      RECT -0.145000 128.100000 12.020000 128.170000 ;
      RECT -0.145000 128.170000 11.950000 128.240000 ;
      RECT -0.145000 128.170000 11.950000 128.240000 ;
      RECT -0.145000 128.240000 11.930000 128.260000 ;
      RECT -0.145000 128.240000 11.930000 128.260000 ;
      RECT -0.145000 128.260000 11.860000 128.330000 ;
      RECT -0.145000 128.260000 11.860000 128.330000 ;
      RECT -0.145000 128.330000 11.790000 128.400000 ;
      RECT -0.145000 128.330000 11.790000 128.400000 ;
      RECT -0.145000 128.400000 11.720000 128.470000 ;
      RECT -0.145000 128.400000 11.720000 128.470000 ;
      RECT -0.145000 128.470000 11.650000 128.540000 ;
      RECT -0.145000 128.470000 11.650000 128.540000 ;
      RECT -0.145000 128.540000 11.580000 128.610000 ;
      RECT -0.145000 128.540000 11.580000 128.610000 ;
      RECT -0.145000 128.610000 11.510000 128.680000 ;
      RECT -0.145000 128.610000 11.510000 128.680000 ;
      RECT -0.145000 128.680000 11.440000 128.750000 ;
      RECT -0.145000 128.680000 11.440000 128.750000 ;
      RECT -0.145000 128.750000 11.370000 128.820000 ;
      RECT -0.145000 128.750000 11.370000 128.820000 ;
      RECT -0.145000 128.820000 11.300000 128.890000 ;
      RECT -0.145000 128.820000 11.300000 128.890000 ;
      RECT -0.145000 128.890000 11.230000 128.960000 ;
      RECT -0.145000 128.890000 11.230000 128.960000 ;
      RECT -0.145000 128.960000 11.160000 129.030000 ;
      RECT -0.145000 128.960000 11.160000 129.030000 ;
      RECT -0.145000 129.030000 11.090000 129.100000 ;
      RECT -0.145000 129.030000 11.090000 129.100000 ;
      RECT -0.145000 129.100000 11.020000 129.170000 ;
      RECT -0.145000 129.100000 11.020000 129.170000 ;
      RECT -0.145000 129.170000 10.950000 129.240000 ;
      RECT -0.145000 129.170000 10.950000 129.240000 ;
      RECT -0.145000 129.240000 10.880000 129.310000 ;
      RECT -0.145000 129.240000 10.880000 129.310000 ;
      RECT -0.145000 129.310000 10.810000 129.380000 ;
      RECT -0.145000 129.310000 10.810000 129.380000 ;
      RECT -0.145000 129.380000 10.740000 129.450000 ;
      RECT -0.145000 129.380000 10.740000 129.450000 ;
      RECT -0.145000 129.450000 10.670000 129.520000 ;
      RECT -0.145000 129.450000 10.670000 129.520000 ;
      RECT -0.145000 129.520000 10.600000 129.590000 ;
      RECT -0.145000 129.520000 10.600000 129.590000 ;
      RECT -0.145000 129.590000 10.530000 129.660000 ;
      RECT -0.145000 129.590000 10.530000 129.660000 ;
      RECT -0.145000 129.660000 10.460000 129.730000 ;
      RECT -0.145000 129.660000 10.460000 129.730000 ;
      RECT -0.145000 129.730000 10.390000 129.800000 ;
      RECT -0.145000 129.730000 10.390000 129.800000 ;
      RECT -0.145000 129.800000 10.320000 129.870000 ;
      RECT -0.145000 129.800000 10.320000 129.870000 ;
      RECT -0.145000 129.870000 10.250000 129.940000 ;
      RECT -0.145000 129.870000 10.250000 129.940000 ;
      RECT -0.145000 129.940000 10.180000 130.010000 ;
      RECT -0.145000 129.940000 10.180000 130.010000 ;
      RECT -0.145000 130.010000 10.110000 130.080000 ;
      RECT -0.145000 130.010000 10.110000 130.080000 ;
      RECT -0.145000 130.080000 10.040000 130.150000 ;
      RECT -0.145000 130.080000 10.040000 130.150000 ;
      RECT -0.145000 130.150000  9.970000 130.220000 ;
      RECT -0.145000 130.150000  9.970000 130.220000 ;
      RECT -0.145000 131.275000  0.940000 131.345000 ;
      RECT -0.145000 131.275000  0.940000 131.345000 ;
      RECT -0.145000 131.345000  1.010000 131.415000 ;
      RECT -0.145000 131.345000  1.010000 131.415000 ;
      RECT -0.145000 131.415000  1.080000 131.485000 ;
      RECT -0.145000 131.415000  1.080000 131.485000 ;
      RECT -0.145000 131.485000  1.150000 131.555000 ;
      RECT -0.145000 131.485000  1.150000 131.555000 ;
      RECT -0.145000 131.555000  1.220000 131.625000 ;
      RECT -0.145000 131.555000  1.220000 131.625000 ;
      RECT -0.145000 131.625000  1.290000 131.695000 ;
      RECT -0.145000 131.625000  1.290000 131.695000 ;
      RECT -0.145000 131.695000  1.360000 131.765000 ;
      RECT -0.145000 131.695000  1.360000 131.765000 ;
      RECT -0.145000 131.765000  1.430000 131.835000 ;
      RECT -0.145000 131.765000  1.430000 131.835000 ;
      RECT -0.145000 131.835000  1.500000 131.905000 ;
      RECT -0.145000 131.835000  1.500000 131.905000 ;
      RECT -0.145000 131.905000  1.570000 131.975000 ;
      RECT -0.145000 131.905000  1.570000 131.975000 ;
      RECT -0.145000 131.975000  1.640000 132.045000 ;
      RECT -0.145000 131.975000  1.640000 132.045000 ;
      RECT -0.145000 132.045000  1.710000 132.115000 ;
      RECT -0.145000 132.045000  1.710000 132.115000 ;
      RECT -0.145000 132.115000  1.780000 132.185000 ;
      RECT -0.145000 132.115000  1.780000 132.185000 ;
      RECT -0.145000 132.185000  1.850000 132.255000 ;
      RECT -0.145000 132.185000  1.850000 132.255000 ;
      RECT -0.145000 132.255000  1.920000 132.325000 ;
      RECT -0.145000 132.255000  1.920000 132.325000 ;
      RECT -0.145000 132.325000  1.990000 132.395000 ;
      RECT -0.145000 132.325000  1.990000 132.395000 ;
      RECT -0.145000 132.395000  2.060000 132.465000 ;
      RECT -0.145000 132.395000  2.060000 132.465000 ;
      RECT -0.145000 132.465000  2.130000 132.535000 ;
      RECT -0.145000 132.465000  2.130000 132.535000 ;
      RECT -0.145000 132.535000  2.200000 132.605000 ;
      RECT -0.145000 132.535000  2.200000 132.605000 ;
      RECT -0.145000 132.605000  2.270000 132.675000 ;
      RECT -0.145000 132.605000  2.270000 132.675000 ;
      RECT -0.145000 132.675000  2.340000 132.740000 ;
      RECT -0.145000 132.675000  2.340000 132.740000 ;
      RECT -0.145000 132.740000  2.405000 132.810000 ;
      RECT -0.145000 132.740000  2.405000 132.810000 ;
      RECT -0.145000 132.810000  2.475000 132.880000 ;
      RECT -0.145000 132.810000  2.475000 132.880000 ;
      RECT -0.145000 132.880000  2.545000 132.950000 ;
      RECT -0.145000 132.880000  2.545000 132.950000 ;
      RECT -0.145000 132.950000  2.615000 133.020000 ;
      RECT -0.145000 132.950000  2.615000 133.020000 ;
      RECT -0.145000 133.020000  2.685000 133.090000 ;
      RECT -0.145000 133.020000  2.685000 133.090000 ;
      RECT -0.145000 133.090000  2.755000 133.160000 ;
      RECT -0.145000 133.090000  2.755000 133.160000 ;
      RECT -0.145000 133.160000  2.825000 133.230000 ;
      RECT -0.145000 133.160000  2.825000 133.230000 ;
      RECT -0.145000 133.230000  2.895000 133.300000 ;
      RECT -0.145000 133.230000  2.895000 133.300000 ;
      RECT -0.145000 133.300000  2.965000 133.370000 ;
      RECT -0.145000 133.300000  2.965000 133.370000 ;
      RECT -0.145000 133.370000  3.035000 133.440000 ;
      RECT -0.145000 133.370000  3.035000 133.440000 ;
      RECT -0.145000 133.440000  3.105000 133.510000 ;
      RECT -0.145000 133.440000  3.105000 133.510000 ;
      RECT -0.145000 133.510000  3.175000 133.580000 ;
      RECT -0.145000 133.510000  3.175000 133.580000 ;
      RECT -0.145000 133.580000  3.245000 133.650000 ;
      RECT -0.145000 133.580000  3.245000 133.650000 ;
      RECT -0.145000 133.650000  3.315000 133.720000 ;
      RECT -0.145000 133.650000  3.315000 133.720000 ;
      RECT -0.145000 133.720000  3.385000 133.790000 ;
      RECT -0.145000 133.720000  3.385000 133.790000 ;
      RECT -0.145000 133.790000  3.455000 133.860000 ;
      RECT -0.145000 133.790000  3.455000 133.860000 ;
      RECT -0.145000 133.860000  3.525000 133.930000 ;
      RECT -0.145000 133.860000  3.525000 133.930000 ;
      RECT -0.145000 133.930000  3.595000 134.000000 ;
      RECT -0.145000 133.930000  3.595000 134.000000 ;
      RECT -0.145000 134.000000  3.665000 134.070000 ;
      RECT -0.145000 134.000000  3.665000 134.070000 ;
      RECT -0.145000 134.070000  3.735000 134.140000 ;
      RECT -0.145000 134.070000  3.735000 134.140000 ;
      RECT -0.145000 134.140000  3.805000 134.180000 ;
      RECT -0.145000 134.140000  3.805000 134.180000 ;
      RECT -0.145000 134.179000  3.773000 134.250000 ;
      RECT -0.145000 134.179000  3.773000 134.250000 ;
      RECT -0.145000 134.250000  3.703000 134.320000 ;
      RECT -0.145000 134.250000  3.703000 134.320000 ;
      RECT -0.145000 134.320000  3.633000 134.390000 ;
      RECT -0.145000 134.320000  3.633000 134.390000 ;
      RECT -0.145000 134.390000  3.562000 134.460000 ;
      RECT -0.145000 134.390000  3.562000 134.460000 ;
      RECT -0.145000 134.460000  3.492000 134.530000 ;
      RECT -0.145000 134.460000  3.492000 134.530000 ;
      RECT -0.145000 134.530000  3.422000 134.600000 ;
      RECT -0.145000 134.530000  3.422000 134.600000 ;
      RECT -0.145000 134.600000  3.352000 134.670000 ;
      RECT -0.145000 134.600000  3.352000 134.670000 ;
      RECT -0.145000 134.670000  3.282000 134.740000 ;
      RECT -0.145000 134.670000  3.282000 134.740000 ;
      RECT -0.145000 134.740000  3.212000 134.810000 ;
      RECT -0.145000 134.740000  3.212000 134.810000 ;
      RECT -0.145000 134.810000  3.141000 134.880000 ;
      RECT -0.145000 134.810000  3.141000 134.880000 ;
      RECT -0.145000 134.880000  3.071000 134.950000 ;
      RECT -0.145000 134.880000  3.071000 134.950000 ;
      RECT -0.145000 134.950000  3.001000 135.020000 ;
      RECT -0.145000 134.950000  3.001000 135.020000 ;
      RECT -0.145000 135.020000  2.931000 135.090000 ;
      RECT -0.145000 135.020000  2.931000 135.090000 ;
      RECT -0.145000 135.090000  2.861000 135.160000 ;
      RECT -0.145000 135.090000  2.861000 135.160000 ;
      RECT -0.145000 135.160000  2.791000 135.230000 ;
      RECT -0.145000 135.160000  2.791000 135.230000 ;
      RECT -0.145000 135.230000  2.720000 135.300000 ;
      RECT -0.145000 135.230000  2.720000 135.300000 ;
      RECT -0.145000 135.300000  2.650000 135.370000 ;
      RECT -0.145000 135.300000  2.650000 135.370000 ;
      RECT -0.145000 135.370000  2.580000 135.440000 ;
      RECT -0.145000 135.370000  2.580000 135.440000 ;
      RECT -0.145000 135.440000  2.550000 135.470000 ;
      RECT -0.145000 135.440000  2.550000 135.470000 ;
      RECT -0.145000 135.470000  2.480000 135.540000 ;
      RECT -0.145000 135.470000  2.480000 135.540000 ;
      RECT -0.145000 135.540000  2.410000 135.610000 ;
      RECT -0.145000 135.540000  2.410000 135.610000 ;
      RECT -0.145000 135.610000  2.339000 135.680000 ;
      RECT -0.145000 135.610000  2.339000 135.680000 ;
      RECT -0.145000 135.680000  2.269000 135.750000 ;
      RECT -0.145000 135.680000  2.269000 135.750000 ;
      RECT -0.145000 135.750000  2.199000 135.820000 ;
      RECT -0.145000 135.750000  2.199000 135.820000 ;
      RECT -0.145000 135.820000  2.129000 135.890000 ;
      RECT -0.145000 135.820000  2.129000 135.890000 ;
      RECT -0.145000 135.890000  2.059000 135.960000 ;
      RECT -0.145000 135.890000  2.059000 135.960000 ;
      RECT -0.145000 135.960000  1.989000 136.030000 ;
      RECT -0.145000 135.960000  1.989000 136.030000 ;
      RECT -0.145000 136.030000  1.918000 136.100000 ;
      RECT -0.145000 136.030000  1.918000 136.100000 ;
      RECT -0.145000 136.100000  1.848000 136.170000 ;
      RECT -0.145000 136.100000  1.848000 136.170000 ;
      RECT -0.145000 136.170000  1.778000 136.240000 ;
      RECT -0.145000 136.170000  1.778000 136.240000 ;
      RECT -0.145000 136.240000  1.708000 136.310000 ;
      RECT -0.145000 136.240000  1.708000 136.310000 ;
      RECT -0.145000 136.310000  1.638000 136.380000 ;
      RECT -0.145000 136.310000  1.638000 136.380000 ;
      RECT -0.145000 136.380000  1.568000 136.450000 ;
      RECT -0.145000 136.380000  1.568000 136.450000 ;
      RECT -0.145000 136.450000  1.497000 136.520000 ;
      RECT -0.145000 136.450000  1.497000 136.520000 ;
      RECT -0.145000 136.520000  1.427000 136.590000 ;
      RECT -0.145000 136.520000  1.427000 136.590000 ;
      RECT -0.145000 136.590000  1.357000 136.660000 ;
      RECT -0.145000 136.590000  1.357000 136.660000 ;
      RECT -0.145000 136.660000  1.287000 136.730000 ;
      RECT -0.145000 136.660000  1.287000 136.730000 ;
      RECT -0.145000 136.730000  1.217000 136.800000 ;
      RECT -0.145000 136.730000  1.217000 136.800000 ;
      RECT -0.145000 136.800000  1.147000 136.870000 ;
      RECT -0.145000 136.800000  1.147000 136.870000 ;
      RECT -0.145000 136.870000  1.076000 136.940000 ;
      RECT -0.145000 136.870000  1.076000 136.940000 ;
      RECT -0.145000 136.940000  1.006000 137.010000 ;
      RECT -0.145000 136.940000  1.006000 137.010000 ;
      RECT -0.145000 137.010000  0.936000 137.080000 ;
      RECT -0.145000 137.010000  0.936000 137.080000 ;
      RECT -0.145000 137.080000  0.866000 137.150000 ;
      RECT -0.145000 137.080000  0.866000 137.150000 ;
      RECT -0.145000 137.150000  0.796000 137.220000 ;
      RECT -0.145000 137.150000  0.796000 137.220000 ;
      RECT -0.145000 137.220000  0.725000 137.290000 ;
      RECT -0.145000 137.220000  0.725000 137.290000 ;
      RECT -0.145000 137.290000  0.655000 137.360000 ;
      RECT -0.145000 137.290000  0.655000 137.360000 ;
      RECT -0.145000 137.360000  0.585000 137.430000 ;
      RECT -0.145000 137.360000  0.585000 137.430000 ;
      RECT -0.145000 137.430000  0.515000 137.500000 ;
      RECT -0.145000 137.430000  0.515000 137.500000 ;
      RECT -0.145000 137.500000  0.445000 137.570000 ;
      RECT -0.145000 137.500000  0.445000 137.570000 ;
      RECT -0.145000 137.570000  0.374000 137.640000 ;
      RECT -0.145000 137.570000  0.374000 137.640000 ;
      RECT -0.145000 137.640000  0.304000 137.710000 ;
      RECT -0.145000 137.640000  0.304000 137.710000 ;
      RECT -0.145000 137.710000  0.234000 137.780000 ;
      RECT -0.145000 137.710000  0.234000 137.780000 ;
      RECT -0.145000 137.780000  0.164000 137.850000 ;
      RECT -0.145000 137.780000  0.164000 137.850000 ;
      RECT -0.145000 137.850000  0.094000 137.920000 ;
      RECT -0.145000 137.850000  0.094000 137.920000 ;
      RECT -0.145000 137.920000  0.023000 137.990000 ;
      RECT -0.145000 137.920000  0.023000 137.990000 ;
      RECT -0.145000 137.990000 -0.047000 138.060000 ;
      RECT -0.145000 137.990000 -0.047000 138.060000 ;
      RECT -0.145000 138.060000 -0.117000 138.130000 ;
      RECT -0.145000 138.060000 -0.117000 138.130000 ;
      RECT -0.145000 138.158000  0.940000 139.015000 ;
      RECT -0.145000 139.015000  0.940000 139.085000 ;
      RECT -0.145000 139.085000  1.010000 139.155000 ;
      RECT -0.145000 139.155000  1.080000 139.225000 ;
      RECT -0.145000 139.225000  1.150000 139.295000 ;
      RECT -0.145000 139.295000  1.220000 139.365000 ;
      RECT -0.145000 139.365000  1.290000 139.435000 ;
      RECT -0.145000 139.435000  1.360000 139.505000 ;
      RECT -0.145000 139.505000 11.105000 139.540000 ;
      RECT -0.145000 139.540000 11.140000 139.575000 ;
      RECT -0.145000 139.575000 69.715000 139.645000 ;
      RECT -0.145000 139.645000 69.785000 139.715000 ;
      RECT -0.145000 139.715000 69.855000 139.785000 ;
      RECT -0.145000 139.785000 69.925000 139.850000 ;
      RECT -0.145000 139.850000  1.385000 139.920000 ;
      RECT -0.145000 139.920000  1.315000 139.990000 ;
      RECT -0.145000 139.990000  1.245000 140.060000 ;
      RECT -0.145000 140.060000  1.175000 140.130000 ;
      RECT -0.145000 140.130000  1.105000 140.200000 ;
      RECT -0.145000 140.200000  1.035000 140.270000 ;
      RECT -0.145000 140.270000  0.965000 140.340000 ;
      RECT -0.145000 140.340000  0.940000 140.365000 ;
      RECT -0.145000 140.365000  0.940000 143.640000 ;
      RECT -0.145000 143.640000  0.940000 143.710000 ;
      RECT -0.145000 143.710000  1.010000 143.780000 ;
      RECT -0.145000 143.780000  1.080000 143.850000 ;
      RECT -0.145000 143.850000  1.150000 143.920000 ;
      RECT -0.145000 143.920000  1.220000 143.990000 ;
      RECT -0.145000 143.990000  1.290000 144.060000 ;
      RECT -0.145000 144.060000  1.360000 144.130000 ;
      RECT -0.145000 144.130000  1.430000 144.200000 ;
      RECT -0.145000 144.200000  1.500000 144.270000 ;
      RECT -0.145000 144.270000  1.570000 144.340000 ;
      RECT -0.145000 144.340000  1.640000 144.410000 ;
      RECT -0.145000 144.410000  1.710000 144.480000 ;
      RECT -0.145000 144.480000  1.780000 144.550000 ;
      RECT -0.145000 144.550000  1.850000 144.620000 ;
      RECT -0.145000 144.620000  1.920000 144.690000 ;
      RECT -0.145000 144.690000  1.990000 144.760000 ;
      RECT -0.145000 144.760000  2.060000 144.830000 ;
      RECT -0.145000 144.830000  2.130000 144.900000 ;
      RECT -0.145000 144.900000  2.200000 144.970000 ;
      RECT -0.145000 144.970000  2.270000 145.040000 ;
      RECT -0.145000 145.040000  2.340000 145.110000 ;
      RECT -0.145000 145.110000  2.410000 145.130000 ;
      RECT -0.127000  96.525000  3.310000  96.545000 ;
      RECT -0.127000  96.525000  3.310000  96.545000 ;
      RECT -0.117000 138.130000  0.940000 138.160000 ;
      RECT -0.057000  96.455000  3.240000  96.525000 ;
      RECT -0.057000  96.455000  3.240000  96.525000 ;
      RECT -0.047000 138.060000  0.940000 138.130000 ;
      RECT  0.000000   0.000000  0.705000  84.591000 ;
      RECT  0.000000   0.000000 12.145000   6.437000 ;
      RECT  0.000000   6.437000 11.777000   6.805000 ;
      RECT  0.000000   6.805000 12.230000   6.983000 ;
      RECT  0.000000   6.983000 12.555000   7.308000 ;
      RECT  0.000000   7.308000 12.555000  10.370000 ;
      RECT  0.000000  10.370000 12.660000  10.445000 ;
      RECT  0.000000  10.445000 14.415000  12.398000 ;
      RECT  0.000000  12.398000 18.077000  16.060000 ;
      RECT  0.000000  16.060000 24.085000  18.668000 ;
      RECT  0.000000  18.668000 24.085000  25.413000 ;
      RECT  0.000000  25.413000 24.675000  26.003000 ;
      RECT  0.000000  26.003000 24.675000  42.682000 ;
      RECT  0.000000  42.682000 24.212000  43.145000 ;
      RECT  0.000000  43.145000  5.925000  43.685000 ;
      RECT  0.000000  43.685000 75.000000 200.000000 ;
      RECT  0.000000  84.591000  0.705000  84.660000 ;
      RECT  0.000000  84.660000  0.774000  84.730000 ;
      RECT  0.000000  84.730000  0.844000  84.800000 ;
      RECT  0.000000  84.800000  0.914000  84.825000 ;
      RECT  0.000000  84.826000  0.940000  95.064000 ;
      RECT  0.000000  95.064000  0.869000  95.135000 ;
      RECT  0.000000  95.135000  0.799000  95.205000 ;
      RECT  0.000000  95.205000  0.729000  95.275000 ;
      RECT  0.000000  95.275000  0.659000  95.345000 ;
      RECT  0.000000  95.345000  0.589000  95.415000 ;
      RECT  0.000000  95.415000  0.519000  95.485000 ;
      RECT  0.000000  95.485000  0.449000  95.555000 ;
      RECT  0.000000  95.555000  0.389000  95.615000 ;
      RECT  0.000000 101.700000 73.490000 104.845000 ;
      RECT  0.000000 104.845000 74.035000 125.160000 ;
      RECT  0.000000 130.500000 10.016000 130.570000 ;
      RECT  0.000000 130.570000  9.946000 130.640000 ;
      RECT  0.000000 130.640000  9.876000 130.710000 ;
      RECT  0.000000 130.710000  9.806000 130.780000 ;
      RECT  0.000000 130.780000  9.736000 130.850000 ;
      RECT  0.000000 130.850000  9.666000 130.920000 ;
      RECT  0.000000 130.920000  9.596000 130.990000 ;
      RECT  0.000000 130.990000  9.591000 130.995000 ;
      RECT  0.000000 145.410000  2.595000 146.420000 ;
      RECT  0.000000 146.420000 59.500000 199.490000 ;
      RECT  0.000000 146.420000 70.525000 146.425000 ;
      RECT  0.000000 146.420000 70.525000 195.970000 ;
      RECT  0.000000 146.425000 73.405000 195.970000 ;
      RECT  0.000000 146.425000 75.000000 174.220000 ;
      RECT  0.000000 174.220000 73.405000 175.420000 ;
      RECT  0.000000 175.420000 75.000000 195.970000 ;
      RECT  0.000000 195.970000 59.500000 199.490000 ;
      RECT  0.000000 199.490000 59.500000 200.000000 ;
      RECT  0.014000  96.385000  3.170000  96.455000 ;
      RECT  0.014000  96.385000  3.170000  96.455000 ;
      RECT  0.023000 137.990000  0.940000 138.060000 ;
      RECT  0.084000  96.315000  3.100000  96.385000 ;
      RECT  0.084000  96.315000  3.100000  96.385000 ;
      RECT  0.094000 137.920000  0.940000 137.990000 ;
      RECT  0.154000  96.245000  3.030000  96.315000 ;
      RECT  0.154000  96.245000  3.030000  96.315000 ;
      RECT  0.164000 137.850000  0.940000 137.920000 ;
      RECT  0.225000  96.175000  2.960000  96.245000 ;
      RECT  0.225000  96.175000  2.960000  96.245000 ;
      RECT  0.234000 137.780000  0.940000 137.850000 ;
      RECT  0.295000  96.105000  2.890000  96.175000 ;
      RECT  0.295000  96.105000  2.890000  96.175000 ;
      RECT  0.304000 137.710000  0.940000 137.780000 ;
      RECT  0.365000  96.035000  2.820000  96.105000 ;
      RECT  0.365000  96.035000  2.820000  96.105000 ;
      RECT  0.374000 137.640000  0.940000 137.710000 ;
      RECT  0.436000  95.965000  2.750000  96.035000 ;
      RECT  0.436000  95.965000  2.750000  96.035000 ;
      RECT  0.445000 137.570000  0.940000 137.640000 ;
      RECT  0.506000  95.895000  2.680000  95.965000 ;
      RECT  0.506000  95.895000  2.680000  95.965000 ;
      RECT  0.515000 137.500000  0.940000 137.570000 ;
      RECT  0.520000  95.880000  2.665000  95.895000 ;
      RECT  0.521000  95.880000  2.665000  95.895000 ;
      RECT  0.521000  95.880000  2.665000  95.895000 ;
      RECT  0.535000  95.865000  2.650000  95.880000 ;
      RECT  0.536000  95.865000  2.650000  95.880000 ;
      RECT  0.536000  95.865000  2.650000  95.880000 ;
      RECT  0.585000 137.430000  0.940000 137.500000 ;
      RECT  0.590000  95.810000  2.650000  95.865000 ;
      RECT  0.591000  95.810000  2.595000  95.865000 ;
      RECT  0.591000  95.810000  2.595000  95.865000 ;
      RECT  0.655000 137.360000  0.940000 137.430000 ;
      RECT  0.660000  95.740000  2.650000  95.810000 ;
      RECT  0.662000  95.740000  2.525000  95.810000 ;
      RECT  0.662000  95.740000  2.525000  95.810000 ;
      RECT  0.725000 137.290000  0.940000 137.360000 ;
      RECT  0.730000  95.670000  2.650000  95.740000 ;
      RECT  0.732000  95.670000  2.455000  95.740000 ;
      RECT  0.732000  95.670000  2.455000  95.740000 ;
      RECT  0.796000 137.220000  0.940000 137.290000 ;
      RECT  0.800000  95.600000  2.650000  95.670000 ;
      RECT  0.802000  95.600000  2.385000  95.670000 ;
      RECT  0.802000  95.600000  2.385000  95.670000 ;
      RECT  0.866000 137.150000  0.940000 137.220000 ;
      RECT  0.870000  95.530000  2.650000  95.600000 ;
      RECT  0.872000  95.530000  2.315000  95.600000 ;
      RECT  0.872000  95.530000  2.315000  95.600000 ;
      RECT  0.936000 137.080000  0.940000 137.150000 ;
      RECT  0.940000  95.460000  2.650000  95.530000 ;
      RECT  0.943000  95.460000  2.245000  95.530000 ;
      RECT  0.943000  95.460000  2.245000  95.530000 ;
      RECT  0.985000   0.240000 11.975000   0.590000 ;
      RECT  0.985000   0.590000  3.300000   0.660000 ;
      RECT  0.985000   0.660000  3.230000   0.730000 ;
      RECT  0.985000   0.730000  3.160000   0.800000 ;
      RECT  0.985000   0.800000  3.090000   0.870000 ;
      RECT  0.985000   0.870000  3.020000   0.940000 ;
      RECT  0.985000   0.940000  2.950000   1.010000 ;
      RECT  0.985000   1.010000  2.880000   1.080000 ;
      RECT  0.985000   1.080000  2.810000   1.150000 ;
      RECT  0.985000   1.150000  2.740000   1.220000 ;
      RECT  0.985000   1.220000  2.670000   1.290000 ;
      RECT  0.985000   1.290000  2.600000   1.360000 ;
      RECT  0.985000   1.360000  2.530000   1.430000 ;
      RECT  0.985000   1.430000  2.460000   1.500000 ;
      RECT  0.985000   1.500000  2.415000   1.545000 ;
      RECT  0.985000   1.545000  2.415000   3.150000 ;
      RECT  0.985000   3.150000  2.415000   3.220000 ;
      RECT  0.985000   3.220000  2.485000   3.290000 ;
      RECT  0.985000   3.290000  2.555000   3.360000 ;
      RECT  0.985000   3.360000  2.625000   3.430000 ;
      RECT  0.985000   3.430000  2.695000   3.500000 ;
      RECT  0.985000   3.500000  2.765000   3.570000 ;
      RECT  0.985000   3.570000  2.835000   3.640000 ;
      RECT  0.985000   3.640000  2.905000   3.710000 ;
      RECT  0.985000   3.710000  2.975000   3.780000 ;
      RECT  0.985000   3.780000  3.045000   3.850000 ;
      RECT  0.985000   3.850000  3.115000   3.920000 ;
      RECT  0.985000   3.920000  3.185000   3.990000 ;
      RECT  0.985000   3.990000  3.255000   4.060000 ;
      RECT  0.985000   4.060000  3.325000   4.105000 ;
      RECT  0.985000   4.105000  4.515000  71.340000 ;
      RECT  0.985000  71.910000 19.260000  79.760000 ;
      RECT  0.985000  80.435000 30.155000  84.475000 ;
      RECT  1.010000  95.390000  2.650000  95.460000 ;
      RECT  1.013000  95.390000  2.175000  95.460000 ;
      RECT  1.013000  95.390000  2.175000  95.460000 ;
      RECT  1.055000  84.475000  3.865000  84.545000 ;
      RECT  1.055000  84.475000  3.865000  84.545000 ;
      RECT  1.080000  95.320000  2.650000  95.390000 ;
      RECT  1.083000  95.320000  2.105000  95.390000 ;
      RECT  1.083000  95.320000  2.105000  95.390000 ;
      RECT  1.125000  84.545000  3.795000  84.615000 ;
      RECT  1.125000  84.545000  3.795000  84.615000 ;
      RECT  1.126000 130.995000 72.380000 131.065000 ;
      RECT  1.150000  95.250000  2.650000  95.320000 ;
      RECT  1.154000  95.250000  2.035000  95.320000 ;
      RECT  1.154000  95.250000  2.035000  95.320000 ;
      RECT  1.195000  84.615000  3.725000  84.685000 ;
      RECT  1.195000  84.615000  3.725000  84.685000 ;
      RECT  1.196000 131.065000 72.380000 131.135000 ;
      RECT  1.220000  81.705000  2.650000  85.760000 ;
      RECT  1.220000  84.685000  3.700000  84.710000 ;
      RECT  1.220000  84.685000  3.700000  84.710000 ;
      RECT  1.220000  84.710000  3.630000  84.780000 ;
      RECT  1.220000  84.780000  3.560000  84.850000 ;
      RECT  1.220000  84.850000  3.490000  84.920000 ;
      RECT  1.220000  84.920000  3.420000  84.990000 ;
      RECT  1.220000  84.990000  3.350000  85.060000 ;
      RECT  1.220000  85.060000  3.280000  85.130000 ;
      RECT  1.220000  85.130000  3.210000  85.200000 ;
      RECT  1.220000  85.200000  3.140000  85.270000 ;
      RECT  1.220000  85.270000  3.070000  85.340000 ;
      RECT  1.220000  85.340000  3.000000  85.410000 ;
      RECT  1.220000  85.410000  2.930000  85.480000 ;
      RECT  1.220000  85.480000  2.860000  85.550000 ;
      RECT  1.220000  85.550000  2.790000  85.620000 ;
      RECT  1.220000  85.620000  2.720000  85.690000 ;
      RECT  1.220000  85.690000  2.650000  85.760000 ;
      RECT  1.220000  85.760000  2.580000  85.830000 ;
      RECT  1.220000  85.760000  2.580000  85.830000 ;
      RECT  1.220000  85.830000  2.510000  85.900000 ;
      RECT  1.220000  85.830000  2.510000  85.900000 ;
      RECT  1.220000  85.900000  2.440000  85.970000 ;
      RECT  1.220000  85.900000  2.440000  85.970000 ;
      RECT  1.220000  85.970000  2.370000  86.040000 ;
      RECT  1.220000  85.970000  2.370000  86.040000 ;
      RECT  1.220000  86.040000  2.300000  86.110000 ;
      RECT  1.220000  86.040000  2.300000  86.110000 ;
      RECT  1.220000  86.110000  2.230000  86.180000 ;
      RECT  1.220000  86.110000  2.230000  86.180000 ;
      RECT  1.220000  86.180000  2.160000  86.250000 ;
      RECT  1.220000  86.180000  2.160000  86.250000 ;
      RECT  1.220000  86.250000  2.090000  86.320000 ;
      RECT  1.220000  86.250000  2.090000  86.320000 ;
      RECT  1.220000  86.320000  2.020000  86.390000 ;
      RECT  1.220000  86.320000  2.020000  86.390000 ;
      RECT  1.220000  86.390000  1.950000  86.460000 ;
      RECT  1.220000  86.390000  1.950000  86.460000 ;
      RECT  1.220000  86.460000  1.880000  86.530000 ;
      RECT  1.220000  86.460000  1.880000  86.530000 ;
      RECT  1.220000  86.530000  1.810000  86.600000 ;
      RECT  1.220000  86.530000  1.810000  86.600000 ;
      RECT  1.220000  86.600000  1.740000  86.670000 ;
      RECT  1.220000  86.600000  1.740000  86.670000 ;
      RECT  1.220000  86.670000  1.670000  86.740000 ;
      RECT  1.220000  86.670000  1.670000  86.740000 ;
      RECT  1.220000  86.740000  1.600000  86.810000 ;
      RECT  1.220000  86.740000  1.600000  86.810000 ;
      RECT  1.220000  86.810000  1.530000  86.880000 ;
      RECT  1.220000  86.810000  1.530000  86.880000 ;
      RECT  1.220000  86.880000  1.460000  86.950000 ;
      RECT  1.220000  86.880000  1.460000  86.950000 ;
      RECT  1.220000  86.950000  1.390000  87.020000 ;
      RECT  1.220000  86.950000  1.390000  87.020000 ;
      RECT  1.220000  87.020000  1.320000  87.090000 ;
      RECT  1.220000  87.020000  1.320000  87.090000 ;
      RECT  1.220000  87.090000  1.250000  87.160000 ;
      RECT  1.220000  87.090000  1.250000  87.160000 ;
      RECT  1.220000  87.190000  2.650000  94.810000 ;
      RECT  1.220000  94.810000  1.525000  94.880000 ;
      RECT  1.220000  94.880000  1.455000  94.950000 ;
      RECT  1.220000  94.950000  1.384000  95.020000 ;
      RECT  1.220000  95.020000  1.314000  95.090000 ;
      RECT  1.220000  95.090000  1.244000  95.160000 ;
      RECT  1.220000  95.160000  1.224000  95.180000 ;
      RECT  1.220000  95.180000  2.650000  95.250000 ;
      RECT  1.220000 135.750000 14.920000 139.225000 ;
      RECT  1.220000 137.196000 70.399000 137.265000 ;
      RECT  1.220000 137.196000 70.399000 137.265000 ;
      RECT  1.220000 137.265000 70.329000 137.335000 ;
      RECT  1.220000 137.265000 70.329000 137.335000 ;
      RECT  1.220000 137.335000 70.259000 137.405000 ;
      RECT  1.220000 137.335000 70.259000 137.405000 ;
      RECT  1.220000 137.405000 70.189000 137.475000 ;
      RECT  1.220000 137.405000 70.189000 137.475000 ;
      RECT  1.220000 137.475000 70.119000 137.545000 ;
      RECT  1.220000 137.475000 70.119000 137.545000 ;
      RECT  1.220000 137.545000 70.049000 137.615000 ;
      RECT  1.220000 137.545000 70.049000 137.615000 ;
      RECT  1.220000 137.615000 69.979000 137.685000 ;
      RECT  1.220000 137.615000 69.979000 137.685000 ;
      RECT  1.220000 137.685000 69.909000 137.755000 ;
      RECT  1.220000 137.685000 69.909000 137.755000 ;
      RECT  1.220000 137.755000 69.839000 137.825000 ;
      RECT  1.220000 137.755000 69.839000 137.825000 ;
      RECT  1.220000 137.825000 69.769000 137.895000 ;
      RECT  1.220000 137.825000 69.769000 137.895000 ;
      RECT  1.220000 137.895000 69.699000 137.965000 ;
      RECT  1.220000 137.895000 69.699000 137.965000 ;
      RECT  1.220000 137.965000 69.629000 138.035000 ;
      RECT  1.220000 137.965000 69.629000 138.035000 ;
      RECT  1.220000 138.035000 69.559000 138.105000 ;
      RECT  1.220000 138.035000 69.559000 138.105000 ;
      RECT  1.220000 138.105000 69.489000 138.175000 ;
      RECT  1.220000 138.105000 69.489000 138.175000 ;
      RECT  1.220000 138.175000 69.419000 138.245000 ;
      RECT  1.220000 138.175000 69.419000 138.245000 ;
      RECT  1.220000 138.245000 69.349000 138.315000 ;
      RECT  1.220000 138.245000 69.349000 138.315000 ;
      RECT  1.220000 138.315000 69.279000 138.385000 ;
      RECT  1.220000 138.315000 69.279000 138.385000 ;
      RECT  1.220000 138.385000 69.209000 138.455000 ;
      RECT  1.220000 138.385000 69.209000 138.455000 ;
      RECT  1.220000 138.455000 69.139000 138.525000 ;
      RECT  1.220000 138.455000 69.139000 138.525000 ;
      RECT  1.220000 138.525000 69.069000 138.595000 ;
      RECT  1.220000 138.525000 69.069000 138.595000 ;
      RECT  1.220000 138.595000 68.999000 138.665000 ;
      RECT  1.220000 138.595000 68.999000 138.665000 ;
      RECT  1.220000 138.665000 16.789000 138.685000 ;
      RECT  1.220000 138.665000 16.789000 138.685000 ;
      RECT  1.220000 138.685000 16.769000 138.705000 ;
      RECT  1.220000 138.685000 16.769000 138.705000 ;
      RECT  1.220000 138.705000 16.764000 138.710000 ;
      RECT  1.220000 138.705000 16.764000 138.710000 ;
      RECT  1.220000 138.710000 14.920000 138.899000 ;
      RECT  1.220000 140.481000 70.225000 140.550000 ;
      RECT  1.220000 140.550000 70.294000 140.620000 ;
      RECT  1.220000 140.620000 70.364000 140.690000 ;
      RECT  1.220000 140.690000 70.434000 140.760000 ;
      RECT  1.220000 140.760000 70.504000 140.780000 ;
      RECT  1.220000 140.781000 70.525000 141.095000 ;
      RECT  1.224000  95.180000  1.965000  95.250000 ;
      RECT  1.224000  95.180000  1.965000  95.250000 ;
      RECT  1.244000  95.160000  1.945000  95.180000 ;
      RECT  1.244000  95.160000  1.945000  95.180000 ;
      RECT  1.266000 131.135000 72.380000 131.205000 ;
      RECT  1.266000 137.150000 70.469000 137.195000 ;
      RECT  1.266000 137.150000 70.469000 137.195000 ;
      RECT  1.291000 138.899000 14.920000 138.970000 ;
      RECT  1.291000 138.899000 14.920000 138.970000 ;
      RECT  1.291000 140.410000 70.154000 140.480000 ;
      RECT  1.314000  95.090000  1.875000  95.160000 ;
      RECT  1.314000  95.090000  1.875000  95.160000 ;
      RECT  1.336000 131.205000 72.380000 131.275000 ;
      RECT  1.336000 137.080000 70.514000 137.150000 ;
      RECT  1.336000 137.080000 70.514000 137.150000 ;
      RECT  1.340000 141.375000 69.645000 143.595000 ;
      RECT  1.361000 138.970000 14.920000 139.040000 ;
      RECT  1.361000 138.970000 14.920000 139.040000 ;
      RECT  1.361000 140.340000 70.084000 140.410000 ;
      RECT  1.384000  95.020000  1.805000  95.090000 ;
      RECT  1.384000  95.020000  1.805000  95.090000 ;
      RECT  1.406000 131.275000 72.380000 131.345000 ;
      RECT  1.406000 137.010000 70.584000 137.080000 ;
      RECT  1.406000 137.010000 70.584000 137.080000 ;
      RECT  1.431000 139.040000 14.920000 139.110000 ;
      RECT  1.431000 139.040000 14.920000 139.110000 ;
      RECT  1.431000 140.270000 70.014000 140.340000 ;
      RECT  1.455000  94.950000  1.735000  95.020000 ;
      RECT  1.455000  94.950000  1.735000  95.020000 ;
      RECT  1.476000 131.345000 72.380000 131.415000 ;
      RECT  1.476000 136.940000 70.654000 137.010000 ;
      RECT  1.476000 136.940000 70.654000 137.010000 ;
      RECT  1.501000 139.110000 14.920000 139.180000 ;
      RECT  1.501000 139.110000 14.920000 139.180000 ;
      RECT  1.501000 140.200000 69.944000 140.270000 ;
      RECT  1.525000  94.880000  1.665000  94.950000 ;
      RECT  1.525000  94.880000  1.665000  94.950000 ;
      RECT  1.546000 131.415000 72.380000 131.485000 ;
      RECT  1.546000 136.870000 70.724000 136.940000 ;
      RECT  1.546000 136.870000 70.724000 136.940000 ;
      RECT  1.546000 139.180000 14.920000 139.225000 ;
      RECT  1.546000 139.180000 14.920000 139.225000 ;
      RECT  1.571000 140.130000 69.874000 140.200000 ;
      RECT  1.616000 131.485000 72.380000 131.555000 ;
      RECT  1.616000 136.800000 70.794000 136.870000 ;
      RECT  1.616000 136.800000 70.794000 136.870000 ;
      RECT  1.641000 143.875000 70.525000 143.945000 ;
      RECT  1.665000  94.810000  2.650000  94.880000 ;
      RECT  1.686000 131.555000 72.380000 131.625000 ;
      RECT  1.686000 136.730000 70.864000 136.800000 ;
      RECT  1.686000 136.730000 70.864000 136.800000 ;
      RECT  1.711000 143.945000 70.525000 144.015000 ;
      RECT  1.735000  94.880000  2.650000  94.950000 ;
      RECT  1.756000 131.625000 72.380000 131.695000 ;
      RECT  1.756000 136.660000 70.934000 136.730000 ;
      RECT  1.756000 136.660000 70.934000 136.730000 ;
      RECT  1.781000 144.015000 70.525000 144.085000 ;
      RECT  1.805000  94.950000  2.650000  95.020000 ;
      RECT  1.826000 131.695000 72.380000 131.765000 ;
      RECT  1.826000 136.590000 71.004000 136.660000 ;
      RECT  1.826000 136.590000 71.004000 136.660000 ;
      RECT  1.851000 144.085000 70.525000 144.155000 ;
      RECT  1.875000  95.020000  2.650000  95.090000 ;
      RECT  1.896000 131.765000 72.380000 131.835000 ;
      RECT  1.896000 136.520000 71.074000 136.590000 ;
      RECT  1.896000 136.520000 71.074000 136.590000 ;
      RECT  1.921000 144.155000 70.525000 144.225000 ;
      RECT  1.945000  95.090000  2.650000  95.160000 ;
      RECT  1.965000  95.160000  2.650000  95.180000 ;
      RECT  1.966000 131.835000 72.380000 131.905000 ;
      RECT  1.966000 136.450000 71.144000 136.520000 ;
      RECT  1.966000 136.450000 71.144000 136.520000 ;
      RECT  1.981000 144.225000 70.525000 144.285000 ;
      RECT  2.036000 131.905000 72.380000 131.975000 ;
      RECT  2.036000 136.380000 71.214000 136.450000 ;
      RECT  2.036000 136.380000 71.214000 136.450000 ;
      RECT  2.051000 144.284000 70.454000 144.355000 ;
      RECT  2.106000 131.975000 72.380000 132.045000 ;
      RECT  2.106000 136.310000 71.284000 136.380000 ;
      RECT  2.106000 136.310000 71.284000 136.380000 ;
      RECT  2.121000 144.355000 70.384000 144.425000 ;
      RECT  2.176000 132.045000 72.380000 132.115000 ;
      RECT  2.176000 136.240000 71.354000 136.310000 ;
      RECT  2.176000 136.240000 71.354000 136.310000 ;
      RECT  2.191000 144.425000 70.314000 144.495000 ;
      RECT  2.246000 132.115000 72.380000 132.185000 ;
      RECT  2.246000 136.170000 71.424000 136.240000 ;
      RECT  2.246000 136.170000 71.424000 136.240000 ;
      RECT  2.261000 144.495000 70.244000 144.565000 ;
      RECT  2.316000 132.185000 72.380000 132.255000 ;
      RECT  2.316000 136.100000 71.494000 136.170000 ;
      RECT  2.316000 136.100000 71.494000 136.170000 ;
      RECT  2.331000 144.565000 70.174000 144.635000 ;
      RECT  2.386000 132.255000 72.380000 132.325000 ;
      RECT  2.386000 136.030000 71.564000 136.100000 ;
      RECT  2.386000 136.030000 71.564000 136.100000 ;
      RECT  2.401000 144.635000 70.104000 144.705000 ;
      RECT  2.456000 132.325000 72.380000 132.395000 ;
      RECT  2.456000 135.960000 71.634000 136.030000 ;
      RECT  2.456000 135.960000 71.634000 136.030000 ;
      RECT  2.471000 144.705000 70.034000 144.775000 ;
      RECT  2.475000 132.740000 13.110000 132.810000 ;
      RECT  2.521000 132.395000 72.380000 132.460000 ;
      RECT  2.526000 135.890000 71.704000 135.960000 ;
      RECT  2.526000 135.890000 71.704000 135.960000 ;
      RECT  2.541000 144.775000 69.964000 144.845000 ;
      RECT  2.545000 132.810000 13.110000 132.880000 ;
      RECT  2.546000 144.845000 69.959000 144.850000 ;
      RECT  2.580000 135.440000 13.110000 135.470000 ;
      RECT  2.596000 135.820000 71.774000 135.890000 ;
      RECT  2.596000 135.820000 71.774000 135.890000 ;
      RECT  2.615000 132.880000 13.110000 132.950000 ;
      RECT  2.650000 135.370000 13.110000 135.440000 ;
      RECT  2.666000 135.750000 71.844000 135.820000 ;
      RECT  2.666000 135.750000 71.844000 135.820000 ;
      RECT  2.685000 132.950000 13.110000 133.020000 ;
      RECT  2.695000   1.661000  3.625000   3.034000 ;
      RECT  2.716000   1.640000  3.625000   1.660000 ;
      RECT  2.720000 135.300000 13.110000 135.370000 ;
      RECT  2.755000 133.020000 13.110000 133.090000 ;
      RECT  2.766000   3.034000  3.625000   3.105000 ;
      RECT  2.786000   1.570000  3.625000   1.640000 ;
      RECT  2.791000 135.230000 13.110000 135.300000 ;
      RECT  2.825000 133.090000 13.110000 133.160000 ;
      RECT  2.836000   3.105000  3.625000   3.175000 ;
      RECT  2.856000   1.500000  3.625000   1.570000 ;
      RECT  2.861000 135.160000 13.110000 135.230000 ;
      RECT  2.875000 145.130000  5.945000 146.140000 ;
      RECT  2.895000 133.160000 13.110000 133.230000 ;
      RECT  2.906000   3.175000  3.625000   3.245000 ;
      RECT  2.926000   1.430000  3.625000   1.500000 ;
      RECT  2.930000  85.876000 71.475000  94.750000 ;
      RECT  2.930000  94.750000 75.000000  95.615000 ;
      RECT  2.930000  95.615000 73.544000  95.680000 ;
      RECT  2.930000  95.680000 73.479000  95.745000 ;
      RECT  2.930000  95.745000 73.474000  95.750000 ;
      RECT  2.931000 135.090000 13.110000 135.160000 ;
      RECT  2.965000 133.230000 13.110000 133.300000 ;
      RECT  2.971000  85.835000 71.475000  85.875000 ;
      RECT  2.971000  85.835000 71.475000  85.875000 ;
      RECT  2.976000   3.245000  3.625000   3.315000 ;
      RECT  2.996000   1.360000  3.625000   1.430000 ;
      RECT  3.001000  95.749000 71.475000  95.820000 ;
      RECT  3.001000  95.749000 71.475000  95.820000 ;
      RECT  3.001000  95.749000 73.404000  95.820000 ;
      RECT  3.001000 135.020000 13.110000 135.090000 ;
      RECT  3.035000 133.300000 13.110000 133.370000 ;
      RECT  3.041000  85.765000 71.475000  85.835000 ;
      RECT  3.041000  85.765000 71.475000  85.835000 ;
      RECT  3.046000   3.315000  3.625000   3.385000 ;
      RECT  3.066000   1.290000  3.625000   1.360000 ;
      RECT  3.071000  95.820000 71.475000  95.890000 ;
      RECT  3.071000  95.820000 71.475000  95.890000 ;
      RECT  3.071000  95.820000 73.334000  95.890000 ;
      RECT  3.071000 134.950000 13.110000 135.020000 ;
      RECT  3.091000   3.385000  3.625000   3.430000 ;
      RECT  3.105000 133.370000 13.110000 133.440000 ;
      RECT  3.111000  85.695000 71.475000  85.765000 ;
      RECT  3.111000  85.695000 71.475000  85.765000 ;
      RECT  3.136000   1.220000  3.625000   1.290000 ;
      RECT  3.141000  95.890000 71.475000  95.960000 ;
      RECT  3.141000  95.890000 71.475000  95.960000 ;
      RECT  3.141000  95.890000 73.264000  95.960000 ;
      RECT  3.141000 134.880000 13.110000 134.950000 ;
      RECT  3.161000   3.430000 12.005000   3.500000 ;
      RECT  3.175000 133.440000 13.110000 133.510000 ;
      RECT  3.181000  85.625000 71.475000  85.695000 ;
      RECT  3.181000  85.625000 71.475000  85.695000 ;
      RECT  3.206000   1.150000  3.625000   1.220000 ;
      RECT  3.211000  95.960000 71.475000  96.030000 ;
      RECT  3.211000  95.960000 71.475000  96.030000 ;
      RECT  3.211000  95.960000 73.194000  96.030000 ;
      RECT  3.212000 134.810000 13.110000 134.880000 ;
      RECT  3.231000   3.500000 12.005000   3.570000 ;
      RECT  3.245000 133.510000 13.110000 133.580000 ;
      RECT  3.251000  85.555000 71.475000  85.625000 ;
      RECT  3.251000  85.555000 71.475000  85.625000 ;
      RECT  3.261000  85.545000 71.475000  85.555000 ;
      RECT  3.261000  85.545000 71.475000  85.555000 ;
      RECT  3.261000  85.545000 75.000000  85.555000 ;
      RECT  3.276000   1.080000  3.625000   1.150000 ;
      RECT  3.281000  96.030000 71.475000  96.100000 ;
      RECT  3.281000  96.030000 71.475000  96.100000 ;
      RECT  3.281000  96.030000 73.124000  96.100000 ;
      RECT  3.282000 134.740000 13.110000 134.810000 ;
      RECT  3.301000   3.570000 12.005000   3.640000 ;
      RECT  3.315000 133.580000 13.110000 133.650000 ;
      RECT  3.331000  85.475000 71.475000  85.545000 ;
      RECT  3.331000  85.475000 71.475000  85.545000 ;
      RECT  3.331000  85.475000 75.000000  85.545000 ;
      RECT  3.346000   1.010000  3.625000   1.080000 ;
      RECT  3.351000  96.100000 71.475000  96.170000 ;
      RECT  3.351000  96.100000 71.475000  96.170000 ;
      RECT  3.351000  96.100000 73.054000  96.170000 ;
      RECT  3.352000 134.670000 13.110000 134.740000 ;
      RECT  3.371000   3.640000 12.005000   3.710000 ;
      RECT  3.385000 133.650000 13.110000 133.720000 ;
      RECT  3.401000  85.405000 71.475000  85.475000 ;
      RECT  3.401000  85.405000 71.475000  85.475000 ;
      RECT  3.401000  85.405000 75.000000  85.475000 ;
      RECT  3.416000   0.940000  3.625000   1.010000 ;
      RECT  3.421000  96.170000 71.475000  96.240000 ;
      RECT  3.421000  96.170000 71.475000  96.240000 ;
      RECT  3.421000  96.170000 72.984000  96.240000 ;
      RECT  3.422000 134.600000 13.110000 134.670000 ;
      RECT  3.441000   3.710000 12.005000   3.780000 ;
      RECT  3.455000 133.720000 13.110000 133.790000 ;
      RECT  3.471000  85.335000 71.475000  85.405000 ;
      RECT  3.471000  85.335000 71.475000  85.405000 ;
      RECT  3.471000  85.335000 75.000000  85.405000 ;
      RECT  3.486000   0.870000  3.625000   0.940000 ;
      RECT  3.486000   3.780000 12.005000   3.825000 ;
      RECT  3.491000  85.315000 33.105000  85.335000 ;
      RECT  3.491000  85.315000 33.105000  85.335000 ;
      RECT  3.491000  96.240000 71.475000  96.310000 ;
      RECT  3.491000  96.240000 71.475000  96.310000 ;
      RECT  3.491000  96.240000 72.914000  96.310000 ;
      RECT  3.492000 134.530000 13.110000 134.600000 ;
      RECT  3.525000 133.790000 13.110000 133.860000 ;
      RECT  3.561000  85.245000 33.105000  85.315000 ;
      RECT  3.561000  85.245000 33.105000  85.315000 ;
      RECT  3.561000  96.310000 71.475000  96.380000 ;
      RECT  3.561000  96.310000 71.475000  96.380000 ;
      RECT  3.561000  96.310000 72.844000  96.380000 ;
      RECT  3.562000 134.460000 13.110000 134.530000 ;
      RECT  3.595000 133.860000 13.110000 133.930000 ;
      RECT  3.631000  85.175000 33.105000  85.245000 ;
      RECT  3.631000  85.175000 33.105000  85.245000 ;
      RECT  3.631000  96.380000 71.475000  96.450000 ;
      RECT  3.631000  96.380000 71.475000  96.450000 ;
      RECT  3.631000  96.380000 72.774000  96.450000 ;
      RECT  3.633000 134.390000 13.110000 134.460000 ;
      RECT  3.665000 133.930000 13.110000 134.000000 ;
      RECT  3.701000  85.105000 33.105000  85.175000 ;
      RECT  3.701000  85.105000 33.105000  85.175000 ;
      RECT  3.701000  96.450000 71.475000  96.520000 ;
      RECT  3.701000  96.450000 71.475000  96.520000 ;
      RECT  3.701000  96.450000 72.704000  96.520000 ;
      RECT  3.703000 134.320000 13.110000 134.390000 ;
      RECT  3.735000 134.000000 13.110000 134.070000 ;
      RECT  3.771000  85.035000 33.105000  85.105000 ;
      RECT  3.771000  85.035000 33.105000  85.105000 ;
      RECT  3.771000  96.520000 71.475000  96.590000 ;
      RECT  3.771000  96.520000 71.475000  96.590000 ;
      RECT  3.771000  96.520000 72.634000  96.590000 ;
      RECT  3.773000 134.250000 13.110000 134.320000 ;
      RECT  3.805000 134.070000 13.110000 134.140000 ;
      RECT  3.841000  84.965000 33.105000  85.035000 ;
      RECT  3.841000  84.965000 33.105000  85.035000 ;
      RECT  3.841000  96.590000 71.475000  96.660000 ;
      RECT  3.841000  96.590000 71.475000  96.660000 ;
      RECT  3.841000  96.590000 72.564000  96.660000 ;
      RECT  3.844000 134.179000 13.110000 134.250000 ;
      RECT  3.845000 134.140000 13.110000 134.180000 ;
      RECT  3.905000   1.140000  5.710000   3.150000 ;
      RECT  3.911000  84.895000 33.105000  84.965000 ;
      RECT  3.911000  84.895000 33.105000  84.965000 ;
      RECT  3.911000  96.660000 71.475000  96.730000 ;
      RECT  3.911000  96.660000 71.475000  96.730000 ;
      RECT  3.911000  96.660000 72.494000  96.730000 ;
      RECT  3.981000  84.825000 33.105000  84.895000 ;
      RECT  3.981000  84.825000 33.105000  84.895000 ;
      RECT  3.981000  96.730000 71.475000  96.800000 ;
      RECT  3.981000  96.730000 71.475000  96.800000 ;
      RECT  3.981000  96.730000 72.424000  96.800000 ;
      RECT  4.051000  84.755000 33.105000  84.825000 ;
      RECT  4.051000  84.755000 33.105000  84.825000 ;
      RECT  4.051000  96.800000 71.475000  96.870000 ;
      RECT  4.051000  96.800000 71.475000  96.870000 ;
      RECT  4.051000  96.800000 72.354000  96.870000 ;
      RECT  4.121000  96.870000 71.475000  96.940000 ;
      RECT  4.121000  96.870000 71.475000  96.940000 ;
      RECT  4.121000  96.870000 72.284000  96.940000 ;
      RECT  4.191000  96.940000 71.475000  97.010000 ;
      RECT  4.191000  96.940000 71.475000  97.010000 ;
      RECT  4.191000  96.940000 72.214000  97.010000 ;
      RECT  4.261000  97.010000 71.475000  97.080000 ;
      RECT  4.261000  97.010000 71.475000  97.080000 ;
      RECT  4.261000  97.010000 72.144000  97.080000 ;
      RECT  4.331000  97.080000 71.475000  97.150000 ;
      RECT  4.331000  97.080000 71.475000  97.150000 ;
      RECT  4.331000  97.080000 72.074000  97.150000 ;
      RECT  4.401000  97.150000 71.475000  97.220000 ;
      RECT  4.401000  97.150000 71.475000  97.220000 ;
      RECT  4.401000  97.150000 72.004000  97.220000 ;
      RECT  4.431000  97.220000 71.475000  97.250000 ;
      RECT  4.431000  97.220000 71.475000  97.250000 ;
      RECT  4.431000  97.220000 71.974000  97.250000 ;
      RECT  4.795000   3.430000 12.005000   3.825000 ;
      RECT  4.795000   3.825000 12.005000   6.379000 ;
      RECT  4.795000   6.379000 11.934000   6.450000 ;
      RECT  4.795000   6.379000 11.934000   6.450000 ;
      RECT  4.795000   6.450000 11.864000   6.520000 ;
      RECT  4.795000   6.450000 11.864000   6.520000 ;
      RECT  4.795000   6.520000 11.794000   6.590000 ;
      RECT  4.795000   6.520000 11.794000   6.590000 ;
      RECT  4.795000   6.590000 11.724000   6.660000 ;
      RECT  4.795000   6.590000 11.724000   6.660000 ;
      RECT  4.795000   6.660000 11.654000   6.730000 ;
      RECT  4.795000   6.660000 11.654000   6.730000 ;
      RECT  4.795000   6.730000 11.584000   6.800000 ;
      RECT  4.795000   6.730000 11.584000   6.800000 ;
      RECT  4.795000   6.800000 11.514000   6.870000 ;
      RECT  4.795000   6.800000 11.514000   6.870000 ;
      RECT  4.795000   6.870000 11.444000   6.940000 ;
      RECT  4.795000   6.870000 11.444000   6.940000 ;
      RECT  4.795000   6.940000 11.439000   6.945000 ;
      RECT  4.795000   6.940000 11.439000   6.945000 ;
      RECT  4.795000   6.945000 12.090000   7.041000 ;
      RECT  4.795000   7.041000 12.090000   7.110000 ;
      RECT  4.795000   7.041000 12.090000   7.110000 ;
      RECT  4.795000   7.110000 12.159000   7.180000 ;
      RECT  4.795000   7.110000 12.159000   7.180000 ;
      RECT  4.795000   7.180000 12.229000   7.250000 ;
      RECT  4.795000   7.180000 12.229000   7.250000 ;
      RECT  4.795000   7.250000 12.299000   7.320000 ;
      RECT  4.795000   7.250000 12.299000   7.320000 ;
      RECT  4.795000   7.320000 12.369000   7.365000 ;
      RECT  4.795000   7.320000 12.369000   7.365000 ;
      RECT  4.795000   7.366000 12.415000  10.510000 ;
      RECT  4.795000   7.366000 12.415000  12.456000 ;
      RECT  4.795000   7.366000 12.415000  12.456000 ;
      RECT  4.795000  10.510000 12.520000  10.585000 ;
      RECT  4.795000  10.585000 14.275000  12.456000 ;
      RECT  4.795000  10.585000 14.275000  16.200000 ;
      RECT  4.795000  12.456000 14.275000  12.525000 ;
      RECT  4.795000  12.456000 14.275000  12.525000 ;
      RECT  4.795000  12.525000 14.344000  12.595000 ;
      RECT  4.795000  12.525000 14.344000  12.595000 ;
      RECT  4.795000  12.595000 14.414000  12.665000 ;
      RECT  4.795000  12.595000 14.414000  12.665000 ;
      RECT  4.795000  12.665000 14.484000  12.735000 ;
      RECT  4.795000  12.665000 14.484000  12.735000 ;
      RECT  4.795000  12.735000 14.554000  12.805000 ;
      RECT  4.795000  12.735000 14.554000  12.805000 ;
      RECT  4.795000  12.805000 14.624000  12.875000 ;
      RECT  4.795000  12.805000 14.624000  12.875000 ;
      RECT  4.795000  12.875000 14.694000  12.945000 ;
      RECT  4.795000  12.875000 14.694000  12.945000 ;
      RECT  4.795000  12.945000 14.764000  13.015000 ;
      RECT  4.795000  12.945000 14.764000  13.015000 ;
      RECT  4.795000  13.015000 14.834000  13.085000 ;
      RECT  4.795000  13.015000 14.834000  13.085000 ;
      RECT  4.795000  13.085000 14.904000  13.155000 ;
      RECT  4.795000  13.085000 14.904000  13.155000 ;
      RECT  4.795000  13.155000 14.974000  13.225000 ;
      RECT  4.795000  13.155000 14.974000  13.225000 ;
      RECT  4.795000  13.225000 15.044000  13.295000 ;
      RECT  4.795000  13.225000 15.044000  13.295000 ;
      RECT  4.795000  13.295000 15.114000  13.365000 ;
      RECT  4.795000  13.295000 15.114000  13.365000 ;
      RECT  4.795000  13.365000 15.184000  13.435000 ;
      RECT  4.795000  13.365000 15.184000  13.435000 ;
      RECT  4.795000  13.435000 15.254000  13.505000 ;
      RECT  4.795000  13.435000 15.254000  13.505000 ;
      RECT  4.795000  13.505000 15.324000  13.575000 ;
      RECT  4.795000  13.505000 15.324000  13.575000 ;
      RECT  4.795000  13.575000 15.394000  13.645000 ;
      RECT  4.795000  13.575000 15.394000  13.645000 ;
      RECT  4.795000  13.645000 15.464000  13.715000 ;
      RECT  4.795000  13.645000 15.464000  13.715000 ;
      RECT  4.795000  13.715000 15.534000  13.785000 ;
      RECT  4.795000  13.715000 15.534000  13.785000 ;
      RECT  4.795000  13.785000 15.604000  13.855000 ;
      RECT  4.795000  13.785000 15.604000  13.855000 ;
      RECT  4.795000  13.855000 15.674000  13.925000 ;
      RECT  4.795000  13.855000 15.674000  13.925000 ;
      RECT  4.795000  13.925000 15.744000  13.995000 ;
      RECT  4.795000  13.925000 15.744000  13.995000 ;
      RECT  4.795000  13.995000 15.814000  14.065000 ;
      RECT  4.795000  13.995000 15.814000  14.065000 ;
      RECT  4.795000  14.065000 15.884000  14.135000 ;
      RECT  4.795000  14.065000 15.884000  14.135000 ;
      RECT  4.795000  14.135000 15.954000  14.205000 ;
      RECT  4.795000  14.135000 15.954000  14.205000 ;
      RECT  4.795000  14.205000 16.024000  14.275000 ;
      RECT  4.795000  14.205000 16.024000  14.275000 ;
      RECT  4.795000  14.275000 16.094000  14.345000 ;
      RECT  4.795000  14.275000 16.094000  14.345000 ;
      RECT  4.795000  14.345000 16.164000  14.415000 ;
      RECT  4.795000  14.345000 16.164000  14.415000 ;
      RECT  4.795000  14.415000 16.234000  14.485000 ;
      RECT  4.795000  14.415000 16.234000  14.485000 ;
      RECT  4.795000  14.485000 16.304000  14.555000 ;
      RECT  4.795000  14.485000 16.304000  14.555000 ;
      RECT  4.795000  14.555000 16.374000  14.625000 ;
      RECT  4.795000  14.555000 16.374000  14.625000 ;
      RECT  4.795000  14.625000 16.444000  14.695000 ;
      RECT  4.795000  14.625000 16.444000  14.695000 ;
      RECT  4.795000  14.695000 16.514000  14.765000 ;
      RECT  4.795000  14.695000 16.514000  14.765000 ;
      RECT  4.795000  14.765000 16.584000  14.835000 ;
      RECT  4.795000  14.765000 16.584000  14.835000 ;
      RECT  4.795000  14.835000 16.654000  14.905000 ;
      RECT  4.795000  14.835000 16.654000  14.905000 ;
      RECT  4.795000  14.905000 16.724000  14.975000 ;
      RECT  4.795000  14.905000 16.724000  14.975000 ;
      RECT  4.795000  14.975000 16.794000  15.045000 ;
      RECT  4.795000  14.975000 16.794000  15.045000 ;
      RECT  4.795000  15.045000 16.864000  15.115000 ;
      RECT  4.795000  15.045000 16.864000  15.115000 ;
      RECT  4.795000  15.115000 16.934000  15.185000 ;
      RECT  4.795000  15.115000 16.934000  15.185000 ;
      RECT  4.795000  15.185000 17.004000  15.255000 ;
      RECT  4.795000  15.185000 17.004000  15.255000 ;
      RECT  4.795000  15.255000 17.074000  15.325000 ;
      RECT  4.795000  15.255000 17.074000  15.325000 ;
      RECT  4.795000  15.325000 17.144000  15.395000 ;
      RECT  4.795000  15.325000 17.144000  15.395000 ;
      RECT  4.795000  15.395000 17.214000  15.465000 ;
      RECT  4.795000  15.395000 17.214000  15.465000 ;
      RECT  4.795000  15.465000 17.284000  15.535000 ;
      RECT  4.795000  15.465000 17.284000  15.535000 ;
      RECT  4.795000  15.535000 17.354000  15.605000 ;
      RECT  4.795000  15.535000 17.354000  15.605000 ;
      RECT  4.795000  15.605000 17.424000  15.675000 ;
      RECT  4.795000  15.605000 17.424000  15.675000 ;
      RECT  4.795000  15.675000 17.494000  15.745000 ;
      RECT  4.795000  15.675000 17.494000  15.745000 ;
      RECT  4.795000  15.745000 17.564000  15.815000 ;
      RECT  4.795000  15.745000 17.564000  15.815000 ;
      RECT  4.795000  15.815000 17.634000  15.885000 ;
      RECT  4.795000  15.815000 17.634000  15.885000 ;
      RECT  4.795000  15.885000 17.704000  15.955000 ;
      RECT  4.795000  15.885000 17.704000  15.955000 ;
      RECT  4.795000  15.955000 17.774000  16.025000 ;
      RECT  4.795000  15.955000 17.774000  16.025000 ;
      RECT  4.795000  16.025000 17.844000  16.095000 ;
      RECT  4.795000  16.025000 17.844000  16.095000 ;
      RECT  4.795000  16.095000 17.914000  16.165000 ;
      RECT  4.795000  16.095000 17.914000  16.165000 ;
      RECT  4.795000  16.165000 17.984000  16.200000 ;
      RECT  4.795000  16.165000 17.984000  16.200000 ;
      RECT  4.795000  16.200000 21.419000  16.270000 ;
      RECT  4.795000  16.200000 21.419000  16.270000 ;
      RECT  4.795000  16.270000 21.489000  16.340000 ;
      RECT  4.795000  16.270000 21.489000  16.340000 ;
      RECT  4.795000  16.340000 21.559000  16.410000 ;
      RECT  4.795000  16.340000 21.559000  16.410000 ;
      RECT  4.795000  16.410000 21.629000  16.480000 ;
      RECT  4.795000  16.410000 21.629000  16.480000 ;
      RECT  4.795000  16.480000 21.699000  16.550000 ;
      RECT  4.795000  16.480000 21.699000  16.550000 ;
      RECT  4.795000  16.550000 21.769000  16.620000 ;
      RECT  4.795000  16.550000 21.769000  16.620000 ;
      RECT  4.795000  16.620000 21.839000  16.690000 ;
      RECT  4.795000  16.620000 21.839000  16.690000 ;
      RECT  4.795000  16.690000 21.909000  16.760000 ;
      RECT  4.795000  16.690000 21.909000  16.760000 ;
      RECT  4.795000  16.760000 21.979000  16.830000 ;
      RECT  4.795000  16.760000 21.979000  16.830000 ;
      RECT  4.795000  16.830000 22.049000  16.900000 ;
      RECT  4.795000  16.830000 22.049000  16.900000 ;
      RECT  4.795000  16.900000 22.119000  16.970000 ;
      RECT  4.795000  16.900000 22.119000  16.970000 ;
      RECT  4.795000  16.970000 22.189000  17.040000 ;
      RECT  4.795000  16.970000 22.189000  17.040000 ;
      RECT  4.795000  17.040000 22.259000  17.110000 ;
      RECT  4.795000  17.040000 22.259000  17.110000 ;
      RECT  4.795000  17.110000 22.329000  17.180000 ;
      RECT  4.795000  17.110000 22.329000  17.180000 ;
      RECT  4.795000  17.180000 22.399000  17.250000 ;
      RECT  4.795000  17.180000 22.399000  17.250000 ;
      RECT  4.795000  17.250000 22.469000  17.320000 ;
      RECT  4.795000  17.250000 22.469000  17.320000 ;
      RECT  4.795000  17.320000 22.539000  17.390000 ;
      RECT  4.795000  17.320000 22.539000  17.390000 ;
      RECT  4.795000  17.390000 22.609000  17.460000 ;
      RECT  4.795000  17.390000 22.609000  17.460000 ;
      RECT  4.795000  17.460000 22.679000  17.530000 ;
      RECT  4.795000  17.460000 22.679000  17.530000 ;
      RECT  4.795000  17.530000 22.749000  17.600000 ;
      RECT  4.795000  17.530000 22.749000  17.600000 ;
      RECT  4.795000  17.600000 22.819000  17.670000 ;
      RECT  4.795000  17.600000 22.819000  17.670000 ;
      RECT  4.795000  17.670000 22.889000  17.740000 ;
      RECT  4.795000  17.670000 22.889000  17.740000 ;
      RECT  4.795000  17.740000 22.959000  17.810000 ;
      RECT  4.795000  17.740000 22.959000  17.810000 ;
      RECT  4.795000  17.810000 23.029000  17.880000 ;
      RECT  4.795000  17.810000 23.029000  17.880000 ;
      RECT  4.795000  17.880000 23.099000  17.950000 ;
      RECT  4.795000  17.880000 23.099000  17.950000 ;
      RECT  4.795000  17.950000 23.169000  18.020000 ;
      RECT  4.795000  17.950000 23.169000  18.020000 ;
      RECT  4.795000  18.020000 23.239000  18.090000 ;
      RECT  4.795000  18.020000 23.239000  18.090000 ;
      RECT  4.795000  18.090000 23.309000  18.160000 ;
      RECT  4.795000  18.090000 23.309000  18.160000 ;
      RECT  4.795000  18.160000 23.379000  18.230000 ;
      RECT  4.795000  18.160000 23.379000  18.230000 ;
      RECT  4.795000  18.230000 23.449000  18.300000 ;
      RECT  4.795000  18.230000 23.449000  18.300000 ;
      RECT  4.795000  18.300000 23.519000  18.370000 ;
      RECT  4.795000  18.300000 23.519000  18.370000 ;
      RECT  4.795000  18.370000 23.589000  18.440000 ;
      RECT  4.795000  18.370000 23.589000  18.440000 ;
      RECT  4.795000  18.440000 23.659000  18.510000 ;
      RECT  4.795000  18.440000 23.659000  18.510000 ;
      RECT  4.795000  18.510000 23.729000  18.580000 ;
      RECT  4.795000  18.510000 23.729000  18.580000 ;
      RECT  4.795000  18.580000 23.799000  18.650000 ;
      RECT  4.795000  18.580000 23.799000  18.650000 ;
      RECT  4.795000  18.650000 23.869000  18.720000 ;
      RECT  4.795000  18.650000 23.869000  18.720000 ;
      RECT  4.795000  18.720000 23.939000  18.725000 ;
      RECT  4.795000  18.720000 23.939000  18.725000 ;
      RECT  4.795000  18.726000 23.945000  25.471000 ;
      RECT  4.795000  18.726000 23.945000  26.061000 ;
      RECT  4.795000  25.471000 23.945000  25.540000 ;
      RECT  4.795000  25.471000 23.945000  25.540000 ;
      RECT  4.795000  25.540000 24.014000  25.610000 ;
      RECT  4.795000  25.540000 24.014000  25.610000 ;
      RECT  4.795000  25.610000 24.084000  25.680000 ;
      RECT  4.795000  25.610000 24.084000  25.680000 ;
      RECT  4.795000  25.680000 24.154000  25.750000 ;
      RECT  4.795000  25.680000 24.154000  25.750000 ;
      RECT  4.795000  25.750000 24.224000  25.820000 ;
      RECT  4.795000  25.750000 24.224000  25.820000 ;
      RECT  4.795000  25.820000 24.294000  25.890000 ;
      RECT  4.795000  25.820000 24.294000  25.890000 ;
      RECT  4.795000  25.890000 24.364000  25.960000 ;
      RECT  4.795000  25.890000 24.364000  25.960000 ;
      RECT  4.795000  25.960000 24.434000  26.030000 ;
      RECT  4.795000  25.960000 24.434000  26.030000 ;
      RECT  4.795000  26.030000 24.504000  26.060000 ;
      RECT  4.795000  26.030000 24.504000  26.060000 ;
      RECT  4.795000  26.061000 24.535000  42.624000 ;
      RECT  4.795000  42.624000 24.464000  42.695000 ;
      RECT  4.795000  42.624000 24.464000  42.695000 ;
      RECT  4.795000  42.695000 24.394000  42.765000 ;
      RECT  4.795000  42.695000 24.394000  42.765000 ;
      RECT  4.795000  42.765000 24.324000  42.835000 ;
      RECT  4.795000  42.765000 24.324000  42.835000 ;
      RECT  4.795000  42.835000 24.254000  42.905000 ;
      RECT  4.795000  42.835000 24.254000  42.905000 ;
      RECT  4.795000  42.905000 24.184000  42.975000 ;
      RECT  4.795000  42.905000 24.184000  42.975000 ;
      RECT  4.795000  42.975000 24.154000  43.005000 ;
      RECT  4.795000  42.975000 24.154000  43.005000 ;
      RECT  4.795000  43.005000  5.785000  43.825000 ;
      RECT  4.795000  43.825000 73.380000  71.630000 ;
      RECT  5.990000   0.870000 12.005000   3.430000 ;
      RECT  6.225000 143.875000 70.525000 144.284000 ;
      RECT  6.225000 144.284000 70.454000 144.355000 ;
      RECT  6.225000 144.284000 70.454000 144.355000 ;
      RECT  6.225000 144.355000 70.384000 144.425000 ;
      RECT  6.225000 144.355000 70.384000 144.425000 ;
      RECT  6.225000 144.425000 70.314000 144.495000 ;
      RECT  6.225000 144.425000 70.314000 144.495000 ;
      RECT  6.225000 144.495000 70.244000 144.565000 ;
      RECT  6.225000 144.495000 70.244000 144.565000 ;
      RECT  6.225000 144.565000 70.174000 144.635000 ;
      RECT  6.225000 144.565000 70.174000 144.635000 ;
      RECT  6.225000 144.635000 70.104000 144.705000 ;
      RECT  6.225000 144.635000 70.104000 144.705000 ;
      RECT  6.225000 144.705000 70.034000 144.775000 ;
      RECT  6.225000 144.705000 70.034000 144.775000 ;
      RECT  6.225000 144.775000 69.964000 144.845000 ;
      RECT  6.225000 144.775000 69.964000 144.845000 ;
      RECT  6.225000 144.845000 69.959000 144.850000 ;
      RECT  6.225000 144.845000 69.959000 144.850000 ;
      RECT  6.225000 144.850000 69.889000 144.920000 ;
      RECT  6.225000 144.850000 69.889000 144.920000 ;
      RECT  6.225000 144.920000 69.819000 144.990000 ;
      RECT  6.225000 144.920000 69.819000 144.990000 ;
      RECT  6.225000 144.990000 69.749000 145.060000 ;
      RECT  6.225000 144.990000 69.749000 145.060000 ;
      RECT  6.225000 145.060000 69.679000 145.130000 ;
      RECT  6.225000 145.060000 69.679000 145.130000 ;
      RECT  6.225000 145.130000 69.609000 145.200000 ;
      RECT  6.225000 145.130000 69.609000 145.200000 ;
      RECT  6.225000 145.200000 69.539000 145.270000 ;
      RECT  6.225000 145.200000 69.539000 145.270000 ;
      RECT  6.225000 145.270000 69.469000 145.340000 ;
      RECT  6.225000 145.270000 69.469000 145.340000 ;
      RECT  6.225000 145.340000 69.399000 145.410000 ;
      RECT  6.225000 145.340000 69.399000 145.410000 ;
      RECT  6.225000 145.410000 70.525000 146.420000 ;
      RECT  6.225000 145.410000 70.525000 195.970000 ;
      RECT  8.191000 132.395000 72.380000 132.460000 ;
      RECT  8.191000 132.395000 72.380000 132.460000 ;
      RECT  8.261000 132.325000 72.380000 132.395000 ;
      RECT  8.261000 132.325000 72.380000 132.395000 ;
      RECT  8.331000 132.255000 72.380000 132.325000 ;
      RECT  8.331000 132.255000 72.380000 132.325000 ;
      RECT  8.401000 132.185000 72.380000 132.255000 ;
      RECT  8.401000 132.185000 72.380000 132.255000 ;
      RECT  8.471000 132.115000 72.380000 132.185000 ;
      RECT  8.471000 132.115000 72.380000 132.185000 ;
      RECT  8.541000 132.045000 72.380000 132.115000 ;
      RECT  8.541000 132.045000 72.380000 132.115000 ;
      RECT  8.611000 131.975000 72.380000 132.045000 ;
      RECT  8.611000 131.975000 72.380000 132.045000 ;
      RECT  8.681000 131.905000 72.380000 131.975000 ;
      RECT  8.681000 131.905000 72.380000 131.975000 ;
      RECT  8.751000 131.835000 72.380000 131.905000 ;
      RECT  8.751000 131.835000 72.380000 131.905000 ;
      RECT  8.821000 131.765000 72.380000 131.835000 ;
      RECT  8.821000 131.765000 72.380000 131.835000 ;
      RECT  8.891000 131.695000 72.380000 131.765000 ;
      RECT  8.891000 131.695000 72.380000 131.765000 ;
      RECT  8.961000 131.625000 72.380000 131.695000 ;
      RECT  8.961000 131.625000 72.380000 131.695000 ;
      RECT  9.031000 131.555000 72.380000 131.625000 ;
      RECT  9.031000 131.555000 72.380000 131.625000 ;
      RECT  9.101000 131.485000 72.380000 131.555000 ;
      RECT  9.101000 131.485000 72.380000 131.555000 ;
      RECT  9.171000 131.415000 72.380000 131.485000 ;
      RECT  9.171000 131.415000 72.380000 131.485000 ;
      RECT  9.241000 131.345000 72.380000 131.415000 ;
      RECT  9.241000 131.345000 72.380000 131.415000 ;
      RECT  9.311000 131.275000 72.380000 131.345000 ;
      RECT  9.311000 131.275000 72.380000 131.345000 ;
      RECT  9.381000 131.205000 72.380000 131.275000 ;
      RECT  9.381000 131.205000 72.380000 131.275000 ;
      RECT  9.451000 131.135000 72.380000 131.205000 ;
      RECT  9.451000 131.135000 72.380000 131.205000 ;
      RECT  9.521000 131.065000 72.380000 131.135000 ;
      RECT  9.521000 131.065000 72.380000 131.135000 ;
      RECT  9.591000 130.995000 72.380000 131.065000 ;
      RECT  9.591000 130.995000 72.380000 131.065000 ;
      RECT  9.596000 130.990000 72.380000 130.995000 ;
      RECT  9.596000 130.990000 72.380000 130.995000 ;
      RECT  9.666000 130.920000 72.380000 130.990000 ;
      RECT  9.666000 130.920000 72.380000 130.990000 ;
      RECT  9.736000 130.850000 72.380000 130.920000 ;
      RECT  9.736000 130.850000 72.380000 130.920000 ;
      RECT  9.806000 130.780000 72.380000 130.850000 ;
      RECT  9.806000 130.780000 72.380000 130.850000 ;
      RECT  9.876000 130.710000 72.380000 130.780000 ;
      RECT  9.876000 130.710000 72.380000 130.780000 ;
      RECT  9.946000 130.640000 72.380000 130.710000 ;
      RECT  9.946000 130.640000 72.380000 130.710000 ;
      RECT 10.016000 130.570000 72.380000 130.640000 ;
      RECT 10.016000 130.570000 72.380000 130.640000 ;
      RECT 10.086000 130.500000 72.380000 130.570000 ;
      RECT 10.086000 130.500000 72.380000 130.570000 ;
      RECT 10.156000 130.430000 64.844000 130.500000 ;
      RECT 10.156000 130.430000 64.844000 130.500000 ;
      RECT 10.226000 130.360000 64.774000 130.430000 ;
      RECT 10.226000 130.360000 64.774000 130.430000 ;
      RECT 10.296000 130.290000 64.704000 130.360000 ;
      RECT 10.296000 130.290000 64.704000 130.360000 ;
      RECT 10.366000 130.220000 64.634000 130.290000 ;
      RECT 10.366000 130.220000 64.634000 130.290000 ;
      RECT 10.436000 130.150000 64.564000 130.220000 ;
      RECT 10.436000 130.150000 64.564000 130.220000 ;
      RECT 10.506000 130.080000 64.494000 130.150000 ;
      RECT 10.506000 130.080000 64.494000 130.150000 ;
      RECT 10.576000 130.010000 64.424000 130.080000 ;
      RECT 10.576000 130.010000 64.424000 130.080000 ;
      RECT 10.646000 129.940000 64.354000 130.010000 ;
      RECT 10.646000 129.940000 64.354000 130.010000 ;
      RECT 10.716000 129.870000 64.284000 129.940000 ;
      RECT 10.716000 129.870000 64.284000 129.940000 ;
      RECT 10.786000 129.800000 64.214000 129.870000 ;
      RECT 10.786000 129.800000 64.214000 129.870000 ;
      RECT 10.856000 129.730000 64.144000 129.800000 ;
      RECT 10.856000 129.730000 64.144000 129.800000 ;
      RECT 10.926000 129.660000 64.074000 129.730000 ;
      RECT 10.926000 129.660000 64.074000 129.730000 ;
      RECT 10.996000 129.590000 64.004000 129.660000 ;
      RECT 10.996000 129.590000 64.004000 129.660000 ;
      RECT 11.066000 129.520000 63.934000 129.590000 ;
      RECT 11.066000 129.520000 63.934000 129.590000 ;
      RECT 11.136000 129.450000 63.864000 129.520000 ;
      RECT 11.136000 129.450000 63.864000 129.520000 ;
      RECT 11.206000 129.380000 63.794000 129.450000 ;
      RECT 11.206000 129.380000 63.794000 129.450000 ;
      RECT 11.256000 139.225000 14.920000 139.260000 ;
      RECT 11.256000 139.225000 14.920000 139.260000 ;
      RECT 11.276000 129.310000 63.724000 129.380000 ;
      RECT 11.276000 129.310000 63.724000 129.380000 ;
      RECT 11.291000 139.260000 14.920000 139.295000 ;
      RECT 11.291000 139.260000 14.920000 139.295000 ;
      RECT 11.346000 129.240000 63.654000 129.310000 ;
      RECT 11.346000 129.240000 63.654000 129.310000 ;
      RECT 11.416000 129.170000 63.584000 129.240000 ;
      RECT 11.416000 129.170000 63.584000 129.240000 ;
      RECT 11.486000 129.100000 63.514000 129.170000 ;
      RECT 11.486000 129.100000 63.514000 129.170000 ;
      RECT 11.556000 129.030000 63.444000 129.100000 ;
      RECT 11.556000 129.030000 63.444000 129.100000 ;
      RECT 11.626000 128.960000 63.374000 129.030000 ;
      RECT 11.626000 128.960000 63.374000 129.030000 ;
      RECT 11.696000 128.890000 63.304000 128.960000 ;
      RECT 11.696000 128.890000 63.304000 128.960000 ;
      RECT 11.766000 128.820000 63.234000 128.890000 ;
      RECT 11.766000 128.820000 63.234000 128.890000 ;
      RECT 11.836000 128.750000 63.164000 128.820000 ;
      RECT 11.836000 128.750000 63.164000 128.820000 ;
      RECT 11.906000 128.680000 63.094000 128.750000 ;
      RECT 11.906000 128.680000 63.094000 128.750000 ;
      RECT 11.950000 128.240000 63.050000 128.260000 ;
      RECT 11.976000 128.610000 63.024000 128.680000 ;
      RECT 11.976000 128.610000 63.024000 128.680000 ;
      RECT 12.020000 128.170000 62.980000 128.240000 ;
      RECT 12.046000 128.540000 62.954000 128.610000 ;
      RECT 12.046000 128.540000 62.954000 128.610000 ;
      RECT 12.090000 128.100000 62.910000 128.170000 ;
      RECT 12.160000 128.030000 62.840000 128.100000 ;
      RECT 12.230000 127.960000 62.770000 128.030000 ;
      RECT 12.300000 127.890000 62.700000 127.960000 ;
      RECT 12.370000 127.820000 62.630000 127.890000 ;
      RECT 12.440000 127.750000 62.560000 127.820000 ;
      RECT 12.510000 127.680000 62.490000 127.750000 ;
      RECT 12.580000 127.610000 62.420000 127.680000 ;
      RECT 12.650000 127.540000 62.350000 127.610000 ;
      RECT 12.685000   0.000000 14.415000   6.717000 ;
      RECT 12.685000   6.717000 14.415000   7.072000 ;
      RECT 12.720000 127.470000 62.280000 127.540000 ;
      RECT 12.790000 127.400000 62.210000 127.470000 ;
      RECT 12.825000   3.550000 14.275000   6.659000 ;
      RECT 12.860000 127.330000 62.140000 127.400000 ;
      RECT 12.896000   6.659000 14.275000   6.730000 ;
      RECT 12.920000   0.240000 13.915000   3.270000 ;
      RECT 12.930000 127.260000 62.070000 127.330000 ;
      RECT 12.966000   6.730000 14.275000   6.800000 ;
      RECT 12.971000  10.555000 14.275000  10.585000 ;
      RECT 13.000000 127.190000 62.000000 127.260000 ;
      RECT 13.036000   6.800000 14.275000   6.870000 ;
      RECT 13.040000   7.072000 14.415000  10.288000 ;
      RECT 13.040000  10.288000 14.415000  10.445000 ;
      RECT 13.041000  10.485000 14.275000  10.555000 ;
      RECT 13.070000 127.120000 61.930000 127.190000 ;
      RECT 13.106000   6.870000 14.275000   6.940000 ;
      RECT 13.111000  10.415000 14.275000  10.485000 ;
      RECT 13.140000 127.050000 61.860000 127.120000 ;
      RECT 13.176000   6.940000 14.275000   7.010000 ;
      RECT 13.180000   7.014000 14.275000  10.346000 ;
      RECT 13.180000  10.346000 14.275000  10.415000 ;
      RECT 13.181000   7.010000 14.275000   7.015000 ;
      RECT 13.210000 126.980000 61.790000 127.050000 ;
      RECT 13.280000 126.910000 61.720000 126.980000 ;
      RECT 13.350000 126.840000 61.650000 126.910000 ;
      RECT 13.390000 130.500000 72.380000 135.750000 ;
      RECT 13.390000 132.460000 72.380000 135.284000 ;
      RECT 13.390000 135.284000 72.309000 135.355000 ;
      RECT 13.390000 135.284000 72.309000 135.355000 ;
      RECT 13.390000 135.355000 72.239000 135.425000 ;
      RECT 13.390000 135.355000 72.239000 135.425000 ;
      RECT 13.390000 135.425000 72.169000 135.495000 ;
      RECT 13.390000 135.425000 72.169000 135.495000 ;
      RECT 13.390000 135.495000 72.099000 135.565000 ;
      RECT 13.390000 135.495000 72.099000 135.565000 ;
      RECT 13.390000 135.565000 72.029000 135.635000 ;
      RECT 13.390000 135.565000 72.029000 135.635000 ;
      RECT 13.390000 135.635000 71.959000 135.705000 ;
      RECT 13.390000 135.635000 71.959000 135.705000 ;
      RECT 13.390000 135.705000 71.914000 135.750000 ;
      RECT 13.390000 135.705000 71.914000 135.750000 ;
      RECT 13.420000 126.770000 61.580000 126.840000 ;
      RECT 13.490000 126.700000 61.510000 126.770000 ;
      RECT 13.560000 126.630000 61.440000 126.700000 ;
      RECT 13.630000 126.560000 61.370000 126.630000 ;
      RECT 13.700000 126.490000 61.300000 126.560000 ;
      RECT 13.770000 126.420000 61.230000 126.490000 ;
      RECT 13.840000 126.350000 61.160000 126.420000 ;
      RECT 13.910000 126.280000 61.090000 126.350000 ;
      RECT 13.980000 126.210000 61.020000 126.280000 ;
      RECT 14.050000 126.140000 60.950000 126.210000 ;
      RECT 14.120000 126.070000 60.880000 126.140000 ;
      RECT 14.190000 126.000000 60.810000 126.070000 ;
      RECT 14.260000 125.930000 60.740000 126.000000 ;
      RECT 14.330000 125.860000 60.670000 125.930000 ;
      RECT 14.400000 125.790000 60.600000 125.860000 ;
      RECT 14.470000 125.720000 60.530000 125.790000 ;
      RECT 14.540000 125.650000 60.460000 125.720000 ;
      RECT 14.610000 125.580000 60.390000 125.650000 ;
      RECT 14.680000 125.510000 60.320000 125.580000 ;
      RECT 14.750000 125.440000 60.250000 125.510000 ;
      RECT 15.200000 138.990000 69.130000 139.060000 ;
      RECT 15.200000 139.060000 69.200000 139.130000 ;
      RECT 15.200000 139.130000 69.270000 139.200000 ;
      RECT 15.200000 139.200000 69.340000 139.270000 ;
      RECT 15.200000 139.270000 69.410000 139.340000 ;
      RECT 15.200000 139.340000 69.480000 139.410000 ;
      RECT 15.200000 139.410000 69.550000 139.480000 ;
      RECT 15.200000 139.480000 69.620000 139.550000 ;
      RECT 15.200000 139.550000 69.690000 139.575000 ;
      RECT 15.275000   0.000000 22.220000   1.345000 ;
      RECT 15.275000   1.345000 24.765000  11.280000 ;
      RECT 15.275000  11.280000 16.460000  12.152000 ;
      RECT 15.275000  12.152000 16.460000  12.468000 ;
      RECT 15.415000   0.830000 16.780000   3.430000 ;
      RECT 15.415000   3.430000 24.625000  11.140000 ;
      RECT 15.415000  11.140000 16.320000  12.094000 ;
      RECT 15.486000  12.094000 16.320000  12.165000 ;
      RECT 15.525000   0.200000 21.315000   0.550000 ;
      RECT 15.556000  12.165000 16.320000  12.235000 ;
      RECT 15.591000  12.468000 16.997000  13.005000 ;
      RECT 15.626000  12.235000 16.320000  12.305000 ;
      RECT 15.696000  12.305000 16.320000  12.375000 ;
      RECT 15.766000  12.375000 16.320000  12.445000 ;
      RECT 15.836000  12.445000 16.320000  12.515000 ;
      RECT 15.846000  12.515000 16.320000  12.525000 ;
      RECT 15.916000  12.526000 16.320000  12.595000 ;
      RECT 15.986000  12.595000 16.389000  12.665000 ;
      RECT 16.056000  12.665000 16.459000  12.735000 ;
      RECT 16.126000  12.735000 16.529000  12.805000 ;
      RECT 16.128000  13.005000 25.015000  13.173000 ;
      RECT 16.196000  12.805000 16.599000  12.875000 ;
      RECT 16.266000  12.875000 16.669000  12.945000 ;
      RECT 16.296000  13.173000 25.015000  15.193000 ;
      RECT 16.336000  12.945000 16.739000  13.015000 ;
      RECT 16.406000  13.015000 16.809000  13.085000 ;
      RECT 16.466000  13.085000 16.879000  13.145000 ;
      RECT 16.511000  13.145000 24.789000  13.190000 ;
      RECT 16.551000  13.190000 24.834000  13.230000 ;
      RECT 16.621000  13.231000 24.875000  13.300000 ;
      RECT 16.691000  13.300000 24.875000  13.370000 ;
      RECT 16.761000  13.370000 24.875000  13.440000 ;
      RECT 16.831000  13.440000 24.875000  13.510000 ;
      RECT 16.885000 138.985000 75.145000 138.990000 ;
      RECT 16.901000  13.510000 24.875000  13.580000 ;
      RECT 16.905000 138.965000 75.145000 138.985000 ;
      RECT 16.925000 138.945000 75.145000 138.965000 ;
      RECT 16.970000  11.280000 24.765000  12.252000 ;
      RECT 16.970000  12.252000 24.765000  12.292000 ;
      RECT 16.971000  13.580000 24.875000  13.650000 ;
      RECT 17.010000  12.292000 24.562000  12.495000 ;
      RECT 17.041000  13.650000 24.875000  13.720000 ;
      RECT 17.060000   1.140000 18.910000   3.150000 ;
      RECT 17.110000   3.430000 24.625000  12.194000 ;
      RECT 17.110000  11.140000 24.625000  12.194000 ;
      RECT 17.111000  13.720000 24.875000  13.790000 ;
      RECT 17.131000  12.194000 24.625000  12.215000 ;
      RECT 17.131000  12.194000 24.625000  12.215000 ;
      RECT 17.151000  12.215000 24.625000  12.235000 ;
      RECT 17.151000  12.215000 24.625000  12.235000 ;
      RECT 17.181000  13.790000 24.875000  13.860000 ;
      RECT 17.211000  12.234000 24.564000  12.295000 ;
      RECT 17.211000  12.234000 24.564000  12.295000 ;
      RECT 17.251000  13.860000 24.875000  13.930000 ;
      RECT 17.271000  12.295000 24.504000  12.355000 ;
      RECT 17.271000  12.295000 24.504000  12.355000 ;
      RECT 17.321000  13.930000 24.875000  14.000000 ;
      RECT 17.391000  14.000000 24.875000  14.070000 ;
      RECT 17.461000  14.070000 24.875000  14.140000 ;
      RECT 17.531000  14.140000 24.875000  14.210000 ;
      RECT 17.601000  14.210000 24.875000  14.280000 ;
      RECT 17.671000  14.280000 24.875000  14.350000 ;
      RECT 17.741000  14.350000 24.875000  14.420000 ;
      RECT 17.811000  14.420000 24.875000  14.490000 ;
      RECT 17.881000  14.490000 24.875000  14.560000 ;
      RECT 17.951000  14.560000 24.875000  14.630000 ;
      RECT 18.021000  14.630000 24.875000  14.700000 ;
      RECT 18.091000  14.700000 24.875000  14.770000 ;
      RECT 18.161000  14.770000 24.875000  14.840000 ;
      RECT 18.231000  14.840000 24.875000  14.910000 ;
      RECT 18.301000  14.910000 24.875000  14.980000 ;
      RECT 18.316000  15.193000 25.102000  15.280000 ;
      RECT 18.371000  14.980000 24.875000  15.050000 ;
      RECT 18.441000  15.050000 24.875000  15.120000 ;
      RECT 18.461000  15.120000 24.875000  15.140000 ;
      RECT 18.985000   0.550000 21.315000   0.620000 ;
      RECT 19.055000   0.620000 21.315000   0.690000 ;
      RECT 19.125000   0.690000 21.315000   0.760000 ;
      RECT 19.190000   2.785000 22.899000   2.855000 ;
      RECT 19.190000   2.785000 22.899000   2.855000 ;
      RECT 19.190000   2.855000 22.969000   2.925000 ;
      RECT 19.190000   2.855000 22.969000   2.925000 ;
      RECT 19.190000   2.925000 23.039000   2.995000 ;
      RECT 19.190000   2.925000 23.039000   2.995000 ;
      RECT 19.190000   2.995000 23.109000   3.065000 ;
      RECT 19.190000   2.995000 23.109000   3.065000 ;
      RECT 19.190000   3.065000 23.179000   3.135000 ;
      RECT 19.190000   3.065000 23.179000   3.135000 ;
      RECT 19.190000   3.135000 23.249000   3.205000 ;
      RECT 19.190000   3.135000 23.249000   3.205000 ;
      RECT 19.190000   3.205000 23.319000   3.275000 ;
      RECT 19.190000   3.205000 23.319000   3.275000 ;
      RECT 19.190000   3.275000 23.389000   3.280000 ;
      RECT 19.190000   3.275000 23.389000   3.280000 ;
      RECT 19.190000   3.280000 24.625000   3.430000 ;
      RECT 19.190000   3.280000 24.625000  11.140000 ;
      RECT 19.190000   3.280000 24.625000  11.140000 ;
      RECT 19.195000   0.760000 21.315000   0.830000 ;
      RECT 19.265000   0.830000 21.385000   0.900000 ;
      RECT 19.335000   0.900000 21.455000   0.970000 ;
      RECT 19.405000   0.970000 21.525000   1.040000 ;
      RECT 19.475000   1.040000 21.595000   1.110000 ;
      RECT 19.540000  71.630000 73.380000  80.155000 ;
      RECT 19.545000   1.110000 21.665000   1.180000 ;
      RECT 19.580000   1.180000 21.735000   1.215000 ;
      RECT 19.580000   1.215000 21.770000   1.285000 ;
      RECT 19.580000   1.285000 21.840000   1.355000 ;
      RECT 19.580000   1.355000 21.910000   1.425000 ;
      RECT 19.580000   1.425000 21.980000   1.495000 ;
      RECT 19.580000   1.495000 22.050000   1.565000 ;
      RECT 19.580000   1.565000 22.120000   1.585000 ;
      RECT 19.580000   1.585000 24.585000   2.505000 ;
      RECT 21.595000   0.000000 22.080000   0.644000 ;
      RECT 21.666000   0.644000 22.080000   0.715000 ;
      RECT 21.736000   0.715000 22.080000   0.785000 ;
      RECT 21.803000  15.280000 25.807000  15.985000 ;
      RECT 21.806000   0.785000 22.080000   0.855000 ;
      RECT 21.876000   0.855000 22.080000   0.925000 ;
      RECT 21.916000  15.140000 24.875000  15.195000 ;
      RECT 21.946000   0.925000 22.080000   0.995000 ;
      RECT 21.971000  15.195000 24.875000  15.250000 ;
      RECT 22.016000   0.995000 22.080000   1.065000 ;
      RECT 22.041000  15.251000 24.875000  15.320000 ;
      RECT 22.111000  15.320000 24.944000  15.390000 ;
      RECT 22.181000  15.390000 25.014000  15.460000 ;
      RECT 22.251000  15.460000 25.084000  15.530000 ;
      RECT 22.321000  15.530000 25.154000  15.600000 ;
      RECT 22.391000  15.600000 25.224000  15.670000 ;
      RECT 22.461000  15.670000 25.294000  15.740000 ;
      RECT 22.508000  15.985000 30.665000  16.843000 ;
      RECT 22.531000  15.740000 25.364000  15.810000 ;
      RECT 22.601000  15.810000 25.434000  15.880000 ;
      RECT 22.671000  15.880000 25.504000  15.950000 ;
      RECT 22.741000  15.950000 25.574000  16.020000 ;
      RECT 22.790000   1.560000 24.585000   1.585000 ;
      RECT 22.800000   0.000000 24.765000   1.345000 ;
      RECT 22.811000  16.020000 25.644000  16.090000 ;
      RECT 22.846000  16.090000 25.714000  16.125000 ;
      RECT 22.860000   1.490000 24.585000   1.560000 ;
      RECT 22.916000  16.125000 29.749000  16.195000 ;
      RECT 22.916000  16.125000 29.749000  16.195000 ;
      RECT 22.930000   1.420000 24.585000   1.490000 ;
      RECT 22.940000   0.000000 24.625000   0.390000 ;
      RECT 22.940000   0.390000 23.210000   0.744000 ;
      RECT 22.940000   0.744000 23.139000   0.815000 ;
      RECT 22.940000   0.815000 23.069000   0.885000 ;
      RECT 22.940000   0.885000 22.999000   0.955000 ;
      RECT 22.986000  16.195000 29.819000  16.265000 ;
      RECT 22.986000  16.195000 29.819000  16.265000 ;
      RECT 23.000000   1.350000 24.585000   1.420000 ;
      RECT 23.056000  16.265000 29.889000  16.335000 ;
      RECT 23.056000  16.265000 29.889000  16.335000 ;
      RECT 23.070000   1.280000 24.585000   1.350000 ;
      RECT 23.085000   2.505000 24.585000   2.575000 ;
      RECT 23.126000  16.335000 29.959000  16.405000 ;
      RECT 23.126000  16.335000 29.959000  16.405000 ;
      RECT 23.140000   1.210000 24.585000   1.280000 ;
      RECT 23.155000   2.575000 24.585000   2.645000 ;
      RECT 23.196000  16.405000 30.029000  16.475000 ;
      RECT 23.196000  16.405000 30.029000  16.475000 ;
      RECT 23.210000   1.140000 24.585000   1.210000 ;
      RECT 23.225000   2.645000 24.585000   2.715000 ;
      RECT 23.266000  16.475000 30.099000  16.545000 ;
      RECT 23.266000  16.475000 30.099000  16.545000 ;
      RECT 23.280000   1.070000 24.585000   1.140000 ;
      RECT 23.295000   2.715000 24.585000   2.785000 ;
      RECT 23.336000  16.545000 30.169000  16.615000 ;
      RECT 23.336000  16.545000 30.169000  16.615000 ;
      RECT 23.350000   1.000000 24.585000   1.070000 ;
      RECT 23.365000   2.785000 24.585000   2.855000 ;
      RECT 23.366000  16.843000 30.665000  18.342000 ;
      RECT 23.406000  16.615000 30.239000  16.685000 ;
      RECT 23.406000  16.615000 30.239000  16.685000 ;
      RECT 23.420000   0.930000 24.585000   1.000000 ;
      RECT 23.435000   2.855000 24.585000   2.925000 ;
      RECT 23.476000  16.685000 30.309000  16.755000 ;
      RECT 23.476000  16.685000 30.309000  16.755000 ;
      RECT 23.490000   0.670000 24.585000   0.860000 ;
      RECT 23.490000   0.860000 24.585000   0.930000 ;
      RECT 23.505000   2.925000 24.585000   2.995000 ;
      RECT 23.510000   2.995000 24.585000   3.000000 ;
      RECT 23.546000  16.755000 30.379000  16.825000 ;
      RECT 23.546000  16.755000 30.379000  16.825000 ;
      RECT 23.616000  16.825000 30.449000  16.895000 ;
      RECT 23.616000  16.825000 30.449000  16.895000 ;
      RECT 23.621000  16.895000 30.519000  16.900000 ;
      RECT 23.621000  16.895000 30.519000  16.900000 ;
      RECT 23.691000  16.901000 30.525000  16.970000 ;
      RECT 23.691000  16.901000 30.525000  16.970000 ;
      RECT 23.761000  16.970000 30.525000  17.040000 ;
      RECT 23.761000  16.970000 30.525000  17.040000 ;
      RECT 23.831000  17.040000 30.525000  17.110000 ;
      RECT 23.831000  17.040000 30.525000  17.110000 ;
      RECT 23.901000  17.110000 30.525000  17.180000 ;
      RECT 23.901000  17.110000 30.525000  17.180000 ;
      RECT 23.971000  17.180000 30.525000  17.250000 ;
      RECT 23.971000  17.180000 30.525000  17.250000 ;
      RECT 24.041000  17.250000 30.525000  17.320000 ;
      RECT 24.041000  17.250000 30.525000  17.320000 ;
      RECT 24.111000  17.320000 30.525000  17.390000 ;
      RECT 24.111000  17.320000 30.525000  17.390000 ;
      RECT 24.181000  17.390000 30.525000  17.460000 ;
      RECT 24.181000  17.390000 30.525000  17.460000 ;
      RECT 24.251000  17.460000 30.525000  17.530000 ;
      RECT 24.251000  17.460000 30.525000  17.530000 ;
      RECT 24.321000  17.530000 30.525000  17.600000 ;
      RECT 24.321000  17.530000 30.525000  17.600000 ;
      RECT 24.391000  17.600000 30.525000  17.670000 ;
      RECT 24.391000  17.600000 30.525000  17.670000 ;
      RECT 24.461000  17.670000 30.525000  17.740000 ;
      RECT 24.461000  17.670000 30.525000  17.740000 ;
      RECT 24.531000  17.740000 30.525000  17.810000 ;
      RECT 24.531000  17.740000 30.525000  17.810000 ;
      RECT 24.546000  43.775000 73.380000  43.825000 ;
      RECT 24.546000  43.775000 73.380000  43.825000 ;
      RECT 24.601000  17.810000 30.525000  17.880000 ;
      RECT 24.601000  17.810000 30.525000  17.880000 ;
      RECT 24.616000  43.705000 73.380000  43.775000 ;
      RECT 24.616000  43.705000 73.380000  43.775000 ;
      RECT 24.671000  17.880000 30.525000  17.950000 ;
      RECT 24.671000  17.880000 30.525000  17.950000 ;
      RECT 24.686000  43.635000 73.380000  43.705000 ;
      RECT 24.686000  43.635000 73.380000  43.705000 ;
      RECT 24.741000  17.950000 30.525000  18.020000 ;
      RECT 24.741000  17.950000 30.525000  18.020000 ;
      RECT 24.756000  43.565000 73.380000  43.635000 ;
      RECT 24.756000  43.565000 73.380000  43.635000 ;
      RECT 24.811000  18.020000 30.525000  18.090000 ;
      RECT 24.811000  18.020000 30.525000  18.090000 ;
      RECT 24.826000  43.495000 73.380000  43.565000 ;
      RECT 24.826000  43.495000 73.380000  43.565000 ;
      RECT 24.865000  18.342000 30.665000  19.485000 ;
      RECT 24.865000  19.485000 32.625000  25.087000 ;
      RECT 24.865000  25.087000 32.625000  25.677000 ;
      RECT 24.881000  18.090000 30.525000  18.160000 ;
      RECT 24.881000  18.090000 30.525000  18.160000 ;
      RECT 24.896000  43.425000 73.380000  43.495000 ;
      RECT 24.896000  43.425000 73.380000  43.495000 ;
      RECT 24.951000  18.160000 30.525000  18.230000 ;
      RECT 24.951000  18.160000 30.525000  18.230000 ;
      RECT 24.966000  43.355000 73.380000  43.425000 ;
      RECT 24.966000  43.355000 73.380000  43.425000 ;
      RECT 25.005000  16.901000 30.525000  25.029000 ;
      RECT 25.005000  18.284000 30.525000  19.625000 ;
      RECT 25.005000  19.625000 32.485000  25.029000 ;
      RECT 25.006000  18.230000 30.525000  18.285000 ;
      RECT 25.006000  18.230000 30.525000  18.285000 ;
      RECT 25.036000  43.285000 73.380000  43.355000 ;
      RECT 25.036000  43.285000 73.380000  43.355000 ;
      RECT 25.076000  25.029000 32.485000  25.100000 ;
      RECT 25.076000  25.029000 32.485000  25.100000 ;
      RECT 25.106000  43.215000 73.380000  43.285000 ;
      RECT 25.106000  43.215000 73.380000  43.285000 ;
      RECT 25.146000  25.100000 32.485000  25.170000 ;
      RECT 25.146000  25.100000 32.485000  25.170000 ;
      RECT 25.176000  43.145000 73.380000  43.215000 ;
      RECT 25.176000  43.145000 73.380000  43.215000 ;
      RECT 25.216000  25.170000 32.485000  25.240000 ;
      RECT 25.216000  25.170000 32.485000  25.240000 ;
      RECT 25.246000  43.075000 73.380000  43.145000 ;
      RECT 25.246000  43.075000 73.380000  43.145000 ;
      RECT 25.275000   0.000000 27.440000   3.183000 ;
      RECT 25.275000   3.183000 28.045000   3.788000 ;
      RECT 25.275000   3.788000 28.045000   4.245000 ;
      RECT 25.275000   4.245000 29.312000   4.755000 ;
      RECT 25.275000   4.755000 28.045000   5.685000 ;
      RECT 25.275000   5.685000 32.620000   8.888000 ;
      RECT 25.275000   8.888000 32.625000   8.893000 ;
      RECT 25.275000   8.893000 32.625000  12.417000 ;
      RECT 25.275000  12.417000 32.625000  12.667000 ;
      RECT 25.286000  25.240000 32.485000  25.310000 ;
      RECT 25.286000  25.240000 32.485000  25.310000 ;
      RECT 25.316000  43.005000 73.380000  43.075000 ;
      RECT 25.316000  43.005000 73.380000  43.075000 ;
      RECT 25.356000  25.310000 32.485000  25.380000 ;
      RECT 25.356000  25.310000 32.485000  25.380000 ;
      RECT 25.386000  42.935000 73.380000  43.005000 ;
      RECT 25.386000  42.935000 73.380000  43.005000 ;
      RECT 25.415000   3.515000 27.574000   3.585000 ;
      RECT 25.415000   3.585000 27.644000   3.655000 ;
      RECT 25.415000   3.655000 27.714000   3.725000 ;
      RECT 25.415000   3.725000 27.784000   3.795000 ;
      RECT 25.415000   3.795000 27.854000   3.845000 ;
      RECT 25.415000   3.846000 27.905000   4.385000 ;
      RECT 25.415000   4.385000 29.414000   4.455000 ;
      RECT 25.415000   4.455000 29.344000   4.525000 ;
      RECT 25.415000   4.525000 29.274000   4.595000 ;
      RECT 25.415000   4.595000 29.254000   4.615000 ;
      RECT 25.415000   4.615000 27.905000   5.825000 ;
      RECT 25.415000   5.825000 31.165000   6.800000 ;
      RECT 25.415000   5.825000 31.165000   8.951000 ;
      RECT 25.415000   5.825000 31.165000   8.951000 ;
      RECT 25.415000   5.825000 31.165000   8.951000 ;
      RECT 25.415000   6.800000 32.480000   8.946000 ;
      RECT 25.415000   8.946000 32.480000   8.950000 ;
      RECT 25.415000   8.946000 32.480000   8.950000 ;
      RECT 25.415000   8.951000 32.485000  12.359000 ;
      RECT 25.426000  25.380000 32.485000  25.450000 ;
      RECT 25.426000  25.380000 32.485000  25.450000 ;
      RECT 25.455000  25.677000 32.625000  28.072000 ;
      RECT 25.455000  28.072000 32.487000  28.210000 ;
      RECT 25.455000  28.210000 28.495000  28.482000 ;
      RECT 25.455000  28.482000 28.495000  32.575000 ;
      RECT 25.455000  32.575000 75.000000  42.668000 ;
      RECT 25.455000  42.668000 75.000000  43.685000 ;
      RECT 25.456000  42.865000 73.380000  42.935000 ;
      RECT 25.456000  42.865000 73.380000  42.935000 ;
      RECT 25.486000  12.359000 32.485000  12.430000 ;
      RECT 25.486000  12.359000 32.485000  12.430000 ;
      RECT 25.496000  25.450000 32.485000  25.520000 ;
      RECT 25.496000  25.450000 32.485000  25.520000 ;
      RECT 25.525000  12.667000 32.625000  14.977000 ;
      RECT 25.525000  14.977000 32.625000  15.475000 ;
      RECT 25.526000  42.795000 73.380000  42.865000 ;
      RECT 25.526000  42.795000 73.380000  42.865000 ;
      RECT 25.556000  12.430000 32.485000  12.500000 ;
      RECT 25.556000  12.430000 32.485000  12.500000 ;
      RECT 25.560000   0.185000 27.265000   3.235000 ;
      RECT 25.566000  25.520000 32.485000  25.590000 ;
      RECT 25.566000  25.520000 32.485000  25.590000 ;
      RECT 25.595000  25.619000 32.485000  28.014000 ;
      RECT 25.595000  28.014000 32.459000  28.040000 ;
      RECT 25.595000  28.014000 32.459000  28.040000 ;
      RECT 25.595000  28.040000 32.429000  28.070000 ;
      RECT 25.595000  28.040000 32.429000  28.070000 ;
      RECT 25.595000  28.070000 28.639000  28.140000 ;
      RECT 25.595000  28.070000 28.639000  28.140000 ;
      RECT 25.595000  28.140000 28.569000  28.210000 ;
      RECT 25.595000  28.140000 28.569000  28.210000 ;
      RECT 25.595000  28.210000 28.499000  28.280000 ;
      RECT 25.595000  28.210000 28.499000  28.280000 ;
      RECT 25.595000  28.280000 28.429000  28.350000 ;
      RECT 25.595000  28.280000 28.429000  28.350000 ;
      RECT 25.595000  28.350000 28.359000  28.420000 ;
      RECT 25.595000  28.350000 28.359000  28.420000 ;
      RECT 25.595000  28.420000 28.354000  28.425000 ;
      RECT 25.595000  28.420000 28.354000  28.425000 ;
      RECT 25.595000  28.424000 28.355000  32.715000 ;
      RECT 25.595000  32.715000 73.380000  42.726000 ;
      RECT 25.595000  42.726000 73.380000  42.795000 ;
      RECT 25.595000  42.726000 73.380000  42.795000 ;
      RECT 25.596000  25.590000 32.485000  25.620000 ;
      RECT 25.596000  25.590000 32.485000  25.620000 ;
      RECT 25.626000  12.500000 32.485000  12.570000 ;
      RECT 25.626000  12.500000 32.485000  12.570000 ;
      RECT 25.665000  12.609000 32.485000  14.919000 ;
      RECT 25.666000  12.570000 32.485000  12.610000 ;
      RECT 25.666000  12.570000 32.485000  12.610000 ;
      RECT 25.736000  14.919000 32.485000  14.990000 ;
      RECT 25.736000  14.919000 32.485000  14.990000 ;
      RECT 25.806000  14.990000 32.485000  15.060000 ;
      RECT 25.806000  14.990000 32.485000  15.060000 ;
      RECT 25.876000  15.060000 32.485000  15.130000 ;
      RECT 25.876000  15.060000 32.485000  15.130000 ;
      RECT 25.946000  15.130000 32.485000  15.200000 ;
      RECT 25.946000  15.130000 32.485000  15.200000 ;
      RECT 26.016000  15.200000 32.485000  15.270000 ;
      RECT 26.016000  15.200000 32.485000  15.270000 ;
      RECT 26.081000  15.270000 32.485000  15.335000 ;
      RECT 26.081000  15.270000 32.485000  15.335000 ;
      RECT 28.370000   0.000000 30.365000   2.797000 ;
      RECT 28.370000   2.797000 30.365000   3.402000 ;
      RECT 28.500000   0.185000 30.205000   2.395000 ;
      RECT 28.516000   2.675000 30.225000   2.745000 ;
      RECT 28.586000   2.745000 30.225000   2.815000 ;
      RECT 28.656000   2.815000 30.225000   2.885000 ;
      RECT 28.726000   2.885000 30.225000   2.955000 ;
      RECT 28.796000   2.955000 30.225000   3.025000 ;
      RECT 28.866000   3.025000 30.225000   3.095000 ;
      RECT 28.936000   3.095000 30.225000   3.165000 ;
      RECT 28.975000   3.402000 30.365000   3.702000 ;
      RECT 28.975000   3.702000 29.822000   4.245000 ;
      RECT 29.005000  28.793000 75.000000  32.575000 ;
      RECT 29.006000   3.165000 30.225000   3.235000 ;
      RECT 29.076000   3.235000 30.225000   3.305000 ;
      RECT 29.078000  28.720000 75.000000  28.793000 ;
      RECT 29.115000   3.344000 30.225000   3.644000 ;
      RECT 29.115000   3.644000 30.154000   3.715000 ;
      RECT 29.115000   3.715000 30.084000   3.785000 ;
      RECT 29.115000   3.785000 30.014000   3.855000 ;
      RECT 29.115000   3.855000 29.944000   3.925000 ;
      RECT 29.115000   3.925000 29.874000   3.995000 ;
      RECT 29.115000   3.995000 29.804000   4.065000 ;
      RECT 29.115000   4.065000 29.734000   4.135000 ;
      RECT 29.115000   4.135000 29.664000   4.205000 ;
      RECT 29.115000   4.205000 29.594000   4.275000 ;
      RECT 29.115000   4.275000 29.524000   4.345000 ;
      RECT 29.115000   4.345000 29.484000   4.385000 ;
      RECT 29.116000   3.305000 30.225000   3.345000 ;
      RECT 29.145000  28.860000 73.380000  32.715000 ;
      RECT 29.766000   5.815000 31.165000   5.825000 ;
      RECT 29.836000   5.745000 31.165000   5.815000 ;
      RECT 29.906000   5.675000 31.165000   5.745000 ;
      RECT 29.976000   5.605000 31.165000   5.675000 ;
      RECT 30.023000  15.475000 32.625000  16.627000 ;
      RECT 30.046000   5.535000 31.165000   5.605000 ;
      RECT 30.116000   5.465000 31.165000   5.535000 ;
      RECT 30.151000  15.335000 32.485000  15.405000 ;
      RECT 30.151000  15.335000 32.485000  15.405000 ;
      RECT 30.186000   5.395000 31.165000   5.465000 ;
      RECT 30.221000  15.405000 32.485000  15.475000 ;
      RECT 30.221000  15.405000 32.485000  15.475000 ;
      RECT 30.256000   5.325000 31.165000   5.395000 ;
      RECT 30.291000  15.475000 32.485000  15.545000 ;
      RECT 30.291000  15.475000 32.485000  15.545000 ;
      RECT 30.326000   5.255000 31.165000   5.325000 ;
      RECT 30.361000  15.545000 32.485000  15.615000 ;
      RECT 30.361000  15.545000 32.485000  15.615000 ;
      RECT 30.396000   5.185000 31.165000   5.255000 ;
      RECT 30.431000  15.615000 32.485000  15.685000 ;
      RECT 30.431000  15.615000 32.485000  15.685000 ;
      RECT 30.435000  80.155000 73.380000  84.520000 ;
      RECT 30.435000  84.520000 33.105000  84.755000 ;
      RECT 30.466000   5.115000 31.165000   5.185000 ;
      RECT 30.501000  15.685000 32.485000  15.755000 ;
      RECT 30.501000  15.685000 32.485000  15.755000 ;
      RECT 30.536000   5.045000 31.165000   5.115000 ;
      RECT 30.571000  15.755000 32.485000  15.825000 ;
      RECT 30.571000  15.755000 32.485000  15.825000 ;
      RECT 30.606000   4.975000 31.165000   5.045000 ;
      RECT 30.641000  15.825000 32.485000  15.895000 ;
      RECT 30.641000  15.825000 32.485000  15.895000 ;
      RECT 30.676000   4.905000 31.165000   4.975000 ;
      RECT 30.711000  15.895000 32.485000  15.965000 ;
      RECT 30.711000  15.895000 32.485000  15.965000 ;
      RECT 30.746000   4.835000 31.165000   4.905000 ;
      RECT 30.781000  15.965000 32.485000  16.035000 ;
      RECT 30.781000  15.965000 32.485000  16.035000 ;
      RECT 30.816000   4.765000 31.165000   4.835000 ;
      RECT 30.851000  16.035000 32.485000  16.105000 ;
      RECT 30.851000  16.035000 32.485000  16.105000 ;
      RECT 30.886000   4.695000 31.165000   4.765000 ;
      RECT 30.921000  16.105000 32.485000  16.175000 ;
      RECT 30.921000  16.105000 32.485000  16.175000 ;
      RECT 30.956000   4.625000 31.165000   4.695000 ;
      RECT 30.991000  16.175000 32.485000  16.245000 ;
      RECT 30.991000  16.175000 32.485000  16.245000 ;
      RECT 31.026000   4.555000 31.165000   4.625000 ;
      RECT 31.061000  16.245000 32.485000  16.315000 ;
      RECT 31.061000  16.245000 32.485000  16.315000 ;
      RECT 31.096000   4.485000 31.165000   4.555000 ;
      RECT 31.131000  16.315000 32.485000  16.385000 ;
      RECT 31.131000  16.315000 32.485000  16.385000 ;
      RECT 31.175000  16.627000 32.625000  19.485000 ;
      RECT 31.201000  16.385000 32.485000  16.455000 ;
      RECT 31.201000  16.385000 32.485000  16.455000 ;
      RECT 31.271000  16.455000 32.485000  16.525000 ;
      RECT 31.271000  16.455000 32.485000  16.525000 ;
      RECT 31.295000   0.000000 32.620000   4.088000 ;
      RECT 31.295000   4.088000 32.620000   5.685000 ;
      RECT 31.315000  16.569000 32.485000  19.625000 ;
      RECT 31.316000  16.525000 32.485000  16.570000 ;
      RECT 31.316000  16.525000 32.485000  16.570000 ;
      RECT 31.435000   0.000000 32.480000   0.390000 ;
      RECT 31.445000   0.670000 32.410000   6.520000 ;
      RECT 33.160000   0.000000 75.000000   8.662000 ;
      RECT 33.160000   8.662000 75.000000   8.667000 ;
      RECT 33.165000   8.667000 75.000000  28.720000 ;
      RECT 33.300000   0.000000 75.000000   0.600000 ;
      RECT 33.300000   0.600000 34.820000   0.620000 ;
      RECT 33.300000   0.620000 34.615000   2.160000 ;
      RECT 33.300000   2.160000 39.940000   6.270000 ;
      RECT 33.300000   6.270000 73.109000   6.340000 ;
      RECT 33.300000   6.270000 73.109000   6.340000 ;
      RECT 33.300000   6.340000 73.179000   6.410000 ;
      RECT 33.300000   6.340000 73.179000   6.410000 ;
      RECT 33.300000   6.410000 73.249000   6.480000 ;
      RECT 33.300000   6.410000 73.249000   6.480000 ;
      RECT 33.300000   6.480000 73.319000   6.540000 ;
      RECT 33.300000   6.480000 73.319000   6.540000 ;
      RECT 33.300000   6.541000 73.380000   8.604000 ;
      RECT 33.305000   8.609000 73.380000  28.860000 ;
      RECT 33.305000   8.609000 73.380000  32.715000 ;
      RECT 33.306000   8.604000 73.380000   8.610000 ;
      RECT 33.306000   8.604000 73.380000   8.610000 ;
      RECT 33.385000  84.800000 74.700000  85.055000 ;
      RECT 34.895000   0.900000 38.965000   1.880000 ;
      RECT 35.100000   0.880000 38.920000   0.900000 ;
      RECT 39.200000   0.600000 75.000000   0.620000 ;
      RECT 39.245000   0.620000 75.000000   0.740000 ;
      RECT 39.245000   0.740000 39.940000   2.160000 ;
      RECT 40.220000   1.020000 74.590000   5.990000 ;
      RECT 56.545000 100.330000 72.090000 101.420000 ;
      RECT 56.725000  97.530000 72.090000  97.760000 ;
      RECT 56.825000  98.040000 71.244000  98.110000 ;
      RECT 56.825000  98.110000 71.314000  98.180000 ;
      RECT 56.825000  98.180000 71.384000  98.250000 ;
      RECT 56.825000  98.250000 71.454000  98.320000 ;
      RECT 56.825000  98.320000 71.524000  98.390000 ;
      RECT 56.825000  98.390000 71.594000  98.460000 ;
      RECT 56.825000  98.460000 71.664000  98.530000 ;
      RECT 56.825000  98.530000 71.734000  98.600000 ;
      RECT 56.825000  98.600000 71.804000  98.605000 ;
      RECT 56.825000  98.606000 71.810000  99.404000 ;
      RECT 56.825000  99.404000 71.739000  99.475000 ;
      RECT 56.825000  99.475000 71.669000  99.545000 ;
      RECT 56.825000  99.545000 71.599000  99.615000 ;
      RECT 56.825000  99.615000 71.529000  99.685000 ;
      RECT 56.825000  99.685000 71.459000  99.755000 ;
      RECT 56.825000  99.755000 71.389000  99.825000 ;
      RECT 56.825000  99.825000 71.319000  99.895000 ;
      RECT 56.825000  99.895000 71.249000  99.965000 ;
      RECT 56.825000  99.965000 71.179000 100.035000 ;
      RECT 56.825000 100.035000 71.164000 100.050000 ;
      RECT 59.500000 199.490000 64.600000 200.000000 ;
      RECT 59.780000 196.250000 64.320000 199.210000 ;
      RECT 60.320000 125.440000 75.145000 125.510000 ;
      RECT 60.320000 125.440000 75.145000 125.510000 ;
      RECT 60.390000 125.510000 75.145000 125.580000 ;
      RECT 60.390000 125.510000 75.145000 125.580000 ;
      RECT 60.460000 125.580000 75.145000 125.650000 ;
      RECT 60.460000 125.580000 75.145000 125.650000 ;
      RECT 60.530000 125.650000 75.145000 125.720000 ;
      RECT 60.530000 125.650000 75.145000 125.720000 ;
      RECT 60.600000 125.720000 75.145000 125.790000 ;
      RECT 60.600000 125.720000 75.145000 125.790000 ;
      RECT 60.670000 125.790000 75.145000 125.860000 ;
      RECT 60.670000 125.790000 75.145000 125.860000 ;
      RECT 60.740000 125.860000 75.145000 125.930000 ;
      RECT 60.740000 125.860000 75.145000 125.930000 ;
      RECT 60.810000 125.930000 75.145000 126.000000 ;
      RECT 60.810000 125.930000 75.145000 126.000000 ;
      RECT 60.880000 126.000000 75.145000 126.070000 ;
      RECT 60.880000 126.000000 75.145000 126.070000 ;
      RECT 60.950000 126.070000 75.145000 126.140000 ;
      RECT 60.950000 126.070000 75.145000 126.140000 ;
      RECT 61.020000 126.140000 75.145000 126.210000 ;
      RECT 61.020000 126.140000 75.145000 126.210000 ;
      RECT 61.090000 126.210000 75.145000 126.280000 ;
      RECT 61.090000 126.210000 75.145000 126.280000 ;
      RECT 61.160000 126.280000 75.145000 126.350000 ;
      RECT 61.160000 126.280000 75.145000 126.350000 ;
      RECT 61.230000 126.350000 75.145000 126.420000 ;
      RECT 61.230000 126.350000 75.145000 126.420000 ;
      RECT 61.300000 126.420000 75.145000 126.490000 ;
      RECT 61.300000 126.420000 75.145000 126.490000 ;
      RECT 61.370000 126.490000 75.145000 126.560000 ;
      RECT 61.370000 126.490000 75.145000 126.560000 ;
      RECT 61.440000 126.560000 75.145000 126.630000 ;
      RECT 61.440000 126.560000 75.145000 126.630000 ;
      RECT 61.510000 126.630000 75.145000 126.700000 ;
      RECT 61.510000 126.630000 75.145000 126.700000 ;
      RECT 61.580000 126.700000 75.145000 126.770000 ;
      RECT 61.580000 126.700000 75.145000 126.770000 ;
      RECT 61.650000 126.770000 75.145000 126.840000 ;
      RECT 61.650000 126.770000 75.145000 126.840000 ;
      RECT 61.720000 126.840000 75.145000 126.910000 ;
      RECT 61.720000 126.840000 75.145000 126.910000 ;
      RECT 61.790000 126.910000 75.145000 126.980000 ;
      RECT 61.790000 126.910000 75.145000 126.980000 ;
      RECT 61.860000 126.980000 75.145000 127.050000 ;
      RECT 61.860000 126.980000 75.145000 127.050000 ;
      RECT 61.930000 127.050000 75.145000 127.120000 ;
      RECT 61.930000 127.050000 75.145000 127.120000 ;
      RECT 62.000000 127.120000 75.145000 127.190000 ;
      RECT 62.000000 127.120000 75.145000 127.190000 ;
      RECT 62.070000 127.190000 75.145000 127.260000 ;
      RECT 62.070000 127.190000 75.145000 127.260000 ;
      RECT 62.140000 127.260000 75.145000 127.330000 ;
      RECT 62.140000 127.260000 75.145000 127.330000 ;
      RECT 62.210000 127.330000 75.145000 127.400000 ;
      RECT 62.210000 127.330000 75.145000 127.400000 ;
      RECT 62.280000 127.400000 75.145000 127.470000 ;
      RECT 62.280000 127.400000 75.145000 127.470000 ;
      RECT 62.350000 127.470000 75.145000 127.540000 ;
      RECT 62.350000 127.470000 75.145000 127.540000 ;
      RECT 62.420000 127.540000 75.145000 127.610000 ;
      RECT 62.420000 127.540000 75.145000 127.610000 ;
      RECT 62.490000 127.610000 75.145000 127.680000 ;
      RECT 62.490000 127.610000 75.145000 127.680000 ;
      RECT 62.560000 127.680000 75.145000 127.750000 ;
      RECT 62.560000 127.680000 75.145000 127.750000 ;
      RECT 62.630000 127.750000 75.145000 127.820000 ;
      RECT 62.630000 127.750000 75.145000 127.820000 ;
      RECT 62.700000 127.820000 75.145000 127.890000 ;
      RECT 62.700000 127.820000 75.145000 127.890000 ;
      RECT 62.770000 127.890000 75.145000 127.960000 ;
      RECT 62.770000 127.890000 75.145000 127.960000 ;
      RECT 62.840000 127.960000 75.145000 128.030000 ;
      RECT 62.840000 127.960000 75.145000 128.030000 ;
      RECT 62.910000 128.030000 75.145000 128.100000 ;
      RECT 62.910000 128.030000 75.145000 128.100000 ;
      RECT 62.980000 128.100000 75.145000 128.170000 ;
      RECT 62.980000 128.100000 75.145000 128.170000 ;
      RECT 63.050000 128.170000 75.145000 128.240000 ;
      RECT 63.050000 128.170000 75.145000 128.240000 ;
      RECT 63.070000 128.240000 75.145000 128.260000 ;
      RECT 63.070000 128.240000 75.145000 128.260000 ;
      RECT 63.140000 128.260000 75.145000 128.330000 ;
      RECT 63.140000 128.260000 75.145000 128.330000 ;
      RECT 63.210000 128.330000 75.145000 128.400000 ;
      RECT 63.210000 128.330000 75.145000 128.400000 ;
      RECT 63.280000 128.400000 75.145000 128.470000 ;
      RECT 63.280000 128.400000 75.145000 128.470000 ;
      RECT 63.350000 128.470000 75.145000 128.540000 ;
      RECT 63.350000 128.470000 75.145000 128.540000 ;
      RECT 63.420000 128.540000 75.145000 128.610000 ;
      RECT 63.420000 128.540000 75.145000 128.610000 ;
      RECT 63.490000 128.610000 75.145000 128.680000 ;
      RECT 63.490000 128.610000 75.145000 128.680000 ;
      RECT 63.560000 128.680000 75.145000 128.750000 ;
      RECT 63.560000 128.680000 75.145000 128.750000 ;
      RECT 63.630000 128.750000 75.145000 128.820000 ;
      RECT 63.630000 128.750000 75.145000 128.820000 ;
      RECT 63.700000 128.820000 75.145000 128.890000 ;
      RECT 63.700000 128.820000 75.145000 128.890000 ;
      RECT 63.770000 128.890000 75.145000 128.960000 ;
      RECT 63.770000 128.890000 75.145000 128.960000 ;
      RECT 63.840000 128.960000 75.145000 129.030000 ;
      RECT 63.840000 128.960000 75.145000 129.030000 ;
      RECT 63.910000 129.030000 75.145000 129.100000 ;
      RECT 63.910000 129.030000 75.145000 129.100000 ;
      RECT 63.980000 129.100000 75.145000 129.170000 ;
      RECT 63.980000 129.100000 75.145000 129.170000 ;
      RECT 64.050000 129.170000 75.145000 129.240000 ;
      RECT 64.050000 129.170000 75.145000 129.240000 ;
      RECT 64.120000 129.240000 75.145000 129.310000 ;
      RECT 64.120000 129.240000 75.145000 129.310000 ;
      RECT 64.190000 129.310000 75.145000 129.380000 ;
      RECT 64.190000 129.310000 75.145000 129.380000 ;
      RECT 64.260000 129.380000 75.145000 129.450000 ;
      RECT 64.260000 129.380000 75.145000 129.450000 ;
      RECT 64.330000 129.450000 75.145000 129.520000 ;
      RECT 64.330000 129.450000 75.145000 129.520000 ;
      RECT 64.400000 129.520000 75.145000 129.590000 ;
      RECT 64.400000 129.520000 75.145000 129.590000 ;
      RECT 64.470000 129.590000 75.145000 129.660000 ;
      RECT 64.470000 129.590000 75.145000 129.660000 ;
      RECT 64.540000 129.660000 75.145000 129.730000 ;
      RECT 64.540000 129.660000 75.145000 129.730000 ;
      RECT 64.600000 175.420000 75.000000 200.000000 ;
      RECT 64.600000 195.970000 75.000000 199.490000 ;
      RECT 64.600000 199.490000 75.000000 200.000000 ;
      RECT 64.610000 129.730000 75.145000 129.800000 ;
      RECT 64.610000 129.730000 75.145000 129.800000 ;
      RECT 64.680000 129.800000 75.145000 129.870000 ;
      RECT 64.680000 129.800000 75.145000 129.870000 ;
      RECT 64.750000 129.870000 75.145000 129.940000 ;
      RECT 64.750000 129.870000 75.145000 129.940000 ;
      RECT 64.820000 129.940000 75.145000 130.010000 ;
      RECT 64.820000 129.940000 75.145000 130.010000 ;
      RECT 64.890000 130.010000 75.145000 130.080000 ;
      RECT 64.890000 130.010000 75.145000 130.080000 ;
      RECT 64.960000 130.080000 75.145000 130.150000 ;
      RECT 64.960000 130.080000 75.145000 130.150000 ;
      RECT 65.030000 130.150000 75.145000 130.220000 ;
      RECT 65.030000 130.150000 75.145000 130.220000 ;
      RECT 69.105000 138.955000 75.145000 138.960000 ;
      RECT 69.105000 138.955000 75.145000 138.960000 ;
      RECT 69.110000 138.950000 75.145000 138.955000 ;
      RECT 69.110000 138.950000 75.145000 138.955000 ;
      RECT 69.115000 138.945000 75.145000 138.950000 ;
      RECT 69.115000 138.945000 75.145000 138.950000 ;
      RECT 69.115000 138.960000 75.145000 138.975000 ;
      RECT 69.115000 138.960000 75.145000 138.975000 ;
      RECT 69.130000 138.975000 75.145000 138.990000 ;
      RECT 69.130000 138.975000 75.145000 138.990000 ;
      RECT 69.160000 138.900000 75.145000 138.945000 ;
      RECT 69.160000 138.900000 75.145000 138.945000 ;
      RECT 69.200000 138.990000 75.145000 139.060000 ;
      RECT 69.200000 138.990000 75.145000 139.060000 ;
      RECT 69.230000 138.830000 75.145000 138.900000 ;
      RECT 69.230000 138.830000 75.145000 138.900000 ;
      RECT 69.270000 139.060000 75.145000 139.130000 ;
      RECT 69.270000 139.060000 75.145000 139.130000 ;
      RECT 69.300000 138.760000 75.145000 138.830000 ;
      RECT 69.300000 138.760000 75.145000 138.830000 ;
      RECT 69.340000 139.130000 75.145000 139.200000 ;
      RECT 69.340000 139.130000 75.145000 139.200000 ;
      RECT 69.370000 138.690000 75.145000 138.760000 ;
      RECT 69.370000 138.690000 75.145000 138.760000 ;
      RECT 69.410000 139.200000 75.145000 139.270000 ;
      RECT 69.410000 139.200000 75.145000 139.270000 ;
      RECT 69.440000 138.620000 75.145000 138.690000 ;
      RECT 69.440000 138.620000 75.145000 138.690000 ;
      RECT 69.480000 139.270000 75.145000 139.340000 ;
      RECT 69.480000 139.270000 75.145000 139.340000 ;
      RECT 69.510000 138.550000 75.145000 138.620000 ;
      RECT 69.510000 138.550000 75.145000 138.620000 ;
      RECT 69.550000 139.340000 75.145000 139.410000 ;
      RECT 69.550000 139.340000 75.145000 139.410000 ;
      RECT 69.580000 138.480000 75.145000 138.550000 ;
      RECT 69.580000 138.480000 75.145000 138.550000 ;
      RECT 69.620000 139.410000 75.145000 139.480000 ;
      RECT 69.620000 139.410000 75.145000 139.480000 ;
      RECT 69.650000 138.410000 75.145000 138.480000 ;
      RECT 69.650000 138.410000 75.145000 138.480000 ;
      RECT 69.690000 139.480000 75.145000 139.550000 ;
      RECT 69.690000 139.480000 75.145000 139.550000 ;
      RECT 69.715000 139.550000 75.145000 139.575000 ;
      RECT 69.715000 139.550000 75.145000 139.575000 ;
      RECT 69.720000 138.340000 75.145000 138.410000 ;
      RECT 69.720000 138.340000 75.145000 138.410000 ;
      RECT 69.785000 139.575000 75.145000 139.645000 ;
      RECT 69.785000 139.575000 75.145000 139.645000 ;
      RECT 69.790000 138.270000 75.145000 138.340000 ;
      RECT 69.790000 138.270000 75.145000 138.340000 ;
      RECT 69.855000 139.645000 75.145000 139.715000 ;
      RECT 69.855000 139.645000 75.145000 139.715000 ;
      RECT 69.860000 138.200000 75.145000 138.270000 ;
      RECT 69.860000 138.200000 75.145000 138.270000 ;
      RECT 69.925000 139.715000 75.145000 139.785000 ;
      RECT 69.925000 139.715000 75.145000 139.785000 ;
      RECT 69.925000 141.095000 70.525000 143.875000 ;
      RECT 69.930000 138.130000 75.145000 138.200000 ;
      RECT 69.930000 138.130000 75.145000 138.200000 ;
      RECT 69.990000 139.785000 75.145000 139.850000 ;
      RECT 69.990000 139.785000 75.145000 139.850000 ;
      RECT 70.000000 138.060000 75.145000 138.130000 ;
      RECT 70.000000 138.060000 75.145000 138.130000 ;
      RECT 70.060000 139.850000 75.145000 139.920000 ;
      RECT 70.060000 139.850000 75.145000 139.920000 ;
      RECT 70.070000 137.990000 75.145000 138.060000 ;
      RECT 70.070000 137.990000 75.145000 138.060000 ;
      RECT 70.105000 145.100000 75.145000 145.130000 ;
      RECT 70.130000 139.920000 75.145000 139.990000 ;
      RECT 70.130000 139.920000 75.145000 139.990000 ;
      RECT 70.140000 137.920000 75.145000 137.990000 ;
      RECT 70.140000 137.920000 75.145000 137.990000 ;
      RECT 70.175000 145.030000 75.145000 145.100000 ;
      RECT 70.200000 139.990000 75.145000 140.060000 ;
      RECT 70.200000 139.990000 75.145000 140.060000 ;
      RECT 70.210000 137.850000 75.145000 137.920000 ;
      RECT 70.210000 137.850000 75.145000 137.920000 ;
      RECT 70.245000 144.960000 75.145000 145.030000 ;
      RECT 70.270000 140.060000 75.145000 140.130000 ;
      RECT 70.270000 140.060000 75.145000 140.130000 ;
      RECT 70.280000 137.780000 75.145000 137.850000 ;
      RECT 70.280000 137.780000 75.145000 137.850000 ;
      RECT 70.315000 144.890000 75.145000 144.960000 ;
      RECT 70.340000 140.130000 75.145000 140.200000 ;
      RECT 70.340000 140.130000 75.145000 140.200000 ;
      RECT 70.350000 137.710000 75.145000 137.780000 ;
      RECT 70.350000 137.710000 75.145000 137.780000 ;
      RECT 70.385000 144.820000 75.145000 144.890000 ;
      RECT 70.410000 140.200000 75.145000 140.270000 ;
      RECT 70.410000 140.200000 75.145000 140.270000 ;
      RECT 70.420000 137.640000 75.145000 137.710000 ;
      RECT 70.420000 137.640000 75.145000 137.710000 ;
      RECT 70.455000 144.750000 75.145000 144.820000 ;
      RECT 70.480000 140.270000 75.145000 140.340000 ;
      RECT 70.480000 140.270000 75.145000 140.340000 ;
      RECT 70.490000 137.570000 75.145000 137.640000 ;
      RECT 70.490000 137.570000 75.145000 137.640000 ;
      RECT 70.525000 144.680000 75.145000 144.750000 ;
      RECT 70.550000 140.340000 75.145000 140.410000 ;
      RECT 70.550000 140.340000 75.145000 140.410000 ;
      RECT 70.560000 137.500000 75.145000 137.570000 ;
      RECT 70.560000 137.500000 75.145000 137.570000 ;
      RECT 70.595000 144.610000 75.145000 144.680000 ;
      RECT 70.620000 140.410000 75.145000 140.480000 ;
      RECT 70.620000 140.410000 75.145000 140.480000 ;
      RECT 70.630000 137.430000 75.145000 137.500000 ;
      RECT 70.630000 137.430000 75.145000 137.500000 ;
      RECT 70.665000 144.540000 75.145000 144.610000 ;
      RECT 70.690000 140.480000 75.145000 140.550000 ;
      RECT 70.690000 140.480000 75.145000 140.550000 ;
      RECT 70.700000 137.360000 75.145000 137.430000 ;
      RECT 70.700000 137.360000 75.145000 137.430000 ;
      RECT 70.735000 144.470000 75.145000 144.540000 ;
      RECT 70.760000 140.550000 75.145000 140.620000 ;
      RECT 70.760000 140.550000 75.145000 140.620000 ;
      RECT 70.770000 137.290000 75.145000 137.360000 ;
      RECT 70.770000 137.290000 75.145000 137.360000 ;
      RECT 70.805000 139.850000 75.145000 145.130000 ;
      RECT 70.805000 140.620000 75.145000 140.665000 ;
      RECT 70.805000 140.620000 75.145000 140.665000 ;
      RECT 70.805000 140.665000 75.145000 144.400000 ;
      RECT 70.805000 144.400000 75.145000 144.470000 ;
      RECT 70.805000 144.400000 75.145000 145.130000 ;
      RECT 70.805000 145.130000 73.195000 146.145000 ;
      RECT 70.840000 137.220000 75.145000 137.290000 ;
      RECT 70.840000 137.220000 75.145000 137.290000 ;
      RECT 70.910000 137.150000 75.145000 137.220000 ;
      RECT 70.910000 137.150000 75.145000 137.220000 ;
      RECT 70.980000 137.080000 75.145000 137.150000 ;
      RECT 70.980000 137.080000 75.145000 137.150000 ;
      RECT 71.050000 137.010000 75.145000 137.080000 ;
      RECT 71.050000 137.010000 75.145000 137.080000 ;
      RECT 71.120000 136.940000 75.145000 137.010000 ;
      RECT 71.120000 136.940000 75.145000 137.010000 ;
      RECT 71.190000 136.870000 75.145000 136.940000 ;
      RECT 71.190000 136.870000 75.145000 136.940000 ;
      RECT 71.260000 136.800000 75.145000 136.870000 ;
      RECT 71.260000 136.800000 75.145000 136.870000 ;
      RECT 71.320000 100.290000 75.145000 100.330000 ;
      RECT 71.330000 136.730000 75.145000 136.800000 ;
      RECT 71.330000 136.730000 75.145000 136.800000 ;
      RECT 71.390000 100.220000 75.145000 100.290000 ;
      RECT 71.400000 136.660000 75.145000 136.730000 ;
      RECT 71.400000 136.660000 75.145000 136.730000 ;
      RECT 71.430000  97.760000 75.145000  97.830000 ;
      RECT 71.460000 100.150000 75.145000 100.220000 ;
      RECT 71.470000 136.590000 75.145000 136.660000 ;
      RECT 71.470000 136.590000 75.145000 136.660000 ;
      RECT 71.500000  97.830000 75.145000  97.900000 ;
      RECT 71.530000 100.080000 75.145000 100.150000 ;
      RECT 71.540000 136.520000 75.145000 136.590000 ;
      RECT 71.540000 136.520000 75.145000 136.590000 ;
      RECT 71.570000  97.900000 75.145000  97.970000 ;
      RECT 71.600000 100.010000 75.145000 100.080000 ;
      RECT 71.610000 136.450000 75.145000 136.520000 ;
      RECT 71.610000 136.450000 75.145000 136.520000 ;
      RECT 71.640000  97.970000 75.145000  98.040000 ;
      RECT 71.670000  99.940000 75.145000 100.010000 ;
      RECT 71.680000 136.380000 75.145000 136.450000 ;
      RECT 71.680000 136.380000 75.145000 136.450000 ;
      RECT 71.710000  98.040000 75.145000  98.110000 ;
      RECT 71.740000  99.870000 75.145000  99.940000 ;
      RECT 71.750000 136.310000 75.145000 136.380000 ;
      RECT 71.750000 136.310000 75.145000 136.380000 ;
      RECT 71.755000  85.835000 74.700000  94.470000 ;
      RECT 71.780000  98.110000 75.145000  98.180000 ;
      RECT 71.810000  99.800000 75.145000  99.870000 ;
      RECT 71.820000 136.240000 75.145000 136.310000 ;
      RECT 71.820000 136.240000 75.145000 136.310000 ;
      RECT 71.850000  98.180000 75.145000  98.250000 ;
      RECT 71.880000  99.730000 75.145000  99.800000 ;
      RECT 71.890000 136.170000 75.145000 136.240000 ;
      RECT 71.890000 136.170000 75.145000 136.240000 ;
      RECT 71.920000  98.250000 75.145000  98.320000 ;
      RECT 71.950000  99.660000 75.145000  99.730000 ;
      RECT 71.960000 136.100000 75.145000 136.170000 ;
      RECT 71.960000 136.100000 75.145000 136.170000 ;
      RECT 71.990000  98.320000 75.145000  98.390000 ;
      RECT 72.020000  99.590000 75.145000  99.660000 ;
      RECT 72.030000 136.030000 75.145000 136.100000 ;
      RECT 72.030000 136.030000 75.145000 136.100000 ;
      RECT 72.060000  98.390000 75.145000  98.460000 ;
      RECT 72.090000  97.530000 75.145000 100.765000 ;
      RECT 72.090000  97.760000 75.145000  98.490000 ;
      RECT 72.090000  98.460000 75.145000  98.490000 ;
      RECT 72.090000  98.490000 75.145000  99.520000 ;
      RECT 72.090000  99.520000 75.145000  99.590000 ;
      RECT 72.090000  99.520000 75.145000 100.330000 ;
      RECT 72.090000 100.330000 75.145000 101.420000 ;
      RECT 72.100000 135.960000 75.145000 136.030000 ;
      RECT 72.100000 135.960000 75.145000 136.030000 ;
      RECT 72.115000  97.505000 75.145000  97.530000 ;
      RECT 72.170000 135.890000 75.145000 135.960000 ;
      RECT 72.170000 135.890000 75.145000 135.960000 ;
      RECT 72.185000  97.435000 75.145000  97.505000 ;
      RECT 72.240000 135.820000 75.145000 135.890000 ;
      RECT 72.240000 135.820000 75.145000 135.890000 ;
      RECT 72.255000  97.365000 75.145000  97.435000 ;
      RECT 72.310000 135.750000 75.145000 135.820000 ;
      RECT 72.310000 135.750000 75.145000 135.820000 ;
      RECT 72.325000  97.295000 75.145000  97.365000 ;
      RECT 72.380000 130.500000 75.000000 130.995000 ;
      RECT 72.380000 135.680000 75.145000 135.750000 ;
      RECT 72.380000 135.680000 75.145000 135.750000 ;
      RECT 72.395000  97.225000 75.145000  97.295000 ;
      RECT 72.450000 135.610000 75.145000 135.680000 ;
      RECT 72.450000 135.610000 75.145000 135.680000 ;
      RECT 72.465000  97.155000 75.145000  97.225000 ;
      RECT 72.520000 135.540000 75.145000 135.610000 ;
      RECT 72.520000 135.540000 75.145000 135.610000 ;
      RECT 72.535000  97.085000 75.145000  97.155000 ;
      RECT 72.590000 135.470000 75.145000 135.540000 ;
      RECT 72.590000 135.470000 75.145000 135.540000 ;
      RECT 72.605000  97.015000 75.145000  97.085000 ;
      RECT 72.660000 131.275000 75.145000 132.915000 ;
      RECT 72.660000 135.400000 75.145000 135.470000 ;
      RECT 72.660000 135.400000 75.145000 135.470000 ;
      RECT 72.675000  96.945000 75.145000  97.015000 ;
      RECT 72.695000 135.365000 75.145000 135.400000 ;
      RECT 72.695000 135.365000 75.145000 135.400000 ;
      RECT 72.745000  96.875000 75.145000  96.945000 ;
      RECT 72.765000 135.295000 75.145000 135.365000 ;
      RECT 72.765000 135.295000 75.145000 135.365000 ;
      RECT 72.815000  96.805000 75.145000  96.875000 ;
      RECT 72.835000 135.225000 75.145000 135.295000 ;
      RECT 72.835000 135.225000 75.145000 135.295000 ;
      RECT 72.885000  96.735000 75.145000  96.805000 ;
      RECT 72.905000 135.155000 75.145000 135.225000 ;
      RECT 72.905000 135.155000 75.145000 135.225000 ;
      RECT 72.955000  96.665000 75.145000  96.735000 ;
      RECT 72.975000 135.085000 75.145000 135.155000 ;
      RECT 72.975000 135.085000 75.145000 135.155000 ;
      RECT 73.025000  96.595000 75.145000  96.665000 ;
      RECT 73.045000 135.015000 75.145000 135.085000 ;
      RECT 73.045000 135.015000 75.145000 135.085000 ;
      RECT 73.095000  96.525000 75.145000  96.595000 ;
      RECT 73.115000 134.945000 75.145000 135.015000 ;
      RECT 73.115000 134.945000 75.145000 135.015000 ;
      RECT 73.165000  96.455000 75.145000  96.525000 ;
      RECT 73.185000 134.875000 75.145000 134.945000 ;
      RECT 73.185000 134.875000 75.145000 134.945000 ;
      RECT 73.235000  96.385000 75.145000  96.455000 ;
      RECT 73.255000 134.805000 75.145000 134.875000 ;
      RECT 73.255000 134.805000 75.145000 134.875000 ;
      RECT 73.295000   5.990000 74.590000   6.060000 ;
      RECT 73.305000  96.315000 75.145000  96.385000 ;
      RECT 73.325000 134.735000 75.145000 134.805000 ;
      RECT 73.325000 134.735000 75.145000 134.805000 ;
      RECT 73.365000   6.060000 74.590000   6.130000 ;
      RECT 73.375000  96.245000 75.145000  96.315000 ;
      RECT 73.395000 134.665000 75.145000 134.735000 ;
      RECT 73.395000 134.665000 75.145000 134.735000 ;
      RECT 73.435000   6.130000 74.590000   6.200000 ;
      RECT 73.445000  96.175000 75.145000  96.245000 ;
      RECT 73.465000 134.595000 75.145000 134.665000 ;
      RECT 73.465000 134.595000 75.145000 134.665000 ;
      RECT 73.475000 145.410000 75.000000 146.425000 ;
      RECT 73.505000   6.200000 74.590000   6.270000 ;
      RECT 73.515000  96.105000 75.145000  96.175000 ;
      RECT 73.535000 134.525000 75.145000 134.595000 ;
      RECT 73.535000 134.525000 75.145000 134.595000 ;
      RECT 73.575000   6.270000 74.590000   6.340000 ;
      RECT 73.585000  96.035000 75.145000  96.105000 ;
      RECT 73.605000 134.455000 75.145000 134.525000 ;
      RECT 73.605000 134.455000 75.145000 134.525000 ;
      RECT 73.645000   6.340000 74.590000   6.410000 ;
      RECT 73.655000  95.965000 75.145000  96.035000 ;
      RECT 73.660000   6.410000 74.590000   6.425000 ;
      RECT 73.660000   6.425000 74.590000  79.620000 ;
      RECT 73.660000  79.620000 74.590000  79.675000 ;
      RECT 73.660000  79.675000 74.645000  79.730000 ;
      RECT 73.660000  79.730000 74.700000  84.800000 ;
      RECT 73.675000 134.385000 75.145000 134.455000 ;
      RECT 73.675000 134.385000 75.145000 134.455000 ;
      RECT 73.685000 174.500000 74.745000 175.140000 ;
      RECT 73.725000  95.895000 75.145000  95.965000 ;
      RECT 73.725000  95.895000 75.145000 100.535000 ;
      RECT 73.745000 134.315000 75.145000 134.385000 ;
      RECT 73.745000 134.315000 75.145000 134.385000 ;
      RECT 73.770000 101.420000 74.700000 104.565000 ;
      RECT 73.815000 134.245000 75.145000 134.315000 ;
      RECT 73.815000 134.245000 75.145000 134.315000 ;
      RECT 73.885000 134.175000 75.145000 134.245000 ;
      RECT 73.885000 134.175000 75.145000 134.245000 ;
      RECT 73.955000 134.105000 75.145000 134.175000 ;
      RECT 73.955000 134.105000 75.145000 134.175000 ;
      RECT 74.025000 134.035000 75.145000 134.105000 ;
      RECT 74.025000 134.035000 75.145000 134.105000 ;
      RECT 74.035000 104.845000 75.000000 105.150000 ;
      RECT 74.095000 133.965000 75.145000 134.035000 ;
      RECT 74.095000 133.965000 75.145000 134.035000 ;
      RECT 74.165000 133.895000 75.145000 133.965000 ;
      RECT 74.165000 133.895000 75.145000 133.965000 ;
      RECT 74.235000 133.825000 75.145000 133.895000 ;
      RECT 74.235000 133.825000 75.145000 133.895000 ;
      RECT 74.305000 133.755000 75.145000 133.825000 ;
      RECT 74.305000 133.755000 75.145000 133.825000 ;
      RECT 74.315000 105.430000 74.915000 125.440000 ;
      RECT 74.375000 133.685000 75.145000 133.755000 ;
      RECT 74.375000 133.685000 75.145000 133.755000 ;
      RECT 74.445000 133.615000 75.145000 133.685000 ;
      RECT 74.445000 133.615000 75.145000 133.685000 ;
      RECT 74.515000 133.545000 75.145000 133.615000 ;
      RECT 74.515000 133.545000 75.145000 133.615000 ;
      RECT 74.585000 133.475000 75.145000 133.545000 ;
      RECT 74.585000 133.475000 75.145000 133.545000 ;
      RECT 74.655000 133.405000 75.145000 133.475000 ;
      RECT 74.655000 133.405000 75.145000 133.475000 ;
      RECT 74.725000 133.335000 75.145000 133.405000 ;
      RECT 74.725000 133.335000 75.145000 133.405000 ;
      RECT 74.795000 133.265000 75.145000 133.335000 ;
      RECT 74.795000 133.265000 75.145000 133.335000 ;
      RECT 74.855000 102.200000 74.925000 102.270000 ;
      RECT 74.855000 102.270000 74.995000 102.340000 ;
      RECT 74.855000 102.340000 75.065000 102.410000 ;
      RECT 74.855000 102.410000 75.135000 102.420000 ;
      RECT 74.865000 133.195000 75.145000 133.265000 ;
      RECT 74.865000 133.195000 75.145000 133.265000 ;
      RECT 74.935000 133.125000 75.145000 133.195000 ;
      RECT 74.935000 133.125000 75.145000 133.195000 ;
      RECT 75.005000 133.055000 75.145000 133.125000 ;
      RECT 75.005000 133.055000 75.145000 133.125000 ;
      RECT 75.075000 132.985000 75.145000 133.055000 ;
      RECT 75.075000 132.985000 75.145000 133.055000 ;
    LAYER met2 ;
      RECT  0.000000   0.000000  8.145000   4.404000 ;
      RECT  0.000000   0.000000  8.285000   1.320000 ;
      RECT  0.000000   1.320000 12.145000   1.610000 ;
      RECT  0.000000   1.610000 17.105000   3.275000 ;
      RECT  0.000000   3.155000 10.634000   3.225000 ;
      RECT  0.000000   3.225000 10.564000   3.295000 ;
      RECT  0.000000   3.275000 19.935000   3.295000 ;
      RECT  0.000000   3.295000  9.595000   4.462000 ;
      RECT  0.000000   3.295000 10.494000   3.365000 ;
      RECT  0.000000   3.365000 10.424000   3.435000 ;
      RECT  0.000000   3.435000 10.354000   3.505000 ;
      RECT  0.000000   3.505000 10.284000   3.575000 ;
      RECT  0.000000   3.575000 10.214000   3.645000 ;
      RECT  0.000000   3.645000 10.144000   3.715000 ;
      RECT  0.000000   3.715000 10.074000   3.785000 ;
      RECT  0.000000   3.785000 10.004000   3.855000 ;
      RECT  0.000000   3.855000  9.934000   3.925000 ;
      RECT  0.000000   3.925000  9.864000   3.995000 ;
      RECT  0.000000   3.995000  9.794000   4.065000 ;
      RECT  0.000000   4.065000  9.724000   4.135000 ;
      RECT  0.000000   4.135000  9.654000   4.205000 ;
      RECT  0.000000   4.205000  9.584000   4.275000 ;
      RECT  0.000000   4.275000  9.514000   4.345000 ;
      RECT  0.000000   4.345000  9.454000   4.405000 ;
      RECT  0.000000   4.404000  3.005000  26.494000 ;
      RECT  0.000000   4.462000  9.595000   9.028000 ;
      RECT  0.000000   9.028000 10.725000  10.158000 ;
      RECT  0.000000   9.086000  9.455000   9.155000 ;
      RECT  0.000000   9.155000  9.524000   9.225000 ;
      RECT  0.000000   9.225000  9.594000   9.295000 ;
      RECT  0.000000   9.295000  9.664000   9.365000 ;
      RECT  0.000000   9.365000  9.734000   9.435000 ;
      RECT  0.000000   9.435000  9.804000   9.505000 ;
      RECT  0.000000   9.505000  9.874000   9.575000 ;
      RECT  0.000000   9.575000  9.944000   9.645000 ;
      RECT  0.000000   9.645000 10.014000   9.715000 ;
      RECT  0.000000   9.715000 10.084000   9.785000 ;
      RECT  0.000000   9.785000 10.154000   9.855000 ;
      RECT  0.000000   9.855000 10.224000   9.925000 ;
      RECT  0.000000   9.925000 10.294000   9.995000 ;
      RECT  0.000000   9.995000 10.364000  10.065000 ;
      RECT  0.000000  10.065000 10.434000  10.135000 ;
      RECT  0.000000  10.135000 10.504000  10.205000 ;
      RECT  0.000000  10.158000 10.725000  26.552000 ;
      RECT  0.000000  10.205000 10.574000  10.215000 ;
      RECT  0.000000  26.494000 10.514000  26.565000 ;
      RECT  0.000000  26.552000 10.510000  26.767000 ;
      RECT  0.000000  26.565000 10.444000  26.635000 ;
      RECT  0.000000  26.635000 10.374000  26.705000 ;
      RECT  0.000000  26.705000 10.369000  26.710000 ;
      RECT  0.000000  26.709000  3.005000 196.995000 ;
      RECT  0.000000  26.767000 10.510000  28.468000 ;
      RECT  0.000000  28.468000 10.725000  28.683000 ;
      RECT  0.000000  28.526000 10.370000  28.595000 ;
      RECT  0.000000  28.595000 10.439000  28.665000 ;
      RECT  0.000000  28.665000 10.509000  28.735000 ;
      RECT  0.000000  28.683000 10.725000  31.253000 ;
      RECT  0.000000  28.735000 10.579000  28.740000 ;
      RECT  0.000000  31.253000 11.120000  31.648000 ;
      RECT  0.000000  31.311000 10.585000  31.380000 ;
      RECT  0.000000  31.380000 10.654000  31.450000 ;
      RECT  0.000000  31.450000 10.724000  31.520000 ;
      RECT  0.000000  31.520000 10.794000  31.590000 ;
      RECT  0.000000  31.590000 10.864000  31.660000 ;
      RECT  0.000000  31.648000 11.120000  36.420000 ;
      RECT  0.000000  31.660000 10.934000  31.705000 ;
      RECT  0.000000  36.420000 75.000000 200.000000 ;
      RECT  0.000000 196.995000 75.000000 200.000000 ;
      RECT  3.002000   3.002000  5.143000   4.462000 ;
      RECT  3.002000   4.462000  6.453000  10.330000 ;
      RECT  3.002000  10.330000  6.453000  10.400000 ;
      RECT  3.002000  10.330000  6.453000  10.400000 ;
      RECT  3.002000  10.400000  6.523000  10.470000 ;
      RECT  3.002000  10.400000  6.523000  10.470000 ;
      RECT  3.002000  10.470000  6.593000  10.540000 ;
      RECT  3.002000  10.470000  6.593000  10.540000 ;
      RECT  3.002000  10.540000  6.663000  10.610000 ;
      RECT  3.002000  10.540000  6.663000  10.610000 ;
      RECT  3.002000  10.610000  6.733000  10.680000 ;
      RECT  3.002000  10.610000  6.733000  10.680000 ;
      RECT  3.002000  10.680000  6.803000  10.750000 ;
      RECT  3.002000  10.680000  6.803000  10.750000 ;
      RECT  3.002000  10.750000  6.873000  10.820000 ;
      RECT  3.002000  10.750000  6.873000  10.820000 ;
      RECT  3.002000  10.820000  6.943000  10.890000 ;
      RECT  3.002000  10.820000  6.943000  10.890000 ;
      RECT  3.002000  10.890000  7.013000  10.960000 ;
      RECT  3.002000  10.890000  7.013000  10.960000 ;
      RECT  3.002000  10.960000  7.083000  11.030000 ;
      RECT  3.002000  10.960000  7.083000  11.030000 ;
      RECT  3.002000  11.030000  7.153000  11.100000 ;
      RECT  3.002000  11.030000  7.153000  11.100000 ;
      RECT  3.002000  11.100000  7.223000  11.170000 ;
      RECT  3.002000  11.100000  7.223000  11.170000 ;
      RECT  3.002000  11.170000  7.293000  11.240000 ;
      RECT  3.002000  11.170000  7.293000  11.240000 ;
      RECT  3.002000  11.240000  7.363000  11.310000 ;
      RECT  3.002000  11.240000  7.363000  11.310000 ;
      RECT  3.002000  11.310000  7.433000  11.380000 ;
      RECT  3.002000  11.310000  7.433000  11.380000 ;
      RECT  3.002000  11.380000  7.503000  11.450000 ;
      RECT  3.002000  11.380000  7.503000  11.450000 ;
      RECT  3.002000  11.450000  7.573000  11.460000 ;
      RECT  3.002000  11.450000  7.573000  11.460000 ;
      RECT  3.002000  11.460000  7.583000  25.250000 ;
      RECT  3.002000  25.250000  7.513000  25.320000 ;
      RECT  3.002000  25.250000  7.513000  25.320000 ;
      RECT  3.002000  25.320000  7.443000  25.390000 ;
      RECT  3.002000  25.320000  7.443000  25.390000 ;
      RECT  3.002000  25.390000  7.373000  25.460000 ;
      RECT  3.002000  25.390000  7.373000  25.460000 ;
      RECT  3.002000  25.460000  7.368000  25.465000 ;
      RECT  3.002000  25.460000  7.368000  25.465000 ;
      RECT  3.002000  25.465000  7.368000  29.770000 ;
      RECT  3.002000  29.770000  7.368000  29.840000 ;
      RECT  3.002000  29.770000  7.368000  29.840000 ;
      RECT  3.002000  29.840000  7.438000  29.910000 ;
      RECT  3.002000  29.840000  7.438000  29.910000 ;
      RECT  3.002000  29.910000  7.508000  29.980000 ;
      RECT  3.002000  29.910000  7.508000  29.980000 ;
      RECT  3.002000  29.980000  7.578000  29.985000 ;
      RECT  3.002000  29.980000  7.578000  29.985000 ;
      RECT  3.002000  29.985000  7.583000  32.555000 ;
      RECT  3.002000  32.555000  7.583000  32.625000 ;
      RECT  3.002000  32.555000  7.583000  32.625000 ;
      RECT  3.002000  32.625000  7.653000  32.695000 ;
      RECT  3.002000  32.625000  7.653000  32.695000 ;
      RECT  3.002000  32.695000  7.723000  32.765000 ;
      RECT  3.002000  32.695000  7.723000  32.765000 ;
      RECT  3.002000  32.765000  7.793000  32.835000 ;
      RECT  3.002000  32.765000  7.793000  32.835000 ;
      RECT  3.002000  32.835000  7.863000  32.905000 ;
      RECT  3.002000  32.835000  7.863000  32.905000 ;
      RECT  3.002000  32.905000  7.933000  32.950000 ;
      RECT  3.002000  32.905000  7.933000  32.950000 ;
      RECT  3.002000  32.950000  7.978000  39.562000 ;
      RECT  3.002000  39.562000 71.998000 196.998000 ;
      RECT  5.143000   4.404000  9.455000   7.409000 ;
      RECT  6.450000   1.750000 16.965000   3.155000 ;
      RECT  6.450000   3.155000  9.455000   4.404000 ;
      RECT  6.450000   7.409000  9.455000  10.216000 ;
      RECT  6.453000  10.216000 10.585000  13.221000 ;
      RECT  7.365000  26.709000 10.370000  28.741000 ;
      RECT  7.365000  28.741000 10.585000  31.311000 ;
      RECT  7.368000  23.489000 10.585000  26.494000 ;
      RECT  7.368000  31.311000 10.585000  31.706000 ;
      RECT  7.368000  31.706000 10.980000  31.746000 ;
      RECT  7.580000  13.221000 10.585000  23.489000 ;
      RECT  7.580000  31.746000 10.980000  36.560000 ;
      RECT  7.975000  36.560000 15.435000  39.562000 ;
      RECT  7.978000  39.562000 15.432000  39.565000 ;
      RECT  8.145000   1.460000 12.005000   1.750000 ;
      RECT  9.035000   0.000000 12.145000   1.320000 ;
      RECT  9.175000   0.000000 12.005000   1.460000 ;
      RECT 10.135000   4.688000 15.827000   4.945000 ;
      RECT 10.135000   4.945000 29.180000   5.528000 ;
      RECT 10.135000   5.528000 29.180000   8.802000 ;
      RECT 10.135000   8.802000 29.180000   9.932000 ;
      RECT 10.275000   4.746000 15.430000   4.815000 ;
      RECT 10.275000   4.815000 15.499000   4.885000 ;
      RECT 10.275000   4.885000 15.569000   4.955000 ;
      RECT 10.275000   4.955000 15.639000   5.025000 ;
      RECT 10.275000   5.025000 15.709000   5.085000 ;
      RECT 10.275000   5.085000 28.539000   5.155000 ;
      RECT 10.275000   5.155000 28.609000   5.225000 ;
      RECT 10.275000   5.225000 28.679000   5.295000 ;
      RECT 10.275000   5.295000 28.749000   5.365000 ;
      RECT 10.275000   5.365000 28.819000   5.435000 ;
      RECT 10.275000   5.435000 28.889000   5.505000 ;
      RECT 10.275000   5.505000 28.959000   5.575000 ;
      RECT 10.275000   5.575000 29.029000   5.585000 ;
      RECT 10.275000   5.586000 29.040000   8.591000 ;
      RECT 10.275000   8.591000 14.407000   8.744000 ;
      RECT 10.346000   4.675000 15.359000   4.745000 ;
      RECT 10.346000   8.744000 29.040000   8.815000 ;
      RECT 10.416000   4.605000 15.289000   4.675000 ;
      RECT 10.416000   8.815000 29.040000   8.885000 ;
      RECT 10.486000   4.535000 15.219000   4.605000 ;
      RECT 10.486000   8.885000 29.040000   8.955000 ;
      RECT 10.556000   4.465000 15.149000   4.535000 ;
      RECT 10.556000   8.955000 29.040000   9.025000 ;
      RECT 10.626000   4.395000 15.079000   4.465000 ;
      RECT 10.626000   9.025000 29.040000   9.095000 ;
      RECT 10.696000   4.325000 15.009000   4.395000 ;
      RECT 10.696000   9.095000 29.040000   9.165000 ;
      RECT 10.766000   4.255000 14.939000   4.325000 ;
      RECT 10.766000   9.165000 29.040000   9.235000 ;
      RECT 10.836000   4.185000 14.869000   4.255000 ;
      RECT 10.836000   9.235000 29.040000   9.305000 ;
      RECT 10.906000   4.115000 14.799000   4.185000 ;
      RECT 10.906000   9.305000 29.040000   9.375000 ;
      RECT 10.976000   4.045000 14.729000   4.115000 ;
      RECT 10.976000   9.375000 29.040000   9.445000 ;
      RECT 10.988000   3.835000 15.570000   4.688000 ;
      RECT 11.046000   3.975000 14.659000   4.045000 ;
      RECT 11.046000   9.445000 29.040000   9.515000 ;
      RECT 11.050000  27.358000 75.000000  27.877000 ;
      RECT 11.050000  27.877000 75.000000  28.092000 ;
      RECT 11.116000   9.515000 29.040000   9.585000 ;
      RECT 11.186000   9.585000 29.040000   9.655000 ;
      RECT 11.190000  27.416000 14.805000  27.819000 ;
      RECT 11.196000  27.410000 75.000000  27.415000 ;
      RECT 11.256000   9.655000 29.040000   9.725000 ;
      RECT 11.261000  27.819000 75.000000  27.890000 ;
      RECT 11.265000   9.932000 29.180000  11.143000 ;
      RECT 11.265000  11.143000 29.630000  11.593000 ;
      RECT 11.265000  11.593000 29.630000  15.813000 ;
      RECT 11.265000  15.813000 30.225000  16.408000 ;
      RECT 11.265000  16.408000 30.225000  20.635000 ;
      RECT 11.265000  20.635000 75.000000  27.143000 ;
      RECT 11.265000  27.143000 75.000000  27.358000 ;
      RECT 11.265000  28.092000 75.000000  31.027000 ;
      RECT 11.265000  31.027000 75.000000  31.422000 ;
      RECT 11.266000  27.340000 75.000000  27.410000 ;
      RECT 11.326000   9.725000 29.040000   9.795000 ;
      RECT 11.331000  27.890000 75.000000  27.960000 ;
      RECT 11.336000  27.270000 75.000000  27.340000 ;
      RECT 11.396000   9.795000 29.040000   9.865000 ;
      RECT 11.401000  27.960000 75.000000  28.030000 ;
      RECT 11.405000   9.874000 14.407000  11.201000 ;
      RECT 11.405000  11.201000 29.040000  11.270000 ;
      RECT 11.405000  11.270000 29.109000  11.340000 ;
      RECT 11.405000  11.340000 29.179000  11.410000 ;
      RECT 11.405000  11.410000 29.249000  11.480000 ;
      RECT 11.405000  11.480000 29.319000  11.550000 ;
      RECT 11.405000  11.550000 29.389000  11.620000 ;
      RECT 11.405000  11.620000 29.459000  11.650000 ;
      RECT 11.405000  11.651000 14.410000  15.871000 ;
      RECT 11.405000  15.871000 29.490000  15.940000 ;
      RECT 11.405000  15.940000 29.559000  16.010000 ;
      RECT 11.405000  16.010000 29.629000  16.080000 ;
      RECT 11.405000  16.080000 29.699000  16.150000 ;
      RECT 11.405000  16.150000 29.769000  16.220000 ;
      RECT 11.405000  16.220000 29.839000  16.290000 ;
      RECT 11.405000  16.290000 29.909000  16.360000 ;
      RECT 11.405000  16.360000 29.979000  16.430000 ;
      RECT 11.405000  16.430000 30.049000  16.465000 ;
      RECT 11.405000  16.466000 14.410000  20.775000 ;
      RECT 11.405000  20.775000 14.805000  27.416000 ;
      RECT 11.405000  27.201000 75.000000  27.270000 ;
      RECT 11.405000  27.819000 14.805000  30.969000 ;
      RECT 11.406000   9.865000 29.040000   9.875000 ;
      RECT 11.406000  28.030000 75.000000  28.035000 ;
      RECT 11.476000  30.969000 75.000000  31.040000 ;
      RECT 11.546000  31.040000 75.000000  31.110000 ;
      RECT 11.616000  31.110000 75.000000  31.180000 ;
      RECT 11.660000  31.422000 75.000000  35.880000 ;
      RECT 11.686000  31.180000 75.000000  31.250000 ;
      RECT 11.756000  31.250000 75.000000  31.320000 ;
      RECT 11.800000  30.969000 14.805000  35.740000 ;
      RECT 11.801000  31.320000 75.000000  31.365000 ;
      RECT 12.290000  35.880000 75.000000  36.420000 ;
      RECT 12.430000  20.775000 75.000000  36.560000 ;
      RECT 12.685000   0.000000 14.415000   1.125000 ;
      RECT 12.685000   1.125000 17.105000   1.610000 ;
      RECT 12.795000   1.745000 16.965000   1.750000 ;
      RECT 12.810000   1.730000 16.965000   1.745000 ;
      RECT 12.825000   0.000000 14.275000   1.265000 ;
      RECT 12.825000   1.265000 16.965000   1.715000 ;
      RECT 12.825000   1.715000 16.965000   1.730000 ;
      RECT 13.277000   6.977000 13.415000   7.045000 ;
      RECT 13.277000   6.977000 13.415000   7.045000 ;
      RECT 13.277000   7.045000 13.483000   7.115000 ;
      RECT 13.277000   7.045000 13.483000   7.115000 ;
      RECT 13.277000   7.115000 13.553000   7.185000 ;
      RECT 13.277000   7.115000 13.553000   7.185000 ;
      RECT 13.277000   7.185000 13.623000   7.255000 ;
      RECT 13.277000   7.185000 13.623000   7.255000 ;
      RECT 13.277000   7.255000 13.693000   7.325000 ;
      RECT 13.277000   7.255000 13.693000   7.325000 ;
      RECT 13.277000   7.325000 13.763000   7.395000 ;
      RECT 13.277000   7.325000 13.763000   7.395000 ;
      RECT 13.277000   7.395000 13.833000   7.465000 ;
      RECT 13.277000   7.395000 13.833000   7.465000 ;
      RECT 13.277000   7.465000 13.903000   7.500000 ;
      RECT 13.277000   7.465000 13.903000   7.500000 ;
      RECT 13.347000   7.500000 13.938000   7.570000 ;
      RECT 13.347000   7.500000 13.938000   7.570000 ;
      RECT 13.417000   7.570000 14.008000   7.640000 ;
      RECT 13.417000   7.570000 14.008000   7.640000 ;
      RECT 13.487000   7.640000 14.078000   7.710000 ;
      RECT 13.487000   7.640000 14.078000   7.710000 ;
      RECT 13.557000   7.710000 14.148000   7.780000 ;
      RECT 13.557000   7.710000 14.148000   7.780000 ;
      RECT 13.627000   7.780000 14.218000   7.850000 ;
      RECT 13.627000   7.780000 14.218000   7.850000 ;
      RECT 13.697000   7.850000 14.288000   7.920000 ;
      RECT 13.697000   7.850000 14.288000   7.920000 ;
      RECT 13.767000   7.920000 14.358000   7.990000 ;
      RECT 13.767000   7.920000 14.358000   7.990000 ;
      RECT 13.837000   7.990000 14.428000   8.060000 ;
      RECT 13.837000   7.990000 14.428000   8.060000 ;
      RECT 13.862000   8.060000 14.498000   8.085000 ;
      RECT 13.862000   8.060000 14.498000   8.085000 ;
      RECT 13.932000   8.087000 26.038000   8.155000 ;
      RECT 13.932000   8.087000 26.038000   8.155000 ;
      RECT 14.002000   8.155000 26.038000   8.225000 ;
      RECT 14.002000   8.155000 26.038000   8.225000 ;
      RECT 14.072000   8.225000 26.038000   8.295000 ;
      RECT 14.072000   8.225000 26.038000   8.295000 ;
      RECT 14.142000   8.295000 26.038000   8.365000 ;
      RECT 14.142000   8.295000 26.038000   8.365000 ;
      RECT 14.212000   8.365000 26.038000   8.435000 ;
      RECT 14.212000   8.365000 26.038000   8.435000 ;
      RECT 14.282000   8.435000 26.038000   8.505000 ;
      RECT 14.282000   8.435000 26.038000   8.505000 ;
      RECT 14.352000   8.505000 26.038000   8.575000 ;
      RECT 14.352000   8.505000 26.038000   8.575000 ;
      RECT 14.407000   8.575000 26.038000   8.630000 ;
      RECT 14.407000   8.575000 26.038000   8.630000 ;
      RECT 14.407000   8.630000 26.038000  12.445000 ;
      RECT 14.407000  12.445000 26.038000  12.515000 ;
      RECT 14.407000  12.445000 26.038000  12.515000 ;
      RECT 14.407000  12.515000 26.108000  12.585000 ;
      RECT 14.407000  12.515000 26.108000  12.585000 ;
      RECT 14.407000  12.585000 26.178000  12.655000 ;
      RECT 14.407000  12.585000 26.178000  12.655000 ;
      RECT 14.407000  12.655000 26.248000  12.725000 ;
      RECT 14.407000  12.655000 26.248000  12.725000 ;
      RECT 14.407000  12.725000 26.318000  12.795000 ;
      RECT 14.407000  12.725000 26.318000  12.795000 ;
      RECT 14.407000  12.795000 26.388000  12.865000 ;
      RECT 14.407000  12.795000 26.388000  12.865000 ;
      RECT 14.407000  12.865000 26.458000  12.895000 ;
      RECT 14.407000  12.865000 26.458000  12.895000 ;
      RECT 14.407000  12.895000 26.488000  17.115000 ;
      RECT 14.407000  17.115000 26.488000  17.185000 ;
      RECT 14.407000  17.115000 26.488000  17.185000 ;
      RECT 14.407000  17.185000 26.558000  17.255000 ;
      RECT 14.407000  17.185000 26.558000  17.255000 ;
      RECT 14.407000  17.255000 26.628000  17.325000 ;
      RECT 14.407000  17.255000 26.628000  17.325000 ;
      RECT 14.407000  17.325000 26.698000  17.395000 ;
      RECT 14.407000  17.325000 26.698000  17.395000 ;
      RECT 14.407000  17.395000 26.768000  17.465000 ;
      RECT 14.407000  17.395000 26.768000  17.465000 ;
      RECT 14.407000  17.465000 26.838000  17.535000 ;
      RECT 14.407000  17.465000 26.838000  17.535000 ;
      RECT 14.407000  17.535000 26.908000  17.605000 ;
      RECT 14.407000  17.535000 26.908000  17.605000 ;
      RECT 14.407000  17.605000 26.978000  17.675000 ;
      RECT 14.407000  17.605000 26.978000  17.675000 ;
      RECT 14.407000  17.675000 27.048000  17.710000 ;
      RECT 14.407000  17.675000 27.048000  17.710000 ;
      RECT 14.407000  17.710000 27.083000  23.777000 ;
      RECT 14.407000  23.777000 71.998000  29.725000 ;
      RECT 14.477000  29.725000 71.998000  29.795000 ;
      RECT 14.477000  29.725000 71.998000  29.795000 ;
      RECT 14.547000  29.795000 71.998000  29.865000 ;
      RECT 14.547000  29.795000 71.998000  29.865000 ;
      RECT 14.617000  29.865000 71.998000  29.935000 ;
      RECT 14.617000  29.865000 71.998000  29.935000 ;
      RECT 14.687000  29.935000 71.998000  30.005000 ;
      RECT 14.687000  29.935000 71.998000  30.005000 ;
      RECT 14.757000  30.005000 71.998000  30.075000 ;
      RECT 14.757000  30.005000 71.998000  30.075000 ;
      RECT 14.802000  30.075000 71.998000  30.120000 ;
      RECT 14.802000  30.075000 71.998000  30.120000 ;
      RECT 14.802000  30.120000 71.998000  32.738000 ;
      RECT 14.943000   3.295000 19.935000   3.595000 ;
      RECT 15.071000   3.155000 16.965000   3.225000 ;
      RECT 15.141000   3.225000 16.965000   3.295000 ;
      RECT 15.211000   3.295000 16.965000   3.365000 ;
      RECT 15.243000   3.595000 22.220000   4.187000 ;
      RECT 15.261000   3.365000 16.965000   3.415000 ;
      RECT 15.275000   0.000000 17.105000   1.125000 ;
      RECT 15.331000   3.415000 19.795000   3.485000 ;
      RECT 15.401000   3.485000 19.795000   3.555000 ;
      RECT 15.415000   0.000000 16.965000   1.265000 ;
      RECT 15.432000  32.738000 71.998000  39.562000 ;
      RECT 15.471000   3.555000 19.795000   3.625000 ;
      RECT 15.541000   3.625000 19.795000   3.695000 ;
      RECT 15.581000   3.695000 19.795000   3.735000 ;
      RECT 15.651000   3.735000 22.080000   3.805000 ;
      RECT 15.721000   3.805000 22.080000   3.875000 ;
      RECT 15.791000   3.875000 22.080000   3.945000 ;
      RECT 15.835000   4.187000 22.002000   4.405000 ;
      RECT 15.861000   3.945000 22.080000   4.015000 ;
      RECT 15.931000   4.015000 22.080000   4.085000 ;
      RECT 15.976000   4.085000 22.080000   4.130000 ;
      RECT 16.041000   4.129000 22.014000   4.195000 ;
      RECT 16.111000   4.195000 21.944000   4.265000 ;
      RECT 19.050000   0.000000 19.935000   3.275000 ;
      RECT 19.190000   0.000000 19.795000   3.415000 ;
      RECT 21.365000   0.000000 22.220000   3.595000 ;
      RECT 21.505000   0.000000 22.080000   3.735000 ;
      RECT 22.800000   0.000000 27.440000   0.470000 ;
      RECT 22.800000   0.470000 28.775000   0.475000 ;
      RECT 22.800000   0.475000 32.620000   0.780000 ;
      RECT 22.800000   0.780000 72.075000   0.910000 ;
      RECT 22.800000   0.910000 75.000000   4.202000 ;
      RECT 22.800000   4.202000 75.000000   4.405000 ;
      RECT 22.940000   0.000000 27.300000   0.610000 ;
      RECT 22.940000   0.610000 28.635000   0.615000 ;
      RECT 22.940000   0.615000 32.480000   0.920000 ;
      RECT 22.940000   0.920000 33.300000   3.925000 ;
      RECT 22.940000   3.925000 29.860000   4.144000 ;
      RECT 23.001000   4.144000 75.000000   4.205000 ;
      RECT 23.061000   4.205000 75.000000   4.265000 ;
      RECT 26.035000   8.591000 29.040000   8.744000 ;
      RECT 26.038000   9.874000 29.040000  11.201000 ;
      RECT 26.038000  11.651000 29.490000  14.656000 ;
      RECT 26.485000  14.656000 29.490000  15.871000 ;
      RECT 26.488000  16.466000 30.085000  19.471000 ;
      RECT 27.080000  19.471000 30.085000  20.775000 ;
      RECT 28.370000   0.000000 28.775000   0.470000 ;
      RECT 28.823000   4.405000 75.000000   5.302000 ;
      RECT 28.951000   4.265000 75.000000   4.335000 ;
      RECT 29.021000   4.335000 75.000000   4.405000 ;
      RECT 29.091000   4.405000 75.000000   4.475000 ;
      RECT 29.161000   4.475000 75.000000   4.545000 ;
      RECT 29.231000   4.545000 75.000000   4.615000 ;
      RECT 29.301000   4.615000 75.000000   4.685000 ;
      RECT 29.371000   4.685000 75.000000   4.755000 ;
      RECT 29.441000   4.755000 75.000000   4.825000 ;
      RECT 29.511000   4.825000 75.000000   4.895000 ;
      RECT 29.581000   4.895000 75.000000   4.965000 ;
      RECT 29.651000   4.965000 75.000000   5.035000 ;
      RECT 29.720000   5.302000 75.000000  10.917000 ;
      RECT 29.720000  10.917000 75.000000  11.367000 ;
      RECT 29.721000   5.035000 75.000000   5.105000 ;
      RECT 29.791000   5.105000 75.000000   5.175000 ;
      RECT 29.825000   0.000000 30.365000   0.470000 ;
      RECT 29.825000   0.470000 32.620000   0.475000 ;
      RECT 29.860000   1.050000 75.000000  10.859000 ;
      RECT 29.860000   1.050000 75.000000  10.859000 ;
      RECT 29.861000   5.175000 75.000000   5.245000 ;
      RECT 29.931000  10.859000 75.000000  10.930000 ;
      RECT 29.965000   0.000000 30.225000   0.610000 ;
      RECT 29.965000   0.610000 32.480000   0.615000 ;
      RECT 30.001000  10.930000 75.000000  11.000000 ;
      RECT 30.071000  11.000000 75.000000  11.070000 ;
      RECT 30.141000  11.070000 75.000000  11.140000 ;
      RECT 30.170000  11.367000 75.000000  15.587000 ;
      RECT 30.170000  15.587000 75.000000  16.182000 ;
      RECT 30.211000  11.140000 75.000000  11.210000 ;
      RECT 30.281000  11.210000 75.000000  11.280000 ;
      RECT 30.310000  10.859000 33.315000  12.524000 ;
      RECT 30.310000  12.524000 33.907000  15.529000 ;
      RECT 30.311000  11.280000 75.000000  11.310000 ;
      RECT 30.381000  15.529000 75.000000  15.600000 ;
      RECT 30.451000  15.600000 75.000000  15.670000 ;
      RECT 30.521000  15.670000 75.000000  15.740000 ;
      RECT 30.591000  15.740000 75.000000  15.810000 ;
      RECT 30.661000  15.810000 75.000000  15.880000 ;
      RECT 30.731000  15.880000 75.000000  15.950000 ;
      RECT 30.765000  16.182000 75.000000  20.635000 ;
      RECT 30.801000  15.950000 75.000000  16.020000 ;
      RECT 30.871000  16.020000 75.000000  16.090000 ;
      RECT 30.905000  16.124000 33.910000  20.775000 ;
      RECT 30.906000  16.090000 75.000000  16.125000 ;
      RECT 31.295000   0.000000 32.620000   0.470000 ;
      RECT 31.435000   0.000000 32.480000   0.610000 ;
      RECT 32.822000   3.922000 68.933000   3.960000 ;
      RECT 32.822000   3.922000 68.933000   3.960000 ;
      RECT 32.862000   3.960000 68.933000   4.000000 ;
      RECT 32.862000   3.960000 68.933000   4.000000 ;
      RECT 32.862000   4.000000 68.933000   4.052000 ;
      RECT 32.862000   4.052000 71.998000   9.615000 ;
      RECT 32.932000   9.615000 71.998000   9.685000 ;
      RECT 32.932000   9.615000 71.998000   9.685000 ;
      RECT 33.002000   9.685000 71.998000   9.755000 ;
      RECT 33.002000   9.685000 71.998000   9.755000 ;
      RECT 33.072000   9.755000 71.998000   9.825000 ;
      RECT 33.072000   9.755000 71.998000   9.825000 ;
      RECT 33.142000   9.825000 71.998000   9.895000 ;
      RECT 33.142000   9.825000 71.998000   9.895000 ;
      RECT 33.160000   0.000000 72.075000   0.780000 ;
      RECT 33.212000   9.895000 71.998000   9.965000 ;
      RECT 33.212000   9.895000 71.998000   9.965000 ;
      RECT 33.282000   9.965000 71.998000  10.035000 ;
      RECT 33.282000   9.965000 71.998000  10.035000 ;
      RECT 33.300000   0.000000 71.935000  10.859000 ;
      RECT 33.300000   0.000000 71.935000  10.859000 ;
      RECT 33.312000  10.035000 71.998000  10.065000 ;
      RECT 33.312000  10.035000 71.998000  10.065000 ;
      RECT 33.312000  10.065000 71.998000  14.285000 ;
      RECT 33.382000  14.285000 71.998000  14.355000 ;
      RECT 33.382000  14.285000 71.998000  14.355000 ;
      RECT 33.452000  14.355000 71.998000  14.425000 ;
      RECT 33.452000  14.355000 71.998000  14.425000 ;
      RECT 33.522000  14.425000 71.998000  14.495000 ;
      RECT 33.522000  14.425000 71.998000  14.495000 ;
      RECT 33.592000  14.495000 71.998000  14.565000 ;
      RECT 33.592000  14.495000 71.998000  14.565000 ;
      RECT 33.662000  14.565000 71.998000  14.635000 ;
      RECT 33.662000  14.565000 71.998000  14.635000 ;
      RECT 33.732000  14.635000 71.998000  14.705000 ;
      RECT 33.732000  14.635000 71.998000  14.705000 ;
      RECT 33.802000  14.705000 71.998000  14.775000 ;
      RECT 33.802000  14.705000 71.998000  14.775000 ;
      RECT 33.872000  14.775000 71.998000  14.845000 ;
      RECT 33.872000  14.775000 71.998000  14.845000 ;
      RECT 33.907000  14.845000 71.998000  14.880000 ;
      RECT 33.907000  14.845000 71.998000  14.880000 ;
      RECT 33.907000  14.880000 71.998000  23.777000 ;
      RECT 36.302000   3.002000 68.933000   3.922000 ;
      RECT 71.995000  10.859000 75.000000  15.529000 ;
      RECT 71.995000  16.124000 75.000000  20.775000 ;
      RECT 71.995000  36.560000 75.000000 196.995000 ;
      RECT 73.130000   1.020000 75.000000   1.050000 ;
      RECT 73.375000   0.000000 75.000000   0.910000 ;
      RECT 73.515000   0.000000 75.000000   1.020000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000  8.000000   3.005000 ;
      RECT  0.000000   0.000000  8.100000  15.661000 ;
      RECT  0.000000   3.005000  3.005000  17.244000 ;
      RECT  0.000000  15.619000  7.849000  15.770000 ;
      RECT  0.000000  15.661000  6.475000  17.286000 ;
      RECT  0.000000  15.770000  7.699000  15.920000 ;
      RECT  0.000000  15.920000  7.549000  16.070000 ;
      RECT  0.000000  16.070000  7.399000  16.220000 ;
      RECT  0.000000  16.220000  7.249000  16.370000 ;
      RECT  0.000000  16.370000  7.099000  16.520000 ;
      RECT  0.000000  16.520000  6.949000  16.670000 ;
      RECT  0.000000  16.670000  6.799000  16.820000 ;
      RECT  0.000000  16.820000  6.649000  16.970000 ;
      RECT  0.000000  16.970000  6.499000  17.120000 ;
      RECT  0.000000  17.120000  6.374000  17.245000 ;
      RECT  0.000000  17.244000  6.375000  64.434000 ;
      RECT  0.000000  17.286000  6.475000  31.629000 ;
      RECT  0.000000  31.629000  9.271000  34.425000 ;
      RECT  0.000000  31.671000  6.375000  31.820000 ;
      RECT  0.000000  31.820000  6.524000  31.970000 ;
      RECT  0.000000  31.970000  6.674000  32.120000 ;
      RECT  0.000000  32.120000  6.824000  32.270000 ;
      RECT  0.000000  32.270000  6.974000  32.420000 ;
      RECT  0.000000  32.420000  7.124000  32.570000 ;
      RECT  0.000000  32.570000  7.274000  32.720000 ;
      RECT  0.000000  32.720000  7.424000  32.870000 ;
      RECT  0.000000  32.870000  7.574000  33.020000 ;
      RECT  0.000000  33.020000  7.724000  33.170000 ;
      RECT  0.000000  33.170000  7.874000  33.320000 ;
      RECT  0.000000  33.320000  8.024000  33.470000 ;
      RECT  0.000000  33.470000  8.174000  33.620000 ;
      RECT  0.000000  33.620000  8.324000  33.770000 ;
      RECT  0.000000  33.770000  8.474000  33.920000 ;
      RECT  0.000000  33.920000  8.624000  34.070000 ;
      RECT  0.000000  34.070000  8.774000  34.220000 ;
      RECT  0.000000  34.220000  8.924000  34.370000 ;
      RECT  0.000000  34.370000  9.074000  34.520000 ;
      RECT  0.000000  34.425000 71.890000  64.476000 ;
      RECT  0.000000  34.520000  9.224000  34.525000 ;
      RECT  0.000000  64.434000 71.639000  64.585000 ;
      RECT  0.000000  64.476000 64.560000  71.806000 ;
      RECT  0.000000  64.585000 71.489000  64.735000 ;
      RECT  0.000000  64.735000 71.339000  64.885000 ;
      RECT  0.000000  64.885000 71.189000  65.035000 ;
      RECT  0.000000  65.035000 71.039000  65.185000 ;
      RECT  0.000000  65.185000 70.889000  65.335000 ;
      RECT  0.000000  65.335000 70.739000  65.485000 ;
      RECT  0.000000  65.485000 70.589000  65.635000 ;
      RECT  0.000000  65.635000 70.439000  65.785000 ;
      RECT  0.000000  65.785000 70.289000  65.935000 ;
      RECT  0.000000  65.935000 70.139000  66.085000 ;
      RECT  0.000000  66.085000 69.989000  66.235000 ;
      RECT  0.000000  66.235000 69.839000  66.385000 ;
      RECT  0.000000  66.385000 69.689000  66.535000 ;
      RECT  0.000000  66.535000 69.539000  66.685000 ;
      RECT  0.000000  66.685000 69.389000  66.835000 ;
      RECT  0.000000  66.835000 69.239000  66.985000 ;
      RECT  0.000000  66.985000 69.089000  67.135000 ;
      RECT  0.000000  67.135000 68.939000  67.285000 ;
      RECT  0.000000  67.285000 68.789000  67.435000 ;
      RECT  0.000000  67.435000 68.639000  67.585000 ;
      RECT  0.000000  67.585000 68.489000  67.735000 ;
      RECT  0.000000  67.735000 68.339000  67.885000 ;
      RECT  0.000000  67.885000 68.189000  68.035000 ;
      RECT  0.000000  68.035000 68.039000  68.185000 ;
      RECT  0.000000  68.185000 67.889000  68.335000 ;
      RECT  0.000000  68.335000 67.739000  68.485000 ;
      RECT  0.000000  68.485000 67.589000  68.635000 ;
      RECT  0.000000  68.635000 67.439000  68.785000 ;
      RECT  0.000000  68.785000 67.289000  68.935000 ;
      RECT  0.000000  68.935000 67.139000  69.085000 ;
      RECT  0.000000  69.085000 66.989000  69.235000 ;
      RECT  0.000000  69.235000 66.839000  69.385000 ;
      RECT  0.000000  69.385000 66.689000  69.535000 ;
      RECT  0.000000  69.535000 66.539000  69.685000 ;
      RECT  0.000000  69.685000 66.389000  69.835000 ;
      RECT  0.000000  69.835000 66.239000  69.985000 ;
      RECT  0.000000  69.985000 66.089000  70.135000 ;
      RECT  0.000000  70.135000 65.939000  70.285000 ;
      RECT  0.000000  70.285000 65.789000  70.435000 ;
      RECT  0.000000  70.435000 65.639000  70.585000 ;
      RECT  0.000000  70.585000 65.489000  70.735000 ;
      RECT  0.000000  70.735000 65.339000  70.885000 ;
      RECT  0.000000  70.885000 65.189000  71.035000 ;
      RECT  0.000000  71.035000 65.039000  71.185000 ;
      RECT  0.000000  71.185000 64.889000  71.335000 ;
      RECT  0.000000  71.335000 64.739000  71.485000 ;
      RECT  0.000000  71.485000 64.589000  71.635000 ;
      RECT  0.000000  71.635000 64.459000  71.765000 ;
      RECT  0.000000  71.764000  3.005000 196.995000 ;
      RECT  0.000000  71.806000 64.560000  94.945000 ;
      RECT  0.000000  94.945000 75.000000 200.000000 ;
      RECT  0.000000 196.995000 75.000000 200.000000 ;
      RECT  3.002000   3.002000  4.998000  14.375000 ;
      RECT  3.002000  14.375000  4.848000  14.525000 ;
      RECT  3.002000  14.375000  4.848000  14.525000 ;
      RECT  3.002000  14.525000  4.698000  14.675000 ;
      RECT  3.002000  14.525000  4.698000  14.675000 ;
      RECT  3.002000  14.675000  4.548000  14.825000 ;
      RECT  3.002000  14.675000  4.548000  14.825000 ;
      RECT  3.002000  14.825000  4.398000  14.975000 ;
      RECT  3.002000  14.825000  4.398000  14.975000 ;
      RECT  3.002000  14.975000  4.248000  15.125000 ;
      RECT  3.002000  14.975000  4.248000  15.125000 ;
      RECT  3.002000  15.125000  4.098000  15.275000 ;
      RECT  3.002000  15.125000  4.098000  15.275000 ;
      RECT  3.002000  15.275000  3.948000  15.425000 ;
      RECT  3.002000  15.275000  3.948000  15.425000 ;
      RECT  3.002000  15.425000  3.798000  15.575000 ;
      RECT  3.002000  15.425000  3.798000  15.575000 ;
      RECT  3.002000  15.575000  3.648000  15.725000 ;
      RECT  3.002000  15.575000  3.648000  15.725000 ;
      RECT  3.002000  15.725000  3.498000  15.875000 ;
      RECT  3.002000  15.725000  3.498000  15.875000 ;
      RECT  3.002000  15.875000  3.373000  16.000000 ;
      RECT  3.002000  15.875000  3.373000  16.000000 ;
      RECT  3.002000  16.000000  3.373000  32.915000 ;
      RECT  3.002000  32.915000  3.373000  33.065000 ;
      RECT  3.002000  32.915000  3.373000  33.065000 ;
      RECT  3.002000  33.065000  3.523000  33.215000 ;
      RECT  3.002000  33.065000  3.523000  33.215000 ;
      RECT  3.002000  33.215000  3.673000  33.365000 ;
      RECT  3.002000  33.215000  3.673000  33.365000 ;
      RECT  3.002000  33.365000  3.823000  33.515000 ;
      RECT  3.002000  33.365000  3.823000  33.515000 ;
      RECT  3.002000  33.515000  3.973000  33.665000 ;
      RECT  3.002000  33.515000  3.973000  33.665000 ;
      RECT  3.002000  33.665000  4.123000  33.815000 ;
      RECT  3.002000  33.665000  4.123000  33.815000 ;
      RECT  3.002000  33.815000  4.273000  33.965000 ;
      RECT  3.002000  33.815000  4.273000  33.965000 ;
      RECT  3.002000  33.965000  4.423000  34.115000 ;
      RECT  3.002000  33.965000  4.423000  34.115000 ;
      RECT  3.002000  34.115000  4.573000  34.265000 ;
      RECT  3.002000  34.115000  4.573000  34.265000 ;
      RECT  3.002000  34.265000  4.723000  34.415000 ;
      RECT  3.002000  34.265000  4.723000  34.415000 ;
      RECT  3.002000  34.415000  4.873000  34.565000 ;
      RECT  3.002000  34.415000  4.873000  34.565000 ;
      RECT  3.002000  34.565000  5.023000  34.715000 ;
      RECT  3.002000  34.565000  5.023000  34.715000 ;
      RECT  3.002000  34.715000  5.173000  34.865000 ;
      RECT  3.002000  34.715000  5.173000  34.865000 ;
      RECT  3.002000  34.865000  5.323000  35.015000 ;
      RECT  3.002000  34.865000  5.323000  35.015000 ;
      RECT  3.002000  35.015000  5.473000  35.165000 ;
      RECT  3.002000  35.015000  5.473000  35.165000 ;
      RECT  3.002000  35.165000  5.623000  35.315000 ;
      RECT  3.002000  35.165000  5.623000  35.315000 ;
      RECT  3.002000  35.315000  5.773000  35.465000 ;
      RECT  3.002000  35.315000  5.773000  35.465000 ;
      RECT  3.002000  35.465000  5.923000  35.615000 ;
      RECT  3.002000  35.465000  5.923000  35.615000 ;
      RECT  3.002000  35.615000  6.073000  35.765000 ;
      RECT  3.002000  35.615000  6.073000  35.765000 ;
      RECT  3.002000  35.765000  6.223000  35.915000 ;
      RECT  3.002000  35.765000  6.223000  35.915000 ;
      RECT  3.002000  35.915000  6.373000  36.065000 ;
      RECT  3.002000  35.915000  6.373000  36.065000 ;
      RECT  3.002000  36.065000  6.523000  36.215000 ;
      RECT  3.002000  36.065000  6.523000  36.215000 ;
      RECT  3.002000  36.215000  6.673000  36.365000 ;
      RECT  3.002000  36.215000  6.673000  36.365000 ;
      RECT  3.002000  36.365000  6.823000  36.515000 ;
      RECT  3.002000  36.365000  6.823000  36.515000 ;
      RECT  3.002000  36.515000  6.973000  36.665000 ;
      RECT  3.002000  36.515000  6.973000  36.665000 ;
      RECT  3.002000  36.665000  7.123000  36.815000 ;
      RECT  3.002000  36.665000  7.123000  36.815000 ;
      RECT  3.002000  36.815000  7.273000  36.965000 ;
      RECT  3.002000  36.815000  7.273000  36.965000 ;
      RECT  3.002000  36.965000  7.423000  37.115000 ;
      RECT  3.002000  36.965000  7.423000  37.115000 ;
      RECT  3.002000  37.115000  7.573000  37.265000 ;
      RECT  3.002000  37.115000  7.573000  37.265000 ;
      RECT  3.002000  37.265000  7.723000  37.415000 ;
      RECT  3.002000  37.265000  7.723000  37.415000 ;
      RECT  3.002000  37.415000  7.873000  37.525000 ;
      RECT  3.002000  37.415000  7.873000  37.525000 ;
      RECT  3.002000  37.527000 68.788000  63.190000 ;
      RECT  3.002000  63.190000 68.638000  63.340000 ;
      RECT  3.002000  63.190000 68.638000  63.340000 ;
      RECT  3.002000  63.340000 68.488000  63.490000 ;
      RECT  3.002000  63.340000 68.488000  63.490000 ;
      RECT  3.002000  63.490000 68.338000  63.640000 ;
      RECT  3.002000  63.490000 68.338000  63.640000 ;
      RECT  3.002000  63.640000 68.188000  63.790000 ;
      RECT  3.002000  63.640000 68.188000  63.790000 ;
      RECT  3.002000  63.790000 68.038000  63.940000 ;
      RECT  3.002000  63.790000 68.038000  63.940000 ;
      RECT  3.002000  63.940000 67.888000  64.090000 ;
      RECT  3.002000  63.940000 67.888000  64.090000 ;
      RECT  3.002000  64.090000 67.738000  64.240000 ;
      RECT  3.002000  64.090000 67.738000  64.240000 ;
      RECT  3.002000  64.240000 67.588000  64.390000 ;
      RECT  3.002000  64.240000 67.588000  64.390000 ;
      RECT  3.002000  64.390000 67.438000  64.540000 ;
      RECT  3.002000  64.390000 67.438000  64.540000 ;
      RECT  3.002000  64.540000 67.288000  64.690000 ;
      RECT  3.002000  64.540000 67.288000  64.690000 ;
      RECT  3.002000  64.690000 67.138000  64.840000 ;
      RECT  3.002000  64.690000 67.138000  64.840000 ;
      RECT  3.002000  64.840000 66.988000  64.990000 ;
      RECT  3.002000  64.840000 66.988000  64.990000 ;
      RECT  3.002000  64.990000 66.838000  65.140000 ;
      RECT  3.002000  64.990000 66.838000  65.140000 ;
      RECT  3.002000  65.140000 66.688000  65.290000 ;
      RECT  3.002000  65.140000 66.688000  65.290000 ;
      RECT  3.002000  65.290000 66.538000  65.440000 ;
      RECT  3.002000  65.290000 66.538000  65.440000 ;
      RECT  3.002000  65.440000 66.388000  65.590000 ;
      RECT  3.002000  65.440000 66.388000  65.590000 ;
      RECT  3.002000  65.590000 66.238000  65.740000 ;
      RECT  3.002000  65.590000 66.238000  65.740000 ;
      RECT  3.002000  65.740000 66.088000  65.890000 ;
      RECT  3.002000  65.740000 66.088000  65.890000 ;
      RECT  3.002000  65.890000 65.938000  66.040000 ;
      RECT  3.002000  65.890000 65.938000  66.040000 ;
      RECT  3.002000  66.040000 65.788000  66.190000 ;
      RECT  3.002000  66.040000 65.788000  66.190000 ;
      RECT  3.002000  66.190000 65.638000  66.340000 ;
      RECT  3.002000  66.190000 65.638000  66.340000 ;
      RECT  3.002000  66.340000 65.488000  66.490000 ;
      RECT  3.002000  66.340000 65.488000  66.490000 ;
      RECT  3.002000  66.490000 65.338000  66.640000 ;
      RECT  3.002000  66.490000 65.338000  66.640000 ;
      RECT  3.002000  66.640000 65.188000  66.790000 ;
      RECT  3.002000  66.640000 65.188000  66.790000 ;
      RECT  3.002000  66.790000 65.038000  66.940000 ;
      RECT  3.002000  66.790000 65.038000  66.940000 ;
      RECT  3.002000  66.940000 64.888000  67.090000 ;
      RECT  3.002000  66.940000 64.888000  67.090000 ;
      RECT  3.002000  67.090000 64.738000  67.240000 ;
      RECT  3.002000  67.090000 64.738000  67.240000 ;
      RECT  3.002000  67.240000 64.588000  67.390000 ;
      RECT  3.002000  67.240000 64.588000  67.390000 ;
      RECT  3.002000  67.390000 64.438000  67.540000 ;
      RECT  3.002000  67.390000 64.438000  67.540000 ;
      RECT  3.002000  67.540000 64.288000  67.690000 ;
      RECT  3.002000  67.540000 64.288000  67.690000 ;
      RECT  3.002000  67.690000 64.138000  67.840000 ;
      RECT  3.002000  67.690000 64.138000  67.840000 ;
      RECT  3.002000  67.840000 63.988000  67.990000 ;
      RECT  3.002000  67.840000 63.988000  67.990000 ;
      RECT  3.002000  67.990000 63.838000  68.140000 ;
      RECT  3.002000  67.990000 63.838000  68.140000 ;
      RECT  3.002000  68.140000 63.688000  68.290000 ;
      RECT  3.002000  68.140000 63.688000  68.290000 ;
      RECT  3.002000  68.290000 63.538000  68.440000 ;
      RECT  3.002000  68.290000 63.538000  68.440000 ;
      RECT  3.002000  68.440000 63.388000  68.590000 ;
      RECT  3.002000  68.440000 63.388000  68.590000 ;
      RECT  3.002000  68.590000 63.238000  68.740000 ;
      RECT  3.002000  68.590000 63.238000  68.740000 ;
      RECT  3.002000  68.740000 63.088000  68.890000 ;
      RECT  3.002000  68.740000 63.088000  68.890000 ;
      RECT  3.002000  68.890000 62.938000  69.040000 ;
      RECT  3.002000  68.890000 62.938000  69.040000 ;
      RECT  3.002000  69.040000 62.788000  69.190000 ;
      RECT  3.002000  69.040000 62.788000  69.190000 ;
      RECT  3.002000  69.190000 62.638000  69.340000 ;
      RECT  3.002000  69.190000 62.638000  69.340000 ;
      RECT  3.002000  69.340000 62.488000  69.490000 ;
      RECT  3.002000  69.340000 62.488000  69.490000 ;
      RECT  3.002000  69.490000 62.338000  69.640000 ;
      RECT  3.002000  69.490000 62.338000  69.640000 ;
      RECT  3.002000  69.640000 62.188000  69.790000 ;
      RECT  3.002000  69.640000 62.188000  69.790000 ;
      RECT  3.002000  69.790000 62.038000  69.940000 ;
      RECT  3.002000  69.790000 62.038000  69.940000 ;
      RECT  3.002000  69.940000 61.888000  70.090000 ;
      RECT  3.002000  69.940000 61.888000  70.090000 ;
      RECT  3.002000  70.090000 61.738000  70.240000 ;
      RECT  3.002000  70.090000 61.738000  70.240000 ;
      RECT  3.002000  70.240000 61.588000  70.390000 ;
      RECT  3.002000  70.240000 61.588000  70.390000 ;
      RECT  3.002000  70.390000 61.458000  70.520000 ;
      RECT  3.002000  70.390000 61.458000  70.520000 ;
      RECT  3.002000  70.520000 61.458000  98.047000 ;
      RECT  3.002000  98.047000 71.998000 196.998000 ;
      RECT  3.370000   3.005000  8.000000  15.619000 ;
      RECT  3.370000  15.619000  6.375000  17.244000 ;
      RECT  6.375000  34.525000 25.680000  37.527000 ;
      RECT  6.375000  37.527000 25.677000  37.530000 ;
      RECT  7.595000  17.744000 71.890000  31.171000 ;
      RECT  7.595000  31.171000 71.890000  33.095000 ;
      RECT  7.695000  17.786000 12.325000  28.124000 ;
      RECT  7.695000  28.124000 25.677000  29.993000 ;
      RECT  7.695000  29.993000 25.680000  31.129000 ;
      RECT  7.821000  17.660000 71.790000  17.785000 ;
      RECT  7.846000  31.129000 71.790000  31.280000 ;
      RECT  7.971000  17.510000 71.790000  17.660000 ;
      RECT  7.996000  31.280000 71.790000  31.430000 ;
      RECT  8.121000  17.360000 71.790000  17.510000 ;
      RECT  8.146000  31.430000 71.790000  31.580000 ;
      RECT  8.271000  17.210000 71.790000  17.360000 ;
      RECT  8.296000  31.580000 71.790000  31.730000 ;
      RECT  8.421000  17.060000 71.790000  17.210000 ;
      RECT  8.446000  31.730000 71.790000  31.880000 ;
      RECT  8.571000  16.910000 71.790000  17.060000 ;
      RECT  8.596000  31.880000 71.790000  32.030000 ;
      RECT  8.721000  16.760000 71.790000  16.910000 ;
      RECT  8.746000  32.030000 71.790000  32.180000 ;
      RECT  8.871000  16.610000 71.790000  16.760000 ;
      RECT  8.896000  32.180000 71.790000  32.330000 ;
      RECT  9.021000  16.460000 71.790000  16.610000 ;
      RECT  9.046000  32.330000 71.790000  32.480000 ;
      RECT  9.171000  16.310000 71.790000  16.460000 ;
      RECT  9.196000  32.480000 71.790000  32.630000 ;
      RECT  9.220000   0.000000 16.945000   3.435000 ;
      RECT  9.220000   3.435000 19.775000   7.274000 ;
      RECT  9.220000   7.274000 22.605000  10.104000 ;
      RECT  9.220000  10.104000 22.605000  12.565000 ;
      RECT  9.220000  12.565000 27.870000  15.070000 ;
      RECT  9.220000  15.070000 71.890000  16.119000 ;
      RECT  9.220000  16.119000 71.890000  17.744000 ;
      RECT  9.320000   0.000000 16.845000   7.316000 ;
      RECT  9.320000   0.000000 16.845000  10.146000 ;
      RECT  9.320000   3.535000 19.675000  12.665000 ;
      RECT  9.320000   7.316000 19.675000   7.465000 ;
      RECT  9.320000   7.465000 19.824000   7.615000 ;
      RECT  9.320000   7.615000 19.974000   7.765000 ;
      RECT  9.320000   7.765000 20.124000   7.915000 ;
      RECT  9.320000   7.915000 20.274000   8.065000 ;
      RECT  9.320000   8.065000 20.424000   8.215000 ;
      RECT  9.320000   8.215000 20.574000   8.365000 ;
      RECT  9.320000   8.365000 20.724000   8.515000 ;
      RECT  9.320000   8.515000 20.874000   8.665000 ;
      RECT  9.320000   8.665000 21.024000   8.815000 ;
      RECT  9.320000   8.815000 21.174000   8.965000 ;
      RECT  9.320000   8.965000 21.324000   9.115000 ;
      RECT  9.320000   9.115000 21.474000   9.265000 ;
      RECT  9.320000   9.265000 21.624000   9.415000 ;
      RECT  9.320000   9.415000 21.774000   9.565000 ;
      RECT  9.320000   9.565000 21.924000   9.715000 ;
      RECT  9.320000   9.715000 22.074000   9.865000 ;
      RECT  9.320000   9.865000 22.224000  10.015000 ;
      RECT  9.320000  10.015000 22.374000  10.145000 ;
      RECT  9.320000  12.665000 12.325000  17.786000 ;
      RECT  9.320000  16.161000 71.790000  16.310000 ;
      RECT  9.346000  32.630000 71.790000  32.780000 ;
      RECT  9.496000  32.780000 71.790000  32.930000 ;
      RECT  9.561000  32.930000 71.790000  32.995000 ;
      RECT 10.697000  19.030000 68.788000  29.885000 ;
      RECT 10.752000  29.885000 68.788000  29.940000 ;
      RECT 10.752000  29.885000 68.788000  29.940000 ;
      RECT 10.807000  18.920000 68.788000  19.030000 ;
      RECT 10.807000  18.920000 68.788000  19.030000 ;
      RECT 10.807000  29.940000 68.788000  29.995000 ;
      RECT 10.807000  29.940000 68.788000  29.995000 ;
      RECT 10.957000  18.770000 68.788000  18.920000 ;
      RECT 10.957000  18.770000 68.788000  18.920000 ;
      RECT 11.107000  18.620000 68.788000  18.770000 ;
      RECT 11.107000  18.620000 68.788000  18.770000 ;
      RECT 11.257000  18.470000 68.788000  18.620000 ;
      RECT 11.257000  18.470000 68.788000  18.620000 ;
      RECT 11.407000  18.320000 68.788000  18.470000 ;
      RECT 11.407000  18.320000 68.788000  18.470000 ;
      RECT 11.555000  18.172000 68.788000  18.320000 ;
      RECT 11.555000  18.172000 68.788000  18.320000 ;
      RECT 11.572000  18.155000 24.768000  18.170000 ;
      RECT 11.572000  18.155000 24.768000  18.170000 ;
      RECT 11.722000  18.005000 24.768000  18.155000 ;
      RECT 11.722000  18.005000 24.768000  18.155000 ;
      RECT 11.872000  17.855000 24.768000  18.005000 ;
      RECT 11.872000  17.855000 24.768000  18.005000 ;
      RECT 12.022000  17.705000 24.768000  17.855000 ;
      RECT 12.022000  17.705000 24.768000  17.855000 ;
      RECT 12.172000  17.555000 24.768000  17.705000 ;
      RECT 12.172000  17.555000 24.768000  17.705000 ;
      RECT 12.322000   3.002000 13.843000   6.537000 ;
      RECT 12.322000   6.537000 16.673000   8.560000 ;
      RECT 12.322000   8.560000 16.673000   8.710000 ;
      RECT 12.322000   8.560000 16.673000   8.710000 ;
      RECT 12.322000   8.710000 16.823000   8.860000 ;
      RECT 12.322000   8.710000 16.823000   8.860000 ;
      RECT 12.322000   8.860000 16.973000   9.010000 ;
      RECT 12.322000   8.860000 16.973000   9.010000 ;
      RECT 12.322000   9.010000 17.123000   9.160000 ;
      RECT 12.322000   9.010000 17.123000   9.160000 ;
      RECT 12.322000   9.160000 17.273000   9.310000 ;
      RECT 12.322000   9.160000 17.273000   9.310000 ;
      RECT 12.322000   9.310000 17.423000   9.460000 ;
      RECT 12.322000   9.310000 17.423000   9.460000 ;
      RECT 12.322000   9.460000 17.573000   9.610000 ;
      RECT 12.322000   9.460000 17.573000   9.610000 ;
      RECT 12.322000   9.610000 17.723000   9.760000 ;
      RECT 12.322000   9.610000 17.723000   9.760000 ;
      RECT 12.322000   9.760000 17.873000   9.910000 ;
      RECT 12.322000   9.760000 17.873000   9.910000 ;
      RECT 12.322000   9.910000 18.023000  10.060000 ;
      RECT 12.322000   9.910000 18.023000  10.060000 ;
      RECT 12.322000  10.060000 18.173000  10.210000 ;
      RECT 12.322000  10.060000 18.173000  10.210000 ;
      RECT 12.322000  10.210000 18.323000  10.360000 ;
      RECT 12.322000  10.210000 18.323000  10.360000 ;
      RECT 12.322000  10.360000 18.473000  10.510000 ;
      RECT 12.322000  10.360000 18.473000  10.510000 ;
      RECT 12.322000  10.510000 18.623000  10.660000 ;
      RECT 12.322000  10.510000 18.623000  10.660000 ;
      RECT 12.322000  10.660000 18.773000  10.810000 ;
      RECT 12.322000  10.660000 18.773000  10.810000 ;
      RECT 12.322000  10.810000 18.923000  10.960000 ;
      RECT 12.322000  10.810000 18.923000  10.960000 ;
      RECT 12.322000  10.960000 19.073000  11.110000 ;
      RECT 12.322000  10.960000 19.073000  11.110000 ;
      RECT 12.322000  11.110000 19.223000  11.260000 ;
      RECT 12.322000  11.110000 19.223000  11.260000 ;
      RECT 12.322000  11.260000 19.373000  11.390000 ;
      RECT 12.322000  11.260000 19.373000  11.390000 ;
      RECT 12.322000  11.390000 19.503000  15.667000 ;
      RECT 12.322000  15.667000 24.768000  17.405000 ;
      RECT 12.322000  17.405000 24.768000  17.555000 ;
      RECT 12.322000  17.405000 24.768000  17.555000 ;
      RECT 19.210000   0.000000 19.775000   3.435000 ;
      RECT 19.310000   0.000000 19.675000   3.535000 ;
      RECT 19.500000  10.146000 22.505000  12.665000 ;
      RECT 19.500000  12.665000 27.770000  15.170000 ;
      RECT 19.503000  15.170000 32.305000  18.172000 ;
      RECT 19.503000  18.172000 32.302000  18.175000 ;
      RECT 21.525000   0.000000 28.635000   6.546000 ;
      RECT 21.525000   6.546000 28.635000   9.371000 ;
      RECT 21.625000   0.000000 28.535000   3.005000 ;
      RECT 21.625000   3.005000 24.630000   3.499000 ;
      RECT 21.625000   3.499000 28.535000   6.504000 ;
      RECT 21.776000   6.504000 28.535000   6.655000 ;
      RECT 21.926000   6.655000 28.535000   6.805000 ;
      RECT 22.076000   6.805000 28.535000   6.955000 ;
      RECT 22.226000   6.955000 28.535000   7.105000 ;
      RECT 22.376000   7.105000 28.535000   7.255000 ;
      RECT 22.526000   7.255000 28.535000   7.405000 ;
      RECT 22.575000  33.095000 71.890000  34.425000 ;
      RECT 22.675000  31.129000 25.680000  34.525000 ;
      RECT 22.676000   7.405000 28.535000   7.555000 ;
      RECT 22.826000   7.555000 28.535000   7.705000 ;
      RECT 22.976000   7.705000 28.535000   7.855000 ;
      RECT 23.126000   7.855000 28.535000   8.005000 ;
      RECT 23.276000   8.005000 28.535000   8.155000 ;
      RECT 23.426000   8.155000 28.535000   8.305000 ;
      RECT 23.576000   8.305000 28.535000   8.455000 ;
      RECT 23.726000   8.455000 28.535000   8.605000 ;
      RECT 23.876000   8.605000 28.535000   8.755000 ;
      RECT 24.026000   8.755000 28.535000   8.905000 ;
      RECT 24.176000   8.905000 28.535000   9.055000 ;
      RECT 24.326000   9.055000 28.535000   9.205000 ;
      RECT 24.350000   9.371000 28.635000   9.721000 ;
      RECT 24.350000   9.721000 27.870000  10.486000 ;
      RECT 24.350000  10.486000 27.870000  12.565000 ;
      RECT 24.450000   9.329000 28.535000   9.679000 ;
      RECT 24.450000   9.679000 27.770000  12.665000 ;
      RECT 24.450000   9.679000 28.384000   9.830000 ;
      RECT 24.450000   9.830000 28.234000   9.980000 ;
      RECT 24.450000   9.980000 28.084000  10.130000 ;
      RECT 24.450000  10.130000 27.934000  10.280000 ;
      RECT 24.450000  10.280000 27.784000  10.430000 ;
      RECT 24.450000  10.430000 27.769000  10.445000 ;
      RECT 24.451000   9.205000 28.535000   9.330000 ;
      RECT 24.627000   3.002000 25.533000   5.260000 ;
      RECT 24.627000   3.002000 25.533000   5.260000 ;
      RECT 24.768000  18.175000 32.302000  20.791000 ;
      RECT 25.530000   3.005000 28.535000   3.499000 ;
      RECT 25.677000  29.993000 68.788000  37.527000 ;
      RECT 29.200000  11.034000 71.890000  15.070000 ;
      RECT 29.300000  11.076000 33.067000  14.081000 ;
      RECT 29.300000  14.081000 32.305000  15.170000 ;
      RECT 29.316000  11.060000 71.790000  11.075000 ;
      RECT 29.466000  10.910000 71.790000  11.060000 ;
      RECT 29.616000  10.760000 71.790000  10.910000 ;
      RECT 29.766000  10.610000 71.790000  10.760000 ;
      RECT 29.916000  10.460000 71.790000  10.610000 ;
      RECT 29.965000   0.000000 71.890000  10.269000 ;
      RECT 29.965000  10.269000 71.890000  11.034000 ;
      RECT 30.065000   0.000000 71.790000   3.005000 ;
      RECT 30.065000   3.005000 33.070000  11.076000 ;
      RECT 30.065000  10.311000 71.790000  10.460000 ;
      RECT 32.302000  12.320000 68.788000  18.172000 ;
      RECT 32.317000  12.305000 68.788000  12.320000 ;
      RECT 32.317000  12.305000 68.788000  12.320000 ;
      RECT 32.467000  12.155000 68.788000  12.305000 ;
      RECT 32.467000  12.155000 68.788000  12.305000 ;
      RECT 32.617000  12.005000 68.788000  12.155000 ;
      RECT 32.617000  12.005000 68.788000  12.155000 ;
      RECT 32.767000  11.855000 68.788000  12.005000 ;
      RECT 32.767000  11.855000 68.788000  12.005000 ;
      RECT 32.917000  11.705000 68.788000  11.855000 ;
      RECT 32.917000  11.705000 68.788000  11.855000 ;
      RECT 33.067000   3.002000 68.788000  11.555000 ;
      RECT 33.067000  11.555000 68.788000  11.705000 ;
      RECT 33.067000  11.555000 68.788000  11.705000 ;
      RECT 61.455000  71.764000 64.460000  95.045000 ;
      RECT 61.458000  95.045000 69.392000  98.050000 ;
      RECT 66.290000  72.524000 75.000000  94.945000 ;
      RECT 66.390000  72.566000 70.636000  75.571000 ;
      RECT 66.390000  75.571000 69.395000  95.045000 ;
      RECT 66.526000  72.430000 75.000000  72.565000 ;
      RECT 66.676000  72.280000 75.000000  72.430000 ;
      RECT 66.826000  72.130000 75.000000  72.280000 ;
      RECT 66.976000  71.980000 75.000000  72.130000 ;
      RECT 67.126000  71.830000 75.000000  71.980000 ;
      RECT 67.276000  71.680000 75.000000  71.830000 ;
      RECT 67.426000  71.530000 75.000000  71.680000 ;
      RECT 67.544000  61.429000 71.790000  64.434000 ;
      RECT 67.576000  71.380000 75.000000  71.530000 ;
      RECT 67.726000  71.230000 75.000000  71.380000 ;
      RECT 67.876000  71.080000 75.000000  71.230000 ;
      RECT 68.026000  70.930000 75.000000  71.080000 ;
      RECT 68.176000  70.780000 75.000000  70.930000 ;
      RECT 68.326000  70.630000 75.000000  70.780000 ;
      RECT 68.476000  70.480000 75.000000  70.630000 ;
      RECT 68.626000  70.330000 75.000000  70.480000 ;
      RECT 68.776000  70.180000 75.000000  70.330000 ;
      RECT 68.785000   3.005000 71.790000  61.429000 ;
      RECT 68.926000  70.030000 75.000000  70.180000 ;
      RECT 69.076000  69.880000 75.000000  70.030000 ;
      RECT 69.226000  69.730000 75.000000  69.880000 ;
      RECT 69.376000  69.580000 75.000000  69.730000 ;
      RECT 69.392000  73.810000 71.998000  98.047000 ;
      RECT 69.447000  73.755000 71.998000  73.810000 ;
      RECT 69.447000  73.755000 71.998000  73.810000 ;
      RECT 69.526000  69.430000 75.000000  69.580000 ;
      RECT 69.597000  73.605000 71.998000  73.755000 ;
      RECT 69.597000  73.605000 71.998000  73.755000 ;
      RECT 69.676000  69.280000 75.000000  69.430000 ;
      RECT 69.747000  73.455000 71.998000  73.605000 ;
      RECT 69.747000  73.455000 71.998000  73.605000 ;
      RECT 69.826000  69.130000 75.000000  69.280000 ;
      RECT 69.897000  73.305000 71.998000  73.455000 ;
      RECT 69.897000  73.305000 71.998000  73.455000 ;
      RECT 69.976000  68.980000 75.000000  69.130000 ;
      RECT 70.047000  73.155000 71.998000  73.305000 ;
      RECT 70.047000  73.155000 71.998000  73.305000 ;
      RECT 70.126000  68.830000 75.000000  68.980000 ;
      RECT 70.197000  73.005000 71.998000  73.155000 ;
      RECT 70.197000  73.005000 71.998000  73.155000 ;
      RECT 70.276000  68.680000 75.000000  68.830000 ;
      RECT 70.347000  72.855000 71.998000  73.005000 ;
      RECT 70.347000  72.855000 71.998000  73.005000 ;
      RECT 70.426000  68.530000 75.000000  68.680000 ;
      RECT 70.497000  72.705000 71.998000  72.855000 ;
      RECT 70.497000  72.705000 71.998000  72.855000 ;
      RECT 70.576000  68.380000 75.000000  68.530000 ;
      RECT 70.647000  72.555000 71.998000  72.705000 ;
      RECT 70.647000  72.555000 71.998000  72.705000 ;
      RECT 70.726000  68.230000 75.000000  68.380000 ;
      RECT 70.797000  72.405000 71.998000  72.555000 ;
      RECT 70.797000  72.405000 71.998000  72.555000 ;
      RECT 70.876000  68.080000 75.000000  68.230000 ;
      RECT 70.947000  72.255000 71.998000  72.405000 ;
      RECT 70.947000  72.255000 71.998000  72.405000 ;
      RECT 71.026000  67.930000 75.000000  68.080000 ;
      RECT 71.097000  72.105000 71.998000  72.255000 ;
      RECT 71.097000  72.105000 71.998000  72.255000 ;
      RECT 71.176000  67.780000 75.000000  67.930000 ;
      RECT 71.247000  71.955000 71.998000  72.105000 ;
      RECT 71.247000  71.955000 71.998000  72.105000 ;
      RECT 71.326000  67.630000 75.000000  67.780000 ;
      RECT 71.397000  71.805000 71.998000  71.955000 ;
      RECT 71.397000  71.805000 71.998000  71.955000 ;
      RECT 71.476000  67.480000 75.000000  67.630000 ;
      RECT 71.547000  71.655000 71.998000  71.805000 ;
      RECT 71.547000  71.655000 71.998000  71.805000 ;
      RECT 71.626000  67.330000 75.000000  67.480000 ;
      RECT 71.697000  71.505000 71.998000  71.655000 ;
      RECT 71.697000  71.505000 71.998000  71.655000 ;
      RECT 71.776000  67.180000 75.000000  67.330000 ;
      RECT 71.847000  71.355000 71.998000  71.505000 ;
      RECT 71.847000  71.355000 71.998000  71.505000 ;
      RECT 71.926000  67.030000 75.000000  67.180000 ;
      RECT 71.995000  72.566000 75.000000 196.995000 ;
      RECT 72.076000  66.880000 75.000000  67.030000 ;
      RECT 72.226000  66.730000 75.000000  66.880000 ;
      RECT 72.376000  66.580000 75.000000  66.730000 ;
      RECT 72.526000  66.430000 75.000000  66.580000 ;
      RECT 72.676000  66.280000 75.000000  66.430000 ;
      RECT 72.826000  66.130000 75.000000  66.280000 ;
      RECT 72.976000  65.980000 75.000000  66.130000 ;
      RECT 73.126000  65.830000 75.000000  65.980000 ;
      RECT 73.276000  65.680000 75.000000  65.830000 ;
      RECT 73.426000  65.530000 75.000000  65.680000 ;
      RECT 73.560000   0.000000 75.000000  49.196000 ;
      RECT 73.560000  49.196000 75.000000  49.861000 ;
      RECT 73.576000  65.380000 75.000000  65.530000 ;
      RECT 73.660000   0.000000 75.000000  49.154000 ;
      RECT 73.726000  65.230000 75.000000  65.380000 ;
      RECT 73.811000  49.154000 75.000000  49.305000 ;
      RECT 73.876000  65.080000 75.000000  65.230000 ;
      RECT 73.961000  49.305000 75.000000  49.455000 ;
      RECT 74.026000  64.930000 75.000000  65.080000 ;
      RECT 74.111000  49.455000 75.000000  49.605000 ;
      RECT 74.176000  64.780000 75.000000  64.930000 ;
      RECT 74.225000  49.861000 75.000000  64.589000 ;
      RECT 74.225000  64.589000 75.000000  72.524000 ;
      RECT 74.261000  49.605000 75.000000  49.755000 ;
      RECT 74.325000  49.819000 75.000000  64.631000 ;
      RECT 74.325000  64.631000 75.000000  64.780000 ;
      RECT 74.326000  49.755000 75.000000  49.820000 ;
    LAYER met4 ;
      RECT  0.000000   0.000000  1.670000   1.635000 ;
      RECT  0.000000   0.000000 75.000000   1.635000 ;
      RECT  0.000000   7.885000  1.670000   8.485000 ;
      RECT  0.000000   7.885000 75.000000   8.485000 ;
      RECT  0.000000  13.935000  1.365000  14.535000 ;
      RECT  0.000000  13.935000 75.000000  14.535000 ;
      RECT  0.000000  18.785000  1.365000  19.385000 ;
      RECT  0.000000  18.785000 75.000000  19.385000 ;
      RECT  0.000000  24.835000  1.670000  25.435000 ;
      RECT  0.000000  24.835000 75.000000  25.435000 ;
      RECT  0.000000  30.885000  1.670000  31.485000 ;
      RECT  0.000000  30.885000 75.000000  31.485000 ;
      RECT  0.000000  35.735000  1.670000  36.335000 ;
      RECT  0.000000  35.735000 75.000000  36.335000 ;
      RECT  0.000000  40.585000  1.670000  41.185000 ;
      RECT  0.000000  40.585000 75.000000  41.185000 ;
      RECT  0.000000  46.635000  1.670000  47.335000 ;
      RECT  0.000000  46.635000 75.000000  47.435000 ;
      RECT  0.000000  57.035000 75.000000  57.835000 ;
      RECT  0.000000  57.135000  1.670000  57.835000 ;
      RECT  0.000000  63.085000  1.670000  63.685000 ;
      RECT  0.000000  63.085000 75.000000  63.685000 ;
      RECT  0.000000  68.935000  1.670000  69.635000 ;
      RECT  0.000000  68.935000 75.000000  69.635000 ;
      RECT  0.000000  95.400000 75.000000 175.385000 ;
      RECT  1.365000  13.935000 73.635000  19.385000 ;
      RECT  1.570000  47.435000 73.430000  57.035000 ;
      RECT  1.670000   0.000000 73.330000  13.935000 ;
      RECT  1.670000  19.385000 73.330000  41.230000 ;
      RECT  1.670000  36.335000 73.330000  41.230000 ;
      RECT  1.670000  36.335000 73.330000  41.230000 ;
      RECT  1.670000  41.185000 75.000000  41.255000 ;
      RECT  1.670000  41.230000 73.255000  41.255000 ;
      RECT  1.670000  46.570000 73.255000  46.590000 ;
      RECT  1.670000  46.570000 73.255000  57.135000 ;
      RECT  1.670000  46.570000 75.000000  46.635000 ;
      RECT  1.670000  46.590000 73.330000  57.135000 ;
      RECT  1.670000  46.590000 73.330000  57.135000 ;
      RECT  1.670000  46.590000 73.330000  95.400000 ;
      RECT  1.670000 175.385000 73.330000 200.000000 ;
      RECT  4.120000  41.230000 73.255000  46.570000 ;
      RECT  4.120000  41.255000 73.255000  46.570000 ;
      RECT  4.120000  41.255000 73.255000  57.135000 ;
      RECT  4.120000  41.255000 75.000000  41.285000 ;
      RECT  4.120000  41.285000 73.430000  41.330000 ;
      RECT  4.120000  41.330000 73.355000  46.490000 ;
      RECT  4.120000  46.490000 73.430000  46.535000 ;
      RECT  4.120000  46.535000 75.000000  46.570000 ;
      RECT 73.330000   0.000000 75.000000   1.635000 ;
      RECT 73.330000   7.885000 75.000000   8.485000 ;
      RECT 73.330000  24.835000 75.000000  25.435000 ;
      RECT 73.330000  30.885000 75.000000  31.485000 ;
      RECT 73.330000  35.735000 75.000000  36.335000 ;
      RECT 73.330000  40.585000 75.000000  41.185000 ;
      RECT 73.330000  46.635000 75.000000  47.335000 ;
      RECT 73.330000  57.135000 75.000000  57.835000 ;
      RECT 73.330000  63.085000 75.000000  63.685000 ;
      RECT 73.330000  68.935000 75.000000  69.635000 ;
      RECT 73.635000  13.935000 75.000000  14.535000 ;
      RECT 73.635000  18.785000 75.000000  19.385000 ;
    LAYER met5 ;
      RECT  0.000000   0.000000 75.000000   1.335000 ;
      RECT  0.000000  36.035000 75.000000  36.040000 ;
      RECT  0.000000  95.785000 75.000000 126.315000 ;
      RECT  0.000000 126.315000 28.895000 146.425000 ;
      RECT  0.000000 146.425000 75.000000 174.985000 ;
      RECT  1.765000  14.235000 73.235000  19.085000 ;
      RECT  2.070000   1.335000 72.930000  14.235000 ;
      RECT  2.070000  19.085000 72.930000  95.785000 ;
      RECT  2.070000 174.985000 72.930000 200.000000 ;
      RECT 42.790000 126.315000 75.000000 146.425000 ;
  END
END sky130_fd_io__top_xres4v2
END LIBRARY
