# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__overlay_vccd_lvc
  CLASS BLOCK ;
  FOREIGN sky130_fd_io__overlay_vccd_lvc ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  75.00000 BY  198.0000 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.630000 10.340000 0.950000 10.660000 ;
      LAYER met4 ;
        RECT 0.630000 10.340000 0.950000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 10.770000 0.950000 11.090000 ;
      LAYER met4 ;
        RECT 0.630000 10.770000 0.950000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 11.200000 0.950000 11.520000 ;
      LAYER met4 ;
        RECT 0.630000 11.200000 0.950000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 6.900000 0.950000 7.220000 ;
      LAYER met4 ;
        RECT 0.630000 6.900000 0.950000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 7.330000 0.950000 7.650000 ;
      LAYER met4 ;
        RECT 0.630000 7.330000 0.950000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 7.760000 0.950000 8.080000 ;
      LAYER met4 ;
        RECT 0.630000 7.760000 0.950000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 8.190000 0.950000 8.510000 ;
      LAYER met4 ;
        RECT 0.630000 8.190000 0.950000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 8.620000 0.950000 8.940000 ;
      LAYER met4 ;
        RECT 0.630000 8.620000 0.950000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 9.050000 0.950000 9.370000 ;
      LAYER met4 ;
        RECT 0.630000 9.050000 0.950000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 9.480000 0.950000 9.800000 ;
      LAYER met4 ;
        RECT 0.630000 9.480000 0.950000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 9.910000 0.950000 10.230000 ;
      LAYER met4 ;
        RECT 0.630000 9.910000 0.950000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040000 10.340000 1.360000 10.660000 ;
      LAYER met4 ;
        RECT 1.040000 10.340000 1.360000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040000 10.770000 1.360000 11.090000 ;
      LAYER met4 ;
        RECT 1.040000 10.770000 1.360000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040000 11.200000 1.360000 11.520000 ;
      LAYER met4 ;
        RECT 1.040000 11.200000 1.360000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040000 6.900000 1.360000 7.220000 ;
      LAYER met4 ;
        RECT 1.040000 6.900000 1.360000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040000 7.330000 1.360000 7.650000 ;
      LAYER met4 ;
        RECT 1.040000 7.330000 1.360000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040000 7.760000 1.360000 8.080000 ;
      LAYER met4 ;
        RECT 1.040000 7.760000 1.360000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040000 8.190000 1.360000 8.510000 ;
      LAYER met4 ;
        RECT 1.040000 8.190000 1.360000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040000 8.620000 1.360000 8.940000 ;
      LAYER met4 ;
        RECT 1.040000 8.620000 1.360000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040000 9.050000 1.360000 9.370000 ;
      LAYER met4 ;
        RECT 1.040000 9.050000 1.360000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040000 9.480000 1.360000 9.800000 ;
      LAYER met4 ;
        RECT 1.040000 9.480000 1.360000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040000 9.910000 1.360000 10.230000 ;
      LAYER met4 ;
        RECT 1.040000 9.910000 1.360000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450000 10.340000 1.770000 10.660000 ;
      LAYER met4 ;
        RECT 1.450000 10.340000 1.770000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450000 10.770000 1.770000 11.090000 ;
      LAYER met4 ;
        RECT 1.450000 10.770000 1.770000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450000 11.200000 1.770000 11.520000 ;
      LAYER met4 ;
        RECT 1.450000 11.200000 1.770000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450000 6.900000 1.770000 7.220000 ;
      LAYER met4 ;
        RECT 1.450000 6.900000 1.770000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450000 7.330000 1.770000 7.650000 ;
      LAYER met4 ;
        RECT 1.450000 7.330000 1.770000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450000 7.760000 1.770000 8.080000 ;
      LAYER met4 ;
        RECT 1.450000 7.760000 1.770000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450000 8.190000 1.770000 8.510000 ;
      LAYER met4 ;
        RECT 1.450000 8.190000 1.770000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450000 8.620000 1.770000 8.940000 ;
      LAYER met4 ;
        RECT 1.450000 8.620000 1.770000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450000 9.050000 1.770000 9.370000 ;
      LAYER met4 ;
        RECT 1.450000 9.050000 1.770000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450000 9.480000 1.770000 9.800000 ;
      LAYER met4 ;
        RECT 1.450000 9.480000 1.770000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450000 9.910000 1.770000 10.230000 ;
      LAYER met4 ;
        RECT 1.450000 9.910000 1.770000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860000 10.340000 2.180000 10.660000 ;
      LAYER met4 ;
        RECT 1.860000 10.340000 2.180000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860000 10.770000 2.180000 11.090000 ;
      LAYER met4 ;
        RECT 1.860000 10.770000 2.180000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860000 11.200000 2.180000 11.520000 ;
      LAYER met4 ;
        RECT 1.860000 11.200000 2.180000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860000 6.900000 2.180000 7.220000 ;
      LAYER met4 ;
        RECT 1.860000 6.900000 2.180000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860000 7.330000 2.180000 7.650000 ;
      LAYER met4 ;
        RECT 1.860000 7.330000 2.180000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860000 7.760000 2.180000 8.080000 ;
      LAYER met4 ;
        RECT 1.860000 7.760000 2.180000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860000 8.190000 2.180000 8.510000 ;
      LAYER met4 ;
        RECT 1.860000 8.190000 2.180000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860000 8.620000 2.180000 8.940000 ;
      LAYER met4 ;
        RECT 1.860000 8.620000 2.180000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860000 9.050000 2.180000 9.370000 ;
      LAYER met4 ;
        RECT 1.860000 9.050000 2.180000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860000 9.480000 2.180000 9.800000 ;
      LAYER met4 ;
        RECT 1.860000 9.480000 2.180000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860000 9.910000 2.180000 10.230000 ;
      LAYER met4 ;
        RECT 1.860000 9.910000 2.180000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380000 10.340000 10.700000 10.660000 ;
      LAYER met4 ;
        RECT 10.380000 10.340000 10.700000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380000 10.770000 10.700000 11.090000 ;
      LAYER met4 ;
        RECT 10.380000 10.770000 10.700000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380000 11.200000 10.700000 11.520000 ;
      LAYER met4 ;
        RECT 10.380000 11.200000 10.700000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380000 6.900000 10.700000 7.220000 ;
      LAYER met4 ;
        RECT 10.380000 6.900000 10.700000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380000 7.330000 10.700000 7.650000 ;
      LAYER met4 ;
        RECT 10.380000 7.330000 10.700000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380000 7.760000 10.700000 8.080000 ;
      LAYER met4 ;
        RECT 10.380000 7.760000 10.700000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380000 8.190000 10.700000 8.510000 ;
      LAYER met4 ;
        RECT 10.380000 8.190000 10.700000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380000 8.620000 10.700000 8.940000 ;
      LAYER met4 ;
        RECT 10.380000 8.620000 10.700000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380000 9.050000 10.700000 9.370000 ;
      LAYER met4 ;
        RECT 10.380000 9.050000 10.700000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380000 9.480000 10.700000 9.800000 ;
      LAYER met4 ;
        RECT 10.380000 9.480000 10.700000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380000 9.910000 10.700000 10.230000 ;
      LAYER met4 ;
        RECT 10.380000 9.910000 10.700000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 10.340000 11.105000 10.660000 ;
      LAYER met4 ;
        RECT 10.785000 10.340000 11.105000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 10.770000 11.105000 11.090000 ;
      LAYER met4 ;
        RECT 10.785000 10.770000 11.105000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 11.200000 11.105000 11.520000 ;
      LAYER met4 ;
        RECT 10.785000 11.200000 11.105000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 6.900000 11.105000 7.220000 ;
      LAYER met4 ;
        RECT 10.785000 6.900000 11.105000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 7.330000 11.105000 7.650000 ;
      LAYER met4 ;
        RECT 10.785000 7.330000 11.105000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 7.760000 11.105000 8.080000 ;
      LAYER met4 ;
        RECT 10.785000 7.760000 11.105000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 8.190000 11.105000 8.510000 ;
      LAYER met4 ;
        RECT 10.785000 8.190000 11.105000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 8.620000 11.105000 8.940000 ;
      LAYER met4 ;
        RECT 10.785000 8.620000 11.105000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 9.050000 11.105000 9.370000 ;
      LAYER met4 ;
        RECT 10.785000 9.050000 11.105000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 9.480000 11.105000 9.800000 ;
      LAYER met4 ;
        RECT 10.785000 9.480000 11.105000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 9.910000 11.105000 10.230000 ;
      LAYER met4 ;
        RECT 10.785000 9.910000 11.105000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190000 10.340000 11.510000 10.660000 ;
      LAYER met4 ;
        RECT 11.190000 10.340000 11.510000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190000 10.770000 11.510000 11.090000 ;
      LAYER met4 ;
        RECT 11.190000 10.770000 11.510000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190000 11.200000 11.510000 11.520000 ;
      LAYER met4 ;
        RECT 11.190000 11.200000 11.510000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190000 6.900000 11.510000 7.220000 ;
      LAYER met4 ;
        RECT 11.190000 6.900000 11.510000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190000 7.330000 11.510000 7.650000 ;
      LAYER met4 ;
        RECT 11.190000 7.330000 11.510000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190000 7.760000 11.510000 8.080000 ;
      LAYER met4 ;
        RECT 11.190000 7.760000 11.510000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190000 8.190000 11.510000 8.510000 ;
      LAYER met4 ;
        RECT 11.190000 8.190000 11.510000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190000 8.620000 11.510000 8.940000 ;
      LAYER met4 ;
        RECT 11.190000 8.620000 11.510000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190000 9.050000 11.510000 9.370000 ;
      LAYER met4 ;
        RECT 11.190000 9.050000 11.510000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190000 9.480000 11.510000 9.800000 ;
      LAYER met4 ;
        RECT 11.190000 9.480000 11.510000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190000 9.910000 11.510000 10.230000 ;
      LAYER met4 ;
        RECT 11.190000 9.910000 11.510000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595000 10.340000 11.915000 10.660000 ;
      LAYER met4 ;
        RECT 11.595000 10.340000 11.915000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595000 10.770000 11.915000 11.090000 ;
      LAYER met4 ;
        RECT 11.595000 10.770000 11.915000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595000 11.200000 11.915000 11.520000 ;
      LAYER met4 ;
        RECT 11.595000 11.200000 11.915000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595000 6.900000 11.915000 7.220000 ;
      LAYER met4 ;
        RECT 11.595000 6.900000 11.915000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595000 7.330000 11.915000 7.650000 ;
      LAYER met4 ;
        RECT 11.595000 7.330000 11.915000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595000 7.760000 11.915000 8.080000 ;
      LAYER met4 ;
        RECT 11.595000 7.760000 11.915000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595000 8.190000 11.915000 8.510000 ;
      LAYER met4 ;
        RECT 11.595000 8.190000 11.915000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595000 8.620000 11.915000 8.940000 ;
      LAYER met4 ;
        RECT 11.595000 8.620000 11.915000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595000 9.050000 11.915000 9.370000 ;
      LAYER met4 ;
        RECT 11.595000 9.050000 11.915000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595000 9.480000 11.915000 9.800000 ;
      LAYER met4 ;
        RECT 11.595000 9.480000 11.915000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595000 9.910000 11.915000 10.230000 ;
      LAYER met4 ;
        RECT 11.595000 9.910000 11.915000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000000 10.340000 12.320000 10.660000 ;
      LAYER met4 ;
        RECT 12.000000 10.340000 12.320000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000000 10.770000 12.320000 11.090000 ;
      LAYER met4 ;
        RECT 12.000000 10.770000 12.320000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000000 11.200000 12.320000 11.520000 ;
      LAYER met4 ;
        RECT 12.000000 11.200000 12.320000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000000 6.900000 12.320000 7.220000 ;
      LAYER met4 ;
        RECT 12.000000 6.900000 12.320000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000000 7.330000 12.320000 7.650000 ;
      LAYER met4 ;
        RECT 12.000000 7.330000 12.320000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000000 7.760000 12.320000 8.080000 ;
      LAYER met4 ;
        RECT 12.000000 7.760000 12.320000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000000 8.190000 12.320000 8.510000 ;
      LAYER met4 ;
        RECT 12.000000 8.190000 12.320000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000000 8.620000 12.320000 8.940000 ;
      LAYER met4 ;
        RECT 12.000000 8.620000 12.320000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000000 9.050000 12.320000 9.370000 ;
      LAYER met4 ;
        RECT 12.000000 9.050000 12.320000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000000 9.480000 12.320000 9.800000 ;
      LAYER met4 ;
        RECT 12.000000 9.480000 12.320000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000000 9.910000 12.320000 10.230000 ;
      LAYER met4 ;
        RECT 12.000000 9.910000 12.320000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405000 10.340000 12.725000 10.660000 ;
      LAYER met4 ;
        RECT 12.405000 10.340000 12.725000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405000 10.770000 12.725000 11.090000 ;
      LAYER met4 ;
        RECT 12.405000 10.770000 12.725000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405000 11.200000 12.725000 11.520000 ;
      LAYER met4 ;
        RECT 12.405000 11.200000 12.725000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405000 6.900000 12.725000 7.220000 ;
      LAYER met4 ;
        RECT 12.405000 6.900000 12.725000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405000 7.330000 12.725000 7.650000 ;
      LAYER met4 ;
        RECT 12.405000 7.330000 12.725000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405000 7.760000 12.725000 8.080000 ;
      LAYER met4 ;
        RECT 12.405000 7.760000 12.725000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405000 8.190000 12.725000 8.510000 ;
      LAYER met4 ;
        RECT 12.405000 8.190000 12.725000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405000 8.620000 12.725000 8.940000 ;
      LAYER met4 ;
        RECT 12.405000 8.620000 12.725000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405000 9.050000 12.725000 9.370000 ;
      LAYER met4 ;
        RECT 12.405000 9.050000 12.725000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405000 9.480000 12.725000 9.800000 ;
      LAYER met4 ;
        RECT 12.405000 9.480000 12.725000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405000 9.910000 12.725000 10.230000 ;
      LAYER met4 ;
        RECT 12.405000 9.910000 12.725000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810000 10.340000 13.130000 10.660000 ;
      LAYER met4 ;
        RECT 12.810000 10.340000 13.130000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810000 10.770000 13.130000 11.090000 ;
      LAYER met4 ;
        RECT 12.810000 10.770000 13.130000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810000 11.200000 13.130000 11.520000 ;
      LAYER met4 ;
        RECT 12.810000 11.200000 13.130000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810000 6.900000 13.130000 7.220000 ;
      LAYER met4 ;
        RECT 12.810000 6.900000 13.130000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810000 7.330000 13.130000 7.650000 ;
      LAYER met4 ;
        RECT 12.810000 7.330000 13.130000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810000 7.760000 13.130000 8.080000 ;
      LAYER met4 ;
        RECT 12.810000 7.760000 13.130000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810000 8.190000 13.130000 8.510000 ;
      LAYER met4 ;
        RECT 12.810000 8.190000 13.130000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810000 8.620000 13.130000 8.940000 ;
      LAYER met4 ;
        RECT 12.810000 8.620000 13.130000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810000 9.050000 13.130000 9.370000 ;
      LAYER met4 ;
        RECT 12.810000 9.050000 13.130000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810000 9.480000 13.130000 9.800000 ;
      LAYER met4 ;
        RECT 12.810000 9.480000 13.130000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810000 9.910000 13.130000 10.230000 ;
      LAYER met4 ;
        RECT 12.810000 9.910000 13.130000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215000 10.340000 13.535000 10.660000 ;
      LAYER met4 ;
        RECT 13.215000 10.340000 13.535000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215000 10.770000 13.535000 11.090000 ;
      LAYER met4 ;
        RECT 13.215000 10.770000 13.535000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215000 11.200000 13.535000 11.520000 ;
      LAYER met4 ;
        RECT 13.215000 11.200000 13.535000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215000 6.900000 13.535000 7.220000 ;
      LAYER met4 ;
        RECT 13.215000 6.900000 13.535000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215000 7.330000 13.535000 7.650000 ;
      LAYER met4 ;
        RECT 13.215000 7.330000 13.535000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215000 7.760000 13.535000 8.080000 ;
      LAYER met4 ;
        RECT 13.215000 7.760000 13.535000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215000 8.190000 13.535000 8.510000 ;
      LAYER met4 ;
        RECT 13.215000 8.190000 13.535000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215000 8.620000 13.535000 8.940000 ;
      LAYER met4 ;
        RECT 13.215000 8.620000 13.535000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215000 9.050000 13.535000 9.370000 ;
      LAYER met4 ;
        RECT 13.215000 9.050000 13.535000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215000 9.480000 13.535000 9.800000 ;
      LAYER met4 ;
        RECT 13.215000 9.480000 13.535000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215000 9.910000 13.535000 10.230000 ;
      LAYER met4 ;
        RECT 13.215000 9.910000 13.535000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620000 10.340000 13.940000 10.660000 ;
      LAYER met4 ;
        RECT 13.620000 10.340000 13.940000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620000 10.770000 13.940000 11.090000 ;
      LAYER met4 ;
        RECT 13.620000 10.770000 13.940000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620000 11.200000 13.940000 11.520000 ;
      LAYER met4 ;
        RECT 13.620000 11.200000 13.940000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620000 6.900000 13.940000 7.220000 ;
      LAYER met4 ;
        RECT 13.620000 6.900000 13.940000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620000 7.330000 13.940000 7.650000 ;
      LAYER met4 ;
        RECT 13.620000 7.330000 13.940000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620000 7.760000 13.940000 8.080000 ;
      LAYER met4 ;
        RECT 13.620000 7.760000 13.940000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620000 8.190000 13.940000 8.510000 ;
      LAYER met4 ;
        RECT 13.620000 8.190000 13.940000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620000 8.620000 13.940000 8.940000 ;
      LAYER met4 ;
        RECT 13.620000 8.620000 13.940000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620000 9.050000 13.940000 9.370000 ;
      LAYER met4 ;
        RECT 13.620000 9.050000 13.940000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620000 9.480000 13.940000 9.800000 ;
      LAYER met4 ;
        RECT 13.620000 9.480000 13.940000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620000 9.910000 13.940000 10.230000 ;
      LAYER met4 ;
        RECT 13.620000 9.910000 13.940000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025000 10.340000 14.345000 10.660000 ;
      LAYER met4 ;
        RECT 14.025000 10.340000 14.345000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025000 10.770000 14.345000 11.090000 ;
      LAYER met4 ;
        RECT 14.025000 10.770000 14.345000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025000 11.200000 14.345000 11.520000 ;
      LAYER met4 ;
        RECT 14.025000 11.200000 14.345000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025000 6.900000 14.345000 7.220000 ;
      LAYER met4 ;
        RECT 14.025000 6.900000 14.345000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025000 7.330000 14.345000 7.650000 ;
      LAYER met4 ;
        RECT 14.025000 7.330000 14.345000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025000 7.760000 14.345000 8.080000 ;
      LAYER met4 ;
        RECT 14.025000 7.760000 14.345000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025000 8.190000 14.345000 8.510000 ;
      LAYER met4 ;
        RECT 14.025000 8.190000 14.345000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025000 8.620000 14.345000 8.940000 ;
      LAYER met4 ;
        RECT 14.025000 8.620000 14.345000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025000 9.050000 14.345000 9.370000 ;
      LAYER met4 ;
        RECT 14.025000 9.050000 14.345000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025000 9.480000 14.345000 9.800000 ;
      LAYER met4 ;
        RECT 14.025000 9.480000 14.345000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025000 9.910000 14.345000 10.230000 ;
      LAYER met4 ;
        RECT 14.025000 9.910000 14.345000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430000 10.340000 14.750000 10.660000 ;
      LAYER met4 ;
        RECT 14.430000 10.340000 14.750000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430000 10.770000 14.750000 11.090000 ;
      LAYER met4 ;
        RECT 14.430000 10.770000 14.750000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430000 11.200000 14.750000 11.520000 ;
      LAYER met4 ;
        RECT 14.430000 11.200000 14.750000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430000 6.900000 14.750000 7.220000 ;
      LAYER met4 ;
        RECT 14.430000 6.900000 14.750000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430000 7.330000 14.750000 7.650000 ;
      LAYER met4 ;
        RECT 14.430000 7.330000 14.750000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430000 7.760000 14.750000 8.080000 ;
      LAYER met4 ;
        RECT 14.430000 7.760000 14.750000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430000 8.190000 14.750000 8.510000 ;
      LAYER met4 ;
        RECT 14.430000 8.190000 14.750000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430000 8.620000 14.750000 8.940000 ;
      LAYER met4 ;
        RECT 14.430000 8.620000 14.750000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430000 9.050000 14.750000 9.370000 ;
      LAYER met4 ;
        RECT 14.430000 9.050000 14.750000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430000 9.480000 14.750000 9.800000 ;
      LAYER met4 ;
        RECT 14.430000 9.480000 14.750000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430000 9.910000 14.750000 10.230000 ;
      LAYER met4 ;
        RECT 14.430000 9.910000 14.750000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835000 10.340000 15.155000 10.660000 ;
      LAYER met4 ;
        RECT 14.835000 10.340000 15.155000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835000 10.770000 15.155000 11.090000 ;
      LAYER met4 ;
        RECT 14.835000 10.770000 15.155000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835000 11.200000 15.155000 11.520000 ;
      LAYER met4 ;
        RECT 14.835000 11.200000 15.155000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835000 6.900000 15.155000 7.220000 ;
      LAYER met4 ;
        RECT 14.835000 6.900000 15.155000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835000 7.330000 15.155000 7.650000 ;
      LAYER met4 ;
        RECT 14.835000 7.330000 15.155000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835000 7.760000 15.155000 8.080000 ;
      LAYER met4 ;
        RECT 14.835000 7.760000 15.155000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835000 8.190000 15.155000 8.510000 ;
      LAYER met4 ;
        RECT 14.835000 8.190000 15.155000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835000 8.620000 15.155000 8.940000 ;
      LAYER met4 ;
        RECT 14.835000 8.620000 15.155000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835000 9.050000 15.155000 9.370000 ;
      LAYER met4 ;
        RECT 14.835000 9.050000 15.155000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835000 9.480000 15.155000 9.800000 ;
      LAYER met4 ;
        RECT 14.835000 9.480000 15.155000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835000 9.910000 15.155000 10.230000 ;
      LAYER met4 ;
        RECT 14.835000 9.910000 15.155000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240000 10.340000 15.560000 10.660000 ;
      LAYER met4 ;
        RECT 15.240000 10.340000 15.560000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240000 10.770000 15.560000 11.090000 ;
      LAYER met4 ;
        RECT 15.240000 10.770000 15.560000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240000 11.200000 15.560000 11.520000 ;
      LAYER met4 ;
        RECT 15.240000 11.200000 15.560000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240000 6.900000 15.560000 7.220000 ;
      LAYER met4 ;
        RECT 15.240000 6.900000 15.560000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240000 7.330000 15.560000 7.650000 ;
      LAYER met4 ;
        RECT 15.240000 7.330000 15.560000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240000 7.760000 15.560000 8.080000 ;
      LAYER met4 ;
        RECT 15.240000 7.760000 15.560000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240000 8.190000 15.560000 8.510000 ;
      LAYER met4 ;
        RECT 15.240000 8.190000 15.560000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240000 8.620000 15.560000 8.940000 ;
      LAYER met4 ;
        RECT 15.240000 8.620000 15.560000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240000 9.050000 15.560000 9.370000 ;
      LAYER met4 ;
        RECT 15.240000 9.050000 15.560000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240000 9.480000 15.560000 9.800000 ;
      LAYER met4 ;
        RECT 15.240000 9.480000 15.560000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240000 9.910000 15.560000 10.230000 ;
      LAYER met4 ;
        RECT 15.240000 9.910000 15.560000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645000 10.340000 15.965000 10.660000 ;
      LAYER met4 ;
        RECT 15.645000 10.340000 15.965000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645000 10.770000 15.965000 11.090000 ;
      LAYER met4 ;
        RECT 15.645000 10.770000 15.965000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645000 11.200000 15.965000 11.520000 ;
      LAYER met4 ;
        RECT 15.645000 11.200000 15.965000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645000 6.900000 15.965000 7.220000 ;
      LAYER met4 ;
        RECT 15.645000 6.900000 15.965000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645000 7.330000 15.965000 7.650000 ;
      LAYER met4 ;
        RECT 15.645000 7.330000 15.965000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645000 7.760000 15.965000 8.080000 ;
      LAYER met4 ;
        RECT 15.645000 7.760000 15.965000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645000 8.190000 15.965000 8.510000 ;
      LAYER met4 ;
        RECT 15.645000 8.190000 15.965000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645000 8.620000 15.965000 8.940000 ;
      LAYER met4 ;
        RECT 15.645000 8.620000 15.965000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645000 9.050000 15.965000 9.370000 ;
      LAYER met4 ;
        RECT 15.645000 9.050000 15.965000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645000 9.480000 15.965000 9.800000 ;
      LAYER met4 ;
        RECT 15.645000 9.480000 15.965000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645000 9.910000 15.965000 10.230000 ;
      LAYER met4 ;
        RECT 15.645000 9.910000 15.965000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050000 10.340000 16.370000 10.660000 ;
      LAYER met4 ;
        RECT 16.050000 10.340000 16.370000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050000 10.770000 16.370000 11.090000 ;
      LAYER met4 ;
        RECT 16.050000 10.770000 16.370000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050000 11.200000 16.370000 11.520000 ;
      LAYER met4 ;
        RECT 16.050000 11.200000 16.370000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050000 6.900000 16.370000 7.220000 ;
      LAYER met4 ;
        RECT 16.050000 6.900000 16.370000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050000 7.330000 16.370000 7.650000 ;
      LAYER met4 ;
        RECT 16.050000 7.330000 16.370000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050000 7.760000 16.370000 8.080000 ;
      LAYER met4 ;
        RECT 16.050000 7.760000 16.370000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050000 8.190000 16.370000 8.510000 ;
      LAYER met4 ;
        RECT 16.050000 8.190000 16.370000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050000 8.620000 16.370000 8.940000 ;
      LAYER met4 ;
        RECT 16.050000 8.620000 16.370000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050000 9.050000 16.370000 9.370000 ;
      LAYER met4 ;
        RECT 16.050000 9.050000 16.370000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050000 9.480000 16.370000 9.800000 ;
      LAYER met4 ;
        RECT 16.050000 9.480000 16.370000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050000 9.910000 16.370000 10.230000 ;
      LAYER met4 ;
        RECT 16.050000 9.910000 16.370000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 10.340000 16.775000 10.660000 ;
      LAYER met4 ;
        RECT 16.455000 10.340000 16.775000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 10.770000 16.775000 11.090000 ;
      LAYER met4 ;
        RECT 16.455000 10.770000 16.775000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 11.200000 16.775000 11.520000 ;
      LAYER met4 ;
        RECT 16.455000 11.200000 16.775000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 6.900000 16.775000 7.220000 ;
      LAYER met4 ;
        RECT 16.455000 6.900000 16.775000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 7.330000 16.775000 7.650000 ;
      LAYER met4 ;
        RECT 16.455000 7.330000 16.775000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 7.760000 16.775000 8.080000 ;
      LAYER met4 ;
        RECT 16.455000 7.760000 16.775000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 8.190000 16.775000 8.510000 ;
      LAYER met4 ;
        RECT 16.455000 8.190000 16.775000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 8.620000 16.775000 8.940000 ;
      LAYER met4 ;
        RECT 16.455000 8.620000 16.775000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 9.050000 16.775000 9.370000 ;
      LAYER met4 ;
        RECT 16.455000 9.050000 16.775000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 9.480000 16.775000 9.800000 ;
      LAYER met4 ;
        RECT 16.455000 9.480000 16.775000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 9.910000 16.775000 10.230000 ;
      LAYER met4 ;
        RECT 16.455000 9.910000 16.775000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860000 10.340000 17.180000 10.660000 ;
      LAYER met4 ;
        RECT 16.860000 10.340000 17.180000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860000 10.770000 17.180000 11.090000 ;
      LAYER met4 ;
        RECT 16.860000 10.770000 17.180000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860000 11.200000 17.180000 11.520000 ;
      LAYER met4 ;
        RECT 16.860000 11.200000 17.180000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860000 6.900000 17.180000 7.220000 ;
      LAYER met4 ;
        RECT 16.860000 6.900000 17.180000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860000 7.330000 17.180000 7.650000 ;
      LAYER met4 ;
        RECT 16.860000 7.330000 17.180000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860000 7.760000 17.180000 8.080000 ;
      LAYER met4 ;
        RECT 16.860000 7.760000 17.180000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860000 8.190000 17.180000 8.510000 ;
      LAYER met4 ;
        RECT 16.860000 8.190000 17.180000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860000 8.620000 17.180000 8.940000 ;
      LAYER met4 ;
        RECT 16.860000 8.620000 17.180000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860000 9.050000 17.180000 9.370000 ;
      LAYER met4 ;
        RECT 16.860000 9.050000 17.180000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860000 9.480000 17.180000 9.800000 ;
      LAYER met4 ;
        RECT 16.860000 9.480000 17.180000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860000 9.910000 17.180000 10.230000 ;
      LAYER met4 ;
        RECT 16.860000 9.910000 17.180000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265000 10.340000 17.585000 10.660000 ;
      LAYER met4 ;
        RECT 17.265000 10.340000 17.585000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265000 10.770000 17.585000 11.090000 ;
      LAYER met4 ;
        RECT 17.265000 10.770000 17.585000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265000 11.200000 17.585000 11.520000 ;
      LAYER met4 ;
        RECT 17.265000 11.200000 17.585000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265000 6.900000 17.585000 7.220000 ;
      LAYER met4 ;
        RECT 17.265000 6.900000 17.585000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265000 7.330000 17.585000 7.650000 ;
      LAYER met4 ;
        RECT 17.265000 7.330000 17.585000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265000 7.760000 17.585000 8.080000 ;
      LAYER met4 ;
        RECT 17.265000 7.760000 17.585000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265000 8.190000 17.585000 8.510000 ;
      LAYER met4 ;
        RECT 17.265000 8.190000 17.585000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265000 8.620000 17.585000 8.940000 ;
      LAYER met4 ;
        RECT 17.265000 8.620000 17.585000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265000 9.050000 17.585000 9.370000 ;
      LAYER met4 ;
        RECT 17.265000 9.050000 17.585000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265000 9.480000 17.585000 9.800000 ;
      LAYER met4 ;
        RECT 17.265000 9.480000 17.585000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265000 9.910000 17.585000 10.230000 ;
      LAYER met4 ;
        RECT 17.265000 9.910000 17.585000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670000 10.340000 17.990000 10.660000 ;
      LAYER met4 ;
        RECT 17.670000 10.340000 17.990000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670000 10.770000 17.990000 11.090000 ;
      LAYER met4 ;
        RECT 17.670000 10.770000 17.990000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670000 11.200000 17.990000 11.520000 ;
      LAYER met4 ;
        RECT 17.670000 11.200000 17.990000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670000 6.900000 17.990000 7.220000 ;
      LAYER met4 ;
        RECT 17.670000 6.900000 17.990000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670000 7.330000 17.990000 7.650000 ;
      LAYER met4 ;
        RECT 17.670000 7.330000 17.990000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670000 7.760000 17.990000 8.080000 ;
      LAYER met4 ;
        RECT 17.670000 7.760000 17.990000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670000 8.190000 17.990000 8.510000 ;
      LAYER met4 ;
        RECT 17.670000 8.190000 17.990000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670000 8.620000 17.990000 8.940000 ;
      LAYER met4 ;
        RECT 17.670000 8.620000 17.990000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670000 9.050000 17.990000 9.370000 ;
      LAYER met4 ;
        RECT 17.670000 9.050000 17.990000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670000 9.480000 17.990000 9.800000 ;
      LAYER met4 ;
        RECT 17.670000 9.480000 17.990000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670000 9.910000 17.990000 10.230000 ;
      LAYER met4 ;
        RECT 17.670000 9.910000 17.990000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075000 10.340000 18.395000 10.660000 ;
      LAYER met4 ;
        RECT 18.075000 10.340000 18.395000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075000 10.770000 18.395000 11.090000 ;
      LAYER met4 ;
        RECT 18.075000 10.770000 18.395000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075000 11.200000 18.395000 11.520000 ;
      LAYER met4 ;
        RECT 18.075000 11.200000 18.395000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075000 6.900000 18.395000 7.220000 ;
      LAYER met4 ;
        RECT 18.075000 6.900000 18.395000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075000 7.330000 18.395000 7.650000 ;
      LAYER met4 ;
        RECT 18.075000 7.330000 18.395000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075000 7.760000 18.395000 8.080000 ;
      LAYER met4 ;
        RECT 18.075000 7.760000 18.395000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075000 8.190000 18.395000 8.510000 ;
      LAYER met4 ;
        RECT 18.075000 8.190000 18.395000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075000 8.620000 18.395000 8.940000 ;
      LAYER met4 ;
        RECT 18.075000 8.620000 18.395000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075000 9.050000 18.395000 9.370000 ;
      LAYER met4 ;
        RECT 18.075000 9.050000 18.395000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075000 9.480000 18.395000 9.800000 ;
      LAYER met4 ;
        RECT 18.075000 9.480000 18.395000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075000 9.910000 18.395000 10.230000 ;
      LAYER met4 ;
        RECT 18.075000 9.910000 18.395000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480000 10.340000 18.800000 10.660000 ;
      LAYER met4 ;
        RECT 18.480000 10.340000 18.800000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480000 10.770000 18.800000 11.090000 ;
      LAYER met4 ;
        RECT 18.480000 10.770000 18.800000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480000 11.200000 18.800000 11.520000 ;
      LAYER met4 ;
        RECT 18.480000 11.200000 18.800000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480000 6.900000 18.800000 7.220000 ;
      LAYER met4 ;
        RECT 18.480000 6.900000 18.800000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480000 7.330000 18.800000 7.650000 ;
      LAYER met4 ;
        RECT 18.480000 7.330000 18.800000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480000 7.760000 18.800000 8.080000 ;
      LAYER met4 ;
        RECT 18.480000 7.760000 18.800000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480000 8.190000 18.800000 8.510000 ;
      LAYER met4 ;
        RECT 18.480000 8.190000 18.800000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480000 8.620000 18.800000 8.940000 ;
      LAYER met4 ;
        RECT 18.480000 8.620000 18.800000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480000 9.050000 18.800000 9.370000 ;
      LAYER met4 ;
        RECT 18.480000 9.050000 18.800000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480000 9.480000 18.800000 9.800000 ;
      LAYER met4 ;
        RECT 18.480000 9.480000 18.800000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480000 9.910000 18.800000 10.230000 ;
      LAYER met4 ;
        RECT 18.480000 9.910000 18.800000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885000 10.340000 19.205000 10.660000 ;
      LAYER met4 ;
        RECT 18.885000 10.340000 19.205000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885000 10.770000 19.205000 11.090000 ;
      LAYER met4 ;
        RECT 18.885000 10.770000 19.205000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885000 11.200000 19.205000 11.520000 ;
      LAYER met4 ;
        RECT 18.885000 11.200000 19.205000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885000 6.900000 19.205000 7.220000 ;
      LAYER met4 ;
        RECT 18.885000 6.900000 19.205000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885000 7.330000 19.205000 7.650000 ;
      LAYER met4 ;
        RECT 18.885000 7.330000 19.205000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885000 7.760000 19.205000 8.080000 ;
      LAYER met4 ;
        RECT 18.885000 7.760000 19.205000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885000 8.190000 19.205000 8.510000 ;
      LAYER met4 ;
        RECT 18.885000 8.190000 19.205000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885000 8.620000 19.205000 8.940000 ;
      LAYER met4 ;
        RECT 18.885000 8.620000 19.205000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885000 9.050000 19.205000 9.370000 ;
      LAYER met4 ;
        RECT 18.885000 9.050000 19.205000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885000 9.480000 19.205000 9.800000 ;
      LAYER met4 ;
        RECT 18.885000 9.480000 19.205000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885000 9.910000 19.205000 10.230000 ;
      LAYER met4 ;
        RECT 18.885000 9.910000 19.205000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290000 10.340000 19.610000 10.660000 ;
      LAYER met4 ;
        RECT 19.290000 10.340000 19.610000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290000 10.770000 19.610000 11.090000 ;
      LAYER met4 ;
        RECT 19.290000 10.770000 19.610000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290000 11.200000 19.610000 11.520000 ;
      LAYER met4 ;
        RECT 19.290000 11.200000 19.610000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290000 6.900000 19.610000 7.220000 ;
      LAYER met4 ;
        RECT 19.290000 6.900000 19.610000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290000 7.330000 19.610000 7.650000 ;
      LAYER met4 ;
        RECT 19.290000 7.330000 19.610000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290000 7.760000 19.610000 8.080000 ;
      LAYER met4 ;
        RECT 19.290000 7.760000 19.610000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290000 8.190000 19.610000 8.510000 ;
      LAYER met4 ;
        RECT 19.290000 8.190000 19.610000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290000 8.620000 19.610000 8.940000 ;
      LAYER met4 ;
        RECT 19.290000 8.620000 19.610000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290000 9.050000 19.610000 9.370000 ;
      LAYER met4 ;
        RECT 19.290000 9.050000 19.610000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290000 9.480000 19.610000 9.800000 ;
      LAYER met4 ;
        RECT 19.290000 9.480000 19.610000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290000 9.910000 19.610000 10.230000 ;
      LAYER met4 ;
        RECT 19.290000 9.910000 19.610000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695000 10.340000 20.015000 10.660000 ;
      LAYER met4 ;
        RECT 19.695000 10.340000 20.015000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695000 10.770000 20.015000 11.090000 ;
      LAYER met4 ;
        RECT 19.695000 10.770000 20.015000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695000 11.200000 20.015000 11.520000 ;
      LAYER met4 ;
        RECT 19.695000 11.200000 20.015000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695000 6.900000 20.015000 7.220000 ;
      LAYER met4 ;
        RECT 19.695000 6.900000 20.015000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695000 7.330000 20.015000 7.650000 ;
      LAYER met4 ;
        RECT 19.695000 7.330000 20.015000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695000 7.760000 20.015000 8.080000 ;
      LAYER met4 ;
        RECT 19.695000 7.760000 20.015000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695000 8.190000 20.015000 8.510000 ;
      LAYER met4 ;
        RECT 19.695000 8.190000 20.015000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695000 8.620000 20.015000 8.940000 ;
      LAYER met4 ;
        RECT 19.695000 8.620000 20.015000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695000 9.050000 20.015000 9.370000 ;
      LAYER met4 ;
        RECT 19.695000 9.050000 20.015000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695000 9.480000 20.015000 9.800000 ;
      LAYER met4 ;
        RECT 19.695000 9.480000 20.015000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695000 9.910000 20.015000 10.230000 ;
      LAYER met4 ;
        RECT 19.695000 9.910000 20.015000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270000 10.340000 2.590000 10.660000 ;
      LAYER met4 ;
        RECT 2.270000 10.340000 2.590000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270000 10.770000 2.590000 11.090000 ;
      LAYER met4 ;
        RECT 2.270000 10.770000 2.590000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270000 11.200000 2.590000 11.520000 ;
      LAYER met4 ;
        RECT 2.270000 11.200000 2.590000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270000 6.900000 2.590000 7.220000 ;
      LAYER met4 ;
        RECT 2.270000 6.900000 2.590000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270000 7.330000 2.590000 7.650000 ;
      LAYER met4 ;
        RECT 2.270000 7.330000 2.590000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270000 7.760000 2.590000 8.080000 ;
      LAYER met4 ;
        RECT 2.270000 7.760000 2.590000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270000 8.190000 2.590000 8.510000 ;
      LAYER met4 ;
        RECT 2.270000 8.190000 2.590000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270000 8.620000 2.590000 8.940000 ;
      LAYER met4 ;
        RECT 2.270000 8.620000 2.590000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270000 9.050000 2.590000 9.370000 ;
      LAYER met4 ;
        RECT 2.270000 9.050000 2.590000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270000 9.480000 2.590000 9.800000 ;
      LAYER met4 ;
        RECT 2.270000 9.480000 2.590000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270000 9.910000 2.590000 10.230000 ;
      LAYER met4 ;
        RECT 2.270000 9.910000 2.590000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680000 10.340000 3.000000 10.660000 ;
      LAYER met4 ;
        RECT 2.680000 10.340000 3.000000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680000 10.770000 3.000000 11.090000 ;
      LAYER met4 ;
        RECT 2.680000 10.770000 3.000000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680000 11.200000 3.000000 11.520000 ;
      LAYER met4 ;
        RECT 2.680000 11.200000 3.000000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680000 6.900000 3.000000 7.220000 ;
      LAYER met4 ;
        RECT 2.680000 6.900000 3.000000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680000 7.330000 3.000000 7.650000 ;
      LAYER met4 ;
        RECT 2.680000 7.330000 3.000000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680000 7.760000 3.000000 8.080000 ;
      LAYER met4 ;
        RECT 2.680000 7.760000 3.000000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680000 8.190000 3.000000 8.510000 ;
      LAYER met4 ;
        RECT 2.680000 8.190000 3.000000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680000 8.620000 3.000000 8.940000 ;
      LAYER met4 ;
        RECT 2.680000 8.620000 3.000000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680000 9.050000 3.000000 9.370000 ;
      LAYER met4 ;
        RECT 2.680000 9.050000 3.000000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680000 9.480000 3.000000 9.800000 ;
      LAYER met4 ;
        RECT 2.680000 9.480000 3.000000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680000 9.910000 3.000000 10.230000 ;
      LAYER met4 ;
        RECT 2.680000 9.910000 3.000000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100000 10.340000 20.420000 10.660000 ;
      LAYER met4 ;
        RECT 20.100000 10.340000 20.420000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100000 10.770000 20.420000 11.090000 ;
      LAYER met4 ;
        RECT 20.100000 10.770000 20.420000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100000 11.200000 20.420000 11.520000 ;
      LAYER met4 ;
        RECT 20.100000 11.200000 20.420000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100000 6.900000 20.420000 7.220000 ;
      LAYER met4 ;
        RECT 20.100000 6.900000 20.420000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100000 7.330000 20.420000 7.650000 ;
      LAYER met4 ;
        RECT 20.100000 7.330000 20.420000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100000 7.760000 20.420000 8.080000 ;
      LAYER met4 ;
        RECT 20.100000 7.760000 20.420000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100000 8.190000 20.420000 8.510000 ;
      LAYER met4 ;
        RECT 20.100000 8.190000 20.420000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100000 8.620000 20.420000 8.940000 ;
      LAYER met4 ;
        RECT 20.100000 8.620000 20.420000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100000 9.050000 20.420000 9.370000 ;
      LAYER met4 ;
        RECT 20.100000 9.050000 20.420000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100000 9.480000 20.420000 9.800000 ;
      LAYER met4 ;
        RECT 20.100000 9.480000 20.420000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100000 9.910000 20.420000 10.230000 ;
      LAYER met4 ;
        RECT 20.100000 9.910000 20.420000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505000 10.340000 20.825000 10.660000 ;
      LAYER met4 ;
        RECT 20.505000 10.340000 20.825000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505000 10.770000 20.825000 11.090000 ;
      LAYER met4 ;
        RECT 20.505000 10.770000 20.825000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505000 11.200000 20.825000 11.520000 ;
      LAYER met4 ;
        RECT 20.505000 11.200000 20.825000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505000 6.900000 20.825000 7.220000 ;
      LAYER met4 ;
        RECT 20.505000 6.900000 20.825000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505000 7.330000 20.825000 7.650000 ;
      LAYER met4 ;
        RECT 20.505000 7.330000 20.825000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505000 7.760000 20.825000 8.080000 ;
      LAYER met4 ;
        RECT 20.505000 7.760000 20.825000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505000 8.190000 20.825000 8.510000 ;
      LAYER met4 ;
        RECT 20.505000 8.190000 20.825000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505000 8.620000 20.825000 8.940000 ;
      LAYER met4 ;
        RECT 20.505000 8.620000 20.825000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505000 9.050000 20.825000 9.370000 ;
      LAYER met4 ;
        RECT 20.505000 9.050000 20.825000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505000 9.480000 20.825000 9.800000 ;
      LAYER met4 ;
        RECT 20.505000 9.480000 20.825000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505000 9.910000 20.825000 10.230000 ;
      LAYER met4 ;
        RECT 20.505000 9.910000 20.825000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910000 10.340000 21.230000 10.660000 ;
      LAYER met4 ;
        RECT 20.910000 10.340000 21.230000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910000 10.770000 21.230000 11.090000 ;
      LAYER met4 ;
        RECT 20.910000 10.770000 21.230000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910000 11.200000 21.230000 11.520000 ;
      LAYER met4 ;
        RECT 20.910000 11.200000 21.230000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910000 6.900000 21.230000 7.220000 ;
      LAYER met4 ;
        RECT 20.910000 6.900000 21.230000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910000 7.330000 21.230000 7.650000 ;
      LAYER met4 ;
        RECT 20.910000 7.330000 21.230000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910000 7.760000 21.230000 8.080000 ;
      LAYER met4 ;
        RECT 20.910000 7.760000 21.230000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910000 8.190000 21.230000 8.510000 ;
      LAYER met4 ;
        RECT 20.910000 8.190000 21.230000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910000 8.620000 21.230000 8.940000 ;
      LAYER met4 ;
        RECT 20.910000 8.620000 21.230000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910000 9.050000 21.230000 9.370000 ;
      LAYER met4 ;
        RECT 20.910000 9.050000 21.230000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910000 9.480000 21.230000 9.800000 ;
      LAYER met4 ;
        RECT 20.910000 9.480000 21.230000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910000 9.910000 21.230000 10.230000 ;
      LAYER met4 ;
        RECT 20.910000 9.910000 21.230000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315000 10.340000 21.635000 10.660000 ;
      LAYER met4 ;
        RECT 21.315000 10.340000 21.635000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315000 10.770000 21.635000 11.090000 ;
      LAYER met4 ;
        RECT 21.315000 10.770000 21.635000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315000 11.200000 21.635000 11.520000 ;
      LAYER met4 ;
        RECT 21.315000 11.200000 21.635000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315000 6.900000 21.635000 7.220000 ;
      LAYER met4 ;
        RECT 21.315000 6.900000 21.635000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315000 7.330000 21.635000 7.650000 ;
      LAYER met4 ;
        RECT 21.315000 7.330000 21.635000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315000 7.760000 21.635000 8.080000 ;
      LAYER met4 ;
        RECT 21.315000 7.760000 21.635000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315000 8.190000 21.635000 8.510000 ;
      LAYER met4 ;
        RECT 21.315000 8.190000 21.635000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315000 8.620000 21.635000 8.940000 ;
      LAYER met4 ;
        RECT 21.315000 8.620000 21.635000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315000 9.050000 21.635000 9.370000 ;
      LAYER met4 ;
        RECT 21.315000 9.050000 21.635000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315000 9.480000 21.635000 9.800000 ;
      LAYER met4 ;
        RECT 21.315000 9.480000 21.635000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315000 9.910000 21.635000 10.230000 ;
      LAYER met4 ;
        RECT 21.315000 9.910000 21.635000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720000 10.340000 22.040000 10.660000 ;
      LAYER met4 ;
        RECT 21.720000 10.340000 22.040000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720000 10.770000 22.040000 11.090000 ;
      LAYER met4 ;
        RECT 21.720000 10.770000 22.040000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720000 11.200000 22.040000 11.520000 ;
      LAYER met4 ;
        RECT 21.720000 11.200000 22.040000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720000 6.900000 22.040000 7.220000 ;
      LAYER met4 ;
        RECT 21.720000 6.900000 22.040000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720000 7.330000 22.040000 7.650000 ;
      LAYER met4 ;
        RECT 21.720000 7.330000 22.040000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720000 7.760000 22.040000 8.080000 ;
      LAYER met4 ;
        RECT 21.720000 7.760000 22.040000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720000 8.190000 22.040000 8.510000 ;
      LAYER met4 ;
        RECT 21.720000 8.190000 22.040000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720000 8.620000 22.040000 8.940000 ;
      LAYER met4 ;
        RECT 21.720000 8.620000 22.040000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720000 9.050000 22.040000 9.370000 ;
      LAYER met4 ;
        RECT 21.720000 9.050000 22.040000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720000 9.480000 22.040000 9.800000 ;
      LAYER met4 ;
        RECT 21.720000 9.480000 22.040000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720000 9.910000 22.040000 10.230000 ;
      LAYER met4 ;
        RECT 21.720000 9.910000 22.040000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125000 10.340000 22.445000 10.660000 ;
      LAYER met4 ;
        RECT 22.125000 10.340000 22.445000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125000 10.770000 22.445000 11.090000 ;
      LAYER met4 ;
        RECT 22.125000 10.770000 22.445000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125000 11.200000 22.445000 11.520000 ;
      LAYER met4 ;
        RECT 22.125000 11.200000 22.445000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125000 6.900000 22.445000 7.220000 ;
      LAYER met4 ;
        RECT 22.125000 6.900000 22.445000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125000 7.330000 22.445000 7.650000 ;
      LAYER met4 ;
        RECT 22.125000 7.330000 22.445000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125000 7.760000 22.445000 8.080000 ;
      LAYER met4 ;
        RECT 22.125000 7.760000 22.445000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125000 8.190000 22.445000 8.510000 ;
      LAYER met4 ;
        RECT 22.125000 8.190000 22.445000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125000 8.620000 22.445000 8.940000 ;
      LAYER met4 ;
        RECT 22.125000 8.620000 22.445000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125000 9.050000 22.445000 9.370000 ;
      LAYER met4 ;
        RECT 22.125000 9.050000 22.445000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125000 9.480000 22.445000 9.800000 ;
      LAYER met4 ;
        RECT 22.125000 9.480000 22.445000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125000 9.910000 22.445000 10.230000 ;
      LAYER met4 ;
        RECT 22.125000 9.910000 22.445000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530000 10.340000 22.850000 10.660000 ;
      LAYER met4 ;
        RECT 22.530000 10.340000 22.850000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530000 10.770000 22.850000 11.090000 ;
      LAYER met4 ;
        RECT 22.530000 10.770000 22.850000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530000 11.200000 22.850000 11.520000 ;
      LAYER met4 ;
        RECT 22.530000 11.200000 22.850000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530000 6.900000 22.850000 7.220000 ;
      LAYER met4 ;
        RECT 22.530000 6.900000 22.850000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530000 7.330000 22.850000 7.650000 ;
      LAYER met4 ;
        RECT 22.530000 7.330000 22.850000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530000 7.760000 22.850000 8.080000 ;
      LAYER met4 ;
        RECT 22.530000 7.760000 22.850000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530000 8.190000 22.850000 8.510000 ;
      LAYER met4 ;
        RECT 22.530000 8.190000 22.850000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530000 8.620000 22.850000 8.940000 ;
      LAYER met4 ;
        RECT 22.530000 8.620000 22.850000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530000 9.050000 22.850000 9.370000 ;
      LAYER met4 ;
        RECT 22.530000 9.050000 22.850000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530000 9.480000 22.850000 9.800000 ;
      LAYER met4 ;
        RECT 22.530000 9.480000 22.850000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530000 9.910000 22.850000 10.230000 ;
      LAYER met4 ;
        RECT 22.530000 9.910000 22.850000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935000 10.340000 23.255000 10.660000 ;
      LAYER met4 ;
        RECT 22.935000 10.340000 23.255000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935000 10.770000 23.255000 11.090000 ;
      LAYER met4 ;
        RECT 22.935000 10.770000 23.255000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935000 11.200000 23.255000 11.520000 ;
      LAYER met4 ;
        RECT 22.935000 11.200000 23.255000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935000 6.900000 23.255000 7.220000 ;
      LAYER met4 ;
        RECT 22.935000 6.900000 23.255000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935000 7.330000 23.255000 7.650000 ;
      LAYER met4 ;
        RECT 22.935000 7.330000 23.255000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935000 7.760000 23.255000 8.080000 ;
      LAYER met4 ;
        RECT 22.935000 7.760000 23.255000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935000 8.190000 23.255000 8.510000 ;
      LAYER met4 ;
        RECT 22.935000 8.190000 23.255000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935000 8.620000 23.255000 8.940000 ;
      LAYER met4 ;
        RECT 22.935000 8.620000 23.255000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935000 9.050000 23.255000 9.370000 ;
      LAYER met4 ;
        RECT 22.935000 9.050000 23.255000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935000 9.480000 23.255000 9.800000 ;
      LAYER met4 ;
        RECT 22.935000 9.480000 23.255000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935000 9.910000 23.255000 10.230000 ;
      LAYER met4 ;
        RECT 22.935000 9.910000 23.255000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340000 10.340000 23.660000 10.660000 ;
      LAYER met4 ;
        RECT 23.340000 10.340000 23.660000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340000 10.770000 23.660000 11.090000 ;
      LAYER met4 ;
        RECT 23.340000 10.770000 23.660000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340000 11.200000 23.660000 11.520000 ;
      LAYER met4 ;
        RECT 23.340000 11.200000 23.660000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340000 6.900000 23.660000 7.220000 ;
      LAYER met4 ;
        RECT 23.340000 6.900000 23.660000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340000 7.330000 23.660000 7.650000 ;
      LAYER met4 ;
        RECT 23.340000 7.330000 23.660000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340000 7.760000 23.660000 8.080000 ;
      LAYER met4 ;
        RECT 23.340000 7.760000 23.660000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340000 8.190000 23.660000 8.510000 ;
      LAYER met4 ;
        RECT 23.340000 8.190000 23.660000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340000 8.620000 23.660000 8.940000 ;
      LAYER met4 ;
        RECT 23.340000 8.620000 23.660000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340000 9.050000 23.660000 9.370000 ;
      LAYER met4 ;
        RECT 23.340000 9.050000 23.660000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340000 9.480000 23.660000 9.800000 ;
      LAYER met4 ;
        RECT 23.340000 9.480000 23.660000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340000 9.910000 23.660000 10.230000 ;
      LAYER met4 ;
        RECT 23.340000 9.910000 23.660000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 10.340000 24.065000 10.660000 ;
      LAYER met4 ;
        RECT 23.745000 10.340000 24.065000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 10.770000 24.065000 11.090000 ;
      LAYER met4 ;
        RECT 23.745000 10.770000 24.065000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 11.200000 24.065000 11.520000 ;
      LAYER met4 ;
        RECT 23.745000 11.200000 24.065000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 6.900000 24.065000 7.220000 ;
      LAYER met4 ;
        RECT 23.745000 6.900000 24.065000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 7.330000 24.065000 7.650000 ;
      LAYER met4 ;
        RECT 23.745000 7.330000 24.065000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 7.760000 24.065000 8.080000 ;
      LAYER met4 ;
        RECT 23.745000 7.760000 24.065000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 8.190000 24.065000 8.510000 ;
      LAYER met4 ;
        RECT 23.745000 8.190000 24.065000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 8.620000 24.065000 8.940000 ;
      LAYER met4 ;
        RECT 23.745000 8.620000 24.065000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 9.050000 24.065000 9.370000 ;
      LAYER met4 ;
        RECT 23.745000 9.050000 24.065000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 9.480000 24.065000 9.800000 ;
      LAYER met4 ;
        RECT 23.745000 9.480000 24.065000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 9.910000 24.065000 10.230000 ;
      LAYER met4 ;
        RECT 23.745000 9.910000 24.065000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 10.340000 24.470000 10.660000 ;
      LAYER met4 ;
        RECT 24.150000 10.340000 24.470000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 10.770000 24.470000 11.090000 ;
      LAYER met4 ;
        RECT 24.150000 10.770000 24.470000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 11.200000 24.470000 11.520000 ;
      LAYER met4 ;
        RECT 24.150000 11.200000 24.470000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 6.900000 24.470000 7.220000 ;
      LAYER met4 ;
        RECT 24.150000 6.900000 24.470000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 7.330000 24.470000 7.650000 ;
      LAYER met4 ;
        RECT 24.150000 7.330000 24.470000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 7.760000 24.470000 8.080000 ;
      LAYER met4 ;
        RECT 24.150000 7.760000 24.470000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 8.190000 24.470000 8.510000 ;
      LAYER met4 ;
        RECT 24.150000 8.190000 24.470000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 8.620000 24.470000 8.940000 ;
      LAYER met4 ;
        RECT 24.150000 8.620000 24.470000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 9.050000 24.470000 9.370000 ;
      LAYER met4 ;
        RECT 24.150000 9.050000 24.470000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 9.480000 24.470000 9.800000 ;
      LAYER met4 ;
        RECT 24.150000 9.480000 24.470000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 9.910000 24.470000 10.230000 ;
      LAYER met4 ;
        RECT 24.150000 9.910000 24.470000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090000 10.340000 3.410000 10.660000 ;
      LAYER met4 ;
        RECT 3.090000 10.340000 3.410000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090000 10.770000 3.410000 11.090000 ;
      LAYER met4 ;
        RECT 3.090000 10.770000 3.410000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090000 11.200000 3.410000 11.520000 ;
      LAYER met4 ;
        RECT 3.090000 11.200000 3.410000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090000 6.900000 3.410000 7.220000 ;
      LAYER met4 ;
        RECT 3.090000 6.900000 3.410000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090000 7.330000 3.410000 7.650000 ;
      LAYER met4 ;
        RECT 3.090000 7.330000 3.410000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090000 7.760000 3.410000 8.080000 ;
      LAYER met4 ;
        RECT 3.090000 7.760000 3.410000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090000 8.190000 3.410000 8.510000 ;
      LAYER met4 ;
        RECT 3.090000 8.190000 3.410000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090000 8.620000 3.410000 8.940000 ;
      LAYER met4 ;
        RECT 3.090000 8.620000 3.410000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090000 9.050000 3.410000 9.370000 ;
      LAYER met4 ;
        RECT 3.090000 9.050000 3.410000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090000 9.480000 3.410000 9.800000 ;
      LAYER met4 ;
        RECT 3.090000 9.480000 3.410000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090000 9.910000 3.410000 10.230000 ;
      LAYER met4 ;
        RECT 3.090000 9.910000 3.410000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495000 10.340000 3.815000 10.660000 ;
      LAYER met4 ;
        RECT 3.495000 10.340000 3.815000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495000 10.770000 3.815000 11.090000 ;
      LAYER met4 ;
        RECT 3.495000 10.770000 3.815000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495000 11.200000 3.815000 11.520000 ;
      LAYER met4 ;
        RECT 3.495000 11.200000 3.815000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495000 6.900000 3.815000 7.220000 ;
      LAYER met4 ;
        RECT 3.495000 6.900000 3.815000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495000 7.330000 3.815000 7.650000 ;
      LAYER met4 ;
        RECT 3.495000 7.330000 3.815000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495000 7.760000 3.815000 8.080000 ;
      LAYER met4 ;
        RECT 3.495000 7.760000 3.815000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495000 8.190000 3.815000 8.510000 ;
      LAYER met4 ;
        RECT 3.495000 8.190000 3.815000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495000 8.620000 3.815000 8.940000 ;
      LAYER met4 ;
        RECT 3.495000 8.620000 3.815000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495000 9.050000 3.815000 9.370000 ;
      LAYER met4 ;
        RECT 3.495000 9.050000 3.815000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495000 9.480000 3.815000 9.800000 ;
      LAYER met4 ;
        RECT 3.495000 9.480000 3.815000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495000 9.910000 3.815000 10.230000 ;
      LAYER met4 ;
        RECT 3.495000 9.910000 3.815000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900000 10.340000 4.220000 10.660000 ;
      LAYER met4 ;
        RECT 3.900000 10.340000 4.220000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900000 10.770000 4.220000 11.090000 ;
      LAYER met4 ;
        RECT 3.900000 10.770000 4.220000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900000 11.200000 4.220000 11.520000 ;
      LAYER met4 ;
        RECT 3.900000 11.200000 4.220000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900000 6.900000 4.220000 7.220000 ;
      LAYER met4 ;
        RECT 3.900000 6.900000 4.220000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900000 7.330000 4.220000 7.650000 ;
      LAYER met4 ;
        RECT 3.900000 7.330000 4.220000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900000 7.760000 4.220000 8.080000 ;
      LAYER met4 ;
        RECT 3.900000 7.760000 4.220000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900000 8.190000 4.220000 8.510000 ;
      LAYER met4 ;
        RECT 3.900000 8.190000 4.220000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900000 8.620000 4.220000 8.940000 ;
      LAYER met4 ;
        RECT 3.900000 8.620000 4.220000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900000 9.050000 4.220000 9.370000 ;
      LAYER met4 ;
        RECT 3.900000 9.050000 4.220000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900000 9.480000 4.220000 9.800000 ;
      LAYER met4 ;
        RECT 3.900000 9.480000 4.220000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900000 9.910000 4.220000 10.230000 ;
      LAYER met4 ;
        RECT 3.900000 9.910000 4.220000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305000 10.340000 4.625000 10.660000 ;
      LAYER met4 ;
        RECT 4.305000 10.340000 4.625000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305000 10.770000 4.625000 11.090000 ;
      LAYER met4 ;
        RECT 4.305000 10.770000 4.625000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305000 11.200000 4.625000 11.520000 ;
      LAYER met4 ;
        RECT 4.305000 11.200000 4.625000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305000 6.900000 4.625000 7.220000 ;
      LAYER met4 ;
        RECT 4.305000 6.900000 4.625000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305000 7.330000 4.625000 7.650000 ;
      LAYER met4 ;
        RECT 4.305000 7.330000 4.625000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305000 7.760000 4.625000 8.080000 ;
      LAYER met4 ;
        RECT 4.305000 7.760000 4.625000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305000 8.190000 4.625000 8.510000 ;
      LAYER met4 ;
        RECT 4.305000 8.190000 4.625000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305000 8.620000 4.625000 8.940000 ;
      LAYER met4 ;
        RECT 4.305000 8.620000 4.625000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305000 9.050000 4.625000 9.370000 ;
      LAYER met4 ;
        RECT 4.305000 9.050000 4.625000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305000 9.480000 4.625000 9.800000 ;
      LAYER met4 ;
        RECT 4.305000 9.480000 4.625000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305000 9.910000 4.625000 10.230000 ;
      LAYER met4 ;
        RECT 4.305000 9.910000 4.625000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710000 10.340000 5.030000 10.660000 ;
      LAYER met4 ;
        RECT 4.710000 10.340000 5.030000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710000 10.770000 5.030000 11.090000 ;
      LAYER met4 ;
        RECT 4.710000 10.770000 5.030000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710000 11.200000 5.030000 11.520000 ;
      LAYER met4 ;
        RECT 4.710000 11.200000 5.030000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710000 6.900000 5.030000 7.220000 ;
      LAYER met4 ;
        RECT 4.710000 6.900000 5.030000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710000 7.330000 5.030000 7.650000 ;
      LAYER met4 ;
        RECT 4.710000 7.330000 5.030000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710000 7.760000 5.030000 8.080000 ;
      LAYER met4 ;
        RECT 4.710000 7.760000 5.030000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710000 8.190000 5.030000 8.510000 ;
      LAYER met4 ;
        RECT 4.710000 8.190000 5.030000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710000 8.620000 5.030000 8.940000 ;
      LAYER met4 ;
        RECT 4.710000 8.620000 5.030000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710000 9.050000 5.030000 9.370000 ;
      LAYER met4 ;
        RECT 4.710000 9.050000 5.030000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710000 9.480000 5.030000 9.800000 ;
      LAYER met4 ;
        RECT 4.710000 9.480000 5.030000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710000 9.910000 5.030000 10.230000 ;
      LAYER met4 ;
        RECT 4.710000 9.910000 5.030000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115000 10.340000 5.435000 10.660000 ;
      LAYER met4 ;
        RECT 5.115000 10.340000 5.435000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115000 10.770000 5.435000 11.090000 ;
      LAYER met4 ;
        RECT 5.115000 10.770000 5.435000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115000 11.200000 5.435000 11.520000 ;
      LAYER met4 ;
        RECT 5.115000 11.200000 5.435000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115000 6.900000 5.435000 7.220000 ;
      LAYER met4 ;
        RECT 5.115000 6.900000 5.435000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115000 7.330000 5.435000 7.650000 ;
      LAYER met4 ;
        RECT 5.115000 7.330000 5.435000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115000 7.760000 5.435000 8.080000 ;
      LAYER met4 ;
        RECT 5.115000 7.760000 5.435000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115000 8.190000 5.435000 8.510000 ;
      LAYER met4 ;
        RECT 5.115000 8.190000 5.435000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115000 8.620000 5.435000 8.940000 ;
      LAYER met4 ;
        RECT 5.115000 8.620000 5.435000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115000 9.050000 5.435000 9.370000 ;
      LAYER met4 ;
        RECT 5.115000 9.050000 5.435000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115000 9.480000 5.435000 9.800000 ;
      LAYER met4 ;
        RECT 5.115000 9.480000 5.435000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115000 9.910000 5.435000 10.230000 ;
      LAYER met4 ;
        RECT 5.115000 9.910000 5.435000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520000 10.340000 5.840000 10.660000 ;
      LAYER met4 ;
        RECT 5.520000 10.340000 5.840000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520000 10.770000 5.840000 11.090000 ;
      LAYER met4 ;
        RECT 5.520000 10.770000 5.840000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520000 11.200000 5.840000 11.520000 ;
      LAYER met4 ;
        RECT 5.520000 11.200000 5.840000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520000 6.900000 5.840000 7.220000 ;
      LAYER met4 ;
        RECT 5.520000 6.900000 5.840000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520000 7.330000 5.840000 7.650000 ;
      LAYER met4 ;
        RECT 5.520000 7.330000 5.840000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520000 7.760000 5.840000 8.080000 ;
      LAYER met4 ;
        RECT 5.520000 7.760000 5.840000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520000 8.190000 5.840000 8.510000 ;
      LAYER met4 ;
        RECT 5.520000 8.190000 5.840000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520000 8.620000 5.840000 8.940000 ;
      LAYER met4 ;
        RECT 5.520000 8.620000 5.840000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520000 9.050000 5.840000 9.370000 ;
      LAYER met4 ;
        RECT 5.520000 9.050000 5.840000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520000 9.480000 5.840000 9.800000 ;
      LAYER met4 ;
        RECT 5.520000 9.480000 5.840000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520000 9.910000 5.840000 10.230000 ;
      LAYER met4 ;
        RECT 5.520000 9.910000 5.840000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925000 10.340000 6.245000 10.660000 ;
      LAYER met4 ;
        RECT 5.925000 10.340000 6.245000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925000 10.770000 6.245000 11.090000 ;
      LAYER met4 ;
        RECT 5.925000 10.770000 6.245000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925000 11.200000 6.245000 11.520000 ;
      LAYER met4 ;
        RECT 5.925000 11.200000 6.245000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925000 6.900000 6.245000 7.220000 ;
      LAYER met4 ;
        RECT 5.925000 6.900000 6.245000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925000 7.330000 6.245000 7.650000 ;
      LAYER met4 ;
        RECT 5.925000 7.330000 6.245000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925000 7.760000 6.245000 8.080000 ;
      LAYER met4 ;
        RECT 5.925000 7.760000 6.245000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925000 8.190000 6.245000 8.510000 ;
      LAYER met4 ;
        RECT 5.925000 8.190000 6.245000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925000 8.620000 6.245000 8.940000 ;
      LAYER met4 ;
        RECT 5.925000 8.620000 6.245000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925000 9.050000 6.245000 9.370000 ;
      LAYER met4 ;
        RECT 5.925000 9.050000 6.245000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925000 9.480000 6.245000 9.800000 ;
      LAYER met4 ;
        RECT 5.925000 9.480000 6.245000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925000 9.910000 6.245000 10.230000 ;
      LAYER met4 ;
        RECT 5.925000 9.910000 6.245000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 10.340000 51.105000 10.660000 ;
      LAYER met4 ;
        RECT 50.785000 10.340000 51.105000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 10.770000 51.105000 11.090000 ;
      LAYER met4 ;
        RECT 50.785000 10.770000 51.105000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 11.200000 51.105000 11.520000 ;
      LAYER met4 ;
        RECT 50.785000 11.200000 51.105000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 6.900000 51.105000 7.220000 ;
      LAYER met4 ;
        RECT 50.785000 6.900000 51.105000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 7.330000 51.105000 7.650000 ;
      LAYER met4 ;
        RECT 50.785000 7.330000 51.105000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 7.760000 51.105000 8.080000 ;
      LAYER met4 ;
        RECT 50.785000 7.760000 51.105000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 8.190000 51.105000 8.510000 ;
      LAYER met4 ;
        RECT 50.785000 8.190000 51.105000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 8.620000 51.105000 8.940000 ;
      LAYER met4 ;
        RECT 50.785000 8.620000 51.105000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 9.050000 51.105000 9.370000 ;
      LAYER met4 ;
        RECT 50.785000 9.050000 51.105000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 9.480000 51.105000 9.800000 ;
      LAYER met4 ;
        RECT 50.785000 9.480000 51.105000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 9.910000 51.105000 10.230000 ;
      LAYER met4 ;
        RECT 50.785000 9.910000 51.105000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 10.340000 51.515000 10.660000 ;
      LAYER met4 ;
        RECT 51.195000 10.340000 51.515000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 10.770000 51.515000 11.090000 ;
      LAYER met4 ;
        RECT 51.195000 10.770000 51.515000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 11.200000 51.515000 11.520000 ;
      LAYER met4 ;
        RECT 51.195000 11.200000 51.515000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 6.900000 51.515000 7.220000 ;
      LAYER met4 ;
        RECT 51.195000 6.900000 51.515000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 7.330000 51.515000 7.650000 ;
      LAYER met4 ;
        RECT 51.195000 7.330000 51.515000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 7.760000 51.515000 8.080000 ;
      LAYER met4 ;
        RECT 51.195000 7.760000 51.515000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 8.190000 51.515000 8.510000 ;
      LAYER met4 ;
        RECT 51.195000 8.190000 51.515000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 8.620000 51.515000 8.940000 ;
      LAYER met4 ;
        RECT 51.195000 8.620000 51.515000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 9.050000 51.515000 9.370000 ;
      LAYER met4 ;
        RECT 51.195000 9.050000 51.515000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 9.480000 51.515000 9.800000 ;
      LAYER met4 ;
        RECT 51.195000 9.480000 51.515000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 9.910000 51.515000 10.230000 ;
      LAYER met4 ;
        RECT 51.195000 9.910000 51.515000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 10.340000 51.925000 10.660000 ;
      LAYER met4 ;
        RECT 51.605000 10.340000 51.925000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 10.770000 51.925000 11.090000 ;
      LAYER met4 ;
        RECT 51.605000 10.770000 51.925000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 11.200000 51.925000 11.520000 ;
      LAYER met4 ;
        RECT 51.605000 11.200000 51.925000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 6.900000 51.925000 7.220000 ;
      LAYER met4 ;
        RECT 51.605000 6.900000 51.925000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 7.330000 51.925000 7.650000 ;
      LAYER met4 ;
        RECT 51.605000 7.330000 51.925000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 7.760000 51.925000 8.080000 ;
      LAYER met4 ;
        RECT 51.605000 7.760000 51.925000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 8.190000 51.925000 8.510000 ;
      LAYER met4 ;
        RECT 51.605000 8.190000 51.925000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 8.620000 51.925000 8.940000 ;
      LAYER met4 ;
        RECT 51.605000 8.620000 51.925000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 9.050000 51.925000 9.370000 ;
      LAYER met4 ;
        RECT 51.605000 9.050000 51.925000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 9.480000 51.925000 9.800000 ;
      LAYER met4 ;
        RECT 51.605000 9.480000 51.925000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 9.910000 51.925000 10.230000 ;
      LAYER met4 ;
        RECT 51.605000 9.910000 51.925000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 10.340000 52.335000 10.660000 ;
      LAYER met4 ;
        RECT 52.015000 10.340000 52.335000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 10.770000 52.335000 11.090000 ;
      LAYER met4 ;
        RECT 52.015000 10.770000 52.335000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 11.200000 52.335000 11.520000 ;
      LAYER met4 ;
        RECT 52.015000 11.200000 52.335000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 6.900000 52.335000 7.220000 ;
      LAYER met4 ;
        RECT 52.015000 6.900000 52.335000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 7.330000 52.335000 7.650000 ;
      LAYER met4 ;
        RECT 52.015000 7.330000 52.335000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 7.760000 52.335000 8.080000 ;
      LAYER met4 ;
        RECT 52.015000 7.760000 52.335000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 8.190000 52.335000 8.510000 ;
      LAYER met4 ;
        RECT 52.015000 8.190000 52.335000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 8.620000 52.335000 8.940000 ;
      LAYER met4 ;
        RECT 52.015000 8.620000 52.335000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 9.050000 52.335000 9.370000 ;
      LAYER met4 ;
        RECT 52.015000 9.050000 52.335000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 9.480000 52.335000 9.800000 ;
      LAYER met4 ;
        RECT 52.015000 9.480000 52.335000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 9.910000 52.335000 10.230000 ;
      LAYER met4 ;
        RECT 52.015000 9.910000 52.335000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 10.340000 52.745000 10.660000 ;
      LAYER met4 ;
        RECT 52.425000 10.340000 52.745000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 10.770000 52.745000 11.090000 ;
      LAYER met4 ;
        RECT 52.425000 10.770000 52.745000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 11.200000 52.745000 11.520000 ;
      LAYER met4 ;
        RECT 52.425000 11.200000 52.745000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 6.900000 52.745000 7.220000 ;
      LAYER met4 ;
        RECT 52.425000 6.900000 52.745000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 7.330000 52.745000 7.650000 ;
      LAYER met4 ;
        RECT 52.425000 7.330000 52.745000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 7.760000 52.745000 8.080000 ;
      LAYER met4 ;
        RECT 52.425000 7.760000 52.745000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 8.190000 52.745000 8.510000 ;
      LAYER met4 ;
        RECT 52.425000 8.190000 52.745000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 8.620000 52.745000 8.940000 ;
      LAYER met4 ;
        RECT 52.425000 8.620000 52.745000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 9.050000 52.745000 9.370000 ;
      LAYER met4 ;
        RECT 52.425000 9.050000 52.745000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 9.480000 52.745000 9.800000 ;
      LAYER met4 ;
        RECT 52.425000 9.480000 52.745000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 9.910000 52.745000 10.230000 ;
      LAYER met4 ;
        RECT 52.425000 9.910000 52.745000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 10.340000 53.155000 10.660000 ;
      LAYER met4 ;
        RECT 52.835000 10.340000 53.155000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 10.770000 53.155000 11.090000 ;
      LAYER met4 ;
        RECT 52.835000 10.770000 53.155000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 11.200000 53.155000 11.520000 ;
      LAYER met4 ;
        RECT 52.835000 11.200000 53.155000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 6.900000 53.155000 7.220000 ;
      LAYER met4 ;
        RECT 52.835000 6.900000 53.155000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 7.330000 53.155000 7.650000 ;
      LAYER met4 ;
        RECT 52.835000 7.330000 53.155000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 7.760000 53.155000 8.080000 ;
      LAYER met4 ;
        RECT 52.835000 7.760000 53.155000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 8.190000 53.155000 8.510000 ;
      LAYER met4 ;
        RECT 52.835000 8.190000 53.155000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 8.620000 53.155000 8.940000 ;
      LAYER met4 ;
        RECT 52.835000 8.620000 53.155000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 9.050000 53.155000 9.370000 ;
      LAYER met4 ;
        RECT 52.835000 9.050000 53.155000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 9.480000 53.155000 9.800000 ;
      LAYER met4 ;
        RECT 52.835000 9.480000 53.155000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 9.910000 53.155000 10.230000 ;
      LAYER met4 ;
        RECT 52.835000 9.910000 53.155000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 10.340000 53.565000 10.660000 ;
      LAYER met4 ;
        RECT 53.245000 10.340000 53.565000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 10.770000 53.565000 11.090000 ;
      LAYER met4 ;
        RECT 53.245000 10.770000 53.565000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 11.200000 53.565000 11.520000 ;
      LAYER met4 ;
        RECT 53.245000 11.200000 53.565000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 6.900000 53.565000 7.220000 ;
      LAYER met4 ;
        RECT 53.245000 6.900000 53.565000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 7.330000 53.565000 7.650000 ;
      LAYER met4 ;
        RECT 53.245000 7.330000 53.565000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 7.760000 53.565000 8.080000 ;
      LAYER met4 ;
        RECT 53.245000 7.760000 53.565000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 8.190000 53.565000 8.510000 ;
      LAYER met4 ;
        RECT 53.245000 8.190000 53.565000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 8.620000 53.565000 8.940000 ;
      LAYER met4 ;
        RECT 53.245000 8.620000 53.565000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 9.050000 53.565000 9.370000 ;
      LAYER met4 ;
        RECT 53.245000 9.050000 53.565000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 9.480000 53.565000 9.800000 ;
      LAYER met4 ;
        RECT 53.245000 9.480000 53.565000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 9.910000 53.565000 10.230000 ;
      LAYER met4 ;
        RECT 53.245000 9.910000 53.565000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 10.340000 53.970000 10.660000 ;
      LAYER met4 ;
        RECT 53.650000 10.340000 53.970000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 10.770000 53.970000 11.090000 ;
      LAYER met4 ;
        RECT 53.650000 10.770000 53.970000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 11.200000 53.970000 11.520000 ;
      LAYER met4 ;
        RECT 53.650000 11.200000 53.970000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 6.900000 53.970000 7.220000 ;
      LAYER met4 ;
        RECT 53.650000 6.900000 53.970000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 7.330000 53.970000 7.650000 ;
      LAYER met4 ;
        RECT 53.650000 7.330000 53.970000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 7.760000 53.970000 8.080000 ;
      LAYER met4 ;
        RECT 53.650000 7.760000 53.970000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 8.190000 53.970000 8.510000 ;
      LAYER met4 ;
        RECT 53.650000 8.190000 53.970000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 8.620000 53.970000 8.940000 ;
      LAYER met4 ;
        RECT 53.650000 8.620000 53.970000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 9.050000 53.970000 9.370000 ;
      LAYER met4 ;
        RECT 53.650000 9.050000 53.970000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 9.480000 53.970000 9.800000 ;
      LAYER met4 ;
        RECT 53.650000 9.480000 53.970000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 9.910000 53.970000 10.230000 ;
      LAYER met4 ;
        RECT 53.650000 9.910000 53.970000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 10.340000 54.375000 10.660000 ;
      LAYER met4 ;
        RECT 54.055000 10.340000 54.375000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 10.770000 54.375000 11.090000 ;
      LAYER met4 ;
        RECT 54.055000 10.770000 54.375000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 11.200000 54.375000 11.520000 ;
      LAYER met4 ;
        RECT 54.055000 11.200000 54.375000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 6.900000 54.375000 7.220000 ;
      LAYER met4 ;
        RECT 54.055000 6.900000 54.375000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 7.330000 54.375000 7.650000 ;
      LAYER met4 ;
        RECT 54.055000 7.330000 54.375000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 7.760000 54.375000 8.080000 ;
      LAYER met4 ;
        RECT 54.055000 7.760000 54.375000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 8.190000 54.375000 8.510000 ;
      LAYER met4 ;
        RECT 54.055000 8.190000 54.375000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 8.620000 54.375000 8.940000 ;
      LAYER met4 ;
        RECT 54.055000 8.620000 54.375000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 9.050000 54.375000 9.370000 ;
      LAYER met4 ;
        RECT 54.055000 9.050000 54.375000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 9.480000 54.375000 9.800000 ;
      LAYER met4 ;
        RECT 54.055000 9.480000 54.375000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 9.910000 54.375000 10.230000 ;
      LAYER met4 ;
        RECT 54.055000 9.910000 54.375000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 10.340000 54.780000 10.660000 ;
      LAYER met4 ;
        RECT 54.460000 10.340000 54.780000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 10.770000 54.780000 11.090000 ;
      LAYER met4 ;
        RECT 54.460000 10.770000 54.780000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 11.200000 54.780000 11.520000 ;
      LAYER met4 ;
        RECT 54.460000 11.200000 54.780000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 6.900000 54.780000 7.220000 ;
      LAYER met4 ;
        RECT 54.460000 6.900000 54.780000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 7.330000 54.780000 7.650000 ;
      LAYER met4 ;
        RECT 54.460000 7.330000 54.780000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 7.760000 54.780000 8.080000 ;
      LAYER met4 ;
        RECT 54.460000 7.760000 54.780000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 8.190000 54.780000 8.510000 ;
      LAYER met4 ;
        RECT 54.460000 8.190000 54.780000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 8.620000 54.780000 8.940000 ;
      LAYER met4 ;
        RECT 54.460000 8.620000 54.780000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 9.050000 54.780000 9.370000 ;
      LAYER met4 ;
        RECT 54.460000 9.050000 54.780000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 9.480000 54.780000 9.800000 ;
      LAYER met4 ;
        RECT 54.460000 9.480000 54.780000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 9.910000 54.780000 10.230000 ;
      LAYER met4 ;
        RECT 54.460000 9.910000 54.780000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 10.340000 55.185000 10.660000 ;
      LAYER met4 ;
        RECT 54.865000 10.340000 55.185000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 10.770000 55.185000 11.090000 ;
      LAYER met4 ;
        RECT 54.865000 10.770000 55.185000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 11.200000 55.185000 11.520000 ;
      LAYER met4 ;
        RECT 54.865000 11.200000 55.185000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 6.900000 55.185000 7.220000 ;
      LAYER met4 ;
        RECT 54.865000 6.900000 55.185000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 7.330000 55.185000 7.650000 ;
      LAYER met4 ;
        RECT 54.865000 7.330000 55.185000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 7.760000 55.185000 8.080000 ;
      LAYER met4 ;
        RECT 54.865000 7.760000 55.185000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 8.190000 55.185000 8.510000 ;
      LAYER met4 ;
        RECT 54.865000 8.190000 55.185000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 8.620000 55.185000 8.940000 ;
      LAYER met4 ;
        RECT 54.865000 8.620000 55.185000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 9.050000 55.185000 9.370000 ;
      LAYER met4 ;
        RECT 54.865000 9.050000 55.185000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 9.480000 55.185000 9.800000 ;
      LAYER met4 ;
        RECT 54.865000 9.480000 55.185000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 9.910000 55.185000 10.230000 ;
      LAYER met4 ;
        RECT 54.865000 9.910000 55.185000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 10.340000 55.590000 10.660000 ;
      LAYER met4 ;
        RECT 55.270000 10.340000 55.590000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 10.770000 55.590000 11.090000 ;
      LAYER met4 ;
        RECT 55.270000 10.770000 55.590000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 11.200000 55.590000 11.520000 ;
      LAYER met4 ;
        RECT 55.270000 11.200000 55.590000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 6.900000 55.590000 7.220000 ;
      LAYER met4 ;
        RECT 55.270000 6.900000 55.590000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 7.330000 55.590000 7.650000 ;
      LAYER met4 ;
        RECT 55.270000 7.330000 55.590000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 7.760000 55.590000 8.080000 ;
      LAYER met4 ;
        RECT 55.270000 7.760000 55.590000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 8.190000 55.590000 8.510000 ;
      LAYER met4 ;
        RECT 55.270000 8.190000 55.590000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 8.620000 55.590000 8.940000 ;
      LAYER met4 ;
        RECT 55.270000 8.620000 55.590000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 9.050000 55.590000 9.370000 ;
      LAYER met4 ;
        RECT 55.270000 9.050000 55.590000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 9.480000 55.590000 9.800000 ;
      LAYER met4 ;
        RECT 55.270000 9.480000 55.590000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 9.910000 55.590000 10.230000 ;
      LAYER met4 ;
        RECT 55.270000 9.910000 55.590000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 10.340000 55.995000 10.660000 ;
      LAYER met4 ;
        RECT 55.675000 10.340000 55.995000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 10.770000 55.995000 11.090000 ;
      LAYER met4 ;
        RECT 55.675000 10.770000 55.995000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 11.200000 55.995000 11.520000 ;
      LAYER met4 ;
        RECT 55.675000 11.200000 55.995000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 6.900000 55.995000 7.220000 ;
      LAYER met4 ;
        RECT 55.675000 6.900000 55.995000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 7.330000 55.995000 7.650000 ;
      LAYER met4 ;
        RECT 55.675000 7.330000 55.995000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 7.760000 55.995000 8.080000 ;
      LAYER met4 ;
        RECT 55.675000 7.760000 55.995000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 8.190000 55.995000 8.510000 ;
      LAYER met4 ;
        RECT 55.675000 8.190000 55.995000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 8.620000 55.995000 8.940000 ;
      LAYER met4 ;
        RECT 55.675000 8.620000 55.995000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 9.050000 55.995000 9.370000 ;
      LAYER met4 ;
        RECT 55.675000 9.050000 55.995000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 9.480000 55.995000 9.800000 ;
      LAYER met4 ;
        RECT 55.675000 9.480000 55.995000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 9.910000 55.995000 10.230000 ;
      LAYER met4 ;
        RECT 55.675000 9.910000 55.995000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 10.340000 56.400000 10.660000 ;
      LAYER met4 ;
        RECT 56.080000 10.340000 56.400000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 10.770000 56.400000 11.090000 ;
      LAYER met4 ;
        RECT 56.080000 10.770000 56.400000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 11.200000 56.400000 11.520000 ;
      LAYER met4 ;
        RECT 56.080000 11.200000 56.400000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 6.900000 56.400000 7.220000 ;
      LAYER met4 ;
        RECT 56.080000 6.900000 56.400000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 7.330000 56.400000 7.650000 ;
      LAYER met4 ;
        RECT 56.080000 7.330000 56.400000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 7.760000 56.400000 8.080000 ;
      LAYER met4 ;
        RECT 56.080000 7.760000 56.400000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 8.190000 56.400000 8.510000 ;
      LAYER met4 ;
        RECT 56.080000 8.190000 56.400000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 8.620000 56.400000 8.940000 ;
      LAYER met4 ;
        RECT 56.080000 8.620000 56.400000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 9.050000 56.400000 9.370000 ;
      LAYER met4 ;
        RECT 56.080000 9.050000 56.400000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 9.480000 56.400000 9.800000 ;
      LAYER met4 ;
        RECT 56.080000 9.480000 56.400000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 9.910000 56.400000 10.230000 ;
      LAYER met4 ;
        RECT 56.080000 9.910000 56.400000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 10.340000 56.805000 10.660000 ;
      LAYER met4 ;
        RECT 56.485000 10.340000 56.805000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 10.770000 56.805000 11.090000 ;
      LAYER met4 ;
        RECT 56.485000 10.770000 56.805000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 11.200000 56.805000 11.520000 ;
      LAYER met4 ;
        RECT 56.485000 11.200000 56.805000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 6.900000 56.805000 7.220000 ;
      LAYER met4 ;
        RECT 56.485000 6.900000 56.805000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 7.330000 56.805000 7.650000 ;
      LAYER met4 ;
        RECT 56.485000 7.330000 56.805000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 7.760000 56.805000 8.080000 ;
      LAYER met4 ;
        RECT 56.485000 7.760000 56.805000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 8.190000 56.805000 8.510000 ;
      LAYER met4 ;
        RECT 56.485000 8.190000 56.805000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 8.620000 56.805000 8.940000 ;
      LAYER met4 ;
        RECT 56.485000 8.620000 56.805000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 9.050000 56.805000 9.370000 ;
      LAYER met4 ;
        RECT 56.485000 9.050000 56.805000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 9.480000 56.805000 9.800000 ;
      LAYER met4 ;
        RECT 56.485000 9.480000 56.805000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 9.910000 56.805000 10.230000 ;
      LAYER met4 ;
        RECT 56.485000 9.910000 56.805000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 10.340000 57.210000 10.660000 ;
      LAYER met4 ;
        RECT 56.890000 10.340000 57.210000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 10.770000 57.210000 11.090000 ;
      LAYER met4 ;
        RECT 56.890000 10.770000 57.210000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 11.200000 57.210000 11.520000 ;
      LAYER met4 ;
        RECT 56.890000 11.200000 57.210000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 6.900000 57.210000 7.220000 ;
      LAYER met4 ;
        RECT 56.890000 6.900000 57.210000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 7.330000 57.210000 7.650000 ;
      LAYER met4 ;
        RECT 56.890000 7.330000 57.210000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 7.760000 57.210000 8.080000 ;
      LAYER met4 ;
        RECT 56.890000 7.760000 57.210000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 8.190000 57.210000 8.510000 ;
      LAYER met4 ;
        RECT 56.890000 8.190000 57.210000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 8.620000 57.210000 8.940000 ;
      LAYER met4 ;
        RECT 56.890000 8.620000 57.210000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 9.050000 57.210000 9.370000 ;
      LAYER met4 ;
        RECT 56.890000 9.050000 57.210000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 9.480000 57.210000 9.800000 ;
      LAYER met4 ;
        RECT 56.890000 9.480000 57.210000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 9.910000 57.210000 10.230000 ;
      LAYER met4 ;
        RECT 56.890000 9.910000 57.210000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 10.340000 57.615000 10.660000 ;
      LAYER met4 ;
        RECT 57.295000 10.340000 57.615000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 10.770000 57.615000 11.090000 ;
      LAYER met4 ;
        RECT 57.295000 10.770000 57.615000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 11.200000 57.615000 11.520000 ;
      LAYER met4 ;
        RECT 57.295000 11.200000 57.615000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 6.900000 57.615000 7.220000 ;
      LAYER met4 ;
        RECT 57.295000 6.900000 57.615000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 7.330000 57.615000 7.650000 ;
      LAYER met4 ;
        RECT 57.295000 7.330000 57.615000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 7.760000 57.615000 8.080000 ;
      LAYER met4 ;
        RECT 57.295000 7.760000 57.615000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 8.190000 57.615000 8.510000 ;
      LAYER met4 ;
        RECT 57.295000 8.190000 57.615000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 8.620000 57.615000 8.940000 ;
      LAYER met4 ;
        RECT 57.295000 8.620000 57.615000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 9.050000 57.615000 9.370000 ;
      LAYER met4 ;
        RECT 57.295000 9.050000 57.615000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 9.480000 57.615000 9.800000 ;
      LAYER met4 ;
        RECT 57.295000 9.480000 57.615000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 9.910000 57.615000 10.230000 ;
      LAYER met4 ;
        RECT 57.295000 9.910000 57.615000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 10.340000 58.020000 10.660000 ;
      LAYER met4 ;
        RECT 57.700000 10.340000 58.020000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 10.770000 58.020000 11.090000 ;
      LAYER met4 ;
        RECT 57.700000 10.770000 58.020000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 11.200000 58.020000 11.520000 ;
      LAYER met4 ;
        RECT 57.700000 11.200000 58.020000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 6.900000 58.020000 7.220000 ;
      LAYER met4 ;
        RECT 57.700000 6.900000 58.020000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 7.330000 58.020000 7.650000 ;
      LAYER met4 ;
        RECT 57.700000 7.330000 58.020000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 7.760000 58.020000 8.080000 ;
      LAYER met4 ;
        RECT 57.700000 7.760000 58.020000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 8.190000 58.020000 8.510000 ;
      LAYER met4 ;
        RECT 57.700000 8.190000 58.020000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 8.620000 58.020000 8.940000 ;
      LAYER met4 ;
        RECT 57.700000 8.620000 58.020000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 9.050000 58.020000 9.370000 ;
      LAYER met4 ;
        RECT 57.700000 9.050000 58.020000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 9.480000 58.020000 9.800000 ;
      LAYER met4 ;
        RECT 57.700000 9.480000 58.020000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 9.910000 58.020000 10.230000 ;
      LAYER met4 ;
        RECT 57.700000 9.910000 58.020000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 10.340000 58.425000 10.660000 ;
      LAYER met4 ;
        RECT 58.105000 10.340000 58.425000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 10.770000 58.425000 11.090000 ;
      LAYER met4 ;
        RECT 58.105000 10.770000 58.425000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 11.200000 58.425000 11.520000 ;
      LAYER met4 ;
        RECT 58.105000 11.200000 58.425000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 6.900000 58.425000 7.220000 ;
      LAYER met4 ;
        RECT 58.105000 6.900000 58.425000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 7.330000 58.425000 7.650000 ;
      LAYER met4 ;
        RECT 58.105000 7.330000 58.425000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 7.760000 58.425000 8.080000 ;
      LAYER met4 ;
        RECT 58.105000 7.760000 58.425000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 8.190000 58.425000 8.510000 ;
      LAYER met4 ;
        RECT 58.105000 8.190000 58.425000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 8.620000 58.425000 8.940000 ;
      LAYER met4 ;
        RECT 58.105000 8.620000 58.425000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 9.050000 58.425000 9.370000 ;
      LAYER met4 ;
        RECT 58.105000 9.050000 58.425000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 9.480000 58.425000 9.800000 ;
      LAYER met4 ;
        RECT 58.105000 9.480000 58.425000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 9.910000 58.425000 10.230000 ;
      LAYER met4 ;
        RECT 58.105000 9.910000 58.425000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 10.340000 58.830000 10.660000 ;
      LAYER met4 ;
        RECT 58.510000 10.340000 58.830000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 10.770000 58.830000 11.090000 ;
      LAYER met4 ;
        RECT 58.510000 10.770000 58.830000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 11.200000 58.830000 11.520000 ;
      LAYER met4 ;
        RECT 58.510000 11.200000 58.830000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 6.900000 58.830000 7.220000 ;
      LAYER met4 ;
        RECT 58.510000 6.900000 58.830000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 7.330000 58.830000 7.650000 ;
      LAYER met4 ;
        RECT 58.510000 7.330000 58.830000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 7.760000 58.830000 8.080000 ;
      LAYER met4 ;
        RECT 58.510000 7.760000 58.830000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 8.190000 58.830000 8.510000 ;
      LAYER met4 ;
        RECT 58.510000 8.190000 58.830000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 8.620000 58.830000 8.940000 ;
      LAYER met4 ;
        RECT 58.510000 8.620000 58.830000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 9.050000 58.830000 9.370000 ;
      LAYER met4 ;
        RECT 58.510000 9.050000 58.830000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 9.480000 58.830000 9.800000 ;
      LAYER met4 ;
        RECT 58.510000 9.480000 58.830000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 9.910000 58.830000 10.230000 ;
      LAYER met4 ;
        RECT 58.510000 9.910000 58.830000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 10.340000 59.235000 10.660000 ;
      LAYER met4 ;
        RECT 58.915000 10.340000 59.235000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 10.770000 59.235000 11.090000 ;
      LAYER met4 ;
        RECT 58.915000 10.770000 59.235000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 11.200000 59.235000 11.520000 ;
      LAYER met4 ;
        RECT 58.915000 11.200000 59.235000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 6.900000 59.235000 7.220000 ;
      LAYER met4 ;
        RECT 58.915000 6.900000 59.235000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 7.330000 59.235000 7.650000 ;
      LAYER met4 ;
        RECT 58.915000 7.330000 59.235000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 7.760000 59.235000 8.080000 ;
      LAYER met4 ;
        RECT 58.915000 7.760000 59.235000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 8.190000 59.235000 8.510000 ;
      LAYER met4 ;
        RECT 58.915000 8.190000 59.235000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 8.620000 59.235000 8.940000 ;
      LAYER met4 ;
        RECT 58.915000 8.620000 59.235000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 9.050000 59.235000 9.370000 ;
      LAYER met4 ;
        RECT 58.915000 9.050000 59.235000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 9.480000 59.235000 9.800000 ;
      LAYER met4 ;
        RECT 58.915000 9.480000 59.235000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 9.910000 59.235000 10.230000 ;
      LAYER met4 ;
        RECT 58.915000 9.910000 59.235000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 10.340000 59.640000 10.660000 ;
      LAYER met4 ;
        RECT 59.320000 10.340000 59.640000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 10.770000 59.640000 11.090000 ;
      LAYER met4 ;
        RECT 59.320000 10.770000 59.640000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 11.200000 59.640000 11.520000 ;
      LAYER met4 ;
        RECT 59.320000 11.200000 59.640000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 6.900000 59.640000 7.220000 ;
      LAYER met4 ;
        RECT 59.320000 6.900000 59.640000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 7.330000 59.640000 7.650000 ;
      LAYER met4 ;
        RECT 59.320000 7.330000 59.640000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 7.760000 59.640000 8.080000 ;
      LAYER met4 ;
        RECT 59.320000 7.760000 59.640000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 8.190000 59.640000 8.510000 ;
      LAYER met4 ;
        RECT 59.320000 8.190000 59.640000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 8.620000 59.640000 8.940000 ;
      LAYER met4 ;
        RECT 59.320000 8.620000 59.640000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 9.050000 59.640000 9.370000 ;
      LAYER met4 ;
        RECT 59.320000 9.050000 59.640000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 9.480000 59.640000 9.800000 ;
      LAYER met4 ;
        RECT 59.320000 9.480000 59.640000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 9.910000 59.640000 10.230000 ;
      LAYER met4 ;
        RECT 59.320000 9.910000 59.640000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 10.340000 60.045000 10.660000 ;
      LAYER met4 ;
        RECT 59.725000 10.340000 60.045000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 10.770000 60.045000 11.090000 ;
      LAYER met4 ;
        RECT 59.725000 10.770000 60.045000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 11.200000 60.045000 11.520000 ;
      LAYER met4 ;
        RECT 59.725000 11.200000 60.045000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 6.900000 60.045000 7.220000 ;
      LAYER met4 ;
        RECT 59.725000 6.900000 60.045000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 7.330000 60.045000 7.650000 ;
      LAYER met4 ;
        RECT 59.725000 7.330000 60.045000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 7.760000 60.045000 8.080000 ;
      LAYER met4 ;
        RECT 59.725000 7.760000 60.045000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 8.190000 60.045000 8.510000 ;
      LAYER met4 ;
        RECT 59.725000 8.190000 60.045000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 8.620000 60.045000 8.940000 ;
      LAYER met4 ;
        RECT 59.725000 8.620000 60.045000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 9.050000 60.045000 9.370000 ;
      LAYER met4 ;
        RECT 59.725000 9.050000 60.045000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 9.480000 60.045000 9.800000 ;
      LAYER met4 ;
        RECT 59.725000 9.480000 60.045000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 9.910000 60.045000 10.230000 ;
      LAYER met4 ;
        RECT 59.725000 9.910000 60.045000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330000 10.340000 6.650000 10.660000 ;
      LAYER met4 ;
        RECT 6.330000 10.340000 6.650000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330000 10.770000 6.650000 11.090000 ;
      LAYER met4 ;
        RECT 6.330000 10.770000 6.650000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330000 11.200000 6.650000 11.520000 ;
      LAYER met4 ;
        RECT 6.330000 11.200000 6.650000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330000 6.900000 6.650000 7.220000 ;
      LAYER met4 ;
        RECT 6.330000 6.900000 6.650000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330000 7.330000 6.650000 7.650000 ;
      LAYER met4 ;
        RECT 6.330000 7.330000 6.650000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330000 7.760000 6.650000 8.080000 ;
      LAYER met4 ;
        RECT 6.330000 7.760000 6.650000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330000 8.190000 6.650000 8.510000 ;
      LAYER met4 ;
        RECT 6.330000 8.190000 6.650000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330000 8.620000 6.650000 8.940000 ;
      LAYER met4 ;
        RECT 6.330000 8.620000 6.650000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330000 9.050000 6.650000 9.370000 ;
      LAYER met4 ;
        RECT 6.330000 9.050000 6.650000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330000 9.480000 6.650000 9.800000 ;
      LAYER met4 ;
        RECT 6.330000 9.480000 6.650000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330000 9.910000 6.650000 10.230000 ;
      LAYER met4 ;
        RECT 6.330000 9.910000 6.650000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735000 10.340000 7.055000 10.660000 ;
      LAYER met4 ;
        RECT 6.735000 10.340000 7.055000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735000 10.770000 7.055000 11.090000 ;
      LAYER met4 ;
        RECT 6.735000 10.770000 7.055000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735000 11.200000 7.055000 11.520000 ;
      LAYER met4 ;
        RECT 6.735000 11.200000 7.055000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735000 6.900000 7.055000 7.220000 ;
      LAYER met4 ;
        RECT 6.735000 6.900000 7.055000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735000 7.330000 7.055000 7.650000 ;
      LAYER met4 ;
        RECT 6.735000 7.330000 7.055000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735000 7.760000 7.055000 8.080000 ;
      LAYER met4 ;
        RECT 6.735000 7.760000 7.055000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735000 8.190000 7.055000 8.510000 ;
      LAYER met4 ;
        RECT 6.735000 8.190000 7.055000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735000 8.620000 7.055000 8.940000 ;
      LAYER met4 ;
        RECT 6.735000 8.620000 7.055000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735000 9.050000 7.055000 9.370000 ;
      LAYER met4 ;
        RECT 6.735000 9.050000 7.055000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735000 9.480000 7.055000 9.800000 ;
      LAYER met4 ;
        RECT 6.735000 9.480000 7.055000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735000 9.910000 7.055000 10.230000 ;
      LAYER met4 ;
        RECT 6.735000 9.910000 7.055000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 10.340000 60.450000 10.660000 ;
      LAYER met4 ;
        RECT 60.130000 10.340000 60.450000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 10.770000 60.450000 11.090000 ;
      LAYER met4 ;
        RECT 60.130000 10.770000 60.450000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 11.200000 60.450000 11.520000 ;
      LAYER met4 ;
        RECT 60.130000 11.200000 60.450000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 6.900000 60.450000 7.220000 ;
      LAYER met4 ;
        RECT 60.130000 6.900000 60.450000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 7.330000 60.450000 7.650000 ;
      LAYER met4 ;
        RECT 60.130000 7.330000 60.450000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 7.760000 60.450000 8.080000 ;
      LAYER met4 ;
        RECT 60.130000 7.760000 60.450000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 8.190000 60.450000 8.510000 ;
      LAYER met4 ;
        RECT 60.130000 8.190000 60.450000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 8.620000 60.450000 8.940000 ;
      LAYER met4 ;
        RECT 60.130000 8.620000 60.450000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 9.050000 60.450000 9.370000 ;
      LAYER met4 ;
        RECT 60.130000 9.050000 60.450000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 9.480000 60.450000 9.800000 ;
      LAYER met4 ;
        RECT 60.130000 9.480000 60.450000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 9.910000 60.450000 10.230000 ;
      LAYER met4 ;
        RECT 60.130000 9.910000 60.450000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 10.340000 60.855000 10.660000 ;
      LAYER met4 ;
        RECT 60.535000 10.340000 60.855000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 10.770000 60.855000 11.090000 ;
      LAYER met4 ;
        RECT 60.535000 10.770000 60.855000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 11.200000 60.855000 11.520000 ;
      LAYER met4 ;
        RECT 60.535000 11.200000 60.855000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 6.900000 60.855000 7.220000 ;
      LAYER met4 ;
        RECT 60.535000 6.900000 60.855000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 7.330000 60.855000 7.650000 ;
      LAYER met4 ;
        RECT 60.535000 7.330000 60.855000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 7.760000 60.855000 8.080000 ;
      LAYER met4 ;
        RECT 60.535000 7.760000 60.855000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 8.190000 60.855000 8.510000 ;
      LAYER met4 ;
        RECT 60.535000 8.190000 60.855000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 8.620000 60.855000 8.940000 ;
      LAYER met4 ;
        RECT 60.535000 8.620000 60.855000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 9.050000 60.855000 9.370000 ;
      LAYER met4 ;
        RECT 60.535000 9.050000 60.855000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 9.480000 60.855000 9.800000 ;
      LAYER met4 ;
        RECT 60.535000 9.480000 60.855000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 9.910000 60.855000 10.230000 ;
      LAYER met4 ;
        RECT 60.535000 9.910000 60.855000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 10.340000 61.260000 10.660000 ;
      LAYER met4 ;
        RECT 60.940000 10.340000 61.260000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 10.770000 61.260000 11.090000 ;
      LAYER met4 ;
        RECT 60.940000 10.770000 61.260000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 11.200000 61.260000 11.520000 ;
      LAYER met4 ;
        RECT 60.940000 11.200000 61.260000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 6.900000 61.260000 7.220000 ;
      LAYER met4 ;
        RECT 60.940000 6.900000 61.260000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 7.330000 61.260000 7.650000 ;
      LAYER met4 ;
        RECT 60.940000 7.330000 61.260000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 7.760000 61.260000 8.080000 ;
      LAYER met4 ;
        RECT 60.940000 7.760000 61.260000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 8.190000 61.260000 8.510000 ;
      LAYER met4 ;
        RECT 60.940000 8.190000 61.260000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 8.620000 61.260000 8.940000 ;
      LAYER met4 ;
        RECT 60.940000 8.620000 61.260000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 9.050000 61.260000 9.370000 ;
      LAYER met4 ;
        RECT 60.940000 9.050000 61.260000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 9.480000 61.260000 9.800000 ;
      LAYER met4 ;
        RECT 60.940000 9.480000 61.260000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 9.910000 61.260000 10.230000 ;
      LAYER met4 ;
        RECT 60.940000 9.910000 61.260000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 10.340000 61.665000 10.660000 ;
      LAYER met4 ;
        RECT 61.345000 10.340000 61.665000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 10.770000 61.665000 11.090000 ;
      LAYER met4 ;
        RECT 61.345000 10.770000 61.665000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 11.200000 61.665000 11.520000 ;
      LAYER met4 ;
        RECT 61.345000 11.200000 61.665000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 6.900000 61.665000 7.220000 ;
      LAYER met4 ;
        RECT 61.345000 6.900000 61.665000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 7.330000 61.665000 7.650000 ;
      LAYER met4 ;
        RECT 61.345000 7.330000 61.665000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 7.760000 61.665000 8.080000 ;
      LAYER met4 ;
        RECT 61.345000 7.760000 61.665000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 8.190000 61.665000 8.510000 ;
      LAYER met4 ;
        RECT 61.345000 8.190000 61.665000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 8.620000 61.665000 8.940000 ;
      LAYER met4 ;
        RECT 61.345000 8.620000 61.665000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 9.050000 61.665000 9.370000 ;
      LAYER met4 ;
        RECT 61.345000 9.050000 61.665000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 9.480000 61.665000 9.800000 ;
      LAYER met4 ;
        RECT 61.345000 9.480000 61.665000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 9.910000 61.665000 10.230000 ;
      LAYER met4 ;
        RECT 61.345000 9.910000 61.665000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 10.340000 62.070000 10.660000 ;
      LAYER met4 ;
        RECT 61.750000 10.340000 62.070000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 10.770000 62.070000 11.090000 ;
      LAYER met4 ;
        RECT 61.750000 10.770000 62.070000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 11.200000 62.070000 11.520000 ;
      LAYER met4 ;
        RECT 61.750000 11.200000 62.070000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 6.900000 62.070000 7.220000 ;
      LAYER met4 ;
        RECT 61.750000 6.900000 62.070000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 7.330000 62.070000 7.650000 ;
      LAYER met4 ;
        RECT 61.750000 7.330000 62.070000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 7.760000 62.070000 8.080000 ;
      LAYER met4 ;
        RECT 61.750000 7.760000 62.070000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 8.190000 62.070000 8.510000 ;
      LAYER met4 ;
        RECT 61.750000 8.190000 62.070000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 8.620000 62.070000 8.940000 ;
      LAYER met4 ;
        RECT 61.750000 8.620000 62.070000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 9.050000 62.070000 9.370000 ;
      LAYER met4 ;
        RECT 61.750000 9.050000 62.070000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 9.480000 62.070000 9.800000 ;
      LAYER met4 ;
        RECT 61.750000 9.480000 62.070000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 9.910000 62.070000 10.230000 ;
      LAYER met4 ;
        RECT 61.750000 9.910000 62.070000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 10.340000 62.475000 10.660000 ;
      LAYER met4 ;
        RECT 62.155000 10.340000 62.475000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 10.770000 62.475000 11.090000 ;
      LAYER met4 ;
        RECT 62.155000 10.770000 62.475000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 11.200000 62.475000 11.520000 ;
      LAYER met4 ;
        RECT 62.155000 11.200000 62.475000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 6.900000 62.475000 7.220000 ;
      LAYER met4 ;
        RECT 62.155000 6.900000 62.475000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 7.330000 62.475000 7.650000 ;
      LAYER met4 ;
        RECT 62.155000 7.330000 62.475000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 7.760000 62.475000 8.080000 ;
      LAYER met4 ;
        RECT 62.155000 7.760000 62.475000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 8.190000 62.475000 8.510000 ;
      LAYER met4 ;
        RECT 62.155000 8.190000 62.475000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 8.620000 62.475000 8.940000 ;
      LAYER met4 ;
        RECT 62.155000 8.620000 62.475000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 9.050000 62.475000 9.370000 ;
      LAYER met4 ;
        RECT 62.155000 9.050000 62.475000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 9.480000 62.475000 9.800000 ;
      LAYER met4 ;
        RECT 62.155000 9.480000 62.475000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 9.910000 62.475000 10.230000 ;
      LAYER met4 ;
        RECT 62.155000 9.910000 62.475000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 10.340000 62.880000 10.660000 ;
      LAYER met4 ;
        RECT 62.560000 10.340000 62.880000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 10.770000 62.880000 11.090000 ;
      LAYER met4 ;
        RECT 62.560000 10.770000 62.880000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 11.200000 62.880000 11.520000 ;
      LAYER met4 ;
        RECT 62.560000 11.200000 62.880000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 6.900000 62.880000 7.220000 ;
      LAYER met4 ;
        RECT 62.560000 6.900000 62.880000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 7.330000 62.880000 7.650000 ;
      LAYER met4 ;
        RECT 62.560000 7.330000 62.880000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 7.760000 62.880000 8.080000 ;
      LAYER met4 ;
        RECT 62.560000 7.760000 62.880000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 8.190000 62.880000 8.510000 ;
      LAYER met4 ;
        RECT 62.560000 8.190000 62.880000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 8.620000 62.880000 8.940000 ;
      LAYER met4 ;
        RECT 62.560000 8.620000 62.880000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 9.050000 62.880000 9.370000 ;
      LAYER met4 ;
        RECT 62.560000 9.050000 62.880000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 9.480000 62.880000 9.800000 ;
      LAYER met4 ;
        RECT 62.560000 9.480000 62.880000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 9.910000 62.880000 10.230000 ;
      LAYER met4 ;
        RECT 62.560000 9.910000 62.880000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 10.340000 63.285000 10.660000 ;
      LAYER met4 ;
        RECT 62.965000 10.340000 63.285000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 10.770000 63.285000 11.090000 ;
      LAYER met4 ;
        RECT 62.965000 10.770000 63.285000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 11.200000 63.285000 11.520000 ;
      LAYER met4 ;
        RECT 62.965000 11.200000 63.285000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 6.900000 63.285000 7.220000 ;
      LAYER met4 ;
        RECT 62.965000 6.900000 63.285000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 7.330000 63.285000 7.650000 ;
      LAYER met4 ;
        RECT 62.965000 7.330000 63.285000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 7.760000 63.285000 8.080000 ;
      LAYER met4 ;
        RECT 62.965000 7.760000 63.285000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 8.190000 63.285000 8.510000 ;
      LAYER met4 ;
        RECT 62.965000 8.190000 63.285000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 8.620000 63.285000 8.940000 ;
      LAYER met4 ;
        RECT 62.965000 8.620000 63.285000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 9.050000 63.285000 9.370000 ;
      LAYER met4 ;
        RECT 62.965000 9.050000 63.285000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 9.480000 63.285000 9.800000 ;
      LAYER met4 ;
        RECT 62.965000 9.480000 63.285000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 9.910000 63.285000 10.230000 ;
      LAYER met4 ;
        RECT 62.965000 9.910000 63.285000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 10.340000 63.690000 10.660000 ;
      LAYER met4 ;
        RECT 63.370000 10.340000 63.690000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 10.770000 63.690000 11.090000 ;
      LAYER met4 ;
        RECT 63.370000 10.770000 63.690000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 11.200000 63.690000 11.520000 ;
      LAYER met4 ;
        RECT 63.370000 11.200000 63.690000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 6.900000 63.690000 7.220000 ;
      LAYER met4 ;
        RECT 63.370000 6.900000 63.690000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 7.330000 63.690000 7.650000 ;
      LAYER met4 ;
        RECT 63.370000 7.330000 63.690000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 7.760000 63.690000 8.080000 ;
      LAYER met4 ;
        RECT 63.370000 7.760000 63.690000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 8.190000 63.690000 8.510000 ;
      LAYER met4 ;
        RECT 63.370000 8.190000 63.690000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 8.620000 63.690000 8.940000 ;
      LAYER met4 ;
        RECT 63.370000 8.620000 63.690000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 9.050000 63.690000 9.370000 ;
      LAYER met4 ;
        RECT 63.370000 9.050000 63.690000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 9.480000 63.690000 9.800000 ;
      LAYER met4 ;
        RECT 63.370000 9.480000 63.690000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 9.910000 63.690000 10.230000 ;
      LAYER met4 ;
        RECT 63.370000 9.910000 63.690000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 10.340000 64.095000 10.660000 ;
      LAYER met4 ;
        RECT 63.775000 10.340000 64.095000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 10.770000 64.095000 11.090000 ;
      LAYER met4 ;
        RECT 63.775000 10.770000 64.095000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 11.200000 64.095000 11.520000 ;
      LAYER met4 ;
        RECT 63.775000 11.200000 64.095000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 6.900000 64.095000 7.220000 ;
      LAYER met4 ;
        RECT 63.775000 6.900000 64.095000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 7.330000 64.095000 7.650000 ;
      LAYER met4 ;
        RECT 63.775000 7.330000 64.095000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 7.760000 64.095000 8.080000 ;
      LAYER met4 ;
        RECT 63.775000 7.760000 64.095000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 8.190000 64.095000 8.510000 ;
      LAYER met4 ;
        RECT 63.775000 8.190000 64.095000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 8.620000 64.095000 8.940000 ;
      LAYER met4 ;
        RECT 63.775000 8.620000 64.095000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 9.050000 64.095000 9.370000 ;
      LAYER met4 ;
        RECT 63.775000 9.050000 64.095000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 9.480000 64.095000 9.800000 ;
      LAYER met4 ;
        RECT 63.775000 9.480000 64.095000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 9.910000 64.095000 10.230000 ;
      LAYER met4 ;
        RECT 63.775000 9.910000 64.095000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 10.340000 64.500000 10.660000 ;
      LAYER met4 ;
        RECT 64.180000 10.340000 64.500000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 10.770000 64.500000 11.090000 ;
      LAYER met4 ;
        RECT 64.180000 10.770000 64.500000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 11.200000 64.500000 11.520000 ;
      LAYER met4 ;
        RECT 64.180000 11.200000 64.500000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 6.900000 64.500000 7.220000 ;
      LAYER met4 ;
        RECT 64.180000 6.900000 64.500000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 7.330000 64.500000 7.650000 ;
      LAYER met4 ;
        RECT 64.180000 7.330000 64.500000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 7.760000 64.500000 8.080000 ;
      LAYER met4 ;
        RECT 64.180000 7.760000 64.500000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 8.190000 64.500000 8.510000 ;
      LAYER met4 ;
        RECT 64.180000 8.190000 64.500000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 8.620000 64.500000 8.940000 ;
      LAYER met4 ;
        RECT 64.180000 8.620000 64.500000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 9.050000 64.500000 9.370000 ;
      LAYER met4 ;
        RECT 64.180000 9.050000 64.500000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 9.480000 64.500000 9.800000 ;
      LAYER met4 ;
        RECT 64.180000 9.480000 64.500000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 9.910000 64.500000 10.230000 ;
      LAYER met4 ;
        RECT 64.180000 9.910000 64.500000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 10.340000 64.905000 10.660000 ;
      LAYER met4 ;
        RECT 64.585000 10.340000 64.905000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 10.770000 64.905000 11.090000 ;
      LAYER met4 ;
        RECT 64.585000 10.770000 64.905000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 11.200000 64.905000 11.520000 ;
      LAYER met4 ;
        RECT 64.585000 11.200000 64.905000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 6.900000 64.905000 7.220000 ;
      LAYER met4 ;
        RECT 64.585000 6.900000 64.905000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 7.330000 64.905000 7.650000 ;
      LAYER met4 ;
        RECT 64.585000 7.330000 64.905000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 7.760000 64.905000 8.080000 ;
      LAYER met4 ;
        RECT 64.585000 7.760000 64.905000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 8.190000 64.905000 8.510000 ;
      LAYER met4 ;
        RECT 64.585000 8.190000 64.905000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 8.620000 64.905000 8.940000 ;
      LAYER met4 ;
        RECT 64.585000 8.620000 64.905000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 9.050000 64.905000 9.370000 ;
      LAYER met4 ;
        RECT 64.585000 9.050000 64.905000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 9.480000 64.905000 9.800000 ;
      LAYER met4 ;
        RECT 64.585000 9.480000 64.905000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 9.910000 64.905000 10.230000 ;
      LAYER met4 ;
        RECT 64.585000 9.910000 64.905000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 10.340000 65.310000 10.660000 ;
      LAYER met4 ;
        RECT 64.990000 10.340000 65.310000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 10.770000 65.310000 11.090000 ;
      LAYER met4 ;
        RECT 64.990000 10.770000 65.310000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 11.200000 65.310000 11.520000 ;
      LAYER met4 ;
        RECT 64.990000 11.200000 65.310000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 6.900000 65.310000 7.220000 ;
      LAYER met4 ;
        RECT 64.990000 6.900000 65.310000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 7.330000 65.310000 7.650000 ;
      LAYER met4 ;
        RECT 64.990000 7.330000 65.310000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 7.760000 65.310000 8.080000 ;
      LAYER met4 ;
        RECT 64.990000 7.760000 65.310000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 8.190000 65.310000 8.510000 ;
      LAYER met4 ;
        RECT 64.990000 8.190000 65.310000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 8.620000 65.310000 8.940000 ;
      LAYER met4 ;
        RECT 64.990000 8.620000 65.310000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 9.050000 65.310000 9.370000 ;
      LAYER met4 ;
        RECT 64.990000 9.050000 65.310000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 9.480000 65.310000 9.800000 ;
      LAYER met4 ;
        RECT 64.990000 9.480000 65.310000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 9.910000 65.310000 10.230000 ;
      LAYER met4 ;
        RECT 64.990000 9.910000 65.310000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 10.340000 65.715000 10.660000 ;
      LAYER met4 ;
        RECT 65.395000 10.340000 65.715000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 10.770000 65.715000 11.090000 ;
      LAYER met4 ;
        RECT 65.395000 10.770000 65.715000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 11.200000 65.715000 11.520000 ;
      LAYER met4 ;
        RECT 65.395000 11.200000 65.715000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 6.900000 65.715000 7.220000 ;
      LAYER met4 ;
        RECT 65.395000 6.900000 65.715000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 7.330000 65.715000 7.650000 ;
      LAYER met4 ;
        RECT 65.395000 7.330000 65.715000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 7.760000 65.715000 8.080000 ;
      LAYER met4 ;
        RECT 65.395000 7.760000 65.715000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 8.190000 65.715000 8.510000 ;
      LAYER met4 ;
        RECT 65.395000 8.190000 65.715000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 8.620000 65.715000 8.940000 ;
      LAYER met4 ;
        RECT 65.395000 8.620000 65.715000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 9.050000 65.715000 9.370000 ;
      LAYER met4 ;
        RECT 65.395000 9.050000 65.715000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 9.480000 65.715000 9.800000 ;
      LAYER met4 ;
        RECT 65.395000 9.480000 65.715000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 9.910000 65.715000 10.230000 ;
      LAYER met4 ;
        RECT 65.395000 9.910000 65.715000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 10.340000 66.120000 10.660000 ;
      LAYER met4 ;
        RECT 65.800000 10.340000 66.120000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 10.770000 66.120000 11.090000 ;
      LAYER met4 ;
        RECT 65.800000 10.770000 66.120000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 11.200000 66.120000 11.520000 ;
      LAYER met4 ;
        RECT 65.800000 11.200000 66.120000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 6.900000 66.120000 7.220000 ;
      LAYER met4 ;
        RECT 65.800000 6.900000 66.120000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 7.330000 66.120000 7.650000 ;
      LAYER met4 ;
        RECT 65.800000 7.330000 66.120000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 7.760000 66.120000 8.080000 ;
      LAYER met4 ;
        RECT 65.800000 7.760000 66.120000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 8.190000 66.120000 8.510000 ;
      LAYER met4 ;
        RECT 65.800000 8.190000 66.120000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 8.620000 66.120000 8.940000 ;
      LAYER met4 ;
        RECT 65.800000 8.620000 66.120000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 9.050000 66.120000 9.370000 ;
      LAYER met4 ;
        RECT 65.800000 9.050000 66.120000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 9.480000 66.120000 9.800000 ;
      LAYER met4 ;
        RECT 65.800000 9.480000 66.120000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 9.910000 66.120000 10.230000 ;
      LAYER met4 ;
        RECT 65.800000 9.910000 66.120000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 10.340000 66.525000 10.660000 ;
      LAYER met4 ;
        RECT 66.205000 10.340000 66.525000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 10.770000 66.525000 11.090000 ;
      LAYER met4 ;
        RECT 66.205000 10.770000 66.525000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 11.200000 66.525000 11.520000 ;
      LAYER met4 ;
        RECT 66.205000 11.200000 66.525000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 6.900000 66.525000 7.220000 ;
      LAYER met4 ;
        RECT 66.205000 6.900000 66.525000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 7.330000 66.525000 7.650000 ;
      LAYER met4 ;
        RECT 66.205000 7.330000 66.525000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 7.760000 66.525000 8.080000 ;
      LAYER met4 ;
        RECT 66.205000 7.760000 66.525000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 8.190000 66.525000 8.510000 ;
      LAYER met4 ;
        RECT 66.205000 8.190000 66.525000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 8.620000 66.525000 8.940000 ;
      LAYER met4 ;
        RECT 66.205000 8.620000 66.525000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 9.050000 66.525000 9.370000 ;
      LAYER met4 ;
        RECT 66.205000 9.050000 66.525000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 9.480000 66.525000 9.800000 ;
      LAYER met4 ;
        RECT 66.205000 9.480000 66.525000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 9.910000 66.525000 10.230000 ;
      LAYER met4 ;
        RECT 66.205000 9.910000 66.525000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 10.340000 66.930000 10.660000 ;
      LAYER met4 ;
        RECT 66.610000 10.340000 66.930000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 10.770000 66.930000 11.090000 ;
      LAYER met4 ;
        RECT 66.610000 10.770000 66.930000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 11.200000 66.930000 11.520000 ;
      LAYER met4 ;
        RECT 66.610000 11.200000 66.930000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 6.900000 66.930000 7.220000 ;
      LAYER met4 ;
        RECT 66.610000 6.900000 66.930000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 7.330000 66.930000 7.650000 ;
      LAYER met4 ;
        RECT 66.610000 7.330000 66.930000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 7.760000 66.930000 8.080000 ;
      LAYER met4 ;
        RECT 66.610000 7.760000 66.930000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 8.190000 66.930000 8.510000 ;
      LAYER met4 ;
        RECT 66.610000 8.190000 66.930000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 8.620000 66.930000 8.940000 ;
      LAYER met4 ;
        RECT 66.610000 8.620000 66.930000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 9.050000 66.930000 9.370000 ;
      LAYER met4 ;
        RECT 66.610000 9.050000 66.930000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 9.480000 66.930000 9.800000 ;
      LAYER met4 ;
        RECT 66.610000 9.480000 66.930000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 9.910000 66.930000 10.230000 ;
      LAYER met4 ;
        RECT 66.610000 9.910000 66.930000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 10.340000 67.335000 10.660000 ;
      LAYER met4 ;
        RECT 67.015000 10.340000 67.335000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 10.770000 67.335000 11.090000 ;
      LAYER met4 ;
        RECT 67.015000 10.770000 67.335000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 11.200000 67.335000 11.520000 ;
      LAYER met4 ;
        RECT 67.015000 11.200000 67.335000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 6.900000 67.335000 7.220000 ;
      LAYER met4 ;
        RECT 67.015000 6.900000 67.335000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 7.330000 67.335000 7.650000 ;
      LAYER met4 ;
        RECT 67.015000 7.330000 67.335000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 7.760000 67.335000 8.080000 ;
      LAYER met4 ;
        RECT 67.015000 7.760000 67.335000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 8.190000 67.335000 8.510000 ;
      LAYER met4 ;
        RECT 67.015000 8.190000 67.335000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 8.620000 67.335000 8.940000 ;
      LAYER met4 ;
        RECT 67.015000 8.620000 67.335000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 9.050000 67.335000 9.370000 ;
      LAYER met4 ;
        RECT 67.015000 9.050000 67.335000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 9.480000 67.335000 9.800000 ;
      LAYER met4 ;
        RECT 67.015000 9.480000 67.335000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 9.910000 67.335000 10.230000 ;
      LAYER met4 ;
        RECT 67.015000 9.910000 67.335000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 10.340000 67.740000 10.660000 ;
      LAYER met4 ;
        RECT 67.420000 10.340000 67.740000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 10.770000 67.740000 11.090000 ;
      LAYER met4 ;
        RECT 67.420000 10.770000 67.740000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 11.200000 67.740000 11.520000 ;
      LAYER met4 ;
        RECT 67.420000 11.200000 67.740000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 6.900000 67.740000 7.220000 ;
      LAYER met4 ;
        RECT 67.420000 6.900000 67.740000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 7.330000 67.740000 7.650000 ;
      LAYER met4 ;
        RECT 67.420000 7.330000 67.740000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 7.760000 67.740000 8.080000 ;
      LAYER met4 ;
        RECT 67.420000 7.760000 67.740000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 8.190000 67.740000 8.510000 ;
      LAYER met4 ;
        RECT 67.420000 8.190000 67.740000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 8.620000 67.740000 8.940000 ;
      LAYER met4 ;
        RECT 67.420000 8.620000 67.740000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 9.050000 67.740000 9.370000 ;
      LAYER met4 ;
        RECT 67.420000 9.050000 67.740000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 9.480000 67.740000 9.800000 ;
      LAYER met4 ;
        RECT 67.420000 9.480000 67.740000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 9.910000 67.740000 10.230000 ;
      LAYER met4 ;
        RECT 67.420000 9.910000 67.740000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 10.340000 68.145000 10.660000 ;
      LAYER met4 ;
        RECT 67.825000 10.340000 68.145000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 10.770000 68.145000 11.090000 ;
      LAYER met4 ;
        RECT 67.825000 10.770000 68.145000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 11.200000 68.145000 11.520000 ;
      LAYER met4 ;
        RECT 67.825000 11.200000 68.145000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 6.900000 68.145000 7.220000 ;
      LAYER met4 ;
        RECT 67.825000 6.900000 68.145000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 7.330000 68.145000 7.650000 ;
      LAYER met4 ;
        RECT 67.825000 7.330000 68.145000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 7.760000 68.145000 8.080000 ;
      LAYER met4 ;
        RECT 67.825000 7.760000 68.145000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 8.190000 68.145000 8.510000 ;
      LAYER met4 ;
        RECT 67.825000 8.190000 68.145000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 8.620000 68.145000 8.940000 ;
      LAYER met4 ;
        RECT 67.825000 8.620000 68.145000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 9.050000 68.145000 9.370000 ;
      LAYER met4 ;
        RECT 67.825000 9.050000 68.145000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 9.480000 68.145000 9.800000 ;
      LAYER met4 ;
        RECT 67.825000 9.480000 68.145000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 9.910000 68.145000 10.230000 ;
      LAYER met4 ;
        RECT 67.825000 9.910000 68.145000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 10.340000 68.550000 10.660000 ;
      LAYER met4 ;
        RECT 68.230000 10.340000 68.550000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 10.770000 68.550000 11.090000 ;
      LAYER met4 ;
        RECT 68.230000 10.770000 68.550000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 11.200000 68.550000 11.520000 ;
      LAYER met4 ;
        RECT 68.230000 11.200000 68.550000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 6.900000 68.550000 7.220000 ;
      LAYER met4 ;
        RECT 68.230000 6.900000 68.550000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 7.330000 68.550000 7.650000 ;
      LAYER met4 ;
        RECT 68.230000 7.330000 68.550000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 7.760000 68.550000 8.080000 ;
      LAYER met4 ;
        RECT 68.230000 7.760000 68.550000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 8.190000 68.550000 8.510000 ;
      LAYER met4 ;
        RECT 68.230000 8.190000 68.550000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 8.620000 68.550000 8.940000 ;
      LAYER met4 ;
        RECT 68.230000 8.620000 68.550000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 9.050000 68.550000 9.370000 ;
      LAYER met4 ;
        RECT 68.230000 9.050000 68.550000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 9.480000 68.550000 9.800000 ;
      LAYER met4 ;
        RECT 68.230000 9.480000 68.550000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 9.910000 68.550000 10.230000 ;
      LAYER met4 ;
        RECT 68.230000 9.910000 68.550000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 10.340000 68.955000 10.660000 ;
      LAYER met4 ;
        RECT 68.635000 10.340000 68.955000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 10.770000 68.955000 11.090000 ;
      LAYER met4 ;
        RECT 68.635000 10.770000 68.955000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 11.200000 68.955000 11.520000 ;
      LAYER met4 ;
        RECT 68.635000 11.200000 68.955000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 6.900000 68.955000 7.220000 ;
      LAYER met4 ;
        RECT 68.635000 6.900000 68.955000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 7.330000 68.955000 7.650000 ;
      LAYER met4 ;
        RECT 68.635000 7.330000 68.955000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 7.760000 68.955000 8.080000 ;
      LAYER met4 ;
        RECT 68.635000 7.760000 68.955000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 8.190000 68.955000 8.510000 ;
      LAYER met4 ;
        RECT 68.635000 8.190000 68.955000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 8.620000 68.955000 8.940000 ;
      LAYER met4 ;
        RECT 68.635000 8.620000 68.955000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 9.050000 68.955000 9.370000 ;
      LAYER met4 ;
        RECT 68.635000 9.050000 68.955000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 9.480000 68.955000 9.800000 ;
      LAYER met4 ;
        RECT 68.635000 9.480000 68.955000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 9.910000 68.955000 10.230000 ;
      LAYER met4 ;
        RECT 68.635000 9.910000 68.955000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 10.340000 69.360000 10.660000 ;
      LAYER met4 ;
        RECT 69.040000 10.340000 69.360000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 10.770000 69.360000 11.090000 ;
      LAYER met4 ;
        RECT 69.040000 10.770000 69.360000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 11.200000 69.360000 11.520000 ;
      LAYER met4 ;
        RECT 69.040000 11.200000 69.360000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 6.900000 69.360000 7.220000 ;
      LAYER met4 ;
        RECT 69.040000 6.900000 69.360000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 7.330000 69.360000 7.650000 ;
      LAYER met4 ;
        RECT 69.040000 7.330000 69.360000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 7.760000 69.360000 8.080000 ;
      LAYER met4 ;
        RECT 69.040000 7.760000 69.360000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 8.190000 69.360000 8.510000 ;
      LAYER met4 ;
        RECT 69.040000 8.190000 69.360000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 8.620000 69.360000 8.940000 ;
      LAYER met4 ;
        RECT 69.040000 8.620000 69.360000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 9.050000 69.360000 9.370000 ;
      LAYER met4 ;
        RECT 69.040000 9.050000 69.360000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 9.480000 69.360000 9.800000 ;
      LAYER met4 ;
        RECT 69.040000 9.480000 69.360000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 9.910000 69.360000 10.230000 ;
      LAYER met4 ;
        RECT 69.040000 9.910000 69.360000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 10.340000 69.765000 10.660000 ;
      LAYER met4 ;
        RECT 69.445000 10.340000 69.765000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 10.770000 69.765000 11.090000 ;
      LAYER met4 ;
        RECT 69.445000 10.770000 69.765000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 11.200000 69.765000 11.520000 ;
      LAYER met4 ;
        RECT 69.445000 11.200000 69.765000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 6.900000 69.765000 7.220000 ;
      LAYER met4 ;
        RECT 69.445000 6.900000 69.765000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 7.330000 69.765000 7.650000 ;
      LAYER met4 ;
        RECT 69.445000 7.330000 69.765000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 7.760000 69.765000 8.080000 ;
      LAYER met4 ;
        RECT 69.445000 7.760000 69.765000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 8.190000 69.765000 8.510000 ;
      LAYER met4 ;
        RECT 69.445000 8.190000 69.765000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 8.620000 69.765000 8.940000 ;
      LAYER met4 ;
        RECT 69.445000 8.620000 69.765000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 9.050000 69.765000 9.370000 ;
      LAYER met4 ;
        RECT 69.445000 9.050000 69.765000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 9.480000 69.765000 9.800000 ;
      LAYER met4 ;
        RECT 69.445000 9.480000 69.765000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 9.910000 69.765000 10.230000 ;
      LAYER met4 ;
        RECT 69.445000 9.910000 69.765000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 10.340000 70.170000 10.660000 ;
      LAYER met4 ;
        RECT 69.850000 10.340000 70.170000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 10.770000 70.170000 11.090000 ;
      LAYER met4 ;
        RECT 69.850000 10.770000 70.170000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 11.200000 70.170000 11.520000 ;
      LAYER met4 ;
        RECT 69.850000 11.200000 70.170000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 6.900000 70.170000 7.220000 ;
      LAYER met4 ;
        RECT 69.850000 6.900000 70.170000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 7.330000 70.170000 7.650000 ;
      LAYER met4 ;
        RECT 69.850000 7.330000 70.170000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 7.760000 70.170000 8.080000 ;
      LAYER met4 ;
        RECT 69.850000 7.760000 70.170000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 8.190000 70.170000 8.510000 ;
      LAYER met4 ;
        RECT 69.850000 8.190000 70.170000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 8.620000 70.170000 8.940000 ;
      LAYER met4 ;
        RECT 69.850000 8.620000 70.170000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 9.050000 70.170000 9.370000 ;
      LAYER met4 ;
        RECT 69.850000 9.050000 70.170000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 9.480000 70.170000 9.800000 ;
      LAYER met4 ;
        RECT 69.850000 9.480000 70.170000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 9.910000 70.170000 10.230000 ;
      LAYER met4 ;
        RECT 69.850000 9.910000 70.170000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140000 10.340000 7.460000 10.660000 ;
      LAYER met4 ;
        RECT 7.140000 10.340000 7.460000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140000 10.770000 7.460000 11.090000 ;
      LAYER met4 ;
        RECT 7.140000 10.770000 7.460000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140000 11.200000 7.460000 11.520000 ;
      LAYER met4 ;
        RECT 7.140000 11.200000 7.460000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140000 6.900000 7.460000 7.220000 ;
      LAYER met4 ;
        RECT 7.140000 6.900000 7.460000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140000 7.330000 7.460000 7.650000 ;
      LAYER met4 ;
        RECT 7.140000 7.330000 7.460000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140000 7.760000 7.460000 8.080000 ;
      LAYER met4 ;
        RECT 7.140000 7.760000 7.460000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140000 8.190000 7.460000 8.510000 ;
      LAYER met4 ;
        RECT 7.140000 8.190000 7.460000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140000 8.620000 7.460000 8.940000 ;
      LAYER met4 ;
        RECT 7.140000 8.620000 7.460000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140000 9.050000 7.460000 9.370000 ;
      LAYER met4 ;
        RECT 7.140000 9.050000 7.460000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140000 9.480000 7.460000 9.800000 ;
      LAYER met4 ;
        RECT 7.140000 9.480000 7.460000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140000 9.910000 7.460000 10.230000 ;
      LAYER met4 ;
        RECT 7.140000 9.910000 7.460000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545000 10.340000 7.865000 10.660000 ;
      LAYER met4 ;
        RECT 7.545000 10.340000 7.865000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545000 10.770000 7.865000 11.090000 ;
      LAYER met4 ;
        RECT 7.545000 10.770000 7.865000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545000 11.200000 7.865000 11.520000 ;
      LAYER met4 ;
        RECT 7.545000 11.200000 7.865000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545000 6.900000 7.865000 7.220000 ;
      LAYER met4 ;
        RECT 7.545000 6.900000 7.865000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545000 7.330000 7.865000 7.650000 ;
      LAYER met4 ;
        RECT 7.545000 7.330000 7.865000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545000 7.760000 7.865000 8.080000 ;
      LAYER met4 ;
        RECT 7.545000 7.760000 7.865000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545000 8.190000 7.865000 8.510000 ;
      LAYER met4 ;
        RECT 7.545000 8.190000 7.865000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545000 8.620000 7.865000 8.940000 ;
      LAYER met4 ;
        RECT 7.545000 8.620000 7.865000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545000 9.050000 7.865000 9.370000 ;
      LAYER met4 ;
        RECT 7.545000 9.050000 7.865000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545000 9.480000 7.865000 9.800000 ;
      LAYER met4 ;
        RECT 7.545000 9.480000 7.865000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545000 9.910000 7.865000 10.230000 ;
      LAYER met4 ;
        RECT 7.545000 9.910000 7.865000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950000 10.340000 8.270000 10.660000 ;
      LAYER met4 ;
        RECT 7.950000 10.340000 8.270000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950000 10.770000 8.270000 11.090000 ;
      LAYER met4 ;
        RECT 7.950000 10.770000 8.270000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950000 11.200000 8.270000 11.520000 ;
      LAYER met4 ;
        RECT 7.950000 11.200000 8.270000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950000 6.900000 8.270000 7.220000 ;
      LAYER met4 ;
        RECT 7.950000 6.900000 8.270000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950000 7.330000 8.270000 7.650000 ;
      LAYER met4 ;
        RECT 7.950000 7.330000 8.270000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950000 7.760000 8.270000 8.080000 ;
      LAYER met4 ;
        RECT 7.950000 7.760000 8.270000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950000 8.190000 8.270000 8.510000 ;
      LAYER met4 ;
        RECT 7.950000 8.190000 8.270000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950000 8.620000 8.270000 8.940000 ;
      LAYER met4 ;
        RECT 7.950000 8.620000 8.270000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950000 9.050000 8.270000 9.370000 ;
      LAYER met4 ;
        RECT 7.950000 9.050000 8.270000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950000 9.480000 8.270000 9.800000 ;
      LAYER met4 ;
        RECT 7.950000 9.480000 8.270000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950000 9.910000 8.270000 10.230000 ;
      LAYER met4 ;
        RECT 7.950000 9.910000 8.270000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 10.340000 70.575000 10.660000 ;
      LAYER met4 ;
        RECT 70.255000 10.340000 70.575000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 10.770000 70.575000 11.090000 ;
      LAYER met4 ;
        RECT 70.255000 10.770000 70.575000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 11.200000 70.575000 11.520000 ;
      LAYER met4 ;
        RECT 70.255000 11.200000 70.575000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 6.900000 70.575000 7.220000 ;
      LAYER met4 ;
        RECT 70.255000 6.900000 70.575000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 7.330000 70.575000 7.650000 ;
      LAYER met4 ;
        RECT 70.255000 7.330000 70.575000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 7.760000 70.575000 8.080000 ;
      LAYER met4 ;
        RECT 70.255000 7.760000 70.575000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 8.190000 70.575000 8.510000 ;
      LAYER met4 ;
        RECT 70.255000 8.190000 70.575000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 8.620000 70.575000 8.940000 ;
      LAYER met4 ;
        RECT 70.255000 8.620000 70.575000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 9.050000 70.575000 9.370000 ;
      LAYER met4 ;
        RECT 70.255000 9.050000 70.575000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 9.480000 70.575000 9.800000 ;
      LAYER met4 ;
        RECT 70.255000 9.480000 70.575000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 9.910000 70.575000 10.230000 ;
      LAYER met4 ;
        RECT 70.255000 9.910000 70.575000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 10.340000 70.980000 10.660000 ;
      LAYER met4 ;
        RECT 70.660000 10.340000 70.980000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 10.770000 70.980000 11.090000 ;
      LAYER met4 ;
        RECT 70.660000 10.770000 70.980000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 11.200000 70.980000 11.520000 ;
      LAYER met4 ;
        RECT 70.660000 11.200000 70.980000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 6.900000 70.980000 7.220000 ;
      LAYER met4 ;
        RECT 70.660000 6.900000 70.980000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 7.330000 70.980000 7.650000 ;
      LAYER met4 ;
        RECT 70.660000 7.330000 70.980000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 7.760000 70.980000 8.080000 ;
      LAYER met4 ;
        RECT 70.660000 7.760000 70.980000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 8.190000 70.980000 8.510000 ;
      LAYER met4 ;
        RECT 70.660000 8.190000 70.980000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 8.620000 70.980000 8.940000 ;
      LAYER met4 ;
        RECT 70.660000 8.620000 70.980000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 9.050000 70.980000 9.370000 ;
      LAYER met4 ;
        RECT 70.660000 9.050000 70.980000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 9.480000 70.980000 9.800000 ;
      LAYER met4 ;
        RECT 70.660000 9.480000 70.980000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 9.910000 70.980000 10.230000 ;
      LAYER met4 ;
        RECT 70.660000 9.910000 70.980000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 10.340000 71.385000 10.660000 ;
      LAYER met4 ;
        RECT 71.065000 10.340000 71.385000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 10.770000 71.385000 11.090000 ;
      LAYER met4 ;
        RECT 71.065000 10.770000 71.385000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 11.200000 71.385000 11.520000 ;
      LAYER met4 ;
        RECT 71.065000 11.200000 71.385000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 6.900000 71.385000 7.220000 ;
      LAYER met4 ;
        RECT 71.065000 6.900000 71.385000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 7.330000 71.385000 7.650000 ;
      LAYER met4 ;
        RECT 71.065000 7.330000 71.385000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 7.760000 71.385000 8.080000 ;
      LAYER met4 ;
        RECT 71.065000 7.760000 71.385000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 8.190000 71.385000 8.510000 ;
      LAYER met4 ;
        RECT 71.065000 8.190000 71.385000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 8.620000 71.385000 8.940000 ;
      LAYER met4 ;
        RECT 71.065000 8.620000 71.385000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 9.050000 71.385000 9.370000 ;
      LAYER met4 ;
        RECT 71.065000 9.050000 71.385000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 9.480000 71.385000 9.800000 ;
      LAYER met4 ;
        RECT 71.065000 9.480000 71.385000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 9.910000 71.385000 10.230000 ;
      LAYER met4 ;
        RECT 71.065000 9.910000 71.385000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 10.340000 71.790000 10.660000 ;
      LAYER met4 ;
        RECT 71.470000 10.340000 71.790000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 10.770000 71.790000 11.090000 ;
      LAYER met4 ;
        RECT 71.470000 10.770000 71.790000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 11.200000 71.790000 11.520000 ;
      LAYER met4 ;
        RECT 71.470000 11.200000 71.790000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 6.900000 71.790000 7.220000 ;
      LAYER met4 ;
        RECT 71.470000 6.900000 71.790000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 7.330000 71.790000 7.650000 ;
      LAYER met4 ;
        RECT 71.470000 7.330000 71.790000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 7.760000 71.790000 8.080000 ;
      LAYER met4 ;
        RECT 71.470000 7.760000 71.790000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 8.190000 71.790000 8.510000 ;
      LAYER met4 ;
        RECT 71.470000 8.190000 71.790000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 8.620000 71.790000 8.940000 ;
      LAYER met4 ;
        RECT 71.470000 8.620000 71.790000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 9.050000 71.790000 9.370000 ;
      LAYER met4 ;
        RECT 71.470000 9.050000 71.790000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 9.480000 71.790000 9.800000 ;
      LAYER met4 ;
        RECT 71.470000 9.480000 71.790000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 9.910000 71.790000 10.230000 ;
      LAYER met4 ;
        RECT 71.470000 9.910000 71.790000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 10.340000 72.195000 10.660000 ;
      LAYER met4 ;
        RECT 71.875000 10.340000 72.195000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 10.770000 72.195000 11.090000 ;
      LAYER met4 ;
        RECT 71.875000 10.770000 72.195000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 11.200000 72.195000 11.520000 ;
      LAYER met4 ;
        RECT 71.875000 11.200000 72.195000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 6.900000 72.195000 7.220000 ;
      LAYER met4 ;
        RECT 71.875000 6.900000 72.195000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 7.330000 72.195000 7.650000 ;
      LAYER met4 ;
        RECT 71.875000 7.330000 72.195000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 7.760000 72.195000 8.080000 ;
      LAYER met4 ;
        RECT 71.875000 7.760000 72.195000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 8.190000 72.195000 8.510000 ;
      LAYER met4 ;
        RECT 71.875000 8.190000 72.195000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 8.620000 72.195000 8.940000 ;
      LAYER met4 ;
        RECT 71.875000 8.620000 72.195000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 9.050000 72.195000 9.370000 ;
      LAYER met4 ;
        RECT 71.875000 9.050000 72.195000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 9.480000 72.195000 9.800000 ;
      LAYER met4 ;
        RECT 71.875000 9.480000 72.195000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 9.910000 72.195000 10.230000 ;
      LAYER met4 ;
        RECT 71.875000 9.910000 72.195000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 10.340000 72.600000 10.660000 ;
      LAYER met4 ;
        RECT 72.280000 10.340000 72.600000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 10.770000 72.600000 11.090000 ;
      LAYER met4 ;
        RECT 72.280000 10.770000 72.600000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 11.200000 72.600000 11.520000 ;
      LAYER met4 ;
        RECT 72.280000 11.200000 72.600000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 6.900000 72.600000 7.220000 ;
      LAYER met4 ;
        RECT 72.280000 6.900000 72.600000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 7.330000 72.600000 7.650000 ;
      LAYER met4 ;
        RECT 72.280000 7.330000 72.600000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 7.760000 72.600000 8.080000 ;
      LAYER met4 ;
        RECT 72.280000 7.760000 72.600000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 8.190000 72.600000 8.510000 ;
      LAYER met4 ;
        RECT 72.280000 8.190000 72.600000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 8.620000 72.600000 8.940000 ;
      LAYER met4 ;
        RECT 72.280000 8.620000 72.600000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 9.050000 72.600000 9.370000 ;
      LAYER met4 ;
        RECT 72.280000 9.050000 72.600000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 9.480000 72.600000 9.800000 ;
      LAYER met4 ;
        RECT 72.280000 9.480000 72.600000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 9.910000 72.600000 10.230000 ;
      LAYER met4 ;
        RECT 72.280000 9.910000 72.600000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 10.340000 73.005000 10.660000 ;
      LAYER met4 ;
        RECT 72.685000 10.340000 73.005000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 10.770000 73.005000 11.090000 ;
      LAYER met4 ;
        RECT 72.685000 10.770000 73.005000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 11.200000 73.005000 11.520000 ;
      LAYER met4 ;
        RECT 72.685000 11.200000 73.005000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 6.900000 73.005000 7.220000 ;
      LAYER met4 ;
        RECT 72.685000 6.900000 73.005000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 7.330000 73.005000 7.650000 ;
      LAYER met4 ;
        RECT 72.685000 7.330000 73.005000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 7.760000 73.005000 8.080000 ;
      LAYER met4 ;
        RECT 72.685000 7.760000 73.005000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 8.190000 73.005000 8.510000 ;
      LAYER met4 ;
        RECT 72.685000 8.190000 73.005000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 8.620000 73.005000 8.940000 ;
      LAYER met4 ;
        RECT 72.685000 8.620000 73.005000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 9.050000 73.005000 9.370000 ;
      LAYER met4 ;
        RECT 72.685000 9.050000 73.005000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 9.480000 73.005000 9.800000 ;
      LAYER met4 ;
        RECT 72.685000 9.480000 73.005000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 9.910000 73.005000 10.230000 ;
      LAYER met4 ;
        RECT 72.685000 9.910000 73.005000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 10.340000 73.410000 10.660000 ;
      LAYER met4 ;
        RECT 73.090000 10.340000 73.410000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 10.770000 73.410000 11.090000 ;
      LAYER met4 ;
        RECT 73.090000 10.770000 73.410000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 11.200000 73.410000 11.520000 ;
      LAYER met4 ;
        RECT 73.090000 11.200000 73.410000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 6.900000 73.410000 7.220000 ;
      LAYER met4 ;
        RECT 73.090000 6.900000 73.410000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 7.330000 73.410000 7.650000 ;
      LAYER met4 ;
        RECT 73.090000 7.330000 73.410000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 7.760000 73.410000 8.080000 ;
      LAYER met4 ;
        RECT 73.090000 7.760000 73.410000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 8.190000 73.410000 8.510000 ;
      LAYER met4 ;
        RECT 73.090000 8.190000 73.410000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 8.620000 73.410000 8.940000 ;
      LAYER met4 ;
        RECT 73.090000 8.620000 73.410000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 9.050000 73.410000 9.370000 ;
      LAYER met4 ;
        RECT 73.090000 9.050000 73.410000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 9.480000 73.410000 9.800000 ;
      LAYER met4 ;
        RECT 73.090000 9.480000 73.410000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 9.910000 73.410000 10.230000 ;
      LAYER met4 ;
        RECT 73.090000 9.910000 73.410000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 10.340000 73.815000 10.660000 ;
      LAYER met4 ;
        RECT 73.495000 10.340000 73.815000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 10.770000 73.815000 11.090000 ;
      LAYER met4 ;
        RECT 73.495000 10.770000 73.815000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 11.200000 73.815000 11.520000 ;
      LAYER met4 ;
        RECT 73.495000 11.200000 73.815000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 6.900000 73.815000 7.220000 ;
      LAYER met4 ;
        RECT 73.495000 6.900000 73.815000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 7.330000 73.815000 7.650000 ;
      LAYER met4 ;
        RECT 73.495000 7.330000 73.815000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 7.760000 73.815000 8.080000 ;
      LAYER met4 ;
        RECT 73.495000 7.760000 73.815000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 8.190000 73.815000 8.510000 ;
      LAYER met4 ;
        RECT 73.495000 8.190000 73.815000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 8.620000 73.815000 8.940000 ;
      LAYER met4 ;
        RECT 73.495000 8.620000 73.815000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 9.050000 73.815000 9.370000 ;
      LAYER met4 ;
        RECT 73.495000 9.050000 73.815000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 9.480000 73.815000 9.800000 ;
      LAYER met4 ;
        RECT 73.495000 9.480000 73.815000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 9.910000 73.815000 10.230000 ;
      LAYER met4 ;
        RECT 73.495000 9.910000 73.815000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 10.340000 74.220000 10.660000 ;
      LAYER met4 ;
        RECT 73.900000 10.340000 74.220000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 10.770000 74.220000 11.090000 ;
      LAYER met4 ;
        RECT 73.900000 10.770000 74.220000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 11.200000 74.220000 11.520000 ;
      LAYER met4 ;
        RECT 73.900000 11.200000 74.220000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 6.900000 74.220000 7.220000 ;
      LAYER met4 ;
        RECT 73.900000 6.900000 74.220000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 7.330000 74.220000 7.650000 ;
      LAYER met4 ;
        RECT 73.900000 7.330000 74.220000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 7.760000 74.220000 8.080000 ;
      LAYER met4 ;
        RECT 73.900000 7.760000 74.220000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 8.190000 74.220000 8.510000 ;
      LAYER met4 ;
        RECT 73.900000 8.190000 74.220000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 8.620000 74.220000 8.940000 ;
      LAYER met4 ;
        RECT 73.900000 8.620000 74.220000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 9.050000 74.220000 9.370000 ;
      LAYER met4 ;
        RECT 73.900000 9.050000 74.220000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 9.480000 74.220000 9.800000 ;
      LAYER met4 ;
        RECT 73.900000 9.480000 74.220000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 9.910000 74.220000 10.230000 ;
      LAYER met4 ;
        RECT 73.900000 9.910000 74.220000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 10.340000 74.625000 10.660000 ;
      LAYER met4 ;
        RECT 74.305000 10.340000 74.625000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 10.770000 74.625000 11.090000 ;
      LAYER met4 ;
        RECT 74.305000 10.770000 74.625000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 11.200000 74.625000 11.520000 ;
      LAYER met4 ;
        RECT 74.305000 11.200000 74.625000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 6.900000 74.625000 7.220000 ;
      LAYER met4 ;
        RECT 74.305000 6.900000 74.625000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 7.330000 74.625000 7.650000 ;
      LAYER met4 ;
        RECT 74.305000 7.330000 74.625000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 7.760000 74.625000 8.080000 ;
      LAYER met4 ;
        RECT 74.305000 7.760000 74.625000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 8.190000 74.625000 8.510000 ;
      LAYER met4 ;
        RECT 74.305000 8.190000 74.625000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 8.620000 74.625000 8.940000 ;
      LAYER met4 ;
        RECT 74.305000 8.620000 74.625000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 9.050000 74.625000 9.370000 ;
      LAYER met4 ;
        RECT 74.305000 9.050000 74.625000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 9.480000 74.625000 9.800000 ;
      LAYER met4 ;
        RECT 74.305000 9.480000 74.625000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 9.910000 74.625000 10.230000 ;
      LAYER met4 ;
        RECT 74.305000 9.910000 74.625000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355000 10.340000 8.675000 10.660000 ;
      LAYER met4 ;
        RECT 8.355000 10.340000 8.675000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355000 10.770000 8.675000 11.090000 ;
      LAYER met4 ;
        RECT 8.355000 10.770000 8.675000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355000 11.200000 8.675000 11.520000 ;
      LAYER met4 ;
        RECT 8.355000 11.200000 8.675000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355000 6.900000 8.675000 7.220000 ;
      LAYER met4 ;
        RECT 8.355000 6.900000 8.675000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355000 7.330000 8.675000 7.650000 ;
      LAYER met4 ;
        RECT 8.355000 7.330000 8.675000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355000 7.760000 8.675000 8.080000 ;
      LAYER met4 ;
        RECT 8.355000 7.760000 8.675000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355000 8.190000 8.675000 8.510000 ;
      LAYER met4 ;
        RECT 8.355000 8.190000 8.675000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355000 8.620000 8.675000 8.940000 ;
      LAYER met4 ;
        RECT 8.355000 8.620000 8.675000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355000 9.050000 8.675000 9.370000 ;
      LAYER met4 ;
        RECT 8.355000 9.050000 8.675000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355000 9.480000 8.675000 9.800000 ;
      LAYER met4 ;
        RECT 8.355000 9.480000 8.675000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355000 9.910000 8.675000 10.230000 ;
      LAYER met4 ;
        RECT 8.355000 9.910000 8.675000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760000 10.340000 9.080000 10.660000 ;
      LAYER met4 ;
        RECT 8.760000 10.340000 9.080000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760000 10.770000 9.080000 11.090000 ;
      LAYER met4 ;
        RECT 8.760000 10.770000 9.080000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760000 11.200000 9.080000 11.520000 ;
      LAYER met4 ;
        RECT 8.760000 11.200000 9.080000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760000 6.900000 9.080000 7.220000 ;
      LAYER met4 ;
        RECT 8.760000 6.900000 9.080000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760000 7.330000 9.080000 7.650000 ;
      LAYER met4 ;
        RECT 8.760000 7.330000 9.080000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760000 7.760000 9.080000 8.080000 ;
      LAYER met4 ;
        RECT 8.760000 7.760000 9.080000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760000 8.190000 9.080000 8.510000 ;
      LAYER met4 ;
        RECT 8.760000 8.190000 9.080000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760000 8.620000 9.080000 8.940000 ;
      LAYER met4 ;
        RECT 8.760000 8.620000 9.080000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760000 9.050000 9.080000 9.370000 ;
      LAYER met4 ;
        RECT 8.760000 9.050000 9.080000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760000 9.480000 9.080000 9.800000 ;
      LAYER met4 ;
        RECT 8.760000 9.480000 9.080000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760000 9.910000 9.080000 10.230000 ;
      LAYER met4 ;
        RECT 8.760000 9.910000 9.080000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165000 10.340000 9.485000 10.660000 ;
      LAYER met4 ;
        RECT 9.165000 10.340000 9.485000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165000 10.770000 9.485000 11.090000 ;
      LAYER met4 ;
        RECT 9.165000 10.770000 9.485000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165000 11.200000 9.485000 11.520000 ;
      LAYER met4 ;
        RECT 9.165000 11.200000 9.485000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165000 6.900000 9.485000 7.220000 ;
      LAYER met4 ;
        RECT 9.165000 6.900000 9.485000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165000 7.330000 9.485000 7.650000 ;
      LAYER met4 ;
        RECT 9.165000 7.330000 9.485000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165000 7.760000 9.485000 8.080000 ;
      LAYER met4 ;
        RECT 9.165000 7.760000 9.485000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165000 8.190000 9.485000 8.510000 ;
      LAYER met4 ;
        RECT 9.165000 8.190000 9.485000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165000 8.620000 9.485000 8.940000 ;
      LAYER met4 ;
        RECT 9.165000 8.620000 9.485000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165000 9.050000 9.485000 9.370000 ;
      LAYER met4 ;
        RECT 9.165000 9.050000 9.485000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165000 9.480000 9.485000 9.800000 ;
      LAYER met4 ;
        RECT 9.165000 9.480000 9.485000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165000 9.910000 9.485000 10.230000 ;
      LAYER met4 ;
        RECT 9.165000 9.910000 9.485000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570000 10.340000 9.890000 10.660000 ;
      LAYER met4 ;
        RECT 9.570000 10.340000 9.890000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570000 10.770000 9.890000 11.090000 ;
      LAYER met4 ;
        RECT 9.570000 10.770000 9.890000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570000 11.200000 9.890000 11.520000 ;
      LAYER met4 ;
        RECT 9.570000 11.200000 9.890000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570000 6.900000 9.890000 7.220000 ;
      LAYER met4 ;
        RECT 9.570000 6.900000 9.890000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570000 7.330000 9.890000 7.650000 ;
      LAYER met4 ;
        RECT 9.570000 7.330000 9.890000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570000 7.760000 9.890000 8.080000 ;
      LAYER met4 ;
        RECT 9.570000 7.760000 9.890000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570000 8.190000 9.890000 8.510000 ;
      LAYER met4 ;
        RECT 9.570000 8.190000 9.890000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570000 8.620000 9.890000 8.940000 ;
      LAYER met4 ;
        RECT 9.570000 8.620000 9.890000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570000 9.050000 9.890000 9.370000 ;
      LAYER met4 ;
        RECT 9.570000 9.050000 9.890000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570000 9.480000 9.890000 9.800000 ;
      LAYER met4 ;
        RECT 9.570000 9.480000 9.890000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570000 9.910000 9.890000 10.230000 ;
      LAYER met4 ;
        RECT 9.570000 9.910000 9.890000 10.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975000 10.340000 10.295000 10.660000 ;
      LAYER met4 ;
        RECT 9.975000 10.340000 10.295000 10.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975000 10.770000 10.295000 11.090000 ;
      LAYER met4 ;
        RECT 9.975000 10.770000 10.295000 11.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975000 11.200000 10.295000 11.520000 ;
      LAYER met4 ;
        RECT 9.975000 11.200000 10.295000 11.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975000 6.900000 10.295000 7.220000 ;
      LAYER met4 ;
        RECT 9.975000 6.900000 10.295000 7.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975000 7.330000 10.295000 7.650000 ;
      LAYER met4 ;
        RECT 9.975000 7.330000 10.295000 7.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975000 7.760000 10.295000 8.080000 ;
      LAYER met4 ;
        RECT 9.975000 7.760000 10.295000 8.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975000 8.190000 10.295000 8.510000 ;
      LAYER met4 ;
        RECT 9.975000 8.190000 10.295000 8.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975000 8.620000 10.295000 8.940000 ;
      LAYER met4 ;
        RECT 9.975000 8.620000 10.295000 8.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975000 9.050000 10.295000 9.370000 ;
      LAYER met4 ;
        RECT 9.975000 9.050000 10.295000 9.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975000 9.480000 10.295000 9.800000 ;
      LAYER met4 ;
        RECT 9.975000 9.480000 10.295000 9.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975000 9.910000 10.295000 10.230000 ;
      LAYER met4 ;
        RECT 9.975000 9.910000 10.295000 10.230000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met3 ;
      RECT 0.600000 6.890000 74.655000 11.530000 ;
    LAYER met4 ;
      RECT 0.000000  0.035000 75.000000  45.965000 ;
      RECT 0.000000 49.745000 75.000000  50.725000 ;
      RECT 0.000000 54.505000 75.000000 198.000000 ;
    LAYER met5 ;
      RECT 0.000000  0.135000 72.130000   6.985000 ;
      RECT 0.000000  6.985000 75.000000  11.435000 ;
      RECT 0.000000 11.435000 72.435000  17.885000 ;
      RECT 0.000000 17.885000 75.000000  22.335000 ;
      RECT 0.000000 22.335000 72.130000  34.835000 ;
      RECT 0.000000 34.835000 75.000000  38.085000 ;
      RECT 0.000000 38.085000 72.130000  94.585000 ;
      RECT 0.000000 94.585000 75.000000 198.000000 ;
  END
END sky130_fd_io__overlay_vccd_lvc
END LIBRARY
