/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_IO__TOP_SIO_SYMBOL_V
`define SKY130_FD_IO__TOP_SIO_SYMBOL_V

/**
 * top_sio: Special I/O PAD that provides additionally a
 *          regulated output buffer and a differential input buffer.
 *          SIO cells are ONLY available IN pairs (see top_sio_macro).
 *
 * Verilog stub (without power pins) for graphical symbol definition
 * generation.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_io__top_sio (
           //# {{data|Data Signals}}
           input        SLOW         ,
           output       IN           ,
           input        INP_DIS      ,
           output       IN_H         ,
           input        OUT          ,
           inout        PAD          ,
           inout        PAD_A_ESD_0_H,
           inout        PAD_A_ESD_1_H,
           inout        PAD_A_NOESD_H,

           //# {{control|Control Signals}}
           input  [2:0] DM           ,
           input        ENABLE_H     ,
           input        HLD_H_N      ,
           input        HLD_OVR      ,
           input        IBUF_SEL     ,
           input        OE_N         ,

           //# {{power|Power}}
           input        VREG_EN      ,
           input        VTRIP_SEL    ,
           input        REFLEAK_BIAS ,
           input        VINREF       ,
           input        VOUTREF      ,
           output       TIE_LO_ESD
       );

// Voltage supply signals
supply0 VSSIO  ;
supply0 VSSIO_Q;
supply0 VSSD   ;
supply1 VCCD   ;
supply1 VDDIO  ;
supply1 VCCHIB ;
supply1 VDDIO_Q;

endmodule

`default_nettype wire
`endif  // SKY130_FD_IO__TOP_SIO_SYMBOL_V
