# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__overlay_vdda_hvc
  CLASS BLOCK ;
  FOREIGN sky130_fd_io__overlay_vdda_hvc ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  75.00000 BY  200.0000 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.525000 14.960000 0.845000 15.280000 ;
      LAYER met4 ;
        RECT 0.525000 14.960000 0.845000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 15.400000 0.845000 15.720000 ;
      LAYER met4 ;
        RECT 0.525000 15.400000 0.845000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 15.840000 0.845000 16.160000 ;
      LAYER met4 ;
        RECT 0.525000 15.840000 0.845000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 16.280000 0.845000 16.600000 ;
      LAYER met4 ;
        RECT 0.525000 16.280000 0.845000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 16.720000 0.845000 17.040000 ;
      LAYER met4 ;
        RECT 0.525000 16.720000 0.845000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 17.160000 0.845000 17.480000 ;
      LAYER met4 ;
        RECT 0.525000 17.160000 0.845000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 17.600000 0.845000 17.920000 ;
      LAYER met4 ;
        RECT 0.525000 17.600000 0.845000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 18.040000 0.845000 18.360000 ;
      LAYER met4 ;
        RECT 0.525000 18.040000 0.845000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 14.960000 1.255000 15.280000 ;
      LAYER met4 ;
        RECT 0.935000 14.960000 1.255000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 15.400000 1.255000 15.720000 ;
      LAYER met4 ;
        RECT 0.935000 15.400000 1.255000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 15.840000 1.255000 16.160000 ;
      LAYER met4 ;
        RECT 0.935000 15.840000 1.255000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 16.280000 1.255000 16.600000 ;
      LAYER met4 ;
        RECT 0.935000 16.280000 1.255000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 16.720000 1.255000 17.040000 ;
      LAYER met4 ;
        RECT 0.935000 16.720000 1.255000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 17.160000 1.255000 17.480000 ;
      LAYER met4 ;
        RECT 0.935000 17.160000 1.255000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 17.600000 1.255000 17.920000 ;
      LAYER met4 ;
        RECT 0.935000 17.600000 1.255000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 18.040000 1.255000 18.360000 ;
      LAYER met4 ;
        RECT 0.935000 18.040000 1.255000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 14.960000 1.665000 15.280000 ;
      LAYER met4 ;
        RECT 1.345000 14.960000 1.665000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 15.400000 1.665000 15.720000 ;
      LAYER met4 ;
        RECT 1.345000 15.400000 1.665000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 15.840000 1.665000 16.160000 ;
      LAYER met4 ;
        RECT 1.345000 15.840000 1.665000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 16.280000 1.665000 16.600000 ;
      LAYER met4 ;
        RECT 1.345000 16.280000 1.665000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 16.720000 1.665000 17.040000 ;
      LAYER met4 ;
        RECT 1.345000 16.720000 1.665000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 17.160000 1.665000 17.480000 ;
      LAYER met4 ;
        RECT 1.345000 17.160000 1.665000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 17.600000 1.665000 17.920000 ;
      LAYER met4 ;
        RECT 1.345000 17.600000 1.665000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 18.040000 1.665000 18.360000 ;
      LAYER met4 ;
        RECT 1.345000 18.040000 1.665000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 14.960000 2.075000 15.280000 ;
      LAYER met4 ;
        RECT 1.755000 14.960000 2.075000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 15.400000 2.075000 15.720000 ;
      LAYER met4 ;
        RECT 1.755000 15.400000 2.075000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 15.840000 2.075000 16.160000 ;
      LAYER met4 ;
        RECT 1.755000 15.840000 2.075000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 16.280000 2.075000 16.600000 ;
      LAYER met4 ;
        RECT 1.755000 16.280000 2.075000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 16.720000 2.075000 17.040000 ;
      LAYER met4 ;
        RECT 1.755000 16.720000 2.075000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 17.160000 2.075000 17.480000 ;
      LAYER met4 ;
        RECT 1.755000 17.160000 2.075000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 17.600000 2.075000 17.920000 ;
      LAYER met4 ;
        RECT 1.755000 17.600000 2.075000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 18.040000 2.075000 18.360000 ;
      LAYER met4 ;
        RECT 1.755000 18.040000 2.075000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 14.960000 10.595000 15.280000 ;
      LAYER met4 ;
        RECT 10.275000 14.960000 10.595000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 15.400000 10.595000 15.720000 ;
      LAYER met4 ;
        RECT 10.275000 15.400000 10.595000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 15.840000 10.595000 16.160000 ;
      LAYER met4 ;
        RECT 10.275000 15.840000 10.595000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 16.280000 10.595000 16.600000 ;
      LAYER met4 ;
        RECT 10.275000 16.280000 10.595000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 16.720000 10.595000 17.040000 ;
      LAYER met4 ;
        RECT 10.275000 16.720000 10.595000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 17.160000 10.595000 17.480000 ;
      LAYER met4 ;
        RECT 10.275000 17.160000 10.595000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 17.600000 10.595000 17.920000 ;
      LAYER met4 ;
        RECT 10.275000 17.600000 10.595000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 18.040000 10.595000 18.360000 ;
      LAYER met4 ;
        RECT 10.275000 18.040000 10.595000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 14.960000 11.000000 15.280000 ;
      LAYER met4 ;
        RECT 10.680000 14.960000 11.000000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 15.400000 11.000000 15.720000 ;
      LAYER met4 ;
        RECT 10.680000 15.400000 11.000000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 15.840000 11.000000 16.160000 ;
      LAYER met4 ;
        RECT 10.680000 15.840000 11.000000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 16.280000 11.000000 16.600000 ;
      LAYER met4 ;
        RECT 10.680000 16.280000 11.000000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 16.720000 11.000000 17.040000 ;
      LAYER met4 ;
        RECT 10.680000 16.720000 11.000000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 17.160000 11.000000 17.480000 ;
      LAYER met4 ;
        RECT 10.680000 17.160000 11.000000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 17.600000 11.000000 17.920000 ;
      LAYER met4 ;
        RECT 10.680000 17.600000 11.000000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 18.040000 11.000000 18.360000 ;
      LAYER met4 ;
        RECT 10.680000 18.040000 11.000000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 14.960000 11.405000 15.280000 ;
      LAYER met4 ;
        RECT 11.085000 14.960000 11.405000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 15.400000 11.405000 15.720000 ;
      LAYER met4 ;
        RECT 11.085000 15.400000 11.405000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 15.840000 11.405000 16.160000 ;
      LAYER met4 ;
        RECT 11.085000 15.840000 11.405000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 16.280000 11.405000 16.600000 ;
      LAYER met4 ;
        RECT 11.085000 16.280000 11.405000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 16.720000 11.405000 17.040000 ;
      LAYER met4 ;
        RECT 11.085000 16.720000 11.405000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 17.160000 11.405000 17.480000 ;
      LAYER met4 ;
        RECT 11.085000 17.160000 11.405000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 17.600000 11.405000 17.920000 ;
      LAYER met4 ;
        RECT 11.085000 17.600000 11.405000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 18.040000 11.405000 18.360000 ;
      LAYER met4 ;
        RECT 11.085000 18.040000 11.405000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 14.960000 11.810000 15.280000 ;
      LAYER met4 ;
        RECT 11.490000 14.960000 11.810000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 15.400000 11.810000 15.720000 ;
      LAYER met4 ;
        RECT 11.490000 15.400000 11.810000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 15.840000 11.810000 16.160000 ;
      LAYER met4 ;
        RECT 11.490000 15.840000 11.810000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 16.280000 11.810000 16.600000 ;
      LAYER met4 ;
        RECT 11.490000 16.280000 11.810000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 16.720000 11.810000 17.040000 ;
      LAYER met4 ;
        RECT 11.490000 16.720000 11.810000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 17.160000 11.810000 17.480000 ;
      LAYER met4 ;
        RECT 11.490000 17.160000 11.810000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 17.600000 11.810000 17.920000 ;
      LAYER met4 ;
        RECT 11.490000 17.600000 11.810000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 18.040000 11.810000 18.360000 ;
      LAYER met4 ;
        RECT 11.490000 18.040000 11.810000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 14.960000 12.215000 15.280000 ;
      LAYER met4 ;
        RECT 11.895000 14.960000 12.215000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 15.400000 12.215000 15.720000 ;
      LAYER met4 ;
        RECT 11.895000 15.400000 12.215000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 15.840000 12.215000 16.160000 ;
      LAYER met4 ;
        RECT 11.895000 15.840000 12.215000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 16.280000 12.215000 16.600000 ;
      LAYER met4 ;
        RECT 11.895000 16.280000 12.215000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 16.720000 12.215000 17.040000 ;
      LAYER met4 ;
        RECT 11.895000 16.720000 12.215000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 17.160000 12.215000 17.480000 ;
      LAYER met4 ;
        RECT 11.895000 17.160000 12.215000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 17.600000 12.215000 17.920000 ;
      LAYER met4 ;
        RECT 11.895000 17.600000 12.215000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 18.040000 12.215000 18.360000 ;
      LAYER met4 ;
        RECT 11.895000 18.040000 12.215000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 14.960000 12.620000 15.280000 ;
      LAYER met4 ;
        RECT 12.300000 14.960000 12.620000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 15.400000 12.620000 15.720000 ;
      LAYER met4 ;
        RECT 12.300000 15.400000 12.620000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 15.840000 12.620000 16.160000 ;
      LAYER met4 ;
        RECT 12.300000 15.840000 12.620000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 16.280000 12.620000 16.600000 ;
      LAYER met4 ;
        RECT 12.300000 16.280000 12.620000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 16.720000 12.620000 17.040000 ;
      LAYER met4 ;
        RECT 12.300000 16.720000 12.620000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 17.160000 12.620000 17.480000 ;
      LAYER met4 ;
        RECT 12.300000 17.160000 12.620000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 17.600000 12.620000 17.920000 ;
      LAYER met4 ;
        RECT 12.300000 17.600000 12.620000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 18.040000 12.620000 18.360000 ;
      LAYER met4 ;
        RECT 12.300000 18.040000 12.620000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 14.960000 13.025000 15.280000 ;
      LAYER met4 ;
        RECT 12.705000 14.960000 13.025000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 15.400000 13.025000 15.720000 ;
      LAYER met4 ;
        RECT 12.705000 15.400000 13.025000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 15.840000 13.025000 16.160000 ;
      LAYER met4 ;
        RECT 12.705000 15.840000 13.025000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 16.280000 13.025000 16.600000 ;
      LAYER met4 ;
        RECT 12.705000 16.280000 13.025000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 16.720000 13.025000 17.040000 ;
      LAYER met4 ;
        RECT 12.705000 16.720000 13.025000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 17.160000 13.025000 17.480000 ;
      LAYER met4 ;
        RECT 12.705000 17.160000 13.025000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 17.600000 13.025000 17.920000 ;
      LAYER met4 ;
        RECT 12.705000 17.600000 13.025000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 18.040000 13.025000 18.360000 ;
      LAYER met4 ;
        RECT 12.705000 18.040000 13.025000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 14.960000 13.430000 15.280000 ;
      LAYER met4 ;
        RECT 13.110000 14.960000 13.430000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 15.400000 13.430000 15.720000 ;
      LAYER met4 ;
        RECT 13.110000 15.400000 13.430000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 15.840000 13.430000 16.160000 ;
      LAYER met4 ;
        RECT 13.110000 15.840000 13.430000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 16.280000 13.430000 16.600000 ;
      LAYER met4 ;
        RECT 13.110000 16.280000 13.430000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 16.720000 13.430000 17.040000 ;
      LAYER met4 ;
        RECT 13.110000 16.720000 13.430000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 17.160000 13.430000 17.480000 ;
      LAYER met4 ;
        RECT 13.110000 17.160000 13.430000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 17.600000 13.430000 17.920000 ;
      LAYER met4 ;
        RECT 13.110000 17.600000 13.430000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 18.040000 13.430000 18.360000 ;
      LAYER met4 ;
        RECT 13.110000 18.040000 13.430000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 14.960000 13.835000 15.280000 ;
      LAYER met4 ;
        RECT 13.515000 14.960000 13.835000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 15.400000 13.835000 15.720000 ;
      LAYER met4 ;
        RECT 13.515000 15.400000 13.835000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 15.840000 13.835000 16.160000 ;
      LAYER met4 ;
        RECT 13.515000 15.840000 13.835000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 16.280000 13.835000 16.600000 ;
      LAYER met4 ;
        RECT 13.515000 16.280000 13.835000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 16.720000 13.835000 17.040000 ;
      LAYER met4 ;
        RECT 13.515000 16.720000 13.835000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 17.160000 13.835000 17.480000 ;
      LAYER met4 ;
        RECT 13.515000 17.160000 13.835000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 17.600000 13.835000 17.920000 ;
      LAYER met4 ;
        RECT 13.515000 17.600000 13.835000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 18.040000 13.835000 18.360000 ;
      LAYER met4 ;
        RECT 13.515000 18.040000 13.835000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 14.960000 14.240000 15.280000 ;
      LAYER met4 ;
        RECT 13.920000 14.960000 14.240000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 15.400000 14.240000 15.720000 ;
      LAYER met4 ;
        RECT 13.920000 15.400000 14.240000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 15.840000 14.240000 16.160000 ;
      LAYER met4 ;
        RECT 13.920000 15.840000 14.240000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 16.280000 14.240000 16.600000 ;
      LAYER met4 ;
        RECT 13.920000 16.280000 14.240000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 16.720000 14.240000 17.040000 ;
      LAYER met4 ;
        RECT 13.920000 16.720000 14.240000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 17.160000 14.240000 17.480000 ;
      LAYER met4 ;
        RECT 13.920000 17.160000 14.240000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 17.600000 14.240000 17.920000 ;
      LAYER met4 ;
        RECT 13.920000 17.600000 14.240000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 18.040000 14.240000 18.360000 ;
      LAYER met4 ;
        RECT 13.920000 18.040000 14.240000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 14.960000 14.645000 15.280000 ;
      LAYER met4 ;
        RECT 14.325000 14.960000 14.645000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 15.400000 14.645000 15.720000 ;
      LAYER met4 ;
        RECT 14.325000 15.400000 14.645000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 15.840000 14.645000 16.160000 ;
      LAYER met4 ;
        RECT 14.325000 15.840000 14.645000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 16.280000 14.645000 16.600000 ;
      LAYER met4 ;
        RECT 14.325000 16.280000 14.645000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 16.720000 14.645000 17.040000 ;
      LAYER met4 ;
        RECT 14.325000 16.720000 14.645000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 17.160000 14.645000 17.480000 ;
      LAYER met4 ;
        RECT 14.325000 17.160000 14.645000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 17.600000 14.645000 17.920000 ;
      LAYER met4 ;
        RECT 14.325000 17.600000 14.645000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 18.040000 14.645000 18.360000 ;
      LAYER met4 ;
        RECT 14.325000 18.040000 14.645000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 14.960000 15.050000 15.280000 ;
      LAYER met4 ;
        RECT 14.730000 14.960000 15.050000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 15.400000 15.050000 15.720000 ;
      LAYER met4 ;
        RECT 14.730000 15.400000 15.050000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 15.840000 15.050000 16.160000 ;
      LAYER met4 ;
        RECT 14.730000 15.840000 15.050000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 16.280000 15.050000 16.600000 ;
      LAYER met4 ;
        RECT 14.730000 16.280000 15.050000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 16.720000 15.050000 17.040000 ;
      LAYER met4 ;
        RECT 14.730000 16.720000 15.050000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 17.160000 15.050000 17.480000 ;
      LAYER met4 ;
        RECT 14.730000 17.160000 15.050000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 17.600000 15.050000 17.920000 ;
      LAYER met4 ;
        RECT 14.730000 17.600000 15.050000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 18.040000 15.050000 18.360000 ;
      LAYER met4 ;
        RECT 14.730000 18.040000 15.050000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 14.960000 15.455000 15.280000 ;
      LAYER met4 ;
        RECT 15.135000 14.960000 15.455000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 15.400000 15.455000 15.720000 ;
      LAYER met4 ;
        RECT 15.135000 15.400000 15.455000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 15.840000 15.455000 16.160000 ;
      LAYER met4 ;
        RECT 15.135000 15.840000 15.455000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 16.280000 15.455000 16.600000 ;
      LAYER met4 ;
        RECT 15.135000 16.280000 15.455000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 16.720000 15.455000 17.040000 ;
      LAYER met4 ;
        RECT 15.135000 16.720000 15.455000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 17.160000 15.455000 17.480000 ;
      LAYER met4 ;
        RECT 15.135000 17.160000 15.455000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 17.600000 15.455000 17.920000 ;
      LAYER met4 ;
        RECT 15.135000 17.600000 15.455000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 18.040000 15.455000 18.360000 ;
      LAYER met4 ;
        RECT 15.135000 18.040000 15.455000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 14.960000 15.860000 15.280000 ;
      LAYER met4 ;
        RECT 15.540000 14.960000 15.860000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 15.400000 15.860000 15.720000 ;
      LAYER met4 ;
        RECT 15.540000 15.400000 15.860000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 15.840000 15.860000 16.160000 ;
      LAYER met4 ;
        RECT 15.540000 15.840000 15.860000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 16.280000 15.860000 16.600000 ;
      LAYER met4 ;
        RECT 15.540000 16.280000 15.860000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 16.720000 15.860000 17.040000 ;
      LAYER met4 ;
        RECT 15.540000 16.720000 15.860000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 17.160000 15.860000 17.480000 ;
      LAYER met4 ;
        RECT 15.540000 17.160000 15.860000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 17.600000 15.860000 17.920000 ;
      LAYER met4 ;
        RECT 15.540000 17.600000 15.860000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 18.040000 15.860000 18.360000 ;
      LAYER met4 ;
        RECT 15.540000 18.040000 15.860000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 14.960000 16.265000 15.280000 ;
      LAYER met4 ;
        RECT 15.945000 14.960000 16.265000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 15.400000 16.265000 15.720000 ;
      LAYER met4 ;
        RECT 15.945000 15.400000 16.265000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 15.840000 16.265000 16.160000 ;
      LAYER met4 ;
        RECT 15.945000 15.840000 16.265000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 16.280000 16.265000 16.600000 ;
      LAYER met4 ;
        RECT 15.945000 16.280000 16.265000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 16.720000 16.265000 17.040000 ;
      LAYER met4 ;
        RECT 15.945000 16.720000 16.265000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 17.160000 16.265000 17.480000 ;
      LAYER met4 ;
        RECT 15.945000 17.160000 16.265000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 17.600000 16.265000 17.920000 ;
      LAYER met4 ;
        RECT 15.945000 17.600000 16.265000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 18.040000 16.265000 18.360000 ;
      LAYER met4 ;
        RECT 15.945000 18.040000 16.265000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 14.960000 16.670000 15.280000 ;
      LAYER met4 ;
        RECT 16.350000 14.960000 16.670000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 15.400000 16.670000 15.720000 ;
      LAYER met4 ;
        RECT 16.350000 15.400000 16.670000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 15.840000 16.670000 16.160000 ;
      LAYER met4 ;
        RECT 16.350000 15.840000 16.670000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 16.280000 16.670000 16.600000 ;
      LAYER met4 ;
        RECT 16.350000 16.280000 16.670000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 16.720000 16.670000 17.040000 ;
      LAYER met4 ;
        RECT 16.350000 16.720000 16.670000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 17.160000 16.670000 17.480000 ;
      LAYER met4 ;
        RECT 16.350000 17.160000 16.670000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 17.600000 16.670000 17.920000 ;
      LAYER met4 ;
        RECT 16.350000 17.600000 16.670000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 18.040000 16.670000 18.360000 ;
      LAYER met4 ;
        RECT 16.350000 18.040000 16.670000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 14.960000 17.075000 15.280000 ;
      LAYER met4 ;
        RECT 16.755000 14.960000 17.075000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 15.400000 17.075000 15.720000 ;
      LAYER met4 ;
        RECT 16.755000 15.400000 17.075000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 15.840000 17.075000 16.160000 ;
      LAYER met4 ;
        RECT 16.755000 15.840000 17.075000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 16.280000 17.075000 16.600000 ;
      LAYER met4 ;
        RECT 16.755000 16.280000 17.075000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 16.720000 17.075000 17.040000 ;
      LAYER met4 ;
        RECT 16.755000 16.720000 17.075000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 17.160000 17.075000 17.480000 ;
      LAYER met4 ;
        RECT 16.755000 17.160000 17.075000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 17.600000 17.075000 17.920000 ;
      LAYER met4 ;
        RECT 16.755000 17.600000 17.075000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 18.040000 17.075000 18.360000 ;
      LAYER met4 ;
        RECT 16.755000 18.040000 17.075000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 14.960000 17.480000 15.280000 ;
      LAYER met4 ;
        RECT 17.160000 14.960000 17.480000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 15.400000 17.480000 15.720000 ;
      LAYER met4 ;
        RECT 17.160000 15.400000 17.480000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 15.840000 17.480000 16.160000 ;
      LAYER met4 ;
        RECT 17.160000 15.840000 17.480000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 16.280000 17.480000 16.600000 ;
      LAYER met4 ;
        RECT 17.160000 16.280000 17.480000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 16.720000 17.480000 17.040000 ;
      LAYER met4 ;
        RECT 17.160000 16.720000 17.480000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 17.160000 17.480000 17.480000 ;
      LAYER met4 ;
        RECT 17.160000 17.160000 17.480000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 17.600000 17.480000 17.920000 ;
      LAYER met4 ;
        RECT 17.160000 17.600000 17.480000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 18.040000 17.480000 18.360000 ;
      LAYER met4 ;
        RECT 17.160000 18.040000 17.480000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 14.960000 17.885000 15.280000 ;
      LAYER met4 ;
        RECT 17.565000 14.960000 17.885000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 15.400000 17.885000 15.720000 ;
      LAYER met4 ;
        RECT 17.565000 15.400000 17.885000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 15.840000 17.885000 16.160000 ;
      LAYER met4 ;
        RECT 17.565000 15.840000 17.885000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 16.280000 17.885000 16.600000 ;
      LAYER met4 ;
        RECT 17.565000 16.280000 17.885000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 16.720000 17.885000 17.040000 ;
      LAYER met4 ;
        RECT 17.565000 16.720000 17.885000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 17.160000 17.885000 17.480000 ;
      LAYER met4 ;
        RECT 17.565000 17.160000 17.885000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 17.600000 17.885000 17.920000 ;
      LAYER met4 ;
        RECT 17.565000 17.600000 17.885000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 18.040000 17.885000 18.360000 ;
      LAYER met4 ;
        RECT 17.565000 18.040000 17.885000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 14.960000 18.290000 15.280000 ;
      LAYER met4 ;
        RECT 17.970000 14.960000 18.290000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 15.400000 18.290000 15.720000 ;
      LAYER met4 ;
        RECT 17.970000 15.400000 18.290000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 15.840000 18.290000 16.160000 ;
      LAYER met4 ;
        RECT 17.970000 15.840000 18.290000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 16.280000 18.290000 16.600000 ;
      LAYER met4 ;
        RECT 17.970000 16.280000 18.290000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 16.720000 18.290000 17.040000 ;
      LAYER met4 ;
        RECT 17.970000 16.720000 18.290000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 17.160000 18.290000 17.480000 ;
      LAYER met4 ;
        RECT 17.970000 17.160000 18.290000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 17.600000 18.290000 17.920000 ;
      LAYER met4 ;
        RECT 17.970000 17.600000 18.290000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 18.040000 18.290000 18.360000 ;
      LAYER met4 ;
        RECT 17.970000 18.040000 18.290000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 14.960000 18.695000 15.280000 ;
      LAYER met4 ;
        RECT 18.375000 14.960000 18.695000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 15.400000 18.695000 15.720000 ;
      LAYER met4 ;
        RECT 18.375000 15.400000 18.695000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 15.840000 18.695000 16.160000 ;
      LAYER met4 ;
        RECT 18.375000 15.840000 18.695000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 16.280000 18.695000 16.600000 ;
      LAYER met4 ;
        RECT 18.375000 16.280000 18.695000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 16.720000 18.695000 17.040000 ;
      LAYER met4 ;
        RECT 18.375000 16.720000 18.695000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 17.160000 18.695000 17.480000 ;
      LAYER met4 ;
        RECT 18.375000 17.160000 18.695000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 17.600000 18.695000 17.920000 ;
      LAYER met4 ;
        RECT 18.375000 17.600000 18.695000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 18.040000 18.695000 18.360000 ;
      LAYER met4 ;
        RECT 18.375000 18.040000 18.695000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 14.960000 19.100000 15.280000 ;
      LAYER met4 ;
        RECT 18.780000 14.960000 19.100000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 15.400000 19.100000 15.720000 ;
      LAYER met4 ;
        RECT 18.780000 15.400000 19.100000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 15.840000 19.100000 16.160000 ;
      LAYER met4 ;
        RECT 18.780000 15.840000 19.100000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 16.280000 19.100000 16.600000 ;
      LAYER met4 ;
        RECT 18.780000 16.280000 19.100000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 16.720000 19.100000 17.040000 ;
      LAYER met4 ;
        RECT 18.780000 16.720000 19.100000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 17.160000 19.100000 17.480000 ;
      LAYER met4 ;
        RECT 18.780000 17.160000 19.100000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 17.600000 19.100000 17.920000 ;
      LAYER met4 ;
        RECT 18.780000 17.600000 19.100000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 18.040000 19.100000 18.360000 ;
      LAYER met4 ;
        RECT 18.780000 18.040000 19.100000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 14.960000 19.505000 15.280000 ;
      LAYER met4 ;
        RECT 19.185000 14.960000 19.505000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 15.400000 19.505000 15.720000 ;
      LAYER met4 ;
        RECT 19.185000 15.400000 19.505000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 15.840000 19.505000 16.160000 ;
      LAYER met4 ;
        RECT 19.185000 15.840000 19.505000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 16.280000 19.505000 16.600000 ;
      LAYER met4 ;
        RECT 19.185000 16.280000 19.505000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 16.720000 19.505000 17.040000 ;
      LAYER met4 ;
        RECT 19.185000 16.720000 19.505000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 17.160000 19.505000 17.480000 ;
      LAYER met4 ;
        RECT 19.185000 17.160000 19.505000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 17.600000 19.505000 17.920000 ;
      LAYER met4 ;
        RECT 19.185000 17.600000 19.505000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 18.040000 19.505000 18.360000 ;
      LAYER met4 ;
        RECT 19.185000 18.040000 19.505000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 14.960000 19.910000 15.280000 ;
      LAYER met4 ;
        RECT 19.590000 14.960000 19.910000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 15.400000 19.910000 15.720000 ;
      LAYER met4 ;
        RECT 19.590000 15.400000 19.910000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 15.840000 19.910000 16.160000 ;
      LAYER met4 ;
        RECT 19.590000 15.840000 19.910000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 16.280000 19.910000 16.600000 ;
      LAYER met4 ;
        RECT 19.590000 16.280000 19.910000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 16.720000 19.910000 17.040000 ;
      LAYER met4 ;
        RECT 19.590000 16.720000 19.910000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 17.160000 19.910000 17.480000 ;
      LAYER met4 ;
        RECT 19.590000 17.160000 19.910000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 17.600000 19.910000 17.920000 ;
      LAYER met4 ;
        RECT 19.590000 17.600000 19.910000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 18.040000 19.910000 18.360000 ;
      LAYER met4 ;
        RECT 19.590000 18.040000 19.910000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 14.960000 20.315000 15.280000 ;
      LAYER met4 ;
        RECT 19.995000 14.960000 20.315000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 15.400000 20.315000 15.720000 ;
      LAYER met4 ;
        RECT 19.995000 15.400000 20.315000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 15.840000 20.315000 16.160000 ;
      LAYER met4 ;
        RECT 19.995000 15.840000 20.315000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 16.280000 20.315000 16.600000 ;
      LAYER met4 ;
        RECT 19.995000 16.280000 20.315000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 16.720000 20.315000 17.040000 ;
      LAYER met4 ;
        RECT 19.995000 16.720000 20.315000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 17.160000 20.315000 17.480000 ;
      LAYER met4 ;
        RECT 19.995000 17.160000 20.315000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 17.600000 20.315000 17.920000 ;
      LAYER met4 ;
        RECT 19.995000 17.600000 20.315000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 18.040000 20.315000 18.360000 ;
      LAYER met4 ;
        RECT 19.995000 18.040000 20.315000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 14.960000 2.485000 15.280000 ;
      LAYER met4 ;
        RECT 2.165000 14.960000 2.485000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 15.400000 2.485000 15.720000 ;
      LAYER met4 ;
        RECT 2.165000 15.400000 2.485000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 15.840000 2.485000 16.160000 ;
      LAYER met4 ;
        RECT 2.165000 15.840000 2.485000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 16.280000 2.485000 16.600000 ;
      LAYER met4 ;
        RECT 2.165000 16.280000 2.485000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 16.720000 2.485000 17.040000 ;
      LAYER met4 ;
        RECT 2.165000 16.720000 2.485000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 17.160000 2.485000 17.480000 ;
      LAYER met4 ;
        RECT 2.165000 17.160000 2.485000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 17.600000 2.485000 17.920000 ;
      LAYER met4 ;
        RECT 2.165000 17.600000 2.485000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 18.040000 2.485000 18.360000 ;
      LAYER met4 ;
        RECT 2.165000 18.040000 2.485000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 14.960000 2.895000 15.280000 ;
      LAYER met4 ;
        RECT 2.575000 14.960000 2.895000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 15.400000 2.895000 15.720000 ;
      LAYER met4 ;
        RECT 2.575000 15.400000 2.895000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 15.840000 2.895000 16.160000 ;
      LAYER met4 ;
        RECT 2.575000 15.840000 2.895000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 16.280000 2.895000 16.600000 ;
      LAYER met4 ;
        RECT 2.575000 16.280000 2.895000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 16.720000 2.895000 17.040000 ;
      LAYER met4 ;
        RECT 2.575000 16.720000 2.895000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 17.160000 2.895000 17.480000 ;
      LAYER met4 ;
        RECT 2.575000 17.160000 2.895000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 17.600000 2.895000 17.920000 ;
      LAYER met4 ;
        RECT 2.575000 17.600000 2.895000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 18.040000 2.895000 18.360000 ;
      LAYER met4 ;
        RECT 2.575000 18.040000 2.895000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 14.960000 3.305000 15.280000 ;
      LAYER met4 ;
        RECT 2.985000 14.960000 3.305000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 15.400000 3.305000 15.720000 ;
      LAYER met4 ;
        RECT 2.985000 15.400000 3.305000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 15.840000 3.305000 16.160000 ;
      LAYER met4 ;
        RECT 2.985000 15.840000 3.305000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 16.280000 3.305000 16.600000 ;
      LAYER met4 ;
        RECT 2.985000 16.280000 3.305000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 16.720000 3.305000 17.040000 ;
      LAYER met4 ;
        RECT 2.985000 16.720000 3.305000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 17.160000 3.305000 17.480000 ;
      LAYER met4 ;
        RECT 2.985000 17.160000 3.305000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 17.600000 3.305000 17.920000 ;
      LAYER met4 ;
        RECT 2.985000 17.600000 3.305000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 18.040000 3.305000 18.360000 ;
      LAYER met4 ;
        RECT 2.985000 18.040000 3.305000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 14.960000 20.720000 15.280000 ;
      LAYER met4 ;
        RECT 20.400000 14.960000 20.720000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 15.400000 20.720000 15.720000 ;
      LAYER met4 ;
        RECT 20.400000 15.400000 20.720000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 15.840000 20.720000 16.160000 ;
      LAYER met4 ;
        RECT 20.400000 15.840000 20.720000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 16.280000 20.720000 16.600000 ;
      LAYER met4 ;
        RECT 20.400000 16.280000 20.720000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 16.720000 20.720000 17.040000 ;
      LAYER met4 ;
        RECT 20.400000 16.720000 20.720000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 17.160000 20.720000 17.480000 ;
      LAYER met4 ;
        RECT 20.400000 17.160000 20.720000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 17.600000 20.720000 17.920000 ;
      LAYER met4 ;
        RECT 20.400000 17.600000 20.720000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 18.040000 20.720000 18.360000 ;
      LAYER met4 ;
        RECT 20.400000 18.040000 20.720000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 14.960000 21.125000 15.280000 ;
      LAYER met4 ;
        RECT 20.805000 14.960000 21.125000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 15.400000 21.125000 15.720000 ;
      LAYER met4 ;
        RECT 20.805000 15.400000 21.125000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 15.840000 21.125000 16.160000 ;
      LAYER met4 ;
        RECT 20.805000 15.840000 21.125000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 16.280000 21.125000 16.600000 ;
      LAYER met4 ;
        RECT 20.805000 16.280000 21.125000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 16.720000 21.125000 17.040000 ;
      LAYER met4 ;
        RECT 20.805000 16.720000 21.125000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 17.160000 21.125000 17.480000 ;
      LAYER met4 ;
        RECT 20.805000 17.160000 21.125000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 17.600000 21.125000 17.920000 ;
      LAYER met4 ;
        RECT 20.805000 17.600000 21.125000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 18.040000 21.125000 18.360000 ;
      LAYER met4 ;
        RECT 20.805000 18.040000 21.125000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 14.960000 21.530000 15.280000 ;
      LAYER met4 ;
        RECT 21.210000 14.960000 21.530000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 15.400000 21.530000 15.720000 ;
      LAYER met4 ;
        RECT 21.210000 15.400000 21.530000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 15.840000 21.530000 16.160000 ;
      LAYER met4 ;
        RECT 21.210000 15.840000 21.530000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 16.280000 21.530000 16.600000 ;
      LAYER met4 ;
        RECT 21.210000 16.280000 21.530000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 16.720000 21.530000 17.040000 ;
      LAYER met4 ;
        RECT 21.210000 16.720000 21.530000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 17.160000 21.530000 17.480000 ;
      LAYER met4 ;
        RECT 21.210000 17.160000 21.530000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 17.600000 21.530000 17.920000 ;
      LAYER met4 ;
        RECT 21.210000 17.600000 21.530000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 18.040000 21.530000 18.360000 ;
      LAYER met4 ;
        RECT 21.210000 18.040000 21.530000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 14.960000 21.935000 15.280000 ;
      LAYER met4 ;
        RECT 21.615000 14.960000 21.935000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 15.400000 21.935000 15.720000 ;
      LAYER met4 ;
        RECT 21.615000 15.400000 21.935000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 15.840000 21.935000 16.160000 ;
      LAYER met4 ;
        RECT 21.615000 15.840000 21.935000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 16.280000 21.935000 16.600000 ;
      LAYER met4 ;
        RECT 21.615000 16.280000 21.935000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 16.720000 21.935000 17.040000 ;
      LAYER met4 ;
        RECT 21.615000 16.720000 21.935000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 17.160000 21.935000 17.480000 ;
      LAYER met4 ;
        RECT 21.615000 17.160000 21.935000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 17.600000 21.935000 17.920000 ;
      LAYER met4 ;
        RECT 21.615000 17.600000 21.935000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 18.040000 21.935000 18.360000 ;
      LAYER met4 ;
        RECT 21.615000 18.040000 21.935000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 14.960000 22.340000 15.280000 ;
      LAYER met4 ;
        RECT 22.020000 14.960000 22.340000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 15.400000 22.340000 15.720000 ;
      LAYER met4 ;
        RECT 22.020000 15.400000 22.340000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 15.840000 22.340000 16.160000 ;
      LAYER met4 ;
        RECT 22.020000 15.840000 22.340000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 16.280000 22.340000 16.600000 ;
      LAYER met4 ;
        RECT 22.020000 16.280000 22.340000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 16.720000 22.340000 17.040000 ;
      LAYER met4 ;
        RECT 22.020000 16.720000 22.340000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 17.160000 22.340000 17.480000 ;
      LAYER met4 ;
        RECT 22.020000 17.160000 22.340000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 17.600000 22.340000 17.920000 ;
      LAYER met4 ;
        RECT 22.020000 17.600000 22.340000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 18.040000 22.340000 18.360000 ;
      LAYER met4 ;
        RECT 22.020000 18.040000 22.340000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 14.960000 22.745000 15.280000 ;
      LAYER met4 ;
        RECT 22.425000 14.960000 22.745000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 15.400000 22.745000 15.720000 ;
      LAYER met4 ;
        RECT 22.425000 15.400000 22.745000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 15.840000 22.745000 16.160000 ;
      LAYER met4 ;
        RECT 22.425000 15.840000 22.745000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 16.280000 22.745000 16.600000 ;
      LAYER met4 ;
        RECT 22.425000 16.280000 22.745000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 16.720000 22.745000 17.040000 ;
      LAYER met4 ;
        RECT 22.425000 16.720000 22.745000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 17.160000 22.745000 17.480000 ;
      LAYER met4 ;
        RECT 22.425000 17.160000 22.745000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 17.600000 22.745000 17.920000 ;
      LAYER met4 ;
        RECT 22.425000 17.600000 22.745000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 18.040000 22.745000 18.360000 ;
      LAYER met4 ;
        RECT 22.425000 18.040000 22.745000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 14.960000 23.150000 15.280000 ;
      LAYER met4 ;
        RECT 22.830000 14.960000 23.150000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 15.400000 23.150000 15.720000 ;
      LAYER met4 ;
        RECT 22.830000 15.400000 23.150000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 15.840000 23.150000 16.160000 ;
      LAYER met4 ;
        RECT 22.830000 15.840000 23.150000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 16.280000 23.150000 16.600000 ;
      LAYER met4 ;
        RECT 22.830000 16.280000 23.150000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 16.720000 23.150000 17.040000 ;
      LAYER met4 ;
        RECT 22.830000 16.720000 23.150000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 17.160000 23.150000 17.480000 ;
      LAYER met4 ;
        RECT 22.830000 17.160000 23.150000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 17.600000 23.150000 17.920000 ;
      LAYER met4 ;
        RECT 22.830000 17.600000 23.150000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 18.040000 23.150000 18.360000 ;
      LAYER met4 ;
        RECT 22.830000 18.040000 23.150000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 14.960000 23.555000 15.280000 ;
      LAYER met4 ;
        RECT 23.235000 14.960000 23.555000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 15.400000 23.555000 15.720000 ;
      LAYER met4 ;
        RECT 23.235000 15.400000 23.555000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 15.840000 23.555000 16.160000 ;
      LAYER met4 ;
        RECT 23.235000 15.840000 23.555000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 16.280000 23.555000 16.600000 ;
      LAYER met4 ;
        RECT 23.235000 16.280000 23.555000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 16.720000 23.555000 17.040000 ;
      LAYER met4 ;
        RECT 23.235000 16.720000 23.555000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 17.160000 23.555000 17.480000 ;
      LAYER met4 ;
        RECT 23.235000 17.160000 23.555000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 17.600000 23.555000 17.920000 ;
      LAYER met4 ;
        RECT 23.235000 17.600000 23.555000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 18.040000 23.555000 18.360000 ;
      LAYER met4 ;
        RECT 23.235000 18.040000 23.555000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 14.960000 23.960000 15.280000 ;
      LAYER met4 ;
        RECT 23.640000 14.960000 23.960000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 15.400000 23.960000 15.720000 ;
      LAYER met4 ;
        RECT 23.640000 15.400000 23.960000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 15.840000 23.960000 16.160000 ;
      LAYER met4 ;
        RECT 23.640000 15.840000 23.960000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 16.280000 23.960000 16.600000 ;
      LAYER met4 ;
        RECT 23.640000 16.280000 23.960000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 16.720000 23.960000 17.040000 ;
      LAYER met4 ;
        RECT 23.640000 16.720000 23.960000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 17.160000 23.960000 17.480000 ;
      LAYER met4 ;
        RECT 23.640000 17.160000 23.960000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 17.600000 23.960000 17.920000 ;
      LAYER met4 ;
        RECT 23.640000 17.600000 23.960000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 18.040000 23.960000 18.360000 ;
      LAYER met4 ;
        RECT 23.640000 18.040000 23.960000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 14.960000 24.365000 15.280000 ;
      LAYER met4 ;
        RECT 24.045000 14.960000 24.365000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 15.400000 24.365000 15.720000 ;
      LAYER met4 ;
        RECT 24.045000 15.400000 24.365000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 15.840000 24.365000 16.160000 ;
      LAYER met4 ;
        RECT 24.045000 15.840000 24.365000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 16.280000 24.365000 16.600000 ;
      LAYER met4 ;
        RECT 24.045000 16.280000 24.365000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 16.720000 24.365000 17.040000 ;
      LAYER met4 ;
        RECT 24.045000 16.720000 24.365000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 17.160000 24.365000 17.480000 ;
      LAYER met4 ;
        RECT 24.045000 17.160000 24.365000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 17.600000 24.365000 17.920000 ;
      LAYER met4 ;
        RECT 24.045000 17.600000 24.365000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 18.040000 24.365000 18.360000 ;
      LAYER met4 ;
        RECT 24.045000 18.040000 24.365000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 14.960000 3.710000 15.280000 ;
      LAYER met4 ;
        RECT 3.390000 14.960000 3.710000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 15.400000 3.710000 15.720000 ;
      LAYER met4 ;
        RECT 3.390000 15.400000 3.710000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 15.840000 3.710000 16.160000 ;
      LAYER met4 ;
        RECT 3.390000 15.840000 3.710000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 16.280000 3.710000 16.600000 ;
      LAYER met4 ;
        RECT 3.390000 16.280000 3.710000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 16.720000 3.710000 17.040000 ;
      LAYER met4 ;
        RECT 3.390000 16.720000 3.710000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 17.160000 3.710000 17.480000 ;
      LAYER met4 ;
        RECT 3.390000 17.160000 3.710000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 17.600000 3.710000 17.920000 ;
      LAYER met4 ;
        RECT 3.390000 17.600000 3.710000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 18.040000 3.710000 18.360000 ;
      LAYER met4 ;
        RECT 3.390000 18.040000 3.710000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 14.960000 4.115000 15.280000 ;
      LAYER met4 ;
        RECT 3.795000 14.960000 4.115000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 15.400000 4.115000 15.720000 ;
      LAYER met4 ;
        RECT 3.795000 15.400000 4.115000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 15.840000 4.115000 16.160000 ;
      LAYER met4 ;
        RECT 3.795000 15.840000 4.115000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 16.280000 4.115000 16.600000 ;
      LAYER met4 ;
        RECT 3.795000 16.280000 4.115000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 16.720000 4.115000 17.040000 ;
      LAYER met4 ;
        RECT 3.795000 16.720000 4.115000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 17.160000 4.115000 17.480000 ;
      LAYER met4 ;
        RECT 3.795000 17.160000 4.115000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 17.600000 4.115000 17.920000 ;
      LAYER met4 ;
        RECT 3.795000 17.600000 4.115000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 18.040000 4.115000 18.360000 ;
      LAYER met4 ;
        RECT 3.795000 18.040000 4.115000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 14.960000 4.520000 15.280000 ;
      LAYER met4 ;
        RECT 4.200000 14.960000 4.520000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 15.400000 4.520000 15.720000 ;
      LAYER met4 ;
        RECT 4.200000 15.400000 4.520000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 15.840000 4.520000 16.160000 ;
      LAYER met4 ;
        RECT 4.200000 15.840000 4.520000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 16.280000 4.520000 16.600000 ;
      LAYER met4 ;
        RECT 4.200000 16.280000 4.520000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 16.720000 4.520000 17.040000 ;
      LAYER met4 ;
        RECT 4.200000 16.720000 4.520000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 17.160000 4.520000 17.480000 ;
      LAYER met4 ;
        RECT 4.200000 17.160000 4.520000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 17.600000 4.520000 17.920000 ;
      LAYER met4 ;
        RECT 4.200000 17.600000 4.520000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 18.040000 4.520000 18.360000 ;
      LAYER met4 ;
        RECT 4.200000 18.040000 4.520000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 14.960000 4.925000 15.280000 ;
      LAYER met4 ;
        RECT 4.605000 14.960000 4.925000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 15.400000 4.925000 15.720000 ;
      LAYER met4 ;
        RECT 4.605000 15.400000 4.925000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 15.840000 4.925000 16.160000 ;
      LAYER met4 ;
        RECT 4.605000 15.840000 4.925000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 16.280000 4.925000 16.600000 ;
      LAYER met4 ;
        RECT 4.605000 16.280000 4.925000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 16.720000 4.925000 17.040000 ;
      LAYER met4 ;
        RECT 4.605000 16.720000 4.925000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 17.160000 4.925000 17.480000 ;
      LAYER met4 ;
        RECT 4.605000 17.160000 4.925000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 17.600000 4.925000 17.920000 ;
      LAYER met4 ;
        RECT 4.605000 17.600000 4.925000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 18.040000 4.925000 18.360000 ;
      LAYER met4 ;
        RECT 4.605000 18.040000 4.925000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 14.960000 5.330000 15.280000 ;
      LAYER met4 ;
        RECT 5.010000 14.960000 5.330000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 15.400000 5.330000 15.720000 ;
      LAYER met4 ;
        RECT 5.010000 15.400000 5.330000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 15.840000 5.330000 16.160000 ;
      LAYER met4 ;
        RECT 5.010000 15.840000 5.330000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 16.280000 5.330000 16.600000 ;
      LAYER met4 ;
        RECT 5.010000 16.280000 5.330000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 16.720000 5.330000 17.040000 ;
      LAYER met4 ;
        RECT 5.010000 16.720000 5.330000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 17.160000 5.330000 17.480000 ;
      LAYER met4 ;
        RECT 5.010000 17.160000 5.330000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 17.600000 5.330000 17.920000 ;
      LAYER met4 ;
        RECT 5.010000 17.600000 5.330000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 18.040000 5.330000 18.360000 ;
      LAYER met4 ;
        RECT 5.010000 18.040000 5.330000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 14.960000 5.735000 15.280000 ;
      LAYER met4 ;
        RECT 5.415000 14.960000 5.735000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 15.400000 5.735000 15.720000 ;
      LAYER met4 ;
        RECT 5.415000 15.400000 5.735000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 15.840000 5.735000 16.160000 ;
      LAYER met4 ;
        RECT 5.415000 15.840000 5.735000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 16.280000 5.735000 16.600000 ;
      LAYER met4 ;
        RECT 5.415000 16.280000 5.735000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 16.720000 5.735000 17.040000 ;
      LAYER met4 ;
        RECT 5.415000 16.720000 5.735000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 17.160000 5.735000 17.480000 ;
      LAYER met4 ;
        RECT 5.415000 17.160000 5.735000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 17.600000 5.735000 17.920000 ;
      LAYER met4 ;
        RECT 5.415000 17.600000 5.735000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 18.040000 5.735000 18.360000 ;
      LAYER met4 ;
        RECT 5.415000 18.040000 5.735000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 14.960000 6.140000 15.280000 ;
      LAYER met4 ;
        RECT 5.820000 14.960000 6.140000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 15.400000 6.140000 15.720000 ;
      LAYER met4 ;
        RECT 5.820000 15.400000 6.140000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 15.840000 6.140000 16.160000 ;
      LAYER met4 ;
        RECT 5.820000 15.840000 6.140000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 16.280000 6.140000 16.600000 ;
      LAYER met4 ;
        RECT 5.820000 16.280000 6.140000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 16.720000 6.140000 17.040000 ;
      LAYER met4 ;
        RECT 5.820000 16.720000 6.140000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 17.160000 6.140000 17.480000 ;
      LAYER met4 ;
        RECT 5.820000 17.160000 6.140000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 17.600000 6.140000 17.920000 ;
      LAYER met4 ;
        RECT 5.820000 17.600000 6.140000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 18.040000 6.140000 18.360000 ;
      LAYER met4 ;
        RECT 5.820000 18.040000 6.140000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 14.960000 50.740000 15.280000 ;
      LAYER met4 ;
        RECT 50.420000 14.960000 50.740000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 15.400000 50.740000 15.720000 ;
      LAYER met4 ;
        RECT 50.420000 15.400000 50.740000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 15.840000 50.740000 16.160000 ;
      LAYER met4 ;
        RECT 50.420000 15.840000 50.740000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 16.280000 50.740000 16.600000 ;
      LAYER met4 ;
        RECT 50.420000 16.280000 50.740000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 16.720000 50.740000 17.040000 ;
      LAYER met4 ;
        RECT 50.420000 16.720000 50.740000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 17.160000 50.740000 17.480000 ;
      LAYER met4 ;
        RECT 50.420000 17.160000 50.740000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 17.600000 50.740000 17.920000 ;
      LAYER met4 ;
        RECT 50.420000 17.600000 50.740000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 18.040000 50.740000 18.360000 ;
      LAYER met4 ;
        RECT 50.420000 18.040000 50.740000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 14.960000 51.150000 15.280000 ;
      LAYER met4 ;
        RECT 50.830000 14.960000 51.150000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 15.400000 51.150000 15.720000 ;
      LAYER met4 ;
        RECT 50.830000 15.400000 51.150000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 15.840000 51.150000 16.160000 ;
      LAYER met4 ;
        RECT 50.830000 15.840000 51.150000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 16.280000 51.150000 16.600000 ;
      LAYER met4 ;
        RECT 50.830000 16.280000 51.150000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 16.720000 51.150000 17.040000 ;
      LAYER met4 ;
        RECT 50.830000 16.720000 51.150000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 17.160000 51.150000 17.480000 ;
      LAYER met4 ;
        RECT 50.830000 17.160000 51.150000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 17.600000 51.150000 17.920000 ;
      LAYER met4 ;
        RECT 50.830000 17.600000 51.150000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 18.040000 51.150000 18.360000 ;
      LAYER met4 ;
        RECT 50.830000 18.040000 51.150000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 14.960000 51.560000 15.280000 ;
      LAYER met4 ;
        RECT 51.240000 14.960000 51.560000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 15.400000 51.560000 15.720000 ;
      LAYER met4 ;
        RECT 51.240000 15.400000 51.560000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 15.840000 51.560000 16.160000 ;
      LAYER met4 ;
        RECT 51.240000 15.840000 51.560000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 16.280000 51.560000 16.600000 ;
      LAYER met4 ;
        RECT 51.240000 16.280000 51.560000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 16.720000 51.560000 17.040000 ;
      LAYER met4 ;
        RECT 51.240000 16.720000 51.560000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 17.160000 51.560000 17.480000 ;
      LAYER met4 ;
        RECT 51.240000 17.160000 51.560000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 17.600000 51.560000 17.920000 ;
      LAYER met4 ;
        RECT 51.240000 17.600000 51.560000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 18.040000 51.560000 18.360000 ;
      LAYER met4 ;
        RECT 51.240000 18.040000 51.560000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 14.960000 51.970000 15.280000 ;
      LAYER met4 ;
        RECT 51.650000 14.960000 51.970000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 15.400000 51.970000 15.720000 ;
      LAYER met4 ;
        RECT 51.650000 15.400000 51.970000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 15.840000 51.970000 16.160000 ;
      LAYER met4 ;
        RECT 51.650000 15.840000 51.970000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 16.280000 51.970000 16.600000 ;
      LAYER met4 ;
        RECT 51.650000 16.280000 51.970000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 16.720000 51.970000 17.040000 ;
      LAYER met4 ;
        RECT 51.650000 16.720000 51.970000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 17.160000 51.970000 17.480000 ;
      LAYER met4 ;
        RECT 51.650000 17.160000 51.970000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 17.600000 51.970000 17.920000 ;
      LAYER met4 ;
        RECT 51.650000 17.600000 51.970000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 18.040000 51.970000 18.360000 ;
      LAYER met4 ;
        RECT 51.650000 18.040000 51.970000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 14.960000 52.380000 15.280000 ;
      LAYER met4 ;
        RECT 52.060000 14.960000 52.380000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 15.400000 52.380000 15.720000 ;
      LAYER met4 ;
        RECT 52.060000 15.400000 52.380000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 15.840000 52.380000 16.160000 ;
      LAYER met4 ;
        RECT 52.060000 15.840000 52.380000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 16.280000 52.380000 16.600000 ;
      LAYER met4 ;
        RECT 52.060000 16.280000 52.380000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 16.720000 52.380000 17.040000 ;
      LAYER met4 ;
        RECT 52.060000 16.720000 52.380000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 17.160000 52.380000 17.480000 ;
      LAYER met4 ;
        RECT 52.060000 17.160000 52.380000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 17.600000 52.380000 17.920000 ;
      LAYER met4 ;
        RECT 52.060000 17.600000 52.380000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 18.040000 52.380000 18.360000 ;
      LAYER met4 ;
        RECT 52.060000 18.040000 52.380000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 14.960000 52.790000 15.280000 ;
      LAYER met4 ;
        RECT 52.470000 14.960000 52.790000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 15.400000 52.790000 15.720000 ;
      LAYER met4 ;
        RECT 52.470000 15.400000 52.790000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 15.840000 52.790000 16.160000 ;
      LAYER met4 ;
        RECT 52.470000 15.840000 52.790000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 16.280000 52.790000 16.600000 ;
      LAYER met4 ;
        RECT 52.470000 16.280000 52.790000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 16.720000 52.790000 17.040000 ;
      LAYER met4 ;
        RECT 52.470000 16.720000 52.790000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 17.160000 52.790000 17.480000 ;
      LAYER met4 ;
        RECT 52.470000 17.160000 52.790000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 17.600000 52.790000 17.920000 ;
      LAYER met4 ;
        RECT 52.470000 17.600000 52.790000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 18.040000 52.790000 18.360000 ;
      LAYER met4 ;
        RECT 52.470000 18.040000 52.790000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 14.960000 53.200000 15.280000 ;
      LAYER met4 ;
        RECT 52.880000 14.960000 53.200000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 15.400000 53.200000 15.720000 ;
      LAYER met4 ;
        RECT 52.880000 15.400000 53.200000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 15.840000 53.200000 16.160000 ;
      LAYER met4 ;
        RECT 52.880000 15.840000 53.200000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 16.280000 53.200000 16.600000 ;
      LAYER met4 ;
        RECT 52.880000 16.280000 53.200000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 16.720000 53.200000 17.040000 ;
      LAYER met4 ;
        RECT 52.880000 16.720000 53.200000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 17.160000 53.200000 17.480000 ;
      LAYER met4 ;
        RECT 52.880000 17.160000 53.200000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 17.600000 53.200000 17.920000 ;
      LAYER met4 ;
        RECT 52.880000 17.600000 53.200000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 18.040000 53.200000 18.360000 ;
      LAYER met4 ;
        RECT 52.880000 18.040000 53.200000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 14.960000 53.605000 15.280000 ;
      LAYER met4 ;
        RECT 53.285000 14.960000 53.605000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 15.400000 53.605000 15.720000 ;
      LAYER met4 ;
        RECT 53.285000 15.400000 53.605000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 15.840000 53.605000 16.160000 ;
      LAYER met4 ;
        RECT 53.285000 15.840000 53.605000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 16.280000 53.605000 16.600000 ;
      LAYER met4 ;
        RECT 53.285000 16.280000 53.605000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 16.720000 53.605000 17.040000 ;
      LAYER met4 ;
        RECT 53.285000 16.720000 53.605000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 17.160000 53.605000 17.480000 ;
      LAYER met4 ;
        RECT 53.285000 17.160000 53.605000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 17.600000 53.605000 17.920000 ;
      LAYER met4 ;
        RECT 53.285000 17.600000 53.605000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 18.040000 53.605000 18.360000 ;
      LAYER met4 ;
        RECT 53.285000 18.040000 53.605000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 14.960000 54.010000 15.280000 ;
      LAYER met4 ;
        RECT 53.690000 14.960000 54.010000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 15.400000 54.010000 15.720000 ;
      LAYER met4 ;
        RECT 53.690000 15.400000 54.010000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 15.840000 54.010000 16.160000 ;
      LAYER met4 ;
        RECT 53.690000 15.840000 54.010000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 16.280000 54.010000 16.600000 ;
      LAYER met4 ;
        RECT 53.690000 16.280000 54.010000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 16.720000 54.010000 17.040000 ;
      LAYER met4 ;
        RECT 53.690000 16.720000 54.010000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 17.160000 54.010000 17.480000 ;
      LAYER met4 ;
        RECT 53.690000 17.160000 54.010000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 17.600000 54.010000 17.920000 ;
      LAYER met4 ;
        RECT 53.690000 17.600000 54.010000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 18.040000 54.010000 18.360000 ;
      LAYER met4 ;
        RECT 53.690000 18.040000 54.010000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 14.960000 54.415000 15.280000 ;
      LAYER met4 ;
        RECT 54.095000 14.960000 54.415000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 15.400000 54.415000 15.720000 ;
      LAYER met4 ;
        RECT 54.095000 15.400000 54.415000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 15.840000 54.415000 16.160000 ;
      LAYER met4 ;
        RECT 54.095000 15.840000 54.415000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 16.280000 54.415000 16.600000 ;
      LAYER met4 ;
        RECT 54.095000 16.280000 54.415000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 16.720000 54.415000 17.040000 ;
      LAYER met4 ;
        RECT 54.095000 16.720000 54.415000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 17.160000 54.415000 17.480000 ;
      LAYER met4 ;
        RECT 54.095000 17.160000 54.415000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 17.600000 54.415000 17.920000 ;
      LAYER met4 ;
        RECT 54.095000 17.600000 54.415000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 18.040000 54.415000 18.360000 ;
      LAYER met4 ;
        RECT 54.095000 18.040000 54.415000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 14.960000 54.820000 15.280000 ;
      LAYER met4 ;
        RECT 54.500000 14.960000 54.820000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 15.400000 54.820000 15.720000 ;
      LAYER met4 ;
        RECT 54.500000 15.400000 54.820000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 15.840000 54.820000 16.160000 ;
      LAYER met4 ;
        RECT 54.500000 15.840000 54.820000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 16.280000 54.820000 16.600000 ;
      LAYER met4 ;
        RECT 54.500000 16.280000 54.820000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 16.720000 54.820000 17.040000 ;
      LAYER met4 ;
        RECT 54.500000 16.720000 54.820000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 17.160000 54.820000 17.480000 ;
      LAYER met4 ;
        RECT 54.500000 17.160000 54.820000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 17.600000 54.820000 17.920000 ;
      LAYER met4 ;
        RECT 54.500000 17.600000 54.820000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 18.040000 54.820000 18.360000 ;
      LAYER met4 ;
        RECT 54.500000 18.040000 54.820000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 14.960000 55.225000 15.280000 ;
      LAYER met4 ;
        RECT 54.905000 14.960000 55.225000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 15.400000 55.225000 15.720000 ;
      LAYER met4 ;
        RECT 54.905000 15.400000 55.225000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 15.840000 55.225000 16.160000 ;
      LAYER met4 ;
        RECT 54.905000 15.840000 55.225000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 16.280000 55.225000 16.600000 ;
      LAYER met4 ;
        RECT 54.905000 16.280000 55.225000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 16.720000 55.225000 17.040000 ;
      LAYER met4 ;
        RECT 54.905000 16.720000 55.225000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 17.160000 55.225000 17.480000 ;
      LAYER met4 ;
        RECT 54.905000 17.160000 55.225000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 17.600000 55.225000 17.920000 ;
      LAYER met4 ;
        RECT 54.905000 17.600000 55.225000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 18.040000 55.225000 18.360000 ;
      LAYER met4 ;
        RECT 54.905000 18.040000 55.225000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 14.960000 55.630000 15.280000 ;
      LAYER met4 ;
        RECT 55.310000 14.960000 55.630000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 15.400000 55.630000 15.720000 ;
      LAYER met4 ;
        RECT 55.310000 15.400000 55.630000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 15.840000 55.630000 16.160000 ;
      LAYER met4 ;
        RECT 55.310000 15.840000 55.630000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 16.280000 55.630000 16.600000 ;
      LAYER met4 ;
        RECT 55.310000 16.280000 55.630000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 16.720000 55.630000 17.040000 ;
      LAYER met4 ;
        RECT 55.310000 16.720000 55.630000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 17.160000 55.630000 17.480000 ;
      LAYER met4 ;
        RECT 55.310000 17.160000 55.630000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 17.600000 55.630000 17.920000 ;
      LAYER met4 ;
        RECT 55.310000 17.600000 55.630000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 18.040000 55.630000 18.360000 ;
      LAYER met4 ;
        RECT 55.310000 18.040000 55.630000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 14.960000 56.035000 15.280000 ;
      LAYER met4 ;
        RECT 55.715000 14.960000 56.035000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 15.400000 56.035000 15.720000 ;
      LAYER met4 ;
        RECT 55.715000 15.400000 56.035000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 15.840000 56.035000 16.160000 ;
      LAYER met4 ;
        RECT 55.715000 15.840000 56.035000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 16.280000 56.035000 16.600000 ;
      LAYER met4 ;
        RECT 55.715000 16.280000 56.035000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 16.720000 56.035000 17.040000 ;
      LAYER met4 ;
        RECT 55.715000 16.720000 56.035000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 17.160000 56.035000 17.480000 ;
      LAYER met4 ;
        RECT 55.715000 17.160000 56.035000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 17.600000 56.035000 17.920000 ;
      LAYER met4 ;
        RECT 55.715000 17.600000 56.035000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 18.040000 56.035000 18.360000 ;
      LAYER met4 ;
        RECT 55.715000 18.040000 56.035000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 14.960000 56.440000 15.280000 ;
      LAYER met4 ;
        RECT 56.120000 14.960000 56.440000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 15.400000 56.440000 15.720000 ;
      LAYER met4 ;
        RECT 56.120000 15.400000 56.440000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 15.840000 56.440000 16.160000 ;
      LAYER met4 ;
        RECT 56.120000 15.840000 56.440000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 16.280000 56.440000 16.600000 ;
      LAYER met4 ;
        RECT 56.120000 16.280000 56.440000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 16.720000 56.440000 17.040000 ;
      LAYER met4 ;
        RECT 56.120000 16.720000 56.440000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 17.160000 56.440000 17.480000 ;
      LAYER met4 ;
        RECT 56.120000 17.160000 56.440000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 17.600000 56.440000 17.920000 ;
      LAYER met4 ;
        RECT 56.120000 17.600000 56.440000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 18.040000 56.440000 18.360000 ;
      LAYER met4 ;
        RECT 56.120000 18.040000 56.440000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 14.960000 56.845000 15.280000 ;
      LAYER met4 ;
        RECT 56.525000 14.960000 56.845000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 15.400000 56.845000 15.720000 ;
      LAYER met4 ;
        RECT 56.525000 15.400000 56.845000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 15.840000 56.845000 16.160000 ;
      LAYER met4 ;
        RECT 56.525000 15.840000 56.845000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 16.280000 56.845000 16.600000 ;
      LAYER met4 ;
        RECT 56.525000 16.280000 56.845000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 16.720000 56.845000 17.040000 ;
      LAYER met4 ;
        RECT 56.525000 16.720000 56.845000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 17.160000 56.845000 17.480000 ;
      LAYER met4 ;
        RECT 56.525000 17.160000 56.845000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 17.600000 56.845000 17.920000 ;
      LAYER met4 ;
        RECT 56.525000 17.600000 56.845000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 18.040000 56.845000 18.360000 ;
      LAYER met4 ;
        RECT 56.525000 18.040000 56.845000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 14.960000 57.250000 15.280000 ;
      LAYER met4 ;
        RECT 56.930000 14.960000 57.250000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 15.400000 57.250000 15.720000 ;
      LAYER met4 ;
        RECT 56.930000 15.400000 57.250000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 15.840000 57.250000 16.160000 ;
      LAYER met4 ;
        RECT 56.930000 15.840000 57.250000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 16.280000 57.250000 16.600000 ;
      LAYER met4 ;
        RECT 56.930000 16.280000 57.250000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 16.720000 57.250000 17.040000 ;
      LAYER met4 ;
        RECT 56.930000 16.720000 57.250000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 17.160000 57.250000 17.480000 ;
      LAYER met4 ;
        RECT 56.930000 17.160000 57.250000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 17.600000 57.250000 17.920000 ;
      LAYER met4 ;
        RECT 56.930000 17.600000 57.250000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 18.040000 57.250000 18.360000 ;
      LAYER met4 ;
        RECT 56.930000 18.040000 57.250000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 14.960000 57.655000 15.280000 ;
      LAYER met4 ;
        RECT 57.335000 14.960000 57.655000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 15.400000 57.655000 15.720000 ;
      LAYER met4 ;
        RECT 57.335000 15.400000 57.655000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 15.840000 57.655000 16.160000 ;
      LAYER met4 ;
        RECT 57.335000 15.840000 57.655000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 16.280000 57.655000 16.600000 ;
      LAYER met4 ;
        RECT 57.335000 16.280000 57.655000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 16.720000 57.655000 17.040000 ;
      LAYER met4 ;
        RECT 57.335000 16.720000 57.655000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 17.160000 57.655000 17.480000 ;
      LAYER met4 ;
        RECT 57.335000 17.160000 57.655000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 17.600000 57.655000 17.920000 ;
      LAYER met4 ;
        RECT 57.335000 17.600000 57.655000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 18.040000 57.655000 18.360000 ;
      LAYER met4 ;
        RECT 57.335000 18.040000 57.655000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 14.960000 58.060000 15.280000 ;
      LAYER met4 ;
        RECT 57.740000 14.960000 58.060000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 15.400000 58.060000 15.720000 ;
      LAYER met4 ;
        RECT 57.740000 15.400000 58.060000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 15.840000 58.060000 16.160000 ;
      LAYER met4 ;
        RECT 57.740000 15.840000 58.060000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 16.280000 58.060000 16.600000 ;
      LAYER met4 ;
        RECT 57.740000 16.280000 58.060000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 16.720000 58.060000 17.040000 ;
      LAYER met4 ;
        RECT 57.740000 16.720000 58.060000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 17.160000 58.060000 17.480000 ;
      LAYER met4 ;
        RECT 57.740000 17.160000 58.060000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 17.600000 58.060000 17.920000 ;
      LAYER met4 ;
        RECT 57.740000 17.600000 58.060000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 18.040000 58.060000 18.360000 ;
      LAYER met4 ;
        RECT 57.740000 18.040000 58.060000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 14.960000 58.465000 15.280000 ;
      LAYER met4 ;
        RECT 58.145000 14.960000 58.465000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 15.400000 58.465000 15.720000 ;
      LAYER met4 ;
        RECT 58.145000 15.400000 58.465000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 15.840000 58.465000 16.160000 ;
      LAYER met4 ;
        RECT 58.145000 15.840000 58.465000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 16.280000 58.465000 16.600000 ;
      LAYER met4 ;
        RECT 58.145000 16.280000 58.465000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 16.720000 58.465000 17.040000 ;
      LAYER met4 ;
        RECT 58.145000 16.720000 58.465000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 17.160000 58.465000 17.480000 ;
      LAYER met4 ;
        RECT 58.145000 17.160000 58.465000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 17.600000 58.465000 17.920000 ;
      LAYER met4 ;
        RECT 58.145000 17.600000 58.465000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 18.040000 58.465000 18.360000 ;
      LAYER met4 ;
        RECT 58.145000 18.040000 58.465000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 14.960000 58.870000 15.280000 ;
      LAYER met4 ;
        RECT 58.550000 14.960000 58.870000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 15.400000 58.870000 15.720000 ;
      LAYER met4 ;
        RECT 58.550000 15.400000 58.870000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 15.840000 58.870000 16.160000 ;
      LAYER met4 ;
        RECT 58.550000 15.840000 58.870000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 16.280000 58.870000 16.600000 ;
      LAYER met4 ;
        RECT 58.550000 16.280000 58.870000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 16.720000 58.870000 17.040000 ;
      LAYER met4 ;
        RECT 58.550000 16.720000 58.870000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 17.160000 58.870000 17.480000 ;
      LAYER met4 ;
        RECT 58.550000 17.160000 58.870000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 17.600000 58.870000 17.920000 ;
      LAYER met4 ;
        RECT 58.550000 17.600000 58.870000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 18.040000 58.870000 18.360000 ;
      LAYER met4 ;
        RECT 58.550000 18.040000 58.870000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 14.960000 59.275000 15.280000 ;
      LAYER met4 ;
        RECT 58.955000 14.960000 59.275000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 15.400000 59.275000 15.720000 ;
      LAYER met4 ;
        RECT 58.955000 15.400000 59.275000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 15.840000 59.275000 16.160000 ;
      LAYER met4 ;
        RECT 58.955000 15.840000 59.275000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 16.280000 59.275000 16.600000 ;
      LAYER met4 ;
        RECT 58.955000 16.280000 59.275000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 16.720000 59.275000 17.040000 ;
      LAYER met4 ;
        RECT 58.955000 16.720000 59.275000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 17.160000 59.275000 17.480000 ;
      LAYER met4 ;
        RECT 58.955000 17.160000 59.275000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 17.600000 59.275000 17.920000 ;
      LAYER met4 ;
        RECT 58.955000 17.600000 59.275000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 18.040000 59.275000 18.360000 ;
      LAYER met4 ;
        RECT 58.955000 18.040000 59.275000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 14.960000 59.680000 15.280000 ;
      LAYER met4 ;
        RECT 59.360000 14.960000 59.680000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 15.400000 59.680000 15.720000 ;
      LAYER met4 ;
        RECT 59.360000 15.400000 59.680000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 15.840000 59.680000 16.160000 ;
      LAYER met4 ;
        RECT 59.360000 15.840000 59.680000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 16.280000 59.680000 16.600000 ;
      LAYER met4 ;
        RECT 59.360000 16.280000 59.680000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 16.720000 59.680000 17.040000 ;
      LAYER met4 ;
        RECT 59.360000 16.720000 59.680000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 17.160000 59.680000 17.480000 ;
      LAYER met4 ;
        RECT 59.360000 17.160000 59.680000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 17.600000 59.680000 17.920000 ;
      LAYER met4 ;
        RECT 59.360000 17.600000 59.680000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 18.040000 59.680000 18.360000 ;
      LAYER met4 ;
        RECT 59.360000 18.040000 59.680000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 14.960000 60.085000 15.280000 ;
      LAYER met4 ;
        RECT 59.765000 14.960000 60.085000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 15.400000 60.085000 15.720000 ;
      LAYER met4 ;
        RECT 59.765000 15.400000 60.085000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 15.840000 60.085000 16.160000 ;
      LAYER met4 ;
        RECT 59.765000 15.840000 60.085000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 16.280000 60.085000 16.600000 ;
      LAYER met4 ;
        RECT 59.765000 16.280000 60.085000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 16.720000 60.085000 17.040000 ;
      LAYER met4 ;
        RECT 59.765000 16.720000 60.085000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 17.160000 60.085000 17.480000 ;
      LAYER met4 ;
        RECT 59.765000 17.160000 60.085000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 17.600000 60.085000 17.920000 ;
      LAYER met4 ;
        RECT 59.765000 17.600000 60.085000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 18.040000 60.085000 18.360000 ;
      LAYER met4 ;
        RECT 59.765000 18.040000 60.085000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 14.960000 6.545000 15.280000 ;
      LAYER met4 ;
        RECT 6.225000 14.960000 6.545000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 15.400000 6.545000 15.720000 ;
      LAYER met4 ;
        RECT 6.225000 15.400000 6.545000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 15.840000 6.545000 16.160000 ;
      LAYER met4 ;
        RECT 6.225000 15.840000 6.545000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 16.280000 6.545000 16.600000 ;
      LAYER met4 ;
        RECT 6.225000 16.280000 6.545000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 16.720000 6.545000 17.040000 ;
      LAYER met4 ;
        RECT 6.225000 16.720000 6.545000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 17.160000 6.545000 17.480000 ;
      LAYER met4 ;
        RECT 6.225000 17.160000 6.545000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 17.600000 6.545000 17.920000 ;
      LAYER met4 ;
        RECT 6.225000 17.600000 6.545000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 18.040000 6.545000 18.360000 ;
      LAYER met4 ;
        RECT 6.225000 18.040000 6.545000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 14.960000 6.950000 15.280000 ;
      LAYER met4 ;
        RECT 6.630000 14.960000 6.950000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 15.400000 6.950000 15.720000 ;
      LAYER met4 ;
        RECT 6.630000 15.400000 6.950000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 15.840000 6.950000 16.160000 ;
      LAYER met4 ;
        RECT 6.630000 15.840000 6.950000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 16.280000 6.950000 16.600000 ;
      LAYER met4 ;
        RECT 6.630000 16.280000 6.950000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 16.720000 6.950000 17.040000 ;
      LAYER met4 ;
        RECT 6.630000 16.720000 6.950000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 17.160000 6.950000 17.480000 ;
      LAYER met4 ;
        RECT 6.630000 17.160000 6.950000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 17.600000 6.950000 17.920000 ;
      LAYER met4 ;
        RECT 6.630000 17.600000 6.950000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 18.040000 6.950000 18.360000 ;
      LAYER met4 ;
        RECT 6.630000 18.040000 6.950000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 14.960000 60.490000 15.280000 ;
      LAYER met4 ;
        RECT 60.170000 14.960000 60.490000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 15.400000 60.490000 15.720000 ;
      LAYER met4 ;
        RECT 60.170000 15.400000 60.490000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 15.840000 60.490000 16.160000 ;
      LAYER met4 ;
        RECT 60.170000 15.840000 60.490000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 16.280000 60.490000 16.600000 ;
      LAYER met4 ;
        RECT 60.170000 16.280000 60.490000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 16.720000 60.490000 17.040000 ;
      LAYER met4 ;
        RECT 60.170000 16.720000 60.490000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 17.160000 60.490000 17.480000 ;
      LAYER met4 ;
        RECT 60.170000 17.160000 60.490000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 17.600000 60.490000 17.920000 ;
      LAYER met4 ;
        RECT 60.170000 17.600000 60.490000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 18.040000 60.490000 18.360000 ;
      LAYER met4 ;
        RECT 60.170000 18.040000 60.490000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 14.960000 60.895000 15.280000 ;
      LAYER met4 ;
        RECT 60.575000 14.960000 60.895000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 15.400000 60.895000 15.720000 ;
      LAYER met4 ;
        RECT 60.575000 15.400000 60.895000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 15.840000 60.895000 16.160000 ;
      LAYER met4 ;
        RECT 60.575000 15.840000 60.895000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 16.280000 60.895000 16.600000 ;
      LAYER met4 ;
        RECT 60.575000 16.280000 60.895000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 16.720000 60.895000 17.040000 ;
      LAYER met4 ;
        RECT 60.575000 16.720000 60.895000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 17.160000 60.895000 17.480000 ;
      LAYER met4 ;
        RECT 60.575000 17.160000 60.895000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 17.600000 60.895000 17.920000 ;
      LAYER met4 ;
        RECT 60.575000 17.600000 60.895000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 18.040000 60.895000 18.360000 ;
      LAYER met4 ;
        RECT 60.575000 18.040000 60.895000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 14.960000 61.300000 15.280000 ;
      LAYER met4 ;
        RECT 60.980000 14.960000 61.300000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 15.400000 61.300000 15.720000 ;
      LAYER met4 ;
        RECT 60.980000 15.400000 61.300000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 15.840000 61.300000 16.160000 ;
      LAYER met4 ;
        RECT 60.980000 15.840000 61.300000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 16.280000 61.300000 16.600000 ;
      LAYER met4 ;
        RECT 60.980000 16.280000 61.300000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 16.720000 61.300000 17.040000 ;
      LAYER met4 ;
        RECT 60.980000 16.720000 61.300000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 17.160000 61.300000 17.480000 ;
      LAYER met4 ;
        RECT 60.980000 17.160000 61.300000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 17.600000 61.300000 17.920000 ;
      LAYER met4 ;
        RECT 60.980000 17.600000 61.300000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 18.040000 61.300000 18.360000 ;
      LAYER met4 ;
        RECT 60.980000 18.040000 61.300000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 14.960000 61.705000 15.280000 ;
      LAYER met4 ;
        RECT 61.385000 14.960000 61.705000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 15.400000 61.705000 15.720000 ;
      LAYER met4 ;
        RECT 61.385000 15.400000 61.705000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 15.840000 61.705000 16.160000 ;
      LAYER met4 ;
        RECT 61.385000 15.840000 61.705000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 16.280000 61.705000 16.600000 ;
      LAYER met4 ;
        RECT 61.385000 16.280000 61.705000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 16.720000 61.705000 17.040000 ;
      LAYER met4 ;
        RECT 61.385000 16.720000 61.705000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 17.160000 61.705000 17.480000 ;
      LAYER met4 ;
        RECT 61.385000 17.160000 61.705000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 17.600000 61.705000 17.920000 ;
      LAYER met4 ;
        RECT 61.385000 17.600000 61.705000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 18.040000 61.705000 18.360000 ;
      LAYER met4 ;
        RECT 61.385000 18.040000 61.705000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 14.960000 62.110000 15.280000 ;
      LAYER met4 ;
        RECT 61.790000 14.960000 62.110000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 15.400000 62.110000 15.720000 ;
      LAYER met4 ;
        RECT 61.790000 15.400000 62.110000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 15.840000 62.110000 16.160000 ;
      LAYER met4 ;
        RECT 61.790000 15.840000 62.110000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 16.280000 62.110000 16.600000 ;
      LAYER met4 ;
        RECT 61.790000 16.280000 62.110000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 16.720000 62.110000 17.040000 ;
      LAYER met4 ;
        RECT 61.790000 16.720000 62.110000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 17.160000 62.110000 17.480000 ;
      LAYER met4 ;
        RECT 61.790000 17.160000 62.110000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 17.600000 62.110000 17.920000 ;
      LAYER met4 ;
        RECT 61.790000 17.600000 62.110000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 18.040000 62.110000 18.360000 ;
      LAYER met4 ;
        RECT 61.790000 18.040000 62.110000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 14.960000 62.515000 15.280000 ;
      LAYER met4 ;
        RECT 62.195000 14.960000 62.515000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 15.400000 62.515000 15.720000 ;
      LAYER met4 ;
        RECT 62.195000 15.400000 62.515000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 15.840000 62.515000 16.160000 ;
      LAYER met4 ;
        RECT 62.195000 15.840000 62.515000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 16.280000 62.515000 16.600000 ;
      LAYER met4 ;
        RECT 62.195000 16.280000 62.515000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 16.720000 62.515000 17.040000 ;
      LAYER met4 ;
        RECT 62.195000 16.720000 62.515000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 17.160000 62.515000 17.480000 ;
      LAYER met4 ;
        RECT 62.195000 17.160000 62.515000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 17.600000 62.515000 17.920000 ;
      LAYER met4 ;
        RECT 62.195000 17.600000 62.515000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 18.040000 62.515000 18.360000 ;
      LAYER met4 ;
        RECT 62.195000 18.040000 62.515000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 14.960000 62.920000 15.280000 ;
      LAYER met4 ;
        RECT 62.600000 14.960000 62.920000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 15.400000 62.920000 15.720000 ;
      LAYER met4 ;
        RECT 62.600000 15.400000 62.920000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 15.840000 62.920000 16.160000 ;
      LAYER met4 ;
        RECT 62.600000 15.840000 62.920000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 16.280000 62.920000 16.600000 ;
      LAYER met4 ;
        RECT 62.600000 16.280000 62.920000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 16.720000 62.920000 17.040000 ;
      LAYER met4 ;
        RECT 62.600000 16.720000 62.920000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 17.160000 62.920000 17.480000 ;
      LAYER met4 ;
        RECT 62.600000 17.160000 62.920000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 17.600000 62.920000 17.920000 ;
      LAYER met4 ;
        RECT 62.600000 17.600000 62.920000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 18.040000 62.920000 18.360000 ;
      LAYER met4 ;
        RECT 62.600000 18.040000 62.920000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 14.960000 63.325000 15.280000 ;
      LAYER met4 ;
        RECT 63.005000 14.960000 63.325000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 15.400000 63.325000 15.720000 ;
      LAYER met4 ;
        RECT 63.005000 15.400000 63.325000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 15.840000 63.325000 16.160000 ;
      LAYER met4 ;
        RECT 63.005000 15.840000 63.325000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 16.280000 63.325000 16.600000 ;
      LAYER met4 ;
        RECT 63.005000 16.280000 63.325000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 16.720000 63.325000 17.040000 ;
      LAYER met4 ;
        RECT 63.005000 16.720000 63.325000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 17.160000 63.325000 17.480000 ;
      LAYER met4 ;
        RECT 63.005000 17.160000 63.325000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 17.600000 63.325000 17.920000 ;
      LAYER met4 ;
        RECT 63.005000 17.600000 63.325000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 18.040000 63.325000 18.360000 ;
      LAYER met4 ;
        RECT 63.005000 18.040000 63.325000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 14.960000 63.730000 15.280000 ;
      LAYER met4 ;
        RECT 63.410000 14.960000 63.730000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 15.400000 63.730000 15.720000 ;
      LAYER met4 ;
        RECT 63.410000 15.400000 63.730000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 15.840000 63.730000 16.160000 ;
      LAYER met4 ;
        RECT 63.410000 15.840000 63.730000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 16.280000 63.730000 16.600000 ;
      LAYER met4 ;
        RECT 63.410000 16.280000 63.730000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 16.720000 63.730000 17.040000 ;
      LAYER met4 ;
        RECT 63.410000 16.720000 63.730000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 17.160000 63.730000 17.480000 ;
      LAYER met4 ;
        RECT 63.410000 17.160000 63.730000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 17.600000 63.730000 17.920000 ;
      LAYER met4 ;
        RECT 63.410000 17.600000 63.730000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 18.040000 63.730000 18.360000 ;
      LAYER met4 ;
        RECT 63.410000 18.040000 63.730000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 14.960000 64.135000 15.280000 ;
      LAYER met4 ;
        RECT 63.815000 14.960000 64.135000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 15.400000 64.135000 15.720000 ;
      LAYER met4 ;
        RECT 63.815000 15.400000 64.135000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 15.840000 64.135000 16.160000 ;
      LAYER met4 ;
        RECT 63.815000 15.840000 64.135000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 16.280000 64.135000 16.600000 ;
      LAYER met4 ;
        RECT 63.815000 16.280000 64.135000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 16.720000 64.135000 17.040000 ;
      LAYER met4 ;
        RECT 63.815000 16.720000 64.135000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 17.160000 64.135000 17.480000 ;
      LAYER met4 ;
        RECT 63.815000 17.160000 64.135000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 17.600000 64.135000 17.920000 ;
      LAYER met4 ;
        RECT 63.815000 17.600000 64.135000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 18.040000 64.135000 18.360000 ;
      LAYER met4 ;
        RECT 63.815000 18.040000 64.135000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 14.960000 64.540000 15.280000 ;
      LAYER met4 ;
        RECT 64.220000 14.960000 64.540000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 15.400000 64.540000 15.720000 ;
      LAYER met4 ;
        RECT 64.220000 15.400000 64.540000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 15.840000 64.540000 16.160000 ;
      LAYER met4 ;
        RECT 64.220000 15.840000 64.540000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 16.280000 64.540000 16.600000 ;
      LAYER met4 ;
        RECT 64.220000 16.280000 64.540000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 16.720000 64.540000 17.040000 ;
      LAYER met4 ;
        RECT 64.220000 16.720000 64.540000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 17.160000 64.540000 17.480000 ;
      LAYER met4 ;
        RECT 64.220000 17.160000 64.540000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 17.600000 64.540000 17.920000 ;
      LAYER met4 ;
        RECT 64.220000 17.600000 64.540000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 18.040000 64.540000 18.360000 ;
      LAYER met4 ;
        RECT 64.220000 18.040000 64.540000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 14.960000 64.945000 15.280000 ;
      LAYER met4 ;
        RECT 64.625000 14.960000 64.945000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 15.400000 64.945000 15.720000 ;
      LAYER met4 ;
        RECT 64.625000 15.400000 64.945000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 15.840000 64.945000 16.160000 ;
      LAYER met4 ;
        RECT 64.625000 15.840000 64.945000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 16.280000 64.945000 16.600000 ;
      LAYER met4 ;
        RECT 64.625000 16.280000 64.945000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 16.720000 64.945000 17.040000 ;
      LAYER met4 ;
        RECT 64.625000 16.720000 64.945000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 17.160000 64.945000 17.480000 ;
      LAYER met4 ;
        RECT 64.625000 17.160000 64.945000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 17.600000 64.945000 17.920000 ;
      LAYER met4 ;
        RECT 64.625000 17.600000 64.945000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 18.040000 64.945000 18.360000 ;
      LAYER met4 ;
        RECT 64.625000 18.040000 64.945000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 14.960000 65.350000 15.280000 ;
      LAYER met4 ;
        RECT 65.030000 14.960000 65.350000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 15.400000 65.350000 15.720000 ;
      LAYER met4 ;
        RECT 65.030000 15.400000 65.350000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 15.840000 65.350000 16.160000 ;
      LAYER met4 ;
        RECT 65.030000 15.840000 65.350000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 16.280000 65.350000 16.600000 ;
      LAYER met4 ;
        RECT 65.030000 16.280000 65.350000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 16.720000 65.350000 17.040000 ;
      LAYER met4 ;
        RECT 65.030000 16.720000 65.350000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 17.160000 65.350000 17.480000 ;
      LAYER met4 ;
        RECT 65.030000 17.160000 65.350000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 17.600000 65.350000 17.920000 ;
      LAYER met4 ;
        RECT 65.030000 17.600000 65.350000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 18.040000 65.350000 18.360000 ;
      LAYER met4 ;
        RECT 65.030000 18.040000 65.350000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 14.960000 65.755000 15.280000 ;
      LAYER met4 ;
        RECT 65.435000 14.960000 65.755000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 15.400000 65.755000 15.720000 ;
      LAYER met4 ;
        RECT 65.435000 15.400000 65.755000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 15.840000 65.755000 16.160000 ;
      LAYER met4 ;
        RECT 65.435000 15.840000 65.755000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 16.280000 65.755000 16.600000 ;
      LAYER met4 ;
        RECT 65.435000 16.280000 65.755000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 16.720000 65.755000 17.040000 ;
      LAYER met4 ;
        RECT 65.435000 16.720000 65.755000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 17.160000 65.755000 17.480000 ;
      LAYER met4 ;
        RECT 65.435000 17.160000 65.755000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 17.600000 65.755000 17.920000 ;
      LAYER met4 ;
        RECT 65.435000 17.600000 65.755000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 18.040000 65.755000 18.360000 ;
      LAYER met4 ;
        RECT 65.435000 18.040000 65.755000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 14.960000 66.160000 15.280000 ;
      LAYER met4 ;
        RECT 65.840000 14.960000 66.160000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 15.400000 66.160000 15.720000 ;
      LAYER met4 ;
        RECT 65.840000 15.400000 66.160000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 15.840000 66.160000 16.160000 ;
      LAYER met4 ;
        RECT 65.840000 15.840000 66.160000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 16.280000 66.160000 16.600000 ;
      LAYER met4 ;
        RECT 65.840000 16.280000 66.160000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 16.720000 66.160000 17.040000 ;
      LAYER met4 ;
        RECT 65.840000 16.720000 66.160000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 17.160000 66.160000 17.480000 ;
      LAYER met4 ;
        RECT 65.840000 17.160000 66.160000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 17.600000 66.160000 17.920000 ;
      LAYER met4 ;
        RECT 65.840000 17.600000 66.160000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 18.040000 66.160000 18.360000 ;
      LAYER met4 ;
        RECT 65.840000 18.040000 66.160000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 14.960000 66.565000 15.280000 ;
      LAYER met4 ;
        RECT 66.245000 14.960000 66.565000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 15.400000 66.565000 15.720000 ;
      LAYER met4 ;
        RECT 66.245000 15.400000 66.565000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 15.840000 66.565000 16.160000 ;
      LAYER met4 ;
        RECT 66.245000 15.840000 66.565000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 16.280000 66.565000 16.600000 ;
      LAYER met4 ;
        RECT 66.245000 16.280000 66.565000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 16.720000 66.565000 17.040000 ;
      LAYER met4 ;
        RECT 66.245000 16.720000 66.565000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 17.160000 66.565000 17.480000 ;
      LAYER met4 ;
        RECT 66.245000 17.160000 66.565000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 17.600000 66.565000 17.920000 ;
      LAYER met4 ;
        RECT 66.245000 17.600000 66.565000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 18.040000 66.565000 18.360000 ;
      LAYER met4 ;
        RECT 66.245000 18.040000 66.565000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 14.960000 66.970000 15.280000 ;
      LAYER met4 ;
        RECT 66.650000 14.960000 66.970000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 15.400000 66.970000 15.720000 ;
      LAYER met4 ;
        RECT 66.650000 15.400000 66.970000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 15.840000 66.970000 16.160000 ;
      LAYER met4 ;
        RECT 66.650000 15.840000 66.970000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 16.280000 66.970000 16.600000 ;
      LAYER met4 ;
        RECT 66.650000 16.280000 66.970000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 16.720000 66.970000 17.040000 ;
      LAYER met4 ;
        RECT 66.650000 16.720000 66.970000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 17.160000 66.970000 17.480000 ;
      LAYER met4 ;
        RECT 66.650000 17.160000 66.970000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 17.600000 66.970000 17.920000 ;
      LAYER met4 ;
        RECT 66.650000 17.600000 66.970000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 18.040000 66.970000 18.360000 ;
      LAYER met4 ;
        RECT 66.650000 18.040000 66.970000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 14.960000 67.375000 15.280000 ;
      LAYER met4 ;
        RECT 67.055000 14.960000 67.375000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 15.400000 67.375000 15.720000 ;
      LAYER met4 ;
        RECT 67.055000 15.400000 67.375000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 15.840000 67.375000 16.160000 ;
      LAYER met4 ;
        RECT 67.055000 15.840000 67.375000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 16.280000 67.375000 16.600000 ;
      LAYER met4 ;
        RECT 67.055000 16.280000 67.375000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 16.720000 67.375000 17.040000 ;
      LAYER met4 ;
        RECT 67.055000 16.720000 67.375000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 17.160000 67.375000 17.480000 ;
      LAYER met4 ;
        RECT 67.055000 17.160000 67.375000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 17.600000 67.375000 17.920000 ;
      LAYER met4 ;
        RECT 67.055000 17.600000 67.375000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 18.040000 67.375000 18.360000 ;
      LAYER met4 ;
        RECT 67.055000 18.040000 67.375000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 14.960000 67.780000 15.280000 ;
      LAYER met4 ;
        RECT 67.460000 14.960000 67.780000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 15.400000 67.780000 15.720000 ;
      LAYER met4 ;
        RECT 67.460000 15.400000 67.780000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 15.840000 67.780000 16.160000 ;
      LAYER met4 ;
        RECT 67.460000 15.840000 67.780000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 16.280000 67.780000 16.600000 ;
      LAYER met4 ;
        RECT 67.460000 16.280000 67.780000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 16.720000 67.780000 17.040000 ;
      LAYER met4 ;
        RECT 67.460000 16.720000 67.780000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 17.160000 67.780000 17.480000 ;
      LAYER met4 ;
        RECT 67.460000 17.160000 67.780000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 17.600000 67.780000 17.920000 ;
      LAYER met4 ;
        RECT 67.460000 17.600000 67.780000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 18.040000 67.780000 18.360000 ;
      LAYER met4 ;
        RECT 67.460000 18.040000 67.780000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 14.960000 68.185000 15.280000 ;
      LAYER met4 ;
        RECT 67.865000 14.960000 68.185000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 15.400000 68.185000 15.720000 ;
      LAYER met4 ;
        RECT 67.865000 15.400000 68.185000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 15.840000 68.185000 16.160000 ;
      LAYER met4 ;
        RECT 67.865000 15.840000 68.185000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 16.280000 68.185000 16.600000 ;
      LAYER met4 ;
        RECT 67.865000 16.280000 68.185000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 16.720000 68.185000 17.040000 ;
      LAYER met4 ;
        RECT 67.865000 16.720000 68.185000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 17.160000 68.185000 17.480000 ;
      LAYER met4 ;
        RECT 67.865000 17.160000 68.185000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 17.600000 68.185000 17.920000 ;
      LAYER met4 ;
        RECT 67.865000 17.600000 68.185000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 18.040000 68.185000 18.360000 ;
      LAYER met4 ;
        RECT 67.865000 18.040000 68.185000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 14.960000 68.590000 15.280000 ;
      LAYER met4 ;
        RECT 68.270000 14.960000 68.590000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 15.400000 68.590000 15.720000 ;
      LAYER met4 ;
        RECT 68.270000 15.400000 68.590000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 15.840000 68.590000 16.160000 ;
      LAYER met4 ;
        RECT 68.270000 15.840000 68.590000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 16.280000 68.590000 16.600000 ;
      LAYER met4 ;
        RECT 68.270000 16.280000 68.590000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 16.720000 68.590000 17.040000 ;
      LAYER met4 ;
        RECT 68.270000 16.720000 68.590000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 17.160000 68.590000 17.480000 ;
      LAYER met4 ;
        RECT 68.270000 17.160000 68.590000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 17.600000 68.590000 17.920000 ;
      LAYER met4 ;
        RECT 68.270000 17.600000 68.590000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 18.040000 68.590000 18.360000 ;
      LAYER met4 ;
        RECT 68.270000 18.040000 68.590000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 14.960000 68.995000 15.280000 ;
      LAYER met4 ;
        RECT 68.675000 14.960000 68.995000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 15.400000 68.995000 15.720000 ;
      LAYER met4 ;
        RECT 68.675000 15.400000 68.995000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 15.840000 68.995000 16.160000 ;
      LAYER met4 ;
        RECT 68.675000 15.840000 68.995000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 16.280000 68.995000 16.600000 ;
      LAYER met4 ;
        RECT 68.675000 16.280000 68.995000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 16.720000 68.995000 17.040000 ;
      LAYER met4 ;
        RECT 68.675000 16.720000 68.995000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 17.160000 68.995000 17.480000 ;
      LAYER met4 ;
        RECT 68.675000 17.160000 68.995000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 17.600000 68.995000 17.920000 ;
      LAYER met4 ;
        RECT 68.675000 17.600000 68.995000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 18.040000 68.995000 18.360000 ;
      LAYER met4 ;
        RECT 68.675000 18.040000 68.995000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 14.960000 69.400000 15.280000 ;
      LAYER met4 ;
        RECT 69.080000 14.960000 69.400000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 15.400000 69.400000 15.720000 ;
      LAYER met4 ;
        RECT 69.080000 15.400000 69.400000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 15.840000 69.400000 16.160000 ;
      LAYER met4 ;
        RECT 69.080000 15.840000 69.400000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 16.280000 69.400000 16.600000 ;
      LAYER met4 ;
        RECT 69.080000 16.280000 69.400000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 16.720000 69.400000 17.040000 ;
      LAYER met4 ;
        RECT 69.080000 16.720000 69.400000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 17.160000 69.400000 17.480000 ;
      LAYER met4 ;
        RECT 69.080000 17.160000 69.400000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 17.600000 69.400000 17.920000 ;
      LAYER met4 ;
        RECT 69.080000 17.600000 69.400000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 18.040000 69.400000 18.360000 ;
      LAYER met4 ;
        RECT 69.080000 18.040000 69.400000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 14.960000 69.805000 15.280000 ;
      LAYER met4 ;
        RECT 69.485000 14.960000 69.805000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 15.400000 69.805000 15.720000 ;
      LAYER met4 ;
        RECT 69.485000 15.400000 69.805000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 15.840000 69.805000 16.160000 ;
      LAYER met4 ;
        RECT 69.485000 15.840000 69.805000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 16.280000 69.805000 16.600000 ;
      LAYER met4 ;
        RECT 69.485000 16.280000 69.805000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 16.720000 69.805000 17.040000 ;
      LAYER met4 ;
        RECT 69.485000 16.720000 69.805000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 17.160000 69.805000 17.480000 ;
      LAYER met4 ;
        RECT 69.485000 17.160000 69.805000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 17.600000 69.805000 17.920000 ;
      LAYER met4 ;
        RECT 69.485000 17.600000 69.805000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 18.040000 69.805000 18.360000 ;
      LAYER met4 ;
        RECT 69.485000 18.040000 69.805000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 14.960000 70.210000 15.280000 ;
      LAYER met4 ;
        RECT 69.890000 14.960000 70.210000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 15.400000 70.210000 15.720000 ;
      LAYER met4 ;
        RECT 69.890000 15.400000 70.210000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 15.840000 70.210000 16.160000 ;
      LAYER met4 ;
        RECT 69.890000 15.840000 70.210000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 16.280000 70.210000 16.600000 ;
      LAYER met4 ;
        RECT 69.890000 16.280000 70.210000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 16.720000 70.210000 17.040000 ;
      LAYER met4 ;
        RECT 69.890000 16.720000 70.210000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 17.160000 70.210000 17.480000 ;
      LAYER met4 ;
        RECT 69.890000 17.160000 70.210000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 17.600000 70.210000 17.920000 ;
      LAYER met4 ;
        RECT 69.890000 17.600000 70.210000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 18.040000 70.210000 18.360000 ;
      LAYER met4 ;
        RECT 69.890000 18.040000 70.210000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 14.960000 7.355000 15.280000 ;
      LAYER met4 ;
        RECT 7.035000 14.960000 7.355000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 15.400000 7.355000 15.720000 ;
      LAYER met4 ;
        RECT 7.035000 15.400000 7.355000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 15.840000 7.355000 16.160000 ;
      LAYER met4 ;
        RECT 7.035000 15.840000 7.355000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 16.280000 7.355000 16.600000 ;
      LAYER met4 ;
        RECT 7.035000 16.280000 7.355000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 16.720000 7.355000 17.040000 ;
      LAYER met4 ;
        RECT 7.035000 16.720000 7.355000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 17.160000 7.355000 17.480000 ;
      LAYER met4 ;
        RECT 7.035000 17.160000 7.355000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 17.600000 7.355000 17.920000 ;
      LAYER met4 ;
        RECT 7.035000 17.600000 7.355000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 18.040000 7.355000 18.360000 ;
      LAYER met4 ;
        RECT 7.035000 18.040000 7.355000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 14.960000 7.760000 15.280000 ;
      LAYER met4 ;
        RECT 7.440000 14.960000 7.760000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 15.400000 7.760000 15.720000 ;
      LAYER met4 ;
        RECT 7.440000 15.400000 7.760000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 15.840000 7.760000 16.160000 ;
      LAYER met4 ;
        RECT 7.440000 15.840000 7.760000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 16.280000 7.760000 16.600000 ;
      LAYER met4 ;
        RECT 7.440000 16.280000 7.760000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 16.720000 7.760000 17.040000 ;
      LAYER met4 ;
        RECT 7.440000 16.720000 7.760000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 17.160000 7.760000 17.480000 ;
      LAYER met4 ;
        RECT 7.440000 17.160000 7.760000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 17.600000 7.760000 17.920000 ;
      LAYER met4 ;
        RECT 7.440000 17.600000 7.760000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 18.040000 7.760000 18.360000 ;
      LAYER met4 ;
        RECT 7.440000 18.040000 7.760000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 14.960000 8.165000 15.280000 ;
      LAYER met4 ;
        RECT 7.845000 14.960000 8.165000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 15.400000 8.165000 15.720000 ;
      LAYER met4 ;
        RECT 7.845000 15.400000 8.165000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 15.840000 8.165000 16.160000 ;
      LAYER met4 ;
        RECT 7.845000 15.840000 8.165000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 16.280000 8.165000 16.600000 ;
      LAYER met4 ;
        RECT 7.845000 16.280000 8.165000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 16.720000 8.165000 17.040000 ;
      LAYER met4 ;
        RECT 7.845000 16.720000 8.165000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 17.160000 8.165000 17.480000 ;
      LAYER met4 ;
        RECT 7.845000 17.160000 8.165000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 17.600000 8.165000 17.920000 ;
      LAYER met4 ;
        RECT 7.845000 17.600000 8.165000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 18.040000 8.165000 18.360000 ;
      LAYER met4 ;
        RECT 7.845000 18.040000 8.165000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 14.960000 70.615000 15.280000 ;
      LAYER met4 ;
        RECT 70.295000 14.960000 70.615000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 15.400000 70.615000 15.720000 ;
      LAYER met4 ;
        RECT 70.295000 15.400000 70.615000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 15.840000 70.615000 16.160000 ;
      LAYER met4 ;
        RECT 70.295000 15.840000 70.615000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 16.280000 70.615000 16.600000 ;
      LAYER met4 ;
        RECT 70.295000 16.280000 70.615000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 16.720000 70.615000 17.040000 ;
      LAYER met4 ;
        RECT 70.295000 16.720000 70.615000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 17.160000 70.615000 17.480000 ;
      LAYER met4 ;
        RECT 70.295000 17.160000 70.615000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 17.600000 70.615000 17.920000 ;
      LAYER met4 ;
        RECT 70.295000 17.600000 70.615000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 18.040000 70.615000 18.360000 ;
      LAYER met4 ;
        RECT 70.295000 18.040000 70.615000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 14.960000 71.020000 15.280000 ;
      LAYER met4 ;
        RECT 70.700000 14.960000 71.020000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 15.400000 71.020000 15.720000 ;
      LAYER met4 ;
        RECT 70.700000 15.400000 71.020000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 15.840000 71.020000 16.160000 ;
      LAYER met4 ;
        RECT 70.700000 15.840000 71.020000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 16.280000 71.020000 16.600000 ;
      LAYER met4 ;
        RECT 70.700000 16.280000 71.020000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 16.720000 71.020000 17.040000 ;
      LAYER met4 ;
        RECT 70.700000 16.720000 71.020000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 17.160000 71.020000 17.480000 ;
      LAYER met4 ;
        RECT 70.700000 17.160000 71.020000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 17.600000 71.020000 17.920000 ;
      LAYER met4 ;
        RECT 70.700000 17.600000 71.020000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 18.040000 71.020000 18.360000 ;
      LAYER met4 ;
        RECT 70.700000 18.040000 71.020000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 14.960000 71.425000 15.280000 ;
      LAYER met4 ;
        RECT 71.105000 14.960000 71.425000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 15.400000 71.425000 15.720000 ;
      LAYER met4 ;
        RECT 71.105000 15.400000 71.425000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 15.840000 71.425000 16.160000 ;
      LAYER met4 ;
        RECT 71.105000 15.840000 71.425000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 16.280000 71.425000 16.600000 ;
      LAYER met4 ;
        RECT 71.105000 16.280000 71.425000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 16.720000 71.425000 17.040000 ;
      LAYER met4 ;
        RECT 71.105000 16.720000 71.425000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 17.160000 71.425000 17.480000 ;
      LAYER met4 ;
        RECT 71.105000 17.160000 71.425000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 17.600000 71.425000 17.920000 ;
      LAYER met4 ;
        RECT 71.105000 17.600000 71.425000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 18.040000 71.425000 18.360000 ;
      LAYER met4 ;
        RECT 71.105000 18.040000 71.425000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 14.960000 71.830000 15.280000 ;
      LAYER met4 ;
        RECT 71.510000 14.960000 71.830000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 15.400000 71.830000 15.720000 ;
      LAYER met4 ;
        RECT 71.510000 15.400000 71.830000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 15.840000 71.830000 16.160000 ;
      LAYER met4 ;
        RECT 71.510000 15.840000 71.830000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 16.280000 71.830000 16.600000 ;
      LAYER met4 ;
        RECT 71.510000 16.280000 71.830000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 16.720000 71.830000 17.040000 ;
      LAYER met4 ;
        RECT 71.510000 16.720000 71.830000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 17.160000 71.830000 17.480000 ;
      LAYER met4 ;
        RECT 71.510000 17.160000 71.830000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 17.600000 71.830000 17.920000 ;
      LAYER met4 ;
        RECT 71.510000 17.600000 71.830000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 18.040000 71.830000 18.360000 ;
      LAYER met4 ;
        RECT 71.510000 18.040000 71.830000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 14.960000 72.235000 15.280000 ;
      LAYER met4 ;
        RECT 71.915000 14.960000 72.235000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 15.400000 72.235000 15.720000 ;
      LAYER met4 ;
        RECT 71.915000 15.400000 72.235000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 15.840000 72.235000 16.160000 ;
      LAYER met4 ;
        RECT 71.915000 15.840000 72.235000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 16.280000 72.235000 16.600000 ;
      LAYER met4 ;
        RECT 71.915000 16.280000 72.235000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 16.720000 72.235000 17.040000 ;
      LAYER met4 ;
        RECT 71.915000 16.720000 72.235000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 17.160000 72.235000 17.480000 ;
      LAYER met4 ;
        RECT 71.915000 17.160000 72.235000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 17.600000 72.235000 17.920000 ;
      LAYER met4 ;
        RECT 71.915000 17.600000 72.235000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 18.040000 72.235000 18.360000 ;
      LAYER met4 ;
        RECT 71.915000 18.040000 72.235000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 14.960000 72.640000 15.280000 ;
      LAYER met4 ;
        RECT 72.320000 14.960000 72.640000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 15.400000 72.640000 15.720000 ;
      LAYER met4 ;
        RECT 72.320000 15.400000 72.640000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 15.840000 72.640000 16.160000 ;
      LAYER met4 ;
        RECT 72.320000 15.840000 72.640000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 16.280000 72.640000 16.600000 ;
      LAYER met4 ;
        RECT 72.320000 16.280000 72.640000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 16.720000 72.640000 17.040000 ;
      LAYER met4 ;
        RECT 72.320000 16.720000 72.640000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 17.160000 72.640000 17.480000 ;
      LAYER met4 ;
        RECT 72.320000 17.160000 72.640000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 17.600000 72.640000 17.920000 ;
      LAYER met4 ;
        RECT 72.320000 17.600000 72.640000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 18.040000 72.640000 18.360000 ;
      LAYER met4 ;
        RECT 72.320000 18.040000 72.640000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 14.960000 73.045000 15.280000 ;
      LAYER met4 ;
        RECT 72.725000 14.960000 73.045000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 15.400000 73.045000 15.720000 ;
      LAYER met4 ;
        RECT 72.725000 15.400000 73.045000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 15.840000 73.045000 16.160000 ;
      LAYER met4 ;
        RECT 72.725000 15.840000 73.045000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 16.280000 73.045000 16.600000 ;
      LAYER met4 ;
        RECT 72.725000 16.280000 73.045000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 16.720000 73.045000 17.040000 ;
      LAYER met4 ;
        RECT 72.725000 16.720000 73.045000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 17.160000 73.045000 17.480000 ;
      LAYER met4 ;
        RECT 72.725000 17.160000 73.045000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 17.600000 73.045000 17.920000 ;
      LAYER met4 ;
        RECT 72.725000 17.600000 73.045000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 18.040000 73.045000 18.360000 ;
      LAYER met4 ;
        RECT 72.725000 18.040000 73.045000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 14.960000 73.450000 15.280000 ;
      LAYER met4 ;
        RECT 73.130000 14.960000 73.450000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 15.400000 73.450000 15.720000 ;
      LAYER met4 ;
        RECT 73.130000 15.400000 73.450000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 15.840000 73.450000 16.160000 ;
      LAYER met4 ;
        RECT 73.130000 15.840000 73.450000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 16.280000 73.450000 16.600000 ;
      LAYER met4 ;
        RECT 73.130000 16.280000 73.450000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 16.720000 73.450000 17.040000 ;
      LAYER met4 ;
        RECT 73.130000 16.720000 73.450000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 17.160000 73.450000 17.480000 ;
      LAYER met4 ;
        RECT 73.130000 17.160000 73.450000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 17.600000 73.450000 17.920000 ;
      LAYER met4 ;
        RECT 73.130000 17.600000 73.450000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 18.040000 73.450000 18.360000 ;
      LAYER met4 ;
        RECT 73.130000 18.040000 73.450000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 14.960000 73.855000 15.280000 ;
      LAYER met4 ;
        RECT 73.535000 14.960000 73.855000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 15.400000 73.855000 15.720000 ;
      LAYER met4 ;
        RECT 73.535000 15.400000 73.855000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 15.840000 73.855000 16.160000 ;
      LAYER met4 ;
        RECT 73.535000 15.840000 73.855000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 16.280000 73.855000 16.600000 ;
      LAYER met4 ;
        RECT 73.535000 16.280000 73.855000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 16.720000 73.855000 17.040000 ;
      LAYER met4 ;
        RECT 73.535000 16.720000 73.855000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 17.160000 73.855000 17.480000 ;
      LAYER met4 ;
        RECT 73.535000 17.160000 73.855000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 17.600000 73.855000 17.920000 ;
      LAYER met4 ;
        RECT 73.535000 17.600000 73.855000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 18.040000 73.855000 18.360000 ;
      LAYER met4 ;
        RECT 73.535000 18.040000 73.855000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 14.960000 74.260000 15.280000 ;
      LAYER met4 ;
        RECT 73.940000 14.960000 74.260000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 15.400000 74.260000 15.720000 ;
      LAYER met4 ;
        RECT 73.940000 15.400000 74.260000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 15.840000 74.260000 16.160000 ;
      LAYER met4 ;
        RECT 73.940000 15.840000 74.260000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 16.280000 74.260000 16.600000 ;
      LAYER met4 ;
        RECT 73.940000 16.280000 74.260000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 16.720000 74.260000 17.040000 ;
      LAYER met4 ;
        RECT 73.940000 16.720000 74.260000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 17.160000 74.260000 17.480000 ;
      LAYER met4 ;
        RECT 73.940000 17.160000 74.260000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 17.600000 74.260000 17.920000 ;
      LAYER met4 ;
        RECT 73.940000 17.600000 74.260000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 18.040000 74.260000 18.360000 ;
      LAYER met4 ;
        RECT 73.940000 18.040000 74.260000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 14.960000 8.570000 15.280000 ;
      LAYER met4 ;
        RECT 8.250000 14.960000 8.570000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 15.400000 8.570000 15.720000 ;
      LAYER met4 ;
        RECT 8.250000 15.400000 8.570000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 15.840000 8.570000 16.160000 ;
      LAYER met4 ;
        RECT 8.250000 15.840000 8.570000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 16.280000 8.570000 16.600000 ;
      LAYER met4 ;
        RECT 8.250000 16.280000 8.570000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 16.720000 8.570000 17.040000 ;
      LAYER met4 ;
        RECT 8.250000 16.720000 8.570000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 17.160000 8.570000 17.480000 ;
      LAYER met4 ;
        RECT 8.250000 17.160000 8.570000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 17.600000 8.570000 17.920000 ;
      LAYER met4 ;
        RECT 8.250000 17.600000 8.570000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 18.040000 8.570000 18.360000 ;
      LAYER met4 ;
        RECT 8.250000 18.040000 8.570000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 14.960000 8.975000 15.280000 ;
      LAYER met4 ;
        RECT 8.655000 14.960000 8.975000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 15.400000 8.975000 15.720000 ;
      LAYER met4 ;
        RECT 8.655000 15.400000 8.975000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 15.840000 8.975000 16.160000 ;
      LAYER met4 ;
        RECT 8.655000 15.840000 8.975000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 16.280000 8.975000 16.600000 ;
      LAYER met4 ;
        RECT 8.655000 16.280000 8.975000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 16.720000 8.975000 17.040000 ;
      LAYER met4 ;
        RECT 8.655000 16.720000 8.975000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 17.160000 8.975000 17.480000 ;
      LAYER met4 ;
        RECT 8.655000 17.160000 8.975000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 17.600000 8.975000 17.920000 ;
      LAYER met4 ;
        RECT 8.655000 17.600000 8.975000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 18.040000 8.975000 18.360000 ;
      LAYER met4 ;
        RECT 8.655000 18.040000 8.975000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 14.960000 9.380000 15.280000 ;
      LAYER met4 ;
        RECT 9.060000 14.960000 9.380000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 15.400000 9.380000 15.720000 ;
      LAYER met4 ;
        RECT 9.060000 15.400000 9.380000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 15.840000 9.380000 16.160000 ;
      LAYER met4 ;
        RECT 9.060000 15.840000 9.380000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 16.280000 9.380000 16.600000 ;
      LAYER met4 ;
        RECT 9.060000 16.280000 9.380000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 16.720000 9.380000 17.040000 ;
      LAYER met4 ;
        RECT 9.060000 16.720000 9.380000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 17.160000 9.380000 17.480000 ;
      LAYER met4 ;
        RECT 9.060000 17.160000 9.380000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 17.600000 9.380000 17.920000 ;
      LAYER met4 ;
        RECT 9.060000 17.600000 9.380000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 18.040000 9.380000 18.360000 ;
      LAYER met4 ;
        RECT 9.060000 18.040000 9.380000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 14.960000 9.785000 15.280000 ;
      LAYER met4 ;
        RECT 9.465000 14.960000 9.785000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 15.400000 9.785000 15.720000 ;
      LAYER met4 ;
        RECT 9.465000 15.400000 9.785000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 15.840000 9.785000 16.160000 ;
      LAYER met4 ;
        RECT 9.465000 15.840000 9.785000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 16.280000 9.785000 16.600000 ;
      LAYER met4 ;
        RECT 9.465000 16.280000 9.785000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 16.720000 9.785000 17.040000 ;
      LAYER met4 ;
        RECT 9.465000 16.720000 9.785000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 17.160000 9.785000 17.480000 ;
      LAYER met4 ;
        RECT 9.465000 17.160000 9.785000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 17.600000 9.785000 17.920000 ;
      LAYER met4 ;
        RECT 9.465000 17.600000 9.785000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 18.040000 9.785000 18.360000 ;
      LAYER met4 ;
        RECT 9.465000 18.040000 9.785000 18.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 14.960000 10.190000 15.280000 ;
      LAYER met4 ;
        RECT 9.870000 14.960000 10.190000 15.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 15.400000 10.190000 15.720000 ;
      LAYER met4 ;
        RECT 9.870000 15.400000 10.190000 15.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 15.840000 10.190000 16.160000 ;
      LAYER met4 ;
        RECT 9.870000 15.840000 10.190000 16.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 16.280000 10.190000 16.600000 ;
      LAYER met4 ;
        RECT 9.870000 16.280000 10.190000 16.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 16.720000 10.190000 17.040000 ;
      LAYER met4 ;
        RECT 9.870000 16.720000 10.190000 17.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 17.160000 10.190000 17.480000 ;
      LAYER met4 ;
        RECT 9.870000 17.160000 10.190000 17.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 17.600000 10.190000 17.920000 ;
      LAYER met4 ;
        RECT 9.870000 17.600000 10.190000 17.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 18.040000 10.190000 18.360000 ;
      LAYER met4 ;
        RECT 9.870000 18.040000 10.190000 18.360000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met3 ;
      RECT 0.495000 14.940000 74.290000 18.380000 ;
    LAYER met4 ;
      RECT 0.000000  2.035000 75.000000  47.965000 ;
      RECT 0.000000 51.745000 75.000000  52.725000 ;
      RECT 0.000000 56.505000 75.000000 200.000000 ;
    LAYER met5 ;
      RECT 0.000000  2.135000 72.130000  15.035000 ;
      RECT 0.000000 15.035000 75.000000  24.335000 ;
      RECT 0.000000 24.335000 72.130000  36.835000 ;
      RECT 0.000000 36.835000 75.000000  40.085000 ;
      RECT 0.000000 40.085000 72.130000  96.585000 ;
      RECT 0.000000 96.585000 75.000000 200.000000 ;
  END
END sky130_fd_io__overlay_vdda_hvc
END LIBRARY
