# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_io__top_ground_lvc_wpad
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 198 ;
  SYMMETRY R90 ;
  PIN AMUXBUS_A
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 1.270000 54.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 1.270000 49.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN G_PAD
    ANTENNAPARTIALMETALSIDEAREA  243.2170 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 31.695000 162.765000 52.340000 167.120000 ;
    END
  END G_PAD
  PIN BDY2_B2B
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 17.630000 5.115000 53.535000 9.540000 ;
        RECT 17.635000 5.110000 53.535000 5.115000 ;
        RECT 17.705000 5.040000 53.535000 5.110000 ;
        RECT 17.775000 4.970000 53.535000 5.040000 ;
        RECT 17.845000 4.900000 53.535000 4.970000 ;
        RECT 17.915000 4.830000 53.535000 4.900000 ;
        RECT 17.985000 4.760000 53.535000 4.830000 ;
        RECT 18.055000 4.690000 53.535000 4.760000 ;
        RECT 18.125000 4.620000 53.535000 4.690000 ;
        RECT 18.195000 4.550000 53.535000 4.620000 ;
        RECT 18.265000 4.480000 53.535000 4.550000 ;
        RECT 18.335000 4.410000 53.535000 4.480000 ;
        RECT 18.405000 4.340000 53.535000 4.410000 ;
        RECT 18.475000 4.270000 53.535000 4.340000 ;
        RECT 18.545000 4.200000 53.535000 4.270000 ;
        RECT 18.615000 4.130000 53.535000 4.200000 ;
        RECT 18.685000 4.060000 53.535000 4.130000 ;
        RECT 18.755000 3.990000 53.535000 4.060000 ;
        RECT 18.825000 3.920000 53.535000 3.990000 ;
        RECT 18.895000 3.850000 53.535000 3.920000 ;
        RECT 18.965000 3.780000 53.535000 3.850000 ;
        RECT 19.035000 3.710000 53.535000 3.780000 ;
        RECT 19.105000 3.640000 53.535000 3.710000 ;
        RECT 19.175000 3.570000 53.535000 3.640000 ;
        RECT 19.245000 3.500000 53.535000 3.570000 ;
        RECT 19.315000 3.430000 53.535000 3.500000 ;
        RECT 19.385000 3.360000 53.535000 3.430000 ;
        RECT 19.455000 3.290000 53.535000 3.360000 ;
        RECT 19.525000 3.220000 53.535000 3.290000 ;
        RECT 19.595000 3.150000 53.535000 3.220000 ;
        RECT 19.665000 3.080000 53.535000 3.150000 ;
        RECT 19.735000 3.010000 53.535000 3.080000 ;
        RECT 19.805000 2.940000 53.535000 3.010000 ;
        RECT 19.875000 2.870000 53.535000 2.940000 ;
        RECT 19.945000 2.800000 53.535000 2.870000 ;
        RECT 20.015000 2.730000 53.535000 2.800000 ;
        RECT 20.085000 2.660000 53.535000 2.730000 ;
        RECT 20.155000 2.590000 53.535000 2.660000 ;
        RECT 20.225000 2.520000 53.535000 2.590000 ;
        RECT 20.295000 2.450000 53.535000 2.520000 ;
        RECT 20.365000 2.380000 53.535000 2.450000 ;
        RECT 20.435000 2.310000 53.535000 2.380000 ;
        RECT 20.505000 2.240000 53.535000 2.310000 ;
        RECT 20.575000 2.170000 53.535000 2.240000 ;
        RECT 20.645000 2.100000 53.535000 2.170000 ;
        RECT 20.715000 2.030000 53.535000 2.100000 ;
        RECT 20.785000 1.960000 53.535000 2.030000 ;
        RECT 20.855000 1.890000 53.535000 1.960000 ;
        RECT 20.925000 0.000000 53.535000 1.820000 ;
        RECT 20.925000 1.820000 53.535000 1.890000 ;
    END
  END BDY2_B2B
  PIN DRN_LVC1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 15.605000  94.310000 23.935000  94.460000 ;
        RECT 15.605000  94.460000 23.785000  94.610000 ;
        RECT 15.605000  94.610000 23.635000  94.760000 ;
        RECT 15.605000  94.760000 23.485000  94.910000 ;
        RECT 15.605000  94.910000 23.335000  95.060000 ;
        RECT 15.605000  95.060000 23.185000  95.210000 ;
        RECT 15.605000  95.210000 23.035000  95.360000 ;
        RECT 15.605000  95.360000 22.885000  95.510000 ;
        RECT 15.605000  95.510000 22.735000  95.660000 ;
        RECT 15.605000  95.660000 22.585000  95.810000 ;
        RECT 15.605000  95.810000 22.435000  95.960000 ;
        RECT 15.605000  95.960000 22.285000  96.110000 ;
        RECT 15.605000  96.110000 22.135000  96.260000 ;
        RECT 15.605000  96.260000 21.985000  96.410000 ;
        RECT 15.605000  96.410000 21.835000  96.560000 ;
        RECT 15.605000  96.560000 21.685000  96.710000 ;
        RECT 15.605000  96.710000 21.605000  96.790000 ;
        RECT 15.605000  96.790000 21.605000 167.100000 ;
        RECT 15.605000 167.100000 21.605000 167.250000 ;
        RECT 15.605000 167.250000 21.755000 167.400000 ;
        RECT 15.605000 167.400000 21.905000 167.550000 ;
        RECT 15.605000 167.550000 22.055000 167.700000 ;
        RECT 15.605000 167.700000 22.205000 167.850000 ;
        RECT 15.605000 167.850000 22.355000 168.000000 ;
        RECT 15.605000 168.000000 22.505000 168.150000 ;
        RECT 15.605000 168.150000 22.655000 168.300000 ;
        RECT 15.605000 168.300000 22.805000 168.450000 ;
        RECT 15.605000 168.450000 22.955000 168.600000 ;
        RECT 15.605000 168.600000 23.105000 168.750000 ;
        RECT 15.605000 168.750000 23.255000 168.900000 ;
        RECT 15.605000 168.900000 23.405000 169.050000 ;
        RECT 15.605000 169.050000 23.555000 169.200000 ;
        RECT 15.605000 169.200000 23.705000 169.350000 ;
        RECT 15.605000 169.350000 23.855000 169.500000 ;
        RECT 15.605000 169.500000 24.005000 169.650000 ;
        RECT 15.605000 169.650000 24.155000 169.800000 ;
        RECT 15.605000 169.800000 24.305000 169.950000 ;
        RECT 15.605000 169.950000 24.455000 170.100000 ;
        RECT 15.605000 170.100000 24.605000 170.250000 ;
        RECT 15.605000 170.250000 24.755000 170.400000 ;
        RECT 15.605000 170.400000 24.905000 170.550000 ;
        RECT 15.605000 170.550000 25.055000 170.610000 ;
        RECT 15.605000 170.610000 25.115000 189.515000 ;
        RECT 15.715000  94.200000 24.085000  94.310000 ;
        RECT 15.865000  94.050000 24.195000  94.200000 ;
        RECT 16.015000  93.900000 24.345000  94.050000 ;
        RECT 16.165000  93.750000 24.495000  93.900000 ;
        RECT 16.315000  93.600000 24.645000  93.750000 ;
        RECT 16.465000  93.450000 24.795000  93.600000 ;
        RECT 16.615000  93.300000 24.945000  93.450000 ;
        RECT 16.765000  93.150000 25.095000  93.300000 ;
        RECT 16.915000  93.000000 25.245000  93.150000 ;
        RECT 17.065000  92.850000 25.395000  93.000000 ;
        RECT 17.215000  92.700000 25.545000  92.850000 ;
        RECT 17.365000  92.550000 25.695000  92.700000 ;
        RECT 17.515000  92.400000 25.845000  92.550000 ;
        RECT 17.665000  92.250000 25.995000  92.400000 ;
        RECT 17.815000  92.100000 26.145000  92.250000 ;
        RECT 17.965000  91.950000 26.295000  92.100000 ;
        RECT 18.115000  91.800000 26.445000  91.950000 ;
        RECT 18.265000  91.650000 26.595000  91.800000 ;
        RECT 18.415000  91.500000 26.745000  91.650000 ;
        RECT 18.565000  91.350000 26.895000  91.500000 ;
        RECT 18.715000  91.200000 27.045000  91.350000 ;
        RECT 18.865000  91.050000 27.195000  91.200000 ;
        RECT 19.015000  90.900000 27.345000  91.050000 ;
        RECT 19.165000  90.750000 27.495000  90.900000 ;
        RECT 19.315000  90.600000 27.645000  90.750000 ;
        RECT 19.465000  90.450000 27.795000  90.600000 ;
        RECT 19.615000  90.300000 27.945000  90.450000 ;
        RECT 19.765000  90.150000 28.095000  90.300000 ;
        RECT 19.915000  90.000000 28.245000  90.150000 ;
        RECT 20.065000  89.850000 28.395000  90.000000 ;
        RECT 20.215000  89.700000 28.545000  89.850000 ;
        RECT 20.365000  89.550000 28.695000  89.700000 ;
        RECT 20.515000  89.400000 28.845000  89.550000 ;
        RECT 20.665000  89.250000 28.995000  89.400000 ;
        RECT 20.815000  89.100000 29.145000  89.250000 ;
        RECT 20.965000  88.950000 29.295000  89.100000 ;
        RECT 21.115000  88.800000 29.445000  88.950000 ;
        RECT 21.265000  88.650000 29.595000  88.800000 ;
        RECT 21.415000  88.500000 29.745000  88.650000 ;
        RECT 21.565000  88.350000 29.895000  88.500000 ;
        RECT 21.715000  88.200000 30.045000  88.350000 ;
        RECT 21.865000  88.050000 30.195000  88.200000 ;
        RECT 22.015000  87.900000 30.345000  88.050000 ;
        RECT 22.165000  87.750000 30.495000  87.900000 ;
        RECT 22.315000  87.600000 30.645000  87.750000 ;
        RECT 22.465000  87.450000 30.795000  87.600000 ;
        RECT 22.615000  87.300000 30.945000  87.450000 ;
        RECT 22.765000  87.150000 31.095000  87.300000 ;
        RECT 22.915000  87.000000 31.245000  87.150000 ;
        RECT 23.065000  86.850000 31.395000  87.000000 ;
        RECT 23.215000  86.700000 31.545000  86.850000 ;
        RECT 23.365000  86.550000 31.695000  86.700000 ;
        RECT 23.515000  86.400000 31.845000  86.550000 ;
        RECT 23.665000  86.250000 31.995000  86.400000 ;
        RECT 23.670000  86.245000 32.145000  86.250000 ;
        RECT 23.760000  86.155000 32.145000  86.245000 ;
        RECT 23.850000  84.650000 32.165000  84.670000 ;
        RECT 23.850000  84.670000 32.145000  84.690000 ;
        RECT 23.850000  84.690000 32.145000  86.065000 ;
        RECT 23.850000  86.065000 32.145000  86.155000 ;
        RECT 23.920000  84.580000 32.185000  84.650000 ;
        RECT 24.070000  84.430000 32.255000  84.580000 ;
        RECT 24.220000  84.280000 32.405000  84.430000 ;
        RECT 24.370000  84.130000 32.555000  84.280000 ;
        RECT 24.520000  83.980000 32.705000  84.130000 ;
        RECT 24.650000  83.850000 48.870000  83.980000 ;
        RECT 24.800000  83.700000 48.870000  83.850000 ;
        RECT 24.950000  83.550000 48.870000  83.700000 ;
        RECT 25.100000  83.400000 48.870000  83.550000 ;
        RECT 25.250000  83.250000 48.870000  83.400000 ;
        RECT 25.400000  83.100000 48.870000  83.250000 ;
        RECT 25.550000  82.950000 48.870000  83.100000 ;
        RECT 25.700000  82.800000 48.870000  82.950000 ;
        RECT 25.850000  82.650000 48.870000  82.800000 ;
        RECT 26.000000   0.000000 36.880000  71.105000 ;
        RECT 26.000000  71.105000 36.880000  71.255000 ;
        RECT 26.000000  71.255000 37.030000  71.405000 ;
        RECT 26.000000  71.405000 37.180000  71.555000 ;
        RECT 26.000000  71.555000 37.330000  71.705000 ;
        RECT 26.000000  71.705000 37.480000  71.855000 ;
        RECT 26.000000  71.855000 37.630000  72.005000 ;
        RECT 26.000000  72.005000 37.780000  72.155000 ;
        RECT 26.000000  72.155000 37.930000  72.305000 ;
        RECT 26.000000  72.305000 38.080000  72.455000 ;
        RECT 26.000000  72.455000 38.230000  72.605000 ;
        RECT 26.000000  72.605000 38.380000  72.755000 ;
        RECT 26.000000  72.755000 38.530000  72.905000 ;
        RECT 26.000000  72.905000 38.680000  73.055000 ;
        RECT 26.000000  73.055000 38.830000  73.205000 ;
        RECT 26.000000  73.205000 38.980000  73.355000 ;
        RECT 26.000000  73.355000 39.130000  73.505000 ;
        RECT 26.000000  73.505000 39.280000  73.655000 ;
        RECT 26.000000  73.655000 39.430000  73.805000 ;
        RECT 26.000000  73.805000 39.580000  73.955000 ;
        RECT 26.000000  73.955000 39.730000  74.105000 ;
        RECT 26.000000  74.105000 39.880000  74.255000 ;
        RECT 26.000000  74.255000 40.030000  74.405000 ;
        RECT 26.000000  74.405000 40.180000  74.555000 ;
        RECT 26.000000  74.555000 40.330000  74.705000 ;
        RECT 26.000000  74.705000 40.480000  74.740000 ;
        RECT 26.000000  74.740000 46.795000  74.890000 ;
        RECT 26.000000  74.890000 46.945000  75.040000 ;
        RECT 26.000000  75.040000 47.095000  75.190000 ;
        RECT 26.000000  75.190000 47.245000  75.340000 ;
        RECT 26.000000  75.340000 47.395000  75.490000 ;
        RECT 26.000000  75.490000 47.545000  75.640000 ;
        RECT 26.000000  75.640000 47.695000  75.790000 ;
        RECT 26.000000  75.790000 47.845000  75.940000 ;
        RECT 26.000000  75.940000 47.995000  76.090000 ;
        RECT 26.000000  76.090000 48.145000  76.240000 ;
        RECT 26.000000  76.240000 48.295000  76.390000 ;
        RECT 26.000000  76.390000 48.445000  76.540000 ;
        RECT 26.000000  76.540000 48.595000  76.690000 ;
        RECT 26.000000  76.690000 48.745000  76.815000 ;
        RECT 26.000000  76.815000 48.870000  82.500000 ;
        RECT 26.000000  82.500000 48.870000  82.650000 ;
        RECT 26.035000  94.500000 32.035000 162.570000 ;
        RECT 26.035000 162.570000 32.035000 162.720000 ;
        RECT 26.035000 162.720000 32.185000 162.870000 ;
        RECT 26.035000 162.870000 32.335000 163.020000 ;
        RECT 26.035000 163.020000 32.485000 163.170000 ;
        RECT 26.035000 163.170000 32.635000 163.320000 ;
        RECT 26.035000 163.320000 32.785000 163.470000 ;
        RECT 26.035000 163.470000 32.935000 163.620000 ;
        RECT 26.035000 163.620000 33.085000 163.770000 ;
        RECT 26.035000 163.770000 33.235000 163.920000 ;
        RECT 26.035000 163.920000 33.385000 164.070000 ;
        RECT 26.035000 164.070000 33.535000 164.220000 ;
        RECT 26.035000 164.220000 33.685000 164.370000 ;
        RECT 26.035000 164.370000 33.835000 164.520000 ;
        RECT 26.035000 164.520000 33.985000 164.670000 ;
        RECT 26.035000 164.670000 34.135000 164.820000 ;
        RECT 26.035000 164.820000 34.285000 164.970000 ;
        RECT 26.035000 164.970000 34.435000 165.120000 ;
        RECT 26.035000 165.120000 34.585000 165.270000 ;
        RECT 26.035000 165.270000 34.735000 165.420000 ;
        RECT 26.035000 165.420000 34.885000 165.570000 ;
        RECT 26.035000 165.570000 35.035000 165.720000 ;
        RECT 26.035000 165.720000 35.185000 165.870000 ;
        RECT 26.035000 165.870000 35.335000 166.020000 ;
        RECT 26.035000 166.020000 35.485000 166.170000 ;
        RECT 26.035000 166.170000 35.635000 166.320000 ;
        RECT 26.035000 166.320000 35.785000 166.470000 ;
        RECT 26.035000 166.470000 35.935000 166.620000 ;
        RECT 26.035000 166.620000 36.085000 166.770000 ;
        RECT 26.035000 166.770000 36.235000 166.920000 ;
        RECT 26.035000 166.920000 36.385000 167.070000 ;
        RECT 26.035000 167.070000 36.535000 167.220000 ;
        RECT 26.035000 167.220000 36.685000 167.370000 ;
        RECT 26.035000 167.370000 36.835000 167.460000 ;
        RECT 26.035000 167.460000 36.925000 189.515000 ;
        RECT 26.095000  94.440000 32.035000  94.500000 ;
        RECT 26.245000  94.290000 32.035000  94.440000 ;
        RECT 26.395000  94.140000 32.035000  94.290000 ;
        RECT 26.545000  93.990000 32.035000  94.140000 ;
        RECT 26.695000  93.840000 32.035000  93.990000 ;
        RECT 26.845000  93.690000 32.035000  93.840000 ;
        RECT 26.995000  93.540000 32.035000  93.690000 ;
        RECT 27.145000  93.390000 32.035000  93.540000 ;
        RECT 27.160000  93.375000 32.035000  93.390000 ;
        RECT 27.310000  93.225000 32.050000  93.375000 ;
        RECT 27.460000  93.075000 32.200000  93.225000 ;
        RECT 27.610000  92.925000 32.350000  93.075000 ;
        RECT 27.760000  92.775000 32.500000  92.925000 ;
        RECT 27.910000  92.625000 32.650000  92.775000 ;
        RECT 28.060000  92.475000 32.800000  92.625000 ;
        RECT 28.210000  92.325000 32.950000  92.475000 ;
        RECT 28.360000  92.175000 33.100000  92.325000 ;
        RECT 28.510000  92.025000 33.250000  92.175000 ;
        RECT 28.660000  91.875000 33.400000  92.025000 ;
        RECT 28.810000  91.725000 33.550000  91.875000 ;
        RECT 28.960000  91.575000 33.700000  91.725000 ;
        RECT 29.110000  91.425000 33.850000  91.575000 ;
        RECT 29.260000  91.275000 34.000000  91.425000 ;
        RECT 29.410000  91.125000 34.150000  91.275000 ;
        RECT 29.560000  90.975000 34.300000  91.125000 ;
        RECT 29.710000  90.825000 34.450000  90.975000 ;
        RECT 29.860000  90.675000 34.600000  90.825000 ;
        RECT 30.010000  90.525000 34.750000  90.675000 ;
        RECT 30.160000  90.375000 34.900000  90.525000 ;
        RECT 30.175000  90.360000 42.385000  90.375000 ;
        RECT 30.325000  90.210000 42.235000  90.360000 ;
        RECT 30.475000  90.060000 42.085000  90.210000 ;
        RECT 30.625000  89.910000 41.935000  90.060000 ;
        RECT 30.775000  89.760000 41.785000  89.910000 ;
        RECT 30.925000  89.610000 41.635000  89.760000 ;
        RECT 31.075000  89.460000 41.485000  89.610000 ;
        RECT 31.225000  89.310000 41.335000  89.460000 ;
        RECT 31.375000  89.160000 41.185000  89.310000 ;
        RECT 31.525000  89.010000 41.035000  89.160000 ;
        RECT 31.675000  88.860000 40.885000  89.010000 ;
        RECT 31.825000  88.710000 40.735000  88.860000 ;
        RECT 31.975000  88.560000 40.585000  88.710000 ;
        RECT 32.125000  88.410000 40.435000  88.560000 ;
        RECT 32.275000  88.260000 40.285000  88.410000 ;
        RECT 32.425000  88.110000 40.135000  88.260000 ;
        RECT 32.575000  87.960000 39.985000  88.110000 ;
        RECT 32.725000  87.810000 39.835000  87.960000 ;
        RECT 32.875000  87.660000 39.685000  87.810000 ;
        RECT 33.025000  87.510000 39.535000  87.660000 ;
        RECT 33.175000  87.360000 39.385000  87.510000 ;
        RECT 33.305000  87.230000 39.385000  87.360000 ;
        RECT 33.455000  87.080000 39.385000  87.230000 ;
        RECT 33.605000  86.930000 39.385000  87.080000 ;
        RECT 33.755000  86.780000 39.385000  86.930000 ;
        RECT 33.905000  86.630000 39.385000  86.780000 ;
        RECT 33.945000  83.980000 39.945000  84.130000 ;
        RECT 34.055000  86.480000 39.385000  86.630000 ;
        RECT 34.095000  84.130000 39.795000  84.280000 ;
        RECT 34.205000  86.330000 39.385000  86.480000 ;
        RECT 34.245000  84.280000 39.645000  84.430000 ;
        RECT 34.355000  86.180000 39.385000  86.330000 ;
        RECT 34.395000  84.430000 39.495000  84.580000 ;
        RECT 34.505000  84.580000 39.385000  84.690000 ;
        RECT 34.505000  84.690000 39.385000  86.030000 ;
        RECT 34.505000  86.030000 39.385000  86.180000 ;
        RECT 37.945000  90.375000 42.400000  90.525000 ;
        RECT 37.945000 169.025000 48.835000 189.515000 ;
        RECT 38.035000 168.935000 48.835000 169.025000 ;
        RECT 38.095000  90.525000 42.550000  90.675000 ;
        RECT 38.185000 168.785000 48.835000 168.935000 ;
        RECT 38.245000  90.675000 42.700000  90.825000 ;
        RECT 38.335000 168.635000 48.835000 168.785000 ;
        RECT 38.395000  90.825000 42.850000  90.975000 ;
        RECT 38.485000 168.485000 48.835000 168.635000 ;
        RECT 38.545000  90.975000 43.000000  91.125000 ;
        RECT 38.635000 168.335000 48.835000 168.485000 ;
        RECT 38.695000  91.125000 43.150000  91.275000 ;
        RECT 38.785000 168.185000 48.835000 168.335000 ;
        RECT 38.845000  91.275000 43.300000  91.425000 ;
        RECT 38.935000 168.035000 48.835000 168.185000 ;
        RECT 38.995000  91.425000 43.450000  91.575000 ;
        RECT 39.085000 167.885000 48.835000 168.035000 ;
        RECT 39.145000  91.575000 43.600000  91.725000 ;
        RECT 39.235000 167.735000 48.835000 167.885000 ;
        RECT 39.295000  91.725000 43.750000  91.875000 ;
        RECT 39.385000 167.585000 48.835000 167.735000 ;
        RECT 39.445000  91.875000 43.900000  92.025000 ;
        RECT 39.535000 167.435000 48.835000 167.585000 ;
        RECT 39.595000  92.025000 44.050000  92.175000 ;
        RECT 39.685000 167.285000 48.835000 167.435000 ;
        RECT 39.745000  92.175000 44.200000  92.325000 ;
        RECT 39.835000 167.135000 48.835000 167.285000 ;
        RECT 39.895000  92.325000 44.350000  92.475000 ;
        RECT 39.985000 166.985000 48.835000 167.135000 ;
        RECT 40.045000  92.475000 44.500000  92.625000 ;
        RECT 40.135000 166.835000 48.835000 166.985000 ;
        RECT 40.195000  92.625000 44.650000  92.775000 ;
        RECT 40.285000 166.685000 48.835000 166.835000 ;
        RECT 40.345000  92.775000 44.800000  92.925000 ;
        RECT 40.435000 166.535000 48.835000 166.685000 ;
        RECT 40.495000  92.925000 44.950000  93.075000 ;
        RECT 40.585000 166.385000 48.835000 166.535000 ;
        RECT 40.645000  93.075000 45.100000  93.225000 ;
        RECT 40.735000 166.235000 48.835000 166.385000 ;
        RECT 40.795000  93.225000 45.250000  93.375000 ;
        RECT 40.885000 166.085000 48.835000 166.235000 ;
        RECT 40.945000  93.375000 45.400000  93.525000 ;
        RECT 41.035000 165.935000 48.835000 166.085000 ;
        RECT 41.050000  83.980000 48.870000  84.130000 ;
        RECT 41.095000  93.525000 45.550000  93.675000 ;
        RECT 41.185000 165.785000 48.835000 165.935000 ;
        RECT 41.200000  84.130000 48.870000  84.280000 ;
        RECT 41.245000  93.675000 45.700000  93.825000 ;
        RECT 41.335000 165.635000 48.835000 165.785000 ;
        RECT 41.350000  84.280000 48.870000  84.430000 ;
        RECT 41.395000  93.825000 45.850000  93.975000 ;
        RECT 41.485000 165.485000 48.835000 165.635000 ;
        RECT 41.500000  84.430000 48.870000  84.580000 ;
        RECT 41.545000  93.975000 46.000000  94.125000 ;
        RECT 41.610000  84.580000 48.870000  84.690000 ;
        RECT 41.610000  84.690000 48.870000  84.810000 ;
        RECT 41.610000  84.810000 48.870000  84.960000 ;
        RECT 41.610000  84.960000 49.020000  85.110000 ;
        RECT 41.610000  85.110000 49.170000  85.260000 ;
        RECT 41.610000  85.260000 49.320000  85.410000 ;
        RECT 41.610000  85.410000 49.470000  85.560000 ;
        RECT 41.610000  85.560000 49.620000  85.710000 ;
        RECT 41.610000  85.710000 49.770000  85.860000 ;
        RECT 41.610000  85.860000 49.920000  86.010000 ;
        RECT 41.610000  86.010000 50.070000  86.160000 ;
        RECT 41.610000  86.160000 50.220000  86.310000 ;
        RECT 41.610000  86.310000 50.370000  86.460000 ;
        RECT 41.610000  86.460000 50.520000  86.610000 ;
        RECT 41.610000  86.610000 50.670000  86.760000 ;
        RECT 41.610000  86.760000 50.820000  86.910000 ;
        RECT 41.610000  86.910000 50.970000  86.960000 ;
        RECT 41.610000  86.960000 51.020000  87.445000 ;
        RECT 41.635000 165.335000 48.835000 165.485000 ;
        RECT 41.695000  94.125000 46.150000  94.275000 ;
        RECT 41.760000  87.445000 51.020000  87.595000 ;
        RECT 41.785000 165.185000 48.835000 165.335000 ;
        RECT 41.845000  94.275000 46.300000  94.425000 ;
        RECT 41.910000  87.595000 51.020000  87.745000 ;
        RECT 41.935000 165.035000 48.835000 165.185000 ;
        RECT 41.995000  94.425000 46.450000  94.575000 ;
        RECT 42.060000  87.745000 51.020000  87.895000 ;
        RECT 42.085000 164.885000 48.835000 165.035000 ;
        RECT 42.145000  94.575000 46.600000  94.725000 ;
        RECT 42.210000  87.895000 51.020000  88.045000 ;
        RECT 42.235000 164.735000 48.835000 164.885000 ;
        RECT 42.295000  94.725000 46.750000  94.875000 ;
        RECT 42.360000  88.045000 51.020000  88.195000 ;
        RECT 42.385000 164.585000 48.835000 164.735000 ;
        RECT 42.445000  94.875000 46.900000  95.025000 ;
        RECT 42.510000  88.195000 51.020000  88.345000 ;
        RECT 42.535000 164.435000 48.835000 164.585000 ;
        RECT 42.540000  88.345000 51.020000  88.375000 ;
        RECT 42.595000  95.025000 47.050000  95.175000 ;
        RECT 42.685000 164.285000 48.835000 164.435000 ;
        RECT 42.690000  88.375000 51.020000  88.525000 ;
        RECT 42.745000  95.175000 47.200000  95.325000 ;
        RECT 42.835000  95.325000 47.350000  95.415000 ;
        RECT 42.835000  95.415000 47.440000  95.565000 ;
        RECT 42.835000  95.565000 47.590000  95.715000 ;
        RECT 42.835000  95.715000 47.740000  95.865000 ;
        RECT 42.835000  95.865000 47.890000  96.015000 ;
        RECT 42.835000  96.015000 48.040000  96.165000 ;
        RECT 42.835000  96.165000 48.190000  96.315000 ;
        RECT 42.835000  96.315000 48.340000  96.465000 ;
        RECT 42.835000  96.465000 48.490000  96.615000 ;
        RECT 42.835000  96.615000 48.640000  96.765000 ;
        RECT 42.835000  96.765000 48.790000  96.810000 ;
        RECT 42.835000  96.810000 48.835000 164.135000 ;
        RECT 42.835000 164.135000 48.835000 164.285000 ;
        RECT 42.840000  88.525000 51.170000  88.675000 ;
        RECT 42.990000  88.675000 51.320000  88.825000 ;
        RECT 43.140000  88.825000 51.470000  88.975000 ;
        RECT 43.290000  88.975000 51.620000  89.125000 ;
        RECT 43.440000  89.125000 51.770000  89.275000 ;
        RECT 43.590000  89.275000 51.920000  89.425000 ;
        RECT 43.740000  89.425000 52.070000  89.575000 ;
        RECT 43.890000  89.575000 52.220000  89.725000 ;
        RECT 44.040000  89.725000 52.370000  89.875000 ;
        RECT 44.190000  89.875000 52.520000  90.025000 ;
        RECT 44.340000  90.025000 52.670000  90.175000 ;
        RECT 44.490000  90.175000 52.820000  90.325000 ;
        RECT 44.640000  90.325000 52.970000  90.475000 ;
        RECT 44.790000  90.475000 53.120000  90.625000 ;
        RECT 44.940000  90.625000 53.270000  90.775000 ;
        RECT 45.090000  90.775000 53.420000  90.925000 ;
        RECT 45.240000  90.925000 53.570000  91.075000 ;
        RECT 45.390000  91.075000 53.720000  91.225000 ;
        RECT 45.540000  91.225000 53.870000  91.375000 ;
        RECT 45.690000  91.375000 54.020000  91.525000 ;
        RECT 45.840000  91.525000 54.170000  91.675000 ;
        RECT 45.990000  91.675000 54.320000  91.825000 ;
        RECT 46.140000  91.825000 54.470000  91.975000 ;
        RECT 46.290000  91.975000 54.620000  92.125000 ;
        RECT 46.440000  92.125000 54.770000  92.275000 ;
        RECT 46.590000  92.275000 54.920000  92.425000 ;
        RECT 46.740000  92.425000 55.070000  92.575000 ;
        RECT 46.890000  92.575000 55.220000  92.725000 ;
        RECT 47.040000  92.725000 55.370000  92.875000 ;
        RECT 47.190000  92.875000 55.520000  93.025000 ;
        RECT 47.340000  93.025000 55.670000  93.175000 ;
        RECT 47.490000  93.175000 55.820000  93.325000 ;
        RECT 47.640000  93.325000 55.970000  93.475000 ;
        RECT 47.790000  93.475000 56.120000  93.625000 ;
        RECT 47.940000  93.625000 56.270000  93.775000 ;
        RECT 48.090000  93.775000 56.420000  93.925000 ;
        RECT 48.240000  93.925000 56.570000  94.075000 ;
        RECT 48.390000  94.075000 56.720000  94.225000 ;
        RECT 48.540000  94.225000 56.870000  94.375000 ;
        RECT 48.690000  94.375000 57.020000  94.525000 ;
        RECT 48.840000  94.525000 57.170000  94.675000 ;
        RECT 48.990000  94.675000 57.320000  94.825000 ;
        RECT 49.140000  94.825000 57.470000  94.975000 ;
        RECT 49.290000  94.975000 57.620000  95.125000 ;
        RECT 49.440000  95.125000 57.770000  95.275000 ;
        RECT 49.590000  95.275000 57.920000  95.425000 ;
        RECT 49.740000  95.425000 58.070000  95.575000 ;
        RECT 49.870000 168.920000 60.330000 189.515000 ;
        RECT 49.890000  95.575000 58.220000  95.725000 ;
        RECT 49.980000 168.810000 60.330000 168.920000 ;
        RECT 50.040000  95.725000 58.370000  95.875000 ;
        RECT 50.130000 168.660000 60.330000 168.810000 ;
        RECT 50.190000  95.875000 58.520000  96.025000 ;
        RECT 50.280000 168.510000 60.330000 168.660000 ;
        RECT 50.340000  96.025000 58.670000  96.175000 ;
        RECT 50.430000 168.360000 60.330000 168.510000 ;
        RECT 50.490000  96.175000 58.820000  96.325000 ;
        RECT 50.580000 168.210000 60.330000 168.360000 ;
        RECT 50.640000  96.325000 58.970000  96.475000 ;
        RECT 50.730000 168.060000 60.330000 168.210000 ;
        RECT 50.790000  96.475000 59.120000  96.625000 ;
        RECT 50.880000 167.910000 60.330000 168.060000 ;
        RECT 50.940000  96.625000 59.270000  96.775000 ;
        RECT 51.030000 167.760000 60.330000 167.910000 ;
        RECT 51.090000  96.775000 59.420000  96.925000 ;
        RECT 51.180000 167.610000 60.330000 167.760000 ;
        RECT 51.240000  96.925000 59.570000  97.075000 ;
        RECT 51.330000 167.460000 60.330000 167.610000 ;
        RECT 51.390000  97.075000 59.720000  97.225000 ;
        RECT 51.480000 167.310000 60.330000 167.460000 ;
        RECT 51.540000  97.225000 59.870000  97.375000 ;
        RECT 51.630000 167.160000 60.330000 167.310000 ;
        RECT 51.690000  97.375000 60.020000  97.525000 ;
        RECT 51.780000 167.010000 60.330000 167.160000 ;
        RECT 51.840000  97.525000 60.170000  97.675000 ;
        RECT 51.850000  97.675000 60.320000  97.685000 ;
        RECT 51.930000 166.860000 60.330000 167.010000 ;
        RECT 52.000000  97.685000 60.330000  97.835000 ;
        RECT 52.080000 166.710000 60.330000 166.860000 ;
        RECT 52.150000  97.835000 60.330000  97.985000 ;
        RECT 52.230000 166.560000 60.330000 166.710000 ;
        RECT 52.300000  97.985000 60.330000  98.135000 ;
        RECT 52.380000 166.410000 60.330000 166.560000 ;
        RECT 52.450000  98.135000 60.330000  98.285000 ;
        RECT 52.530000 166.260000 60.330000 166.410000 ;
        RECT 52.600000  98.285000 60.330000  98.435000 ;
        RECT 52.680000 166.110000 60.330000 166.260000 ;
        RECT 52.750000  98.435000 60.330000  98.585000 ;
        RECT 52.830000 165.960000 60.330000 166.110000 ;
        RECT 52.900000  98.585000 60.330000  98.735000 ;
        RECT 52.980000 165.810000 60.330000 165.960000 ;
        RECT 53.050000  98.735000 60.330000  98.885000 ;
        RECT 53.130000 165.660000 60.330000 165.810000 ;
        RECT 53.200000  98.885000 60.330000  99.035000 ;
        RECT 53.280000 165.510000 60.330000 165.660000 ;
        RECT 53.350000  99.035000 60.330000  99.185000 ;
        RECT 53.430000 165.360000 60.330000 165.510000 ;
        RECT 53.500000  99.185000 60.330000  99.335000 ;
        RECT 53.580000 165.210000 60.330000 165.360000 ;
        RECT 53.650000  99.335000 60.330000  99.485000 ;
        RECT 53.730000 165.060000 60.330000 165.210000 ;
        RECT 53.800000  99.485000 60.330000  99.635000 ;
        RECT 53.880000 164.910000 60.330000 165.060000 ;
        RECT 53.950000  99.635000 60.330000  99.785000 ;
        RECT 54.030000 164.760000 60.330000 164.910000 ;
        RECT 54.100000  99.785000 60.330000  99.935000 ;
        RECT 54.180000 164.610000 60.330000 164.760000 ;
        RECT 54.250000  99.935000 60.330000 100.085000 ;
        RECT 54.330000 100.085000 60.330000 100.165000 ;
        RECT 54.330000 100.165000 60.330000 164.460000 ;
        RECT 54.330000 164.460000 60.330000 164.610000 ;
    END
  END DRN_LVC1
  PIN DRN_LVC2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.380000 0.000000 49.255000 69.490000 ;
    END
  END DRN_LVC2
  PIN G_CORE
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.500000  0.000000 24.500000  82.660000 ;
        RECT 0.500000 82.660000 24.350000  82.810000 ;
        RECT 0.500000 82.810000 24.200000  82.960000 ;
        RECT 0.500000 82.960000 24.050000  83.110000 ;
        RECT 0.500000 83.110000 23.900000  83.260000 ;
        RECT 0.500000 83.260000 23.750000  83.410000 ;
        RECT 0.500000 83.410000 23.600000  83.560000 ;
        RECT 0.500000 83.560000 23.450000  83.710000 ;
        RECT 0.500000 83.710000 23.300000  83.860000 ;
        RECT 0.500000 83.860000 23.150000  84.010000 ;
        RECT 0.500000 84.010000 23.000000  84.160000 ;
        RECT 0.500000 84.160000 22.850000  84.310000 ;
        RECT 0.500000 84.310000 22.700000  84.460000 ;
        RECT 0.500000 84.460000 22.550000  84.610000 ;
        RECT 0.500000 84.610000 22.400000  84.760000 ;
        RECT 0.500000 84.760000 22.250000  84.910000 ;
        RECT 0.500000 84.910000 22.100000  85.060000 ;
        RECT 0.500000 85.060000 21.950000  85.210000 ;
        RECT 0.500000 85.210000 21.800000  85.360000 ;
        RECT 0.500000 85.360000 21.650000  85.510000 ;
        RECT 0.500000 85.510000 21.500000  85.660000 ;
        RECT 0.500000 85.660000 21.350000  85.810000 ;
        RECT 0.500000 85.810000 21.200000  85.960000 ;
        RECT 0.500000 85.960000 21.050000  86.110000 ;
        RECT 0.500000 86.110000 20.900000  86.260000 ;
        RECT 0.500000 86.260000 20.750000  86.410000 ;
        RECT 0.500000 86.410000 20.600000  86.560000 ;
        RECT 0.500000 86.560000 20.450000  86.710000 ;
        RECT 0.500000 86.710000 20.300000  86.860000 ;
        RECT 0.500000 86.860000 20.150000  87.010000 ;
        RECT 0.500000 87.010000 20.000000  87.160000 ;
        RECT 0.500000 87.160000 19.850000  87.310000 ;
        RECT 0.500000 87.310000 19.700000  87.460000 ;
        RECT 0.500000 87.460000 19.550000  87.610000 ;
        RECT 0.500000 87.610000 19.400000  87.760000 ;
        RECT 0.500000 87.760000 19.250000  87.910000 ;
        RECT 0.500000 87.910000 19.100000  88.060000 ;
        RECT 0.500000 88.060000 18.950000  88.210000 ;
        RECT 0.500000 88.210000 18.800000  88.360000 ;
        RECT 0.500000 88.360000 18.650000  88.510000 ;
        RECT 0.500000 88.510000 18.500000  88.660000 ;
        RECT 0.500000 88.660000 18.350000  88.810000 ;
        RECT 0.500000 88.810000 18.200000  88.960000 ;
        RECT 0.500000 88.960000 18.050000  89.110000 ;
        RECT 0.500000 89.110000 17.900000  89.260000 ;
        RECT 0.500000 89.260000 17.750000  89.410000 ;
        RECT 0.500000 89.410000 17.600000  89.560000 ;
        RECT 0.500000 89.560000 17.450000  89.710000 ;
        RECT 0.500000 89.710000 17.300000  89.860000 ;
        RECT 0.500000 89.860000 17.150000  90.010000 ;
        RECT 0.500000 90.010000 17.000000  90.160000 ;
        RECT 0.500000 90.160000 16.850000  90.310000 ;
        RECT 0.500000 90.310000 16.700000  90.460000 ;
        RECT 0.500000 90.460000 16.550000  90.610000 ;
        RECT 0.500000 90.610000 16.400000  90.760000 ;
        RECT 0.500000 90.760000 16.250000  90.910000 ;
        RECT 0.500000 90.910000 16.100000  91.060000 ;
        RECT 0.500000 91.060000 15.950000  91.210000 ;
        RECT 0.500000 91.210000 15.800000  91.360000 ;
        RECT 0.500000 91.360000 15.650000  91.510000 ;
        RECT 0.500000 91.510000 15.500000  91.660000 ;
        RECT 0.500000 91.660000 15.350000  91.810000 ;
        RECT 0.500000 91.810000 15.200000  91.960000 ;
        RECT 0.500000 91.960000 15.050000  92.110000 ;
        RECT 0.500000 92.110000 14.900000  92.260000 ;
        RECT 0.500000 92.260000 14.750000  92.410000 ;
        RECT 0.500000 92.410000 14.600000  92.560000 ;
        RECT 0.500000 92.560000 14.450000  92.710000 ;
        RECT 0.500000 92.710000 14.300000  92.860000 ;
        RECT 0.500000 92.860000 14.150000  93.010000 ;
        RECT 0.500000 93.010000 14.000000  93.160000 ;
        RECT 0.500000 93.160000 13.850000  93.310000 ;
        RECT 0.500000 93.310000 13.700000  93.460000 ;
        RECT 0.500000 93.460000 13.550000  93.610000 ;
        RECT 0.500000 93.610000 13.400000  93.760000 ;
        RECT 0.500000 93.760000 13.250000  93.910000 ;
        RECT 0.500000 93.910000 13.100000  94.060000 ;
        RECT 0.500000 94.060000 12.950000  94.210000 ;
        RECT 0.500000 94.210000 12.900000  94.260000 ;
        RECT 0.500000 94.260000 12.900000 171.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000  0.000000 74.700000  84.465000 ;
        RECT 50.905000 84.465000 74.700000  84.615000 ;
        RECT 51.055000 84.615000 74.700000  84.765000 ;
        RECT 51.205000 84.765000 74.700000  84.915000 ;
        RECT 51.355000 84.915000 74.700000  85.065000 ;
        RECT 51.505000 85.065000 74.700000  85.215000 ;
        RECT 51.655000 85.215000 74.700000  85.365000 ;
        RECT 51.805000 85.365000 74.700000  85.515000 ;
        RECT 51.955000 85.515000 74.700000  85.665000 ;
        RECT 52.105000 85.665000 74.700000  85.815000 ;
        RECT 52.255000 85.815000 74.700000  85.965000 ;
        RECT 52.405000 85.965000 74.700000  86.115000 ;
        RECT 52.555000 86.115000 74.700000  86.265000 ;
        RECT 52.705000 86.265000 74.700000  86.415000 ;
        RECT 52.855000 86.415000 74.700000  86.565000 ;
        RECT 53.005000 86.565000 74.700000  86.715000 ;
        RECT 53.155000 86.715000 74.700000  86.865000 ;
        RECT 53.305000 86.865000 74.700000  87.015000 ;
        RECT 53.455000 87.015000 74.700000  87.165000 ;
        RECT 53.605000 87.165000 74.700000  87.315000 ;
        RECT 53.755000 87.315000 74.700000  87.465000 ;
        RECT 53.905000 87.465000 74.700000  87.615000 ;
        RECT 54.055000 87.615000 74.700000  87.765000 ;
        RECT 54.205000 87.765000 74.700000  87.915000 ;
        RECT 54.355000 87.915000 74.700000  88.065000 ;
        RECT 54.505000 88.065000 74.700000  88.215000 ;
        RECT 54.655000 88.215000 74.700000  88.365000 ;
        RECT 54.805000 88.365000 74.700000  88.515000 ;
        RECT 54.955000 88.515000 74.700000  88.665000 ;
        RECT 55.105000 88.665000 74.700000  88.815000 ;
        RECT 55.255000 88.815000 74.700000  88.965000 ;
        RECT 55.405000 88.965000 74.700000  89.115000 ;
        RECT 55.555000 89.115000 74.700000  89.265000 ;
        RECT 55.705000 89.265000 74.700000  89.415000 ;
        RECT 55.855000 89.415000 74.700000  89.565000 ;
        RECT 56.005000 89.565000 74.700000  89.715000 ;
        RECT 56.155000 89.715000 74.700000  89.865000 ;
        RECT 56.305000 89.865000 74.700000  90.015000 ;
        RECT 56.455000 90.015000 74.700000  90.165000 ;
        RECT 56.605000 90.165000 74.700000  90.315000 ;
        RECT 56.755000 90.315000 74.700000  90.465000 ;
        RECT 56.905000 90.465000 74.700000  90.615000 ;
        RECT 57.055000 90.615000 74.700000  90.765000 ;
        RECT 57.205000 90.765000 74.700000  90.915000 ;
        RECT 57.355000 90.915000 74.700000  91.065000 ;
        RECT 57.505000 91.065000 74.700000  91.215000 ;
        RECT 57.655000 91.215000 74.700000  91.365000 ;
        RECT 57.805000 91.365000 74.700000  91.515000 ;
        RECT 57.955000 91.515000 74.700000  91.665000 ;
        RECT 58.105000 91.665000 74.700000  91.815000 ;
        RECT 58.255000 91.815000 74.700000  91.965000 ;
        RECT 58.405000 91.965000 74.700000  92.115000 ;
        RECT 58.555000 92.115000 74.700000  92.265000 ;
        RECT 58.705000 92.265000 74.700000  92.415000 ;
        RECT 58.855000 92.415000 74.700000  92.565000 ;
        RECT 59.005000 92.565000 74.700000  92.715000 ;
        RECT 59.155000 92.715000 74.700000  92.865000 ;
        RECT 59.305000 92.865000 74.700000  93.015000 ;
        RECT 59.455000 93.015000 74.700000  93.165000 ;
        RECT 59.605000 93.165000 74.700000  93.315000 ;
        RECT 59.755000 93.315000 74.700000  93.465000 ;
        RECT 59.905000 93.465000 74.700000  93.615000 ;
        RECT 60.055000 93.615000 74.700000  93.765000 ;
        RECT 60.205000 93.765000 74.700000  93.915000 ;
        RECT 60.355000 93.915000 74.700000  94.065000 ;
        RECT 60.505000 94.065000 74.700000  94.215000 ;
        RECT 60.655000 94.215000 74.700000  94.365000 ;
        RECT 60.805000 94.365000 74.700000  94.515000 ;
        RECT 60.955000 94.515000 74.700000  94.665000 ;
        RECT 61.105000 94.665000 74.700000  94.815000 ;
        RECT 61.255000 94.815000 74.700000  94.965000 ;
        RECT 61.405000 94.965000 74.700000  95.115000 ;
        RECT 61.555000 95.115000 74.700000  95.265000 ;
        RECT 61.705000 95.265000 74.700000  95.415000 ;
        RECT 61.855000 95.415000 74.700000  95.565000 ;
        RECT 62.005000 95.565000 74.700000  95.715000 ;
        RECT 62.045000 95.715000 74.700000  95.755000 ;
        RECT 62.045000 95.755000 74.700000 172.235000 ;
    END
  END G_CORE
  PIN OGC_LVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 26.210000 0.000000 27.700000 0.170000 ;
    END
  END OGC_LVC
  PIN SRC_BDY_LVC1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT  0.500000   0.000000 20.495000   1.485000 ;
        RECT  0.500000   1.485000 20.425000   1.555000 ;
        RECT  0.500000   1.555000 20.355000   1.625000 ;
        RECT  0.500000   1.625000 20.285000   1.695000 ;
        RECT  0.500000   1.695000 20.215000   1.765000 ;
        RECT  0.500000   1.765000 20.145000   1.835000 ;
        RECT  0.500000   1.835000 20.075000   1.905000 ;
        RECT  0.500000   1.905000 20.005000   1.975000 ;
        RECT  0.500000   1.975000 19.935000   2.045000 ;
        RECT  0.500000   2.045000 19.865000   2.115000 ;
        RECT  0.500000   2.115000 19.795000   2.185000 ;
        RECT  0.500000   2.185000 19.725000   2.255000 ;
        RECT  0.500000   2.255000 19.655000   2.325000 ;
        RECT  0.500000   2.325000 19.585000   2.395000 ;
        RECT  0.500000   2.395000 19.515000   2.465000 ;
        RECT  0.500000   2.465000 19.445000   2.535000 ;
        RECT  0.500000   2.535000 19.375000   2.605000 ;
        RECT  0.500000   2.605000 19.305000   2.675000 ;
        RECT  0.500000   2.675000 19.235000   2.745000 ;
        RECT  0.500000   2.745000 19.165000   2.815000 ;
        RECT  0.500000   2.815000 19.095000   2.885000 ;
        RECT  0.500000   2.885000 19.025000   2.955000 ;
        RECT  0.500000   2.955000 18.955000   3.025000 ;
        RECT  0.500000   3.025000 18.885000   3.095000 ;
        RECT  0.500000   3.095000 18.815000   3.165000 ;
        RECT  0.500000   3.165000 18.745000   3.235000 ;
        RECT  0.500000   3.235000 18.675000   3.305000 ;
        RECT  0.500000   3.305000 18.605000   3.375000 ;
        RECT  0.500000   3.375000 18.535000   3.445000 ;
        RECT  0.500000   3.445000 18.465000   3.515000 ;
        RECT  0.500000   3.515000 18.395000   3.585000 ;
        RECT  0.500000   3.585000 18.325000   3.655000 ;
        RECT  0.500000   3.655000 18.255000   3.725000 ;
        RECT  0.500000   3.725000 18.185000   3.795000 ;
        RECT  0.500000   3.795000 18.115000   3.865000 ;
        RECT  0.500000   3.865000 18.045000   3.935000 ;
        RECT  0.500000   3.935000 17.975000   4.005000 ;
        RECT  0.500000   4.005000 17.905000   4.075000 ;
        RECT  0.500000   4.075000 17.835000   4.145000 ;
        RECT  0.500000   4.145000 17.765000   4.215000 ;
        RECT  0.500000   4.215000 17.695000   4.285000 ;
        RECT  0.500000   4.285000 17.625000   4.355000 ;
        RECT  0.500000   4.355000 17.555000   4.425000 ;
        RECT  0.500000   4.425000 17.485000   4.495000 ;
        RECT  0.500000   4.495000 17.415000   4.565000 ;
        RECT  0.500000   4.565000 17.345000   4.635000 ;
        RECT  0.500000   4.635000 17.275000   4.705000 ;
        RECT  0.500000   4.705000 17.205000   4.775000 ;
        RECT  0.500000   4.775000 17.135000   4.845000 ;
        RECT  0.500000   4.845000 17.065000   4.915000 ;
        RECT  0.500000   4.915000 16.995000   4.985000 ;
        RECT  0.500000   4.985000 16.925000   5.055000 ;
        RECT  0.500000   5.055000 16.860000   5.120000 ;
        RECT  0.500000   5.120000 16.860000   7.655000 ;
        RECT  0.500000   7.655000 10.745000   7.725000 ;
        RECT  0.500000   7.725000 10.675000   7.795000 ;
        RECT  0.500000   7.795000 10.605000   7.865000 ;
        RECT  0.500000   7.865000 10.535000   7.935000 ;
        RECT  0.500000   7.935000 10.465000   8.005000 ;
        RECT  0.500000   8.005000 10.420000   8.050000 ;
        RECT  0.500000   8.050000 10.420000   9.820000 ;
        RECT  0.500000   9.820000 10.420000   9.890000 ;
        RECT  0.500000   9.890000 10.490000   9.960000 ;
        RECT  0.500000   9.960000 10.560000  10.030000 ;
        RECT  0.500000  10.030000 10.630000  10.100000 ;
        RECT  0.500000  10.100000 10.700000  10.170000 ;
        RECT  0.500000  10.170000 10.770000  10.215000 ;
        RECT  0.500000  10.215000 55.595000  17.080000 ;
        RECT  0.500000  17.080000 21.785000  17.150000 ;
        RECT  0.500000  17.150000 21.715000  17.220000 ;
        RECT  0.500000  17.220000 21.645000  17.290000 ;
        RECT  0.500000  17.290000 21.575000  17.360000 ;
        RECT  0.500000  17.360000 21.505000  17.430000 ;
        RECT  0.500000  17.430000 21.435000  17.500000 ;
        RECT  0.500000  17.500000 21.365000  17.570000 ;
        RECT  0.500000  17.570000 21.295000  17.640000 ;
        RECT  0.500000  17.640000 21.225000  17.710000 ;
        RECT  0.500000  17.710000 21.155000  17.780000 ;
        RECT  0.500000  17.780000 21.085000  17.850000 ;
        RECT  0.500000  17.850000 21.015000  17.920000 ;
        RECT  0.500000  17.920000 20.945000  17.990000 ;
        RECT  0.500000  17.990000 20.875000  18.060000 ;
        RECT  0.500000  18.060000 20.805000  18.130000 ;
        RECT  0.500000  18.130000 20.735000  18.200000 ;
        RECT  0.500000  18.200000 20.665000  18.270000 ;
        RECT  0.500000  18.270000 20.595000  18.340000 ;
        RECT  0.500000  18.340000 20.525000  18.410000 ;
        RECT  0.500000  18.410000 20.455000  18.480000 ;
        RECT  0.500000  18.480000 20.385000  18.550000 ;
        RECT  0.500000  18.550000 20.315000  18.620000 ;
        RECT  0.500000  18.620000 20.245000  18.690000 ;
        RECT  0.500000  18.690000 20.175000  18.760000 ;
        RECT  0.500000  18.760000 20.105000  18.830000 ;
        RECT  0.500000  18.830000 20.035000  18.900000 ;
        RECT  0.500000  18.900000 19.965000  18.970000 ;
        RECT  0.500000  18.970000 19.895000  19.040000 ;
        RECT  0.500000  19.040000 19.825000  19.110000 ;
        RECT  0.500000  19.110000 19.755000  19.180000 ;
        RECT  0.500000  19.180000 19.685000  19.250000 ;
        RECT  0.500000  19.250000 19.615000  19.320000 ;
        RECT  0.500000  19.320000 19.545000  19.390000 ;
        RECT  0.500000  19.390000 19.475000  19.460000 ;
        RECT  0.500000  19.460000 19.405000  19.530000 ;
        RECT  0.500000  19.530000 19.335000  19.600000 ;
        RECT  0.500000  19.600000 19.265000  19.670000 ;
        RECT  0.500000  19.670000 19.195000  19.740000 ;
        RECT  0.500000  19.740000 19.125000  19.810000 ;
        RECT  0.500000  19.810000 19.055000  19.880000 ;
        RECT  0.500000  19.880000 18.985000  19.950000 ;
        RECT  0.500000  19.950000 18.915000  20.020000 ;
        RECT  0.500000  20.020000 18.845000  20.090000 ;
        RECT  0.500000  20.090000 18.775000  20.160000 ;
        RECT  0.500000  20.160000 18.705000  20.230000 ;
        RECT  0.500000  20.230000 18.635000  20.300000 ;
        RECT  0.500000  20.300000 18.565000  20.370000 ;
        RECT  0.500000  20.370000 18.495000  20.440000 ;
        RECT  0.500000  20.440000 18.425000  20.510000 ;
        RECT  0.500000  20.510000 18.355000  20.580000 ;
        RECT  0.500000  20.580000 18.285000  20.650000 ;
        RECT  0.500000  20.650000 18.215000  20.720000 ;
        RECT  0.500000  20.720000 18.145000  20.790000 ;
        RECT  0.500000  20.790000 18.075000  20.860000 ;
        RECT  0.500000  20.860000 18.005000  20.930000 ;
        RECT  0.500000  20.930000 17.935000  21.000000 ;
        RECT  0.500000  21.000000 17.865000  21.070000 ;
        RECT  0.500000  21.070000 17.795000  21.140000 ;
        RECT  0.500000  21.140000 17.725000  21.210000 ;
        RECT  0.500000  21.210000 17.655000  21.280000 ;
        RECT  0.500000  21.280000 17.585000  21.350000 ;
        RECT  0.500000  21.350000 17.515000  21.420000 ;
        RECT  0.500000  21.420000 17.445000  21.490000 ;
        RECT  0.500000  21.490000 17.375000  21.560000 ;
        RECT  0.500000  21.560000 17.305000  21.630000 ;
        RECT  0.500000  21.630000 17.235000  21.700000 ;
        RECT  0.500000  21.700000 17.165000  21.770000 ;
        RECT  0.500000  21.770000 17.095000  21.840000 ;
        RECT  0.500000  21.840000 17.025000  21.910000 ;
        RECT  0.500000  21.910000 16.955000  21.980000 ;
        RECT  0.500000  21.980000 16.885000  22.050000 ;
        RECT  0.500000  22.050000 16.815000  22.120000 ;
        RECT  0.500000  22.120000 16.745000  22.190000 ;
        RECT  0.500000  22.190000 16.675000  22.260000 ;
        RECT  0.500000  22.260000 16.605000  22.330000 ;
        RECT  0.500000  22.330000 16.535000  22.400000 ;
        RECT  0.500000  22.400000 16.465000  22.470000 ;
        RECT  0.500000  22.470000 16.395000  22.540000 ;
        RECT  0.500000  22.540000 16.325000  22.610000 ;
        RECT  0.500000  22.610000 16.255000  22.680000 ;
        RECT  0.500000  22.680000 16.185000  22.750000 ;
        RECT  0.500000  22.750000 16.115000  22.820000 ;
        RECT  0.500000  22.820000 16.045000  22.890000 ;
        RECT  0.500000  22.890000 15.975000  22.960000 ;
        RECT  0.500000  22.960000 15.905000  23.030000 ;
        RECT  0.500000  23.030000 15.835000  23.100000 ;
        RECT  0.500000  23.100000 15.765000  23.170000 ;
        RECT  0.500000  23.170000 15.695000  23.240000 ;
        RECT  0.500000  23.240000 15.625000  23.310000 ;
        RECT  0.500000  23.310000 15.555000  23.380000 ;
        RECT  0.500000  23.380000 15.485000  23.450000 ;
        RECT  0.500000  23.450000 15.415000  23.520000 ;
        RECT  0.500000  23.520000 15.345000  23.590000 ;
        RECT  0.500000  23.590000 15.275000  23.660000 ;
        RECT  0.500000  23.660000 15.205000  23.730000 ;
        RECT  0.500000  23.730000 15.135000  23.800000 ;
        RECT  0.500000  23.800000 15.065000  23.870000 ;
        RECT  0.500000  23.870000 14.995000  23.940000 ;
        RECT  0.500000  23.940000 14.925000  24.010000 ;
        RECT  0.500000  24.010000 14.855000  24.080000 ;
        RECT  0.500000  24.080000 14.785000  24.150000 ;
        RECT  0.500000  24.150000 14.715000  24.220000 ;
        RECT  0.500000  24.220000 14.645000  24.290000 ;
        RECT  0.500000  24.290000 14.575000  24.360000 ;
        RECT  0.500000  24.360000 14.505000  24.430000 ;
        RECT  0.500000  24.430000 14.435000  24.500000 ;
        RECT  0.500000  24.500000 14.365000  24.570000 ;
        RECT  0.500000  24.570000 14.295000  24.640000 ;
        RECT  0.500000  24.640000 14.225000  24.710000 ;
        RECT  0.500000  24.710000 14.155000  24.780000 ;
        RECT  0.500000  24.780000 14.085000  24.850000 ;
        RECT  0.500000  24.850000 14.015000  24.920000 ;
        RECT  0.500000  24.920000 13.945000  24.990000 ;
        RECT  0.500000  24.990000 13.875000  25.060000 ;
        RECT  0.500000  25.060000 13.805000  25.130000 ;
        RECT  0.500000  25.130000 13.750000  25.185000 ;
        RECT  0.500000  25.185000 13.750000  74.295000 ;
        RECT  0.500000  74.295000 13.750000  74.365000 ;
        RECT  0.500000  74.365000 13.820000  74.435000 ;
        RECT  0.500000  74.435000 13.890000  74.505000 ;
        RECT  0.500000  74.505000 13.960000 129.935000 ;
        RECT  0.500000 129.935000 13.960000 130.005000 ;
        RECT  0.500000 130.005000 14.030000 130.075000 ;
        RECT  0.500000 130.075000 14.100000 130.145000 ;
        RECT  0.500000 130.145000 14.170000 130.215000 ;
        RECT  0.500000 130.215000 14.240000 130.285000 ;
        RECT  0.500000 130.285000 14.310000 130.355000 ;
        RECT  0.500000 130.355000 14.380000 130.425000 ;
        RECT  0.500000 130.425000 14.450000 130.495000 ;
        RECT  0.500000 130.495000 14.520000 130.565000 ;
        RECT  0.500000 130.565000 14.590000 130.635000 ;
        RECT  0.500000 130.635000 14.660000 130.705000 ;
        RECT  0.500000 130.705000 14.730000 130.775000 ;
        RECT  0.500000 130.775000 14.800000 130.845000 ;
        RECT  0.500000 130.845000 14.870000 130.915000 ;
        RECT  0.500000 130.915000 14.940000 130.985000 ;
        RECT  0.500000 130.985000 68.010000 133.630000 ;
        RECT  0.500000 133.630000 14.940000 133.700000 ;
        RECT  0.500000 133.700000 14.870000 133.770000 ;
        RECT  0.500000 133.770000 14.800000 133.840000 ;
        RECT  0.500000 133.840000 14.730000 133.910000 ;
        RECT  0.500000 133.910000 14.660000 133.980000 ;
        RECT  0.500000 133.980000 14.590000 134.050000 ;
        RECT  0.500000 134.050000 14.520000 134.120000 ;
        RECT  0.500000 134.120000 14.450000 134.190000 ;
        RECT  0.500000 134.190000 14.380000 134.260000 ;
        RECT  0.500000 134.260000 14.310000 134.330000 ;
        RECT  0.500000 134.330000 14.240000 134.400000 ;
        RECT  0.500000 134.400000 14.170000 134.470000 ;
        RECT  0.500000 134.470000 14.100000 134.540000 ;
        RECT  0.500000 134.540000 14.030000 134.610000 ;
        RECT  0.500000 134.610000 13.960000 134.680000 ;
        RECT  0.500000 134.680000 13.960000 139.940000 ;
        RECT  0.500000 139.940000 13.960000 140.010000 ;
        RECT  0.500000 140.010000 14.030000 140.080000 ;
        RECT  0.500000 140.080000 14.100000 140.150000 ;
        RECT  0.500000 140.150000 14.170000 140.220000 ;
        RECT  0.500000 140.220000 14.240000 140.290000 ;
        RECT  0.500000 140.290000 14.310000 140.360000 ;
        RECT  0.500000 140.360000 14.380000 140.430000 ;
        RECT  0.500000 140.430000 14.450000 140.500000 ;
        RECT  0.500000 140.500000 14.520000 140.570000 ;
        RECT  0.500000 140.570000 14.590000 140.640000 ;
        RECT  0.500000 140.640000 14.660000 140.710000 ;
        RECT  0.500000 140.710000 14.730000 140.780000 ;
        RECT  0.500000 140.780000 14.800000 140.850000 ;
        RECT  0.500000 140.850000 14.870000 140.920000 ;
        RECT  0.500000 140.920000 14.940000 140.990000 ;
        RECT  0.500000 140.990000 68.010000 143.630000 ;
        RECT  0.500000 143.630000 14.940000 143.700000 ;
        RECT  0.500000 143.700000 14.870000 143.770000 ;
        RECT  0.500000 143.770000 14.800000 143.840000 ;
        RECT  0.500000 143.840000 14.730000 143.910000 ;
        RECT  0.500000 143.910000 14.660000 143.980000 ;
        RECT  0.500000 143.980000 14.590000 144.050000 ;
        RECT  0.500000 144.050000 14.520000 144.120000 ;
        RECT  0.500000 144.120000 14.450000 144.190000 ;
        RECT  0.500000 144.190000 14.380000 144.260000 ;
        RECT  0.500000 144.260000 14.310000 144.330000 ;
        RECT  0.500000 144.330000 14.240000 144.400000 ;
        RECT  0.500000 144.400000 14.170000 144.470000 ;
        RECT  0.500000 144.470000 14.100000 144.540000 ;
        RECT  0.500000 144.540000 14.030000 144.610000 ;
        RECT  0.500000 144.610000 13.960000 144.680000 ;
        RECT  0.500000 144.680000 13.960000 149.940000 ;
        RECT  0.500000 149.940000 13.960000 150.010000 ;
        RECT  0.500000 150.010000 14.030000 150.080000 ;
        RECT  0.500000 150.080000 14.100000 150.150000 ;
        RECT  0.500000 150.150000 14.170000 150.220000 ;
        RECT  0.500000 150.220000 14.240000 150.290000 ;
        RECT  0.500000 150.290000 14.310000 150.360000 ;
        RECT  0.500000 150.360000 14.380000 150.430000 ;
        RECT  0.500000 150.430000 14.450000 150.500000 ;
        RECT  0.500000 150.500000 14.520000 150.570000 ;
        RECT  0.500000 150.570000 14.590000 150.640000 ;
        RECT  0.500000 150.640000 14.660000 150.710000 ;
        RECT  0.500000 150.710000 14.730000 150.780000 ;
        RECT  0.500000 150.780000 14.800000 150.850000 ;
        RECT  0.500000 150.850000 14.870000 150.920000 ;
        RECT  0.500000 150.920000 14.940000 150.990000 ;
        RECT  0.500000 150.990000 68.010000 153.630000 ;
        RECT  0.500000 153.630000 14.940000 153.700000 ;
        RECT  0.500000 153.700000 14.870000 153.770000 ;
        RECT  0.500000 153.770000 14.800000 153.840000 ;
        RECT  0.500000 153.840000 14.730000 153.910000 ;
        RECT  0.500000 153.910000 14.660000 153.980000 ;
        RECT  0.500000 153.980000 14.590000 154.050000 ;
        RECT  0.500000 154.050000 14.520000 154.120000 ;
        RECT  0.500000 154.120000 14.450000 154.190000 ;
        RECT  0.500000 154.190000 14.380000 154.260000 ;
        RECT  0.500000 154.260000 14.310000 154.330000 ;
        RECT  0.500000 154.330000 14.240000 154.400000 ;
        RECT  0.500000 154.400000 14.170000 154.470000 ;
        RECT  0.500000 154.470000 14.100000 154.540000 ;
        RECT  0.500000 154.540000 14.030000 154.610000 ;
        RECT  0.500000 154.610000 13.960000 154.680000 ;
        RECT  0.500000 154.680000 13.960000 159.940000 ;
        RECT  0.500000 159.940000 13.960000 160.010000 ;
        RECT  0.500000 160.010000 14.030000 160.080000 ;
        RECT  0.500000 160.080000 14.100000 160.150000 ;
        RECT  0.500000 160.150000 14.170000 160.220000 ;
        RECT  0.500000 160.220000 14.240000 160.290000 ;
        RECT  0.500000 160.290000 14.310000 160.360000 ;
        RECT  0.500000 160.360000 14.380000 160.430000 ;
        RECT  0.500000 160.430000 14.450000 160.500000 ;
        RECT  0.500000 160.500000 14.520000 160.570000 ;
        RECT  0.500000 160.570000 14.590000 160.640000 ;
        RECT  0.500000 160.640000 14.660000 160.710000 ;
        RECT  0.500000 160.710000 14.730000 160.780000 ;
        RECT  0.500000 160.780000 14.800000 160.850000 ;
        RECT  0.500000 160.850000 14.870000 160.920000 ;
        RECT  0.500000 160.920000 14.940000 160.990000 ;
        RECT  0.500000 160.990000 68.010000 163.630000 ;
        RECT  0.500000 163.630000 14.940000 163.700000 ;
        RECT  0.500000 163.700000 14.870000 163.770000 ;
        RECT  0.500000 163.770000 14.800000 163.840000 ;
        RECT  0.500000 163.840000 14.730000 163.910000 ;
        RECT  0.500000 163.910000 14.660000 163.980000 ;
        RECT  0.500000 163.980000 14.590000 164.050000 ;
        RECT  0.500000 164.050000 14.520000 164.120000 ;
        RECT  0.500000 164.120000 14.450000 164.190000 ;
        RECT  0.500000 164.190000 14.380000 164.260000 ;
        RECT  0.500000 164.260000 14.310000 164.330000 ;
        RECT  0.500000 164.330000 14.240000 164.400000 ;
        RECT  0.500000 164.400000 14.170000 164.470000 ;
        RECT  0.500000 164.470000 14.100000 164.540000 ;
        RECT  0.500000 164.540000 14.030000 164.610000 ;
        RECT  0.500000 164.610000 13.960000 164.680000 ;
        RECT  0.500000 164.680000 13.960000 169.940000 ;
        RECT  0.500000 169.940000 13.960000 170.010000 ;
        RECT  0.500000 170.010000 14.030000 170.080000 ;
        RECT  0.500000 170.080000 14.100000 170.150000 ;
        RECT  0.500000 170.150000 14.170000 170.220000 ;
        RECT  0.500000 170.220000 14.240000 170.290000 ;
        RECT  0.500000 170.290000 14.310000 170.360000 ;
        RECT  0.500000 170.360000 14.380000 170.430000 ;
        RECT  0.500000 170.430000 14.450000 170.500000 ;
        RECT  0.500000 170.500000 14.520000 170.570000 ;
        RECT  0.500000 170.570000 14.590000 170.640000 ;
        RECT  0.500000 170.640000 14.660000 170.710000 ;
        RECT  0.500000 170.710000 14.730000 170.780000 ;
        RECT  0.500000 170.780000 14.800000 170.850000 ;
        RECT  0.500000 170.850000 14.870000 170.920000 ;
        RECT  0.500000 170.920000 14.940000 170.990000 ;
        RECT  0.500000 170.990000 68.010000 173.630000 ;
        RECT  0.500000 173.630000 14.940000 173.700000 ;
        RECT  0.500000 173.700000 14.870000 173.770000 ;
        RECT  0.500000 173.770000 14.800000 173.840000 ;
        RECT  0.500000 173.840000 14.730000 173.910000 ;
        RECT  0.500000 173.910000 14.660000 173.980000 ;
        RECT  0.500000 173.980000 14.590000 174.050000 ;
        RECT  0.500000 174.050000 14.520000 174.120000 ;
        RECT  0.500000 174.120000 14.450000 174.190000 ;
        RECT  0.500000 174.190000 14.380000 174.260000 ;
        RECT  0.500000 174.260000 14.310000 174.330000 ;
        RECT  0.500000 174.330000 14.240000 174.400000 ;
        RECT  0.500000 174.400000 14.170000 174.470000 ;
        RECT  0.500000 174.470000 14.100000 174.540000 ;
        RECT  0.500000 174.540000 14.030000 174.610000 ;
        RECT  0.500000 174.610000 13.960000 174.680000 ;
        RECT  0.500000 174.680000 13.960000 179.940000 ;
        RECT  0.500000 179.940000 13.960000 180.010000 ;
        RECT  0.500000 180.010000 14.030000 180.080000 ;
        RECT  0.500000 180.080000 14.100000 180.150000 ;
        RECT  0.500000 180.150000 14.170000 180.220000 ;
        RECT  0.500000 180.220000 14.240000 180.290000 ;
        RECT  0.500000 180.290000 14.310000 180.360000 ;
        RECT  0.500000 180.360000 14.380000 180.430000 ;
        RECT  0.500000 180.430000 14.450000 180.500000 ;
        RECT  0.500000 180.500000 14.520000 180.570000 ;
        RECT  0.500000 180.570000 14.590000 180.640000 ;
        RECT  0.500000 180.640000 14.660000 180.710000 ;
        RECT  0.500000 180.710000 14.730000 180.780000 ;
        RECT  0.500000 180.780000 14.800000 180.850000 ;
        RECT  0.500000 180.850000 14.870000 180.920000 ;
        RECT  0.500000 180.920000 14.940000 180.990000 ;
        RECT  0.500000 180.990000 68.010000 183.630000 ;
        RECT  0.500000 183.630000 14.940000 183.700000 ;
        RECT  0.500000 183.700000 14.870000 183.770000 ;
        RECT  0.500000 183.770000 14.800000 183.840000 ;
        RECT  0.500000 183.840000 14.730000 183.910000 ;
        RECT  0.500000 183.910000 14.660000 183.980000 ;
        RECT  0.500000 183.980000 14.590000 184.050000 ;
        RECT  0.500000 184.050000 14.520000 184.120000 ;
        RECT  0.500000 184.120000 14.450000 184.190000 ;
        RECT  0.500000 184.190000 14.380000 184.260000 ;
        RECT  0.500000 184.260000 14.310000 184.330000 ;
        RECT  0.500000 184.330000 14.240000 184.400000 ;
        RECT  0.500000 184.400000 14.170000 184.470000 ;
        RECT  0.500000 184.470000 14.100000 184.540000 ;
        RECT  0.500000 184.540000 14.030000 184.610000 ;
        RECT  0.500000 184.610000 13.960000 184.680000 ;
        RECT  0.500000 184.680000 13.960000 189.940000 ;
        RECT  0.500000 189.940000 13.960000 190.010000 ;
        RECT  0.500000 190.010000 14.030000 190.080000 ;
        RECT  0.500000 190.080000 14.100000 190.150000 ;
        RECT  0.500000 190.150000 14.170000 190.220000 ;
        RECT  0.500000 190.220000 14.240000 190.290000 ;
        RECT  0.500000 190.290000 14.310000 190.360000 ;
        RECT  0.500000 190.360000 14.380000 190.430000 ;
        RECT  0.500000 190.430000 14.450000 190.500000 ;
        RECT  0.500000 190.500000 14.520000 190.570000 ;
        RECT  0.500000 190.570000 14.590000 190.640000 ;
        RECT  0.500000 190.640000 14.660000 190.710000 ;
        RECT  0.500000 190.710000 14.730000 190.780000 ;
        RECT  0.500000 190.780000 14.800000 190.850000 ;
        RECT  0.500000 190.850000 14.870000 190.920000 ;
        RECT  0.500000 190.920000 14.940000 190.990000 ;
        RECT  0.500000 190.990000 68.010000 193.630000 ;
        RECT 11.635000  10.210000 55.595000  10.215000 ;
        RECT 11.695000   7.655000 16.860000   7.725000 ;
        RECT 11.700000  10.145000 55.595000  10.210000 ;
        RECT 11.765000   7.725000 16.860000   7.795000 ;
        RECT 11.765000  10.080000 55.595000  10.145000 ;
        RECT 11.805000  10.040000 17.535000  10.080000 ;
        RECT 11.835000   7.795000 16.860000   7.865000 ;
        RECT 11.875000   9.970000 17.465000  10.040000 ;
        RECT 11.905000   7.865000 16.860000   7.935000 ;
        RECT 11.945000   9.900000 17.395000   9.970000 ;
        RECT 11.975000   7.935000 16.860000   8.005000 ;
        RECT 12.015000   8.005000 16.860000   8.045000 ;
        RECT 12.015000   8.045000 16.860000   9.365000 ;
        RECT 12.015000   9.365000 16.860000   9.435000 ;
        RECT 12.015000   9.435000 16.930000   9.505000 ;
        RECT 12.015000   9.505000 17.000000   9.575000 ;
        RECT 12.015000   9.575000 17.070000   9.645000 ;
        RECT 12.015000   9.645000 17.140000   9.715000 ;
        RECT 12.015000   9.715000 17.210000   9.785000 ;
        RECT 12.015000   9.785000 17.280000   9.830000 ;
        RECT 12.015000   9.830000 17.325000   9.900000 ;
    END
  END SRC_BDY_LVC1
  PIN SRC_BDY_LVC2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 16.135000 31.010000 74.700000 33.650000 ;
        RECT 16.135000 40.990000 74.700000 43.630000 ;
        RECT 16.135000 51.010000 74.700000 53.650000 ;
        RECT 16.135000 60.990000 74.700000 63.630000 ;
        RECT 16.135000 70.990000 74.700000 73.630000 ;
        RECT 54.095000  0.000000 74.700000  7.815000 ;
        RECT 54.095000 19.990000 74.700000 21.695000 ;
        RECT 54.150000 19.935000 74.700000 19.990000 ;
        RECT 54.165000  7.815000 74.700000  7.885000 ;
        RECT 54.220000 19.865000 74.700000 19.935000 ;
        RECT 54.235000  7.885000 74.700000  7.955000 ;
        RECT 54.290000 19.795000 74.700000 19.865000 ;
        RECT 54.305000  7.955000 74.700000  8.025000 ;
        RECT 54.360000 19.725000 74.700000 19.795000 ;
        RECT 54.375000  8.025000 74.700000  8.095000 ;
        RECT 54.430000 19.655000 74.700000 19.725000 ;
        RECT 54.445000  8.095000 74.700000  8.165000 ;
        RECT 54.500000 19.585000 74.700000 19.655000 ;
        RECT 54.515000  8.165000 74.700000  8.235000 ;
        RECT 54.570000 19.515000 74.700000 19.585000 ;
        RECT 54.585000  8.235000 74.700000  8.305000 ;
        RECT 54.640000 19.445000 74.700000 19.515000 ;
        RECT 54.655000  8.305000 74.700000  8.375000 ;
        RECT 54.710000 19.375000 74.700000 19.445000 ;
        RECT 54.725000  8.375000 74.700000  8.445000 ;
        RECT 54.780000 19.305000 74.700000 19.375000 ;
        RECT 54.795000  8.445000 74.700000  8.515000 ;
        RECT 54.850000 19.235000 74.700000 19.305000 ;
        RECT 54.865000  8.515000 74.700000  8.585000 ;
        RECT 54.920000 19.165000 74.700000 19.235000 ;
        RECT 54.935000  8.585000 74.700000  8.655000 ;
        RECT 54.990000 19.095000 74.700000 19.165000 ;
        RECT 55.005000  8.655000 74.700000  8.725000 ;
        RECT 55.060000 19.025000 74.700000 19.095000 ;
        RECT 55.075000  8.725000 74.700000  8.795000 ;
        RECT 55.130000 18.955000 74.700000 19.025000 ;
        RECT 55.145000  8.795000 74.700000  8.865000 ;
        RECT 55.200000 18.885000 74.700000 18.955000 ;
        RECT 55.215000  8.865000 74.700000  8.935000 ;
        RECT 55.270000 18.815000 74.700000 18.885000 ;
        RECT 55.285000  8.935000 74.700000  9.005000 ;
        RECT 55.340000 18.745000 74.700000 18.815000 ;
        RECT 55.355000  9.005000 74.700000  9.075000 ;
        RECT 55.410000 18.675000 74.700000 18.745000 ;
        RECT 55.425000  9.075000 74.700000  9.145000 ;
        RECT 55.480000 18.605000 74.700000 18.675000 ;
        RECT 55.495000  9.145000 74.700000  9.215000 ;
        RECT 55.550000 18.535000 74.700000 18.605000 ;
        RECT 55.565000  9.215000 74.700000  9.285000 ;
        RECT 55.620000 18.465000 74.700000 18.535000 ;
        RECT 55.635000  9.285000 74.700000  9.355000 ;
        RECT 55.690000 18.395000 74.700000 18.465000 ;
        RECT 55.705000  9.355000 74.700000  9.425000 ;
        RECT 55.760000 18.325000 74.700000 18.395000 ;
        RECT 55.775000  9.425000 74.700000  9.495000 ;
        RECT 55.830000 18.255000 74.700000 18.325000 ;
        RECT 55.845000  9.495000 74.700000  9.565000 ;
        RECT 55.900000 18.185000 74.700000 18.255000 ;
        RECT 55.915000  9.565000 74.700000  9.635000 ;
        RECT 55.970000 18.115000 74.700000 18.185000 ;
        RECT 55.985000  9.635000 74.700000  9.705000 ;
        RECT 56.040000 18.045000 74.700000 18.115000 ;
        RECT 56.055000  9.705000 74.700000  9.775000 ;
        RECT 56.110000 17.975000 74.700000 18.045000 ;
        RECT 56.125000  9.775000 74.700000  9.845000 ;
        RECT 56.180000 17.905000 74.700000 17.975000 ;
        RECT 56.195000  9.845000 74.700000  9.915000 ;
        RECT 56.250000  9.915000 74.700000  9.970000 ;
        RECT 56.250000  9.970000 74.700000 17.835000 ;
        RECT 56.250000 17.835000 74.700000 17.905000 ;
        RECT 62.325000 21.695000 74.700000 21.765000 ;
        RECT 62.395000 21.765000 74.700000 21.835000 ;
        RECT 62.465000 21.835000 74.700000 21.905000 ;
        RECT 62.535000 21.905000 74.700000 21.975000 ;
        RECT 62.605000 21.975000 74.700000 22.045000 ;
        RECT 62.675000 22.045000 74.700000 22.115000 ;
        RECT 62.745000 22.115000 74.700000 22.185000 ;
        RECT 62.815000 22.185000 74.700000 22.255000 ;
        RECT 62.885000 22.255000 74.700000 22.325000 ;
        RECT 62.955000 22.325000 74.700000 22.395000 ;
        RECT 63.025000 22.395000 74.700000 22.465000 ;
        RECT 63.095000 22.465000 74.700000 22.535000 ;
        RECT 63.165000 22.535000 74.700000 22.605000 ;
        RECT 63.235000 22.605000 74.700000 22.675000 ;
        RECT 63.305000 22.675000 74.700000 22.745000 ;
        RECT 63.375000 22.745000 74.700000 22.815000 ;
        RECT 63.445000 22.815000 74.700000 22.885000 ;
        RECT 63.515000 22.885000 74.700000 22.955000 ;
        RECT 63.585000 22.955000 74.700000 23.025000 ;
        RECT 63.655000 23.025000 74.700000 23.095000 ;
        RECT 63.725000 23.095000 74.700000 23.165000 ;
        RECT 63.795000 23.165000 74.700000 23.235000 ;
        RECT 63.865000 23.235000 74.700000 23.305000 ;
        RECT 63.935000 23.305000 74.700000 23.375000 ;
        RECT 64.005000 23.375000 74.700000 23.445000 ;
        RECT 64.075000 23.445000 74.700000 23.515000 ;
        RECT 64.145000 23.515000 74.700000 23.585000 ;
        RECT 64.215000 23.585000 74.700000 23.655000 ;
        RECT 64.285000 23.655000 74.700000 23.725000 ;
        RECT 64.355000 23.725000 74.700000 23.795000 ;
        RECT 64.425000 23.795000 74.700000 23.865000 ;
        RECT 64.495000 23.865000 74.700000 23.935000 ;
        RECT 64.565000 23.935000 74.700000 24.005000 ;
        RECT 64.635000 24.005000 74.700000 24.075000 ;
        RECT 64.705000 24.075000 74.700000 24.145000 ;
        RECT 64.775000 24.145000 74.700000 24.215000 ;
        RECT 64.845000 24.215000 74.700000 24.285000 ;
        RECT 64.880000 31.000000 74.700000 31.010000 ;
        RECT 64.915000 24.285000 74.700000 24.355000 ;
        RECT 64.950000 30.930000 74.700000 31.000000 ;
        RECT 64.950000 40.985000 74.700000 40.990000 ;
        RECT 64.950000 51.005000 74.700000 51.010000 ;
        RECT 64.985000 24.355000 74.700000 24.425000 ;
        RECT 65.015000 60.920000 74.700000 60.990000 ;
        RECT 65.015000 63.630000 74.700000 63.700000 ;
        RECT 65.015000 70.920000 74.700000 70.990000 ;
        RECT 65.020000 30.860000 74.700000 30.930000 ;
        RECT 65.020000 40.915000 74.700000 40.985000 ;
        RECT 65.020000 50.935000 74.700000 51.005000 ;
        RECT 65.030000 33.650000 74.700000 33.720000 ;
        RECT 65.030000 43.630000 74.700000 43.700000 ;
        RECT 65.030000 53.650000 74.700000 53.720000 ;
        RECT 65.055000 24.425000 74.700000 24.495000 ;
        RECT 65.085000 60.850000 74.700000 60.920000 ;
        RECT 65.085000 63.700000 74.700000 63.770000 ;
        RECT 65.085000 70.850000 74.700000 70.920000 ;
        RECT 65.090000 30.790000 74.700000 30.860000 ;
        RECT 65.090000 40.845000 74.700000 40.915000 ;
        RECT 65.090000 50.865000 74.700000 50.935000 ;
        RECT 65.100000 33.720000 74.700000 33.790000 ;
        RECT 65.100000 43.700000 74.700000 43.770000 ;
        RECT 65.100000 53.720000 74.700000 53.790000 ;
        RECT 65.125000 24.495000 74.700000 24.565000 ;
        RECT 65.155000 60.780000 74.700000 60.850000 ;
        RECT 65.155000 63.770000 74.700000 63.840000 ;
        RECT 65.155000 70.780000 74.700000 70.850000 ;
        RECT 65.160000 30.720000 74.700000 30.790000 ;
        RECT 65.160000 40.775000 74.700000 40.845000 ;
        RECT 65.160000 50.795000 74.700000 50.865000 ;
        RECT 65.170000 33.790000 74.700000 33.860000 ;
        RECT 65.170000 43.770000 74.700000 43.840000 ;
        RECT 65.170000 53.790000 74.700000 53.860000 ;
        RECT 65.195000 24.565000 74.700000 24.635000 ;
        RECT 65.225000 60.710000 74.700000 60.780000 ;
        RECT 65.225000 63.840000 74.700000 63.910000 ;
        RECT 65.225000 70.710000 74.700000 70.780000 ;
        RECT 65.230000 30.650000 74.700000 30.720000 ;
        RECT 65.230000 40.705000 74.700000 40.775000 ;
        RECT 65.230000 50.725000 74.700000 50.795000 ;
        RECT 65.240000 33.860000 74.700000 33.930000 ;
        RECT 65.240000 43.840000 74.700000 43.910000 ;
        RECT 65.240000 53.860000 74.700000 53.930000 ;
        RECT 65.265000 24.635000 74.700000 24.705000 ;
        RECT 65.270000 73.630000 68.740000 73.700000 ;
        RECT 65.295000 60.640000 74.700000 60.710000 ;
        RECT 65.295000 63.910000 74.700000 63.980000 ;
        RECT 65.295000 70.640000 74.700000 70.710000 ;
        RECT 65.300000 30.580000 74.700000 30.650000 ;
        RECT 65.300000 40.635000 74.700000 40.705000 ;
        RECT 65.300000 50.655000 74.700000 50.725000 ;
        RECT 65.310000 33.930000 74.700000 34.000000 ;
        RECT 65.310000 43.910000 74.700000 43.980000 ;
        RECT 65.310000 53.930000 74.700000 54.000000 ;
        RECT 65.335000 24.705000 74.700000 24.775000 ;
        RECT 65.340000 73.700000 68.670000 73.770000 ;
        RECT 65.365000 60.570000 74.700000 60.640000 ;
        RECT 65.365000 63.980000 74.700000 64.050000 ;
        RECT 65.365000 70.570000 74.700000 70.640000 ;
        RECT 65.370000 30.510000 74.700000 30.580000 ;
        RECT 65.370000 40.565000 74.700000 40.635000 ;
        RECT 65.370000 50.585000 74.700000 50.655000 ;
        RECT 65.380000 34.000000 74.700000 34.070000 ;
        RECT 65.380000 43.980000 74.700000 44.050000 ;
        RECT 65.380000 54.000000 74.700000 54.070000 ;
        RECT 65.405000 24.775000 74.700000 24.845000 ;
        RECT 65.410000 73.770000 68.600000 73.840000 ;
        RECT 65.435000 60.500000 74.700000 60.570000 ;
        RECT 65.435000 64.050000 74.700000 64.120000 ;
        RECT 65.435000 70.500000 74.700000 70.570000 ;
        RECT 65.440000 30.440000 74.700000 30.510000 ;
        RECT 65.440000 40.495000 74.700000 40.565000 ;
        RECT 65.440000 50.515000 74.700000 50.585000 ;
        RECT 65.450000 34.070000 74.700000 34.140000 ;
        RECT 65.450000 44.050000 74.700000 44.120000 ;
        RECT 65.450000 54.070000 74.700000 54.140000 ;
        RECT 65.475000 24.845000 74.700000 24.915000 ;
        RECT 65.480000 73.840000 68.530000 73.910000 ;
        RECT 65.505000 60.430000 74.700000 60.500000 ;
        RECT 65.505000 64.120000 74.700000 64.190000 ;
        RECT 65.505000 70.430000 74.700000 70.500000 ;
        RECT 65.510000 30.370000 74.700000 30.440000 ;
        RECT 65.510000 40.425000 74.700000 40.495000 ;
        RECT 65.510000 50.445000 74.700000 50.515000 ;
        RECT 65.520000 34.140000 74.700000 34.210000 ;
        RECT 65.520000 44.120000 74.700000 44.190000 ;
        RECT 65.520000 54.140000 74.700000 54.210000 ;
        RECT 65.545000 24.915000 74.700000 24.985000 ;
        RECT 65.550000 73.910000 68.460000 73.980000 ;
        RECT 65.575000 60.360000 74.700000 60.430000 ;
        RECT 65.575000 64.190000 74.700000 64.260000 ;
        RECT 65.575000 70.360000 74.700000 70.430000 ;
        RECT 65.580000 30.300000 74.700000 30.370000 ;
        RECT 65.580000 40.355000 74.700000 40.425000 ;
        RECT 65.580000 50.375000 74.700000 50.445000 ;
        RECT 65.590000 34.210000 74.700000 34.280000 ;
        RECT 65.590000 44.190000 74.700000 44.260000 ;
        RECT 65.590000 54.210000 74.700000 54.280000 ;
        RECT 65.615000 24.985000 74.700000 25.055000 ;
        RECT 65.620000 73.980000 68.390000 74.050000 ;
        RECT 65.645000 60.290000 74.700000 60.360000 ;
        RECT 65.645000 64.260000 74.700000 64.330000 ;
        RECT 65.645000 70.290000 74.700000 70.360000 ;
        RECT 65.650000 30.230000 74.700000 30.300000 ;
        RECT 65.650000 40.285000 74.700000 40.355000 ;
        RECT 65.650000 50.305000 74.700000 50.375000 ;
        RECT 65.660000 34.280000 74.700000 34.350000 ;
        RECT 65.660000 44.260000 74.700000 44.330000 ;
        RECT 65.660000 54.280000 74.700000 54.350000 ;
        RECT 65.685000 25.055000 74.700000 25.125000 ;
        RECT 65.690000 74.050000 68.320000 74.120000 ;
        RECT 65.715000 60.220000 74.700000 60.290000 ;
        RECT 65.715000 64.330000 74.700000 64.400000 ;
        RECT 65.715000 70.220000 74.700000 70.290000 ;
        RECT 65.720000 30.160000 74.700000 30.230000 ;
        RECT 65.720000 40.215000 74.700000 40.285000 ;
        RECT 65.720000 50.235000 74.700000 50.305000 ;
        RECT 65.730000 34.350000 74.700000 34.420000 ;
        RECT 65.730000 44.330000 74.700000 44.400000 ;
        RECT 65.730000 54.350000 74.700000 54.420000 ;
        RECT 65.755000 25.125000 74.700000 25.195000 ;
        RECT 65.760000 74.120000 68.250000 74.190000 ;
        RECT 65.785000 60.150000 74.700000 60.220000 ;
        RECT 65.785000 64.400000 74.700000 64.470000 ;
        RECT 65.785000 70.150000 74.700000 70.220000 ;
        RECT 65.790000 30.090000 74.700000 30.160000 ;
        RECT 65.790000 40.145000 74.700000 40.215000 ;
        RECT 65.790000 50.165000 74.700000 50.235000 ;
        RECT 65.800000 34.420000 74.700000 34.490000 ;
        RECT 65.800000 44.400000 74.700000 44.470000 ;
        RECT 65.800000 54.420000 74.700000 54.490000 ;
        RECT 65.825000 25.195000 74.700000 25.265000 ;
        RECT 65.830000 74.190000 68.180000 74.260000 ;
        RECT 65.855000 60.080000 74.700000 60.150000 ;
        RECT 65.855000 64.470000 74.700000 64.540000 ;
        RECT 65.855000 70.080000 74.700000 70.150000 ;
        RECT 65.860000 30.020000 74.700000 30.090000 ;
        RECT 65.860000 40.075000 74.700000 40.145000 ;
        RECT 65.860000 50.095000 74.700000 50.165000 ;
        RECT 65.870000 34.490000 74.700000 34.560000 ;
        RECT 65.870000 44.470000 74.700000 44.540000 ;
        RECT 65.870000 54.490000 74.700000 54.560000 ;
        RECT 65.895000 25.265000 74.700000 25.335000 ;
        RECT 65.900000 74.260000 68.110000 74.330000 ;
        RECT 65.925000 60.010000 74.700000 60.080000 ;
        RECT 65.925000 64.540000 74.700000 64.610000 ;
        RECT 65.925000 70.010000 74.700000 70.080000 ;
        RECT 65.930000 29.950000 74.700000 30.020000 ;
        RECT 65.930000 40.005000 74.700000 40.075000 ;
        RECT 65.930000 50.025000 74.700000 50.095000 ;
        RECT 65.940000 34.560000 74.700000 34.630000 ;
        RECT 65.940000 44.540000 74.700000 44.610000 ;
        RECT 65.940000 54.560000 74.700000 54.630000 ;
        RECT 65.965000 25.335000 74.700000 25.405000 ;
        RECT 65.970000 74.330000 68.040000 74.400000 ;
        RECT 65.995000 54.630000 74.700000 54.685000 ;
        RECT 65.995000 54.685000 74.700000 59.940000 ;
        RECT 65.995000 59.940000 74.700000 60.010000 ;
        RECT 65.995000 64.610000 74.700000 64.680000 ;
        RECT 65.995000 64.680000 74.700000 69.940000 ;
        RECT 65.995000 69.940000 74.700000 70.010000 ;
        RECT 66.000000 25.405000 74.700000 25.440000 ;
        RECT 66.000000 25.440000 74.700000 29.880000 ;
        RECT 66.000000 29.880000 74.700000 29.950000 ;
        RECT 66.000000 34.630000 74.700000 34.690000 ;
        RECT 66.000000 34.690000 74.700000 39.935000 ;
        RECT 66.000000 39.935000 74.700000 40.005000 ;
        RECT 66.000000 44.610000 74.700000 44.670000 ;
        RECT 66.000000 44.670000 74.700000 49.955000 ;
        RECT 66.000000 49.955000 74.700000 50.025000 ;
        RECT 66.000000 74.400000 68.010000 74.430000 ;
        RECT 66.000000 74.430000 68.010000 98.560000 ;
    END
  END SRC_BDY_LVC2
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 6.885000 1.270000 11.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 6.885000 75.000000 11.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 6.985000 1.270000 11.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 0.035000 1.270000 5.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 0.035000 75.000000 5.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 0.135000 1.270000 5.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 12.935000 0.965000 16.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 12.935000 75.000000 16.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 13.035000 0.965000 16.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 17.785000 1.270000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 68.035000 1.270000 93.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 17.785000 75.000000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 68.035000 75.000000 93.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 17.885000 1.270000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 68.035000 1.270000 92.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 17.885000 75.000000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 62.085000 1.270000 66.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 62.085000 75.000000 66.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 62.185000 1.270000 66.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 34.735000 1.270000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 45.735000 1.270000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 49.645000 1.270000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 54.405000 1.270000 54.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 34.735000 75.000000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 45.735000 75.000000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 49.645000 75.000000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 54.405000 75.000000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 34.840000 1.270000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 45.735000 1.270000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 34.840000 75.000000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 39.585000 1.270000 44.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 39.585000 75.000000 44.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 39.685000 1.270000 44.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 23.835000 1.270000 28.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 23.835000 75.000000 28.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 23.935000 1.270000 28.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 56.235000 1.270000 60.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.235000 75.000000 60.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 56.335000 1.270000 60.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 29.885000 1.270000 33.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 29.885000 75.000000 33.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 29.985000 1.270000 33.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT  0.240000  17.210000  2.995000  19.200000 ;
      RECT  1.350000   1.020000  7.110000   1.190000 ;
      RECT  1.350000   1.190000  1.520000  17.040000 ;
      RECT  1.350000  17.040000  7.110000  17.210000 ;
      RECT  1.760000  19.630000  9.385000  20.140000 ;
      RECT  1.760000  20.140000  2.685000  23.060000 ;
      RECT  1.845000   3.220000  2.015000   8.960000 ;
      RECT  1.845000   9.710000  2.015000  16.610000 ;
      RECT  2.070000   1.610000  6.390000   1.780000 ;
      RECT  2.070000   9.260000  6.390000   9.430000 ;
      RECT  2.305000   2.490000  2.475000   8.960000 ;
      RECT  2.305000  10.140000  2.475000  15.440000 ;
      RECT  2.765000   3.220000  2.935000   8.960000 ;
      RECT  2.765000   9.710000  2.935000  16.610000 ;
      RECT  3.225000   2.490000  3.395000   8.960000 ;
      RECT  3.225000  10.140000  3.395000  15.440000 ;
      RECT  3.685000   3.220000  3.855000   8.960000 ;
      RECT  3.685000   9.710000  3.855000  16.610000 ;
      RECT  4.145000   2.490000  4.315000   8.960000 ;
      RECT  4.145000  10.140000  4.315000  15.440000 ;
      RECT  4.605000   3.220000  4.775000   8.960000 ;
      RECT  4.605000   9.710000  4.775000  16.610000 ;
      RECT  4.975000  22.290000 10.650000  23.010000 ;
      RECT  5.065000   2.490000  5.235000   8.960000 ;
      RECT  5.065000  10.140000  5.235000  15.440000 ;
      RECT  5.525000   3.220000  5.695000   8.960000 ;
      RECT  5.525000   9.710000  5.695000  16.610000 ;
      RECT  5.890000  23.010000 10.650000  23.015000 ;
      RECT  5.985000   2.490000  6.155000   8.960000 ;
      RECT  5.985000  10.140000  6.155000  15.440000 ;
      RECT  6.445000   2.060000  6.615000   8.960000 ;
      RECT  6.445000   9.710000  6.615000  16.610000 ;
      RECT  6.940000   1.190000  7.110000  17.040000 ;
      RECT  8.340000 196.360000  8.670000 196.420000 ;
      RECT  8.345000   1.410000 16.655000  18.350000 ;
      RECT  8.420000 195.890000  8.590000 196.360000 ;
      RECT  9.155000 106.965000 10.280000 196.850000 ;
      RECT  9.155000 196.850000 69.720000 197.380000 ;
      RECT  9.185000  23.825000 69.720000  24.355000 ;
      RECT  9.185000  24.355000 10.280000  82.980000 ;
      RECT  9.185000  82.980000 21.740000  83.150000 ;
      RECT  9.185000  83.150000 10.280000  99.490000 ;
      RECT  9.730000  99.490000 10.280000 106.965000 ;
      RECT 10.920000  83.820000 11.830000  84.585000 ;
      RECT 11.065000 168.280000 12.220000 194.935000 ;
      RECT 11.065000 194.935000 68.495000 195.885000 ;
      RECT 11.095000 144.465000 21.490000 145.315000 ;
      RECT 11.095000 145.315000 12.220000 168.280000 ;
      RECT 11.275000  25.065000 68.140000  26.015000 ;
      RECT 11.275000  26.015000 12.220000  34.040000 ;
      RECT 11.275000  36.745000 12.220000  43.620000 ;
      RECT 11.275000  46.905000 12.220000  81.575000 ;
      RECT 11.275000  81.575000 23.280000  82.085000 ;
      RECT 11.370000  34.040000 12.220000  36.745000 ;
      RECT 11.370000  43.620000 12.220000  46.905000 ;
      RECT 12.405000 184.140000 66.575000 186.620000 ;
      RECT 12.430000 184.100000 66.575000 184.140000 ;
      RECT 12.750000  75.785000 12.920000  80.300000 ;
      RECT 12.975000  81.045000 66.655000  81.215000 ;
      RECT 13.060000  44.100000 65.590000  46.620000 ;
      RECT 13.060000  64.100000 65.590000  66.620000 ;
      RECT 13.190000  34.100000 65.590000  36.620000 ;
      RECT 13.190000  54.100000 65.590000  56.620000 ;
      RECT 13.335000 174.100000 65.590000 176.620000 ;
      RECT 13.365000 145.615000 14.305000 145.620000 ;
      RECT 13.365000 145.620000 65.590000 146.620000 ;
      RECT 13.365000 154.100000 65.590000 156.620000 ;
      RECT 13.365000 164.100000 65.590000 166.620000 ;
      RECT 13.395000  26.900000 13.925000  33.570000 ;
      RECT 13.395000  36.900000 13.925000  43.570000 ;
      RECT 13.395000  46.900000 13.925000  53.570000 ;
      RECT 13.395000  56.900000 13.925000  63.570000 ;
      RECT 13.395000  66.900000 13.925000  71.725000 ;
      RECT 13.395000 186.900000 13.925000 193.570000 ;
      RECT 14.360000 194.100000 65.590000 194.270000 ;
      RECT 14.780000  26.900000 15.310000  33.570000 ;
      RECT 14.780000  36.900000 15.310000  43.570000 ;
      RECT 14.780000  46.900000 15.310000  53.570000 ;
      RECT 14.780000  56.900000 15.310000  63.570000 ;
      RECT 14.780000  66.900000 15.310000  71.725000 ;
      RECT 14.780000 186.900000 15.310000 193.570000 ;
      RECT 14.790000  26.840000 15.300000  26.900000 ;
      RECT 14.790000  33.570000 15.300000  33.630000 ;
      RECT 14.790000  36.840000 15.300000  36.900000 ;
      RECT 14.790000  43.570000 15.300000  43.630000 ;
      RECT 14.790000  46.840000 15.300000  46.900000 ;
      RECT 14.790000  53.570000 15.300000  53.630000 ;
      RECT 14.790000  56.840000 15.300000  56.900000 ;
      RECT 14.790000  63.570000 15.300000  63.630000 ;
      RECT 14.790000  66.840000 15.300000  66.900000 ;
      RECT 14.790000 186.840000 15.300000 186.900000 ;
      RECT 14.790000 193.570000 15.300000 193.630000 ;
      RECT 15.865000 146.900000 16.395000 153.570000 ;
      RECT 15.865000 156.900000 16.395000 163.570000 ;
      RECT 15.865000 166.900000 16.395000 173.570000 ;
      RECT 16.165000  26.900000 16.695000  33.570000 ;
      RECT 16.165000  36.900000 16.695000  43.570000 ;
      RECT 16.165000  46.900000 16.695000  53.570000 ;
      RECT 16.165000  56.900000 16.695000  63.570000 ;
      RECT 16.165000  66.900000 16.695000  71.725000 ;
      RECT 16.165000 176.900000 16.695000 183.570000 ;
      RECT 16.165000 186.900000 16.695000 193.570000 ;
      RECT 17.000000  17.580000 56.200000  18.350000 ;
      RECT 17.030000  75.785000 17.200000  80.300000 ;
      RECT 17.550000  26.900000 18.080000  33.570000 ;
      RECT 17.550000  36.900000 18.080000  43.570000 ;
      RECT 17.550000  46.900000 18.080000  53.570000 ;
      RECT 17.550000  56.900000 18.080000  63.570000 ;
      RECT 17.550000  66.900000 18.080000  71.725000 ;
      RECT 17.550000 176.900000 18.080000 183.570000 ;
      RECT 17.550000 186.900000 18.080000 193.570000 ;
      RECT 17.560000  26.840000 18.070000  26.900000 ;
      RECT 17.560000  33.570000 18.070000  33.630000 ;
      RECT 17.560000  36.840000 18.070000  36.900000 ;
      RECT 17.560000  43.570000 18.070000  43.630000 ;
      RECT 17.560000  46.840000 18.070000  46.900000 ;
      RECT 17.560000  53.570000 18.070000  53.630000 ;
      RECT 17.560000  56.840000 18.070000  56.900000 ;
      RECT 17.560000  63.570000 18.070000  63.630000 ;
      RECT 17.560000  66.840000 18.070000  66.900000 ;
      RECT 17.560000 176.840000 18.070000 176.900000 ;
      RECT 17.560000 183.570000 18.070000 183.630000 ;
      RECT 17.560000 186.840000 18.070000 186.900000 ;
      RECT 17.560000 193.570000 18.070000 193.630000 ;
      RECT 17.955000 146.900000 18.485000 153.570000 ;
      RECT 17.955000 156.900000 18.485000 163.570000 ;
      RECT 17.955000 166.900000 18.485000 173.570000 ;
      RECT 17.965000 146.840000 18.475000 146.900000 ;
      RECT 17.965000 153.570000 18.475000 153.630000 ;
      RECT 17.965000 156.840000 18.475000 156.900000 ;
      RECT 17.965000 163.570000 18.475000 163.630000 ;
      RECT 17.965000 166.840000 18.475000 166.900000 ;
      RECT 17.965000 173.570000 18.475000 173.630000 ;
      RECT 18.935000  26.900000 19.465000  33.570000 ;
      RECT 18.935000  36.900000 19.465000  43.570000 ;
      RECT 18.935000  46.900000 19.465000  53.570000 ;
      RECT 18.935000  56.900000 19.465000  63.570000 ;
      RECT 18.935000  66.900000 19.465000  71.725000 ;
      RECT 18.935000 176.900000 19.465000 183.570000 ;
      RECT 18.935000 186.900000 19.465000 193.570000 ;
      RECT 19.495000  83.820000 20.405000  84.585000 ;
      RECT 20.045000 146.900000 20.575000 153.570000 ;
      RECT 20.045000 156.900000 20.575000 163.570000 ;
      RECT 20.045000 166.900000 20.575000 173.570000 ;
      RECT 20.320000  26.900000 20.850000  33.570000 ;
      RECT 20.320000  36.900000 20.850000  43.570000 ;
      RECT 20.320000  46.900000 20.850000  53.570000 ;
      RECT 20.320000  56.900000 20.850000  63.570000 ;
      RECT 20.320000  66.900000 20.850000  71.725000 ;
      RECT 20.320000 176.900000 20.850000 183.570000 ;
      RECT 20.320000 186.900000 20.850000 193.570000 ;
      RECT 20.330000  26.840000 20.840000  26.900000 ;
      RECT 20.330000  33.570000 20.840000  33.630000 ;
      RECT 20.330000  36.840000 20.840000  36.900000 ;
      RECT 20.330000  43.570000 20.840000  43.630000 ;
      RECT 20.330000  46.840000 20.840000  46.900000 ;
      RECT 20.330000  53.570000 20.840000  53.630000 ;
      RECT 20.330000  56.840000 20.840000  56.900000 ;
      RECT 20.330000  63.570000 20.840000  63.630000 ;
      RECT 20.330000  66.840000 20.840000  66.900000 ;
      RECT 20.330000 176.840000 20.840000 176.900000 ;
      RECT 20.330000 183.570000 20.840000 183.630000 ;
      RECT 20.330000 186.840000 20.840000 186.900000 ;
      RECT 20.330000 193.570000 20.840000 193.630000 ;
      RECT 20.640000 100.865000 68.495000 101.035000 ;
      RECT 20.640000 101.035000 21.490000 109.275000 ;
      RECT 20.640000 109.275000 68.495000 109.445000 ;
      RECT 20.640000 109.445000 21.490000 117.770000 ;
      RECT 20.640000 117.770000 68.495000 117.940000 ;
      RECT 20.640000 117.940000 21.490000 144.465000 ;
      RECT 21.570000  83.150000 21.740000  99.925000 ;
      RECT 21.570000  99.925000 69.720000 100.095000 ;
      RECT 21.660000 128.010000 65.590000 128.515000 ;
      RECT 21.690000 134.100000 65.590000 136.620000 ;
      RECT 21.705000  26.900000 22.235000  33.570000 ;
      RECT 21.705000  36.900000 22.235000  43.570000 ;
      RECT 21.705000  46.900000 22.235000  53.570000 ;
      RECT 21.705000  56.900000 22.235000  63.570000 ;
      RECT 21.705000  66.900000 22.235000  71.725000 ;
      RECT 21.705000 176.900000 22.235000 183.570000 ;
      RECT 21.705000 186.900000 22.235000 193.570000 ;
      RECT 22.135000 146.900000 22.665000 153.570000 ;
      RECT 22.135000 156.900000 22.665000 163.570000 ;
      RECT 22.135000 166.900000 22.665000 173.570000 ;
      RECT 22.145000 146.840000 22.655000 146.900000 ;
      RECT 22.145000 153.570000 22.655000 153.630000 ;
      RECT 22.145000 156.840000 22.655000 156.900000 ;
      RECT 22.145000 163.570000 22.655000 163.630000 ;
      RECT 22.145000 166.840000 22.655000 166.900000 ;
      RECT 22.145000 173.570000 22.655000 173.630000 ;
      RECT 22.430000  82.085000 23.280000  82.180000 ;
      RECT 22.430000  82.180000 68.140000  82.350000 ;
      RECT 22.430000  82.350000 23.280000  90.675000 ;
      RECT 22.430000  90.675000 68.140000  90.845000 ;
      RECT 22.430000  90.845000 23.280000  97.890000 ;
      RECT 22.770000  97.890000 23.280000  98.990000 ;
      RECT 22.770000  98.990000 68.140000  99.160000 ;
      RECT 23.090000  26.900000 23.620000  33.570000 ;
      RECT 23.090000  36.900000 23.620000  43.570000 ;
      RECT 23.090000  46.900000 23.620000  53.570000 ;
      RECT 23.090000  56.900000 23.620000  63.570000 ;
      RECT 23.090000  66.900000 23.620000  71.725000 ;
      RECT 23.090000 176.900000 23.620000 183.570000 ;
      RECT 23.090000 186.900000 23.620000 193.570000 ;
      RECT 23.100000  26.840000 23.610000  26.900000 ;
      RECT 23.100000  33.570000 23.610000  33.630000 ;
      RECT 23.100000  36.840000 23.610000  36.900000 ;
      RECT 23.100000  43.570000 23.610000  43.630000 ;
      RECT 23.100000  46.840000 23.610000  46.900000 ;
      RECT 23.100000  53.570000 23.610000  53.630000 ;
      RECT 23.100000  56.840000 23.610000  56.900000 ;
      RECT 23.100000  63.570000 23.610000  63.630000 ;
      RECT 23.100000  66.840000 23.610000  66.900000 ;
      RECT 23.100000 176.840000 23.610000 176.900000 ;
      RECT 23.100000 183.570000 23.610000 183.630000 ;
      RECT 23.100000 186.840000 23.610000 186.900000 ;
      RECT 23.100000 193.570000 23.610000 193.630000 ;
      RECT 23.405000 144.100000 65.590000 145.620000 ;
      RECT 23.635000 101.385000 24.045000 108.175000 ;
      RECT 23.635000 109.880000 24.045000 115.550000 ;
      RECT 23.635000 120.080000 24.045000 125.295000 ;
      RECT 23.685000  82.785000 24.215000  89.575000 ;
      RECT 23.685000  91.280000 24.215000  98.070000 ;
      RECT 23.805000 115.550000 24.045000 116.670000 ;
      RECT 23.805000 118.955000 24.045000 120.080000 ;
      RECT 23.805000 125.295000 24.045000 125.745000 ;
      RECT 24.225000 128.730000 24.755000 133.760000 ;
      RECT 24.225000 136.900000 24.755000 143.570000 ;
      RECT 24.225000 146.900000 24.755000 153.570000 ;
      RECT 24.225000 156.900000 24.755000 163.570000 ;
      RECT 24.225000 166.900000 24.755000 173.570000 ;
      RECT 24.475000  26.900000 25.005000  33.570000 ;
      RECT 24.475000  36.900000 25.005000  43.570000 ;
      RECT 24.475000  46.900000 25.005000  53.570000 ;
      RECT 24.475000  56.900000 25.005000  63.570000 ;
      RECT 24.475000  66.900000 25.005000  71.725000 ;
      RECT 24.475000 176.900000 25.005000 183.570000 ;
      RECT 24.475000 186.900000 25.005000 193.570000 ;
      RECT 24.615000  90.045000 66.655000  90.215000 ;
      RECT 24.615000  98.540000 66.655000  98.710000 ;
      RECT 24.670000 108.645000 66.655000 108.815000 ;
      RECT 24.670000 117.140000 66.655000 117.310000 ;
      RECT 24.670000 118.315000 66.655000 118.485000 ;
      RECT 25.310000  75.785000 25.480000  80.300000 ;
      RECT 25.310000  82.915000 25.480000  89.020000 ;
      RECT 25.310000  91.930000 25.480000  96.925000 ;
      RECT 25.365000 101.385000 25.535000 106.255000 ;
      RECT 25.365000 110.450000 25.535000 115.330000 ;
      RECT 25.365000 120.080000 25.535000 124.860000 ;
      RECT 25.860000  26.900000 26.390000  33.570000 ;
      RECT 25.860000  36.900000 26.390000  43.570000 ;
      RECT 25.860000  46.900000 26.390000  53.570000 ;
      RECT 25.860000  56.900000 26.390000  63.570000 ;
      RECT 25.860000  66.900000 26.390000  71.725000 ;
      RECT 25.860000 176.900000 26.390000 183.570000 ;
      RECT 25.860000 186.900000 26.390000 193.570000 ;
      RECT 25.870000  26.840000 26.380000  26.900000 ;
      RECT 25.870000  33.570000 26.380000  33.630000 ;
      RECT 25.870000  36.840000 26.380000  36.900000 ;
      RECT 25.870000  43.570000 26.380000  43.630000 ;
      RECT 25.870000  46.840000 26.380000  46.900000 ;
      RECT 25.870000  53.570000 26.380000  53.630000 ;
      RECT 25.870000  56.840000 26.380000  56.900000 ;
      RECT 25.870000  63.570000 26.380000  63.630000 ;
      RECT 25.870000  66.840000 26.380000  66.900000 ;
      RECT 25.870000 176.840000 26.380000 176.900000 ;
      RECT 25.870000 183.570000 26.380000 183.630000 ;
      RECT 25.870000 186.840000 26.380000 186.900000 ;
      RECT 25.870000 193.570000 26.380000 193.630000 ;
      RECT 26.315000 128.730000 26.845000 133.715000 ;
      RECT 26.315000 136.900000 26.845000 143.570000 ;
      RECT 26.315000 146.900000 26.845000 153.570000 ;
      RECT 26.315000 156.900000 26.845000 163.570000 ;
      RECT 26.315000 166.900000 26.845000 173.570000 ;
      RECT 26.325000 136.840000 26.835000 136.900000 ;
      RECT 26.325000 143.570000 26.835000 143.630000 ;
      RECT 26.325000 146.840000 26.835000 146.900000 ;
      RECT 26.325000 153.570000 26.835000 153.630000 ;
      RECT 26.325000 156.840000 26.835000 156.900000 ;
      RECT 26.325000 163.570000 26.835000 163.630000 ;
      RECT 26.325000 166.840000 26.835000 166.900000 ;
      RECT 26.325000 173.570000 26.835000 173.630000 ;
      RECT 27.245000  26.900000 27.775000  33.570000 ;
      RECT 27.245000  36.900000 27.775000  43.570000 ;
      RECT 27.245000  46.900000 27.775000  53.570000 ;
      RECT 27.245000  56.900000 27.775000  63.570000 ;
      RECT 27.245000  66.900000 27.775000  71.725000 ;
      RECT 27.245000 176.900000 27.775000 183.570000 ;
      RECT 27.245000 186.900000 27.775000 193.570000 ;
      RECT 28.405000 128.860000 28.935000 133.760000 ;
      RECT 28.405000 136.900000 28.935000 143.570000 ;
      RECT 28.405000 146.900000 28.935000 153.570000 ;
      RECT 28.405000 156.900000 28.935000 163.570000 ;
      RECT 28.405000 166.900000 28.935000 173.570000 ;
      RECT 28.630000  26.900000 29.160000  33.570000 ;
      RECT 28.630000  36.900000 29.160000  43.570000 ;
      RECT 28.630000  46.900000 29.160000  53.570000 ;
      RECT 28.630000  56.900000 29.160000  63.570000 ;
      RECT 28.630000  66.900000 29.160000  71.725000 ;
      RECT 28.630000 176.900000 29.160000 183.570000 ;
      RECT 28.630000 186.900000 29.160000 193.570000 ;
      RECT 28.640000  26.840000 29.150000  26.900000 ;
      RECT 28.640000  33.570000 29.150000  33.630000 ;
      RECT 28.640000  36.840000 29.150000  36.900000 ;
      RECT 28.640000  43.570000 29.150000  43.630000 ;
      RECT 28.640000  46.840000 29.150000  46.900000 ;
      RECT 28.640000  53.570000 29.150000  53.630000 ;
      RECT 28.640000  56.840000 29.150000  56.900000 ;
      RECT 28.640000  63.570000 29.150000  63.630000 ;
      RECT 28.640000  66.840000 29.150000  66.900000 ;
      RECT 28.640000 176.840000 29.150000 176.900000 ;
      RECT 28.640000 183.570000 29.150000 183.630000 ;
      RECT 28.640000 186.840000 29.150000 186.900000 ;
      RECT 28.640000 193.570000 29.150000 193.630000 ;
      RECT 30.015000  26.900000 30.545000  33.570000 ;
      RECT 30.015000  36.900000 30.545000  43.570000 ;
      RECT 30.015000  46.900000 30.545000  53.570000 ;
      RECT 30.015000  56.900000 30.545000  63.570000 ;
      RECT 30.015000  66.900000 30.545000  71.725000 ;
      RECT 30.015000 176.900000 30.545000 183.570000 ;
      RECT 30.015000 186.900000 30.545000 193.570000 ;
      RECT 30.495000 128.730000 31.025000 133.715000 ;
      RECT 30.495000 136.900000 31.025000 143.570000 ;
      RECT 30.495000 146.900000 31.025000 153.570000 ;
      RECT 30.495000 156.900000 31.025000 163.570000 ;
      RECT 30.495000 166.900000 31.025000 173.570000 ;
      RECT 30.505000 136.840000 31.015000 136.900000 ;
      RECT 30.505000 143.570000 31.015000 143.630000 ;
      RECT 30.505000 146.840000 31.015000 146.900000 ;
      RECT 30.505000 153.570000 31.015000 153.630000 ;
      RECT 30.505000 156.840000 31.015000 156.900000 ;
      RECT 30.505000 163.570000 31.015000 163.630000 ;
      RECT 30.505000 166.840000 31.015000 166.900000 ;
      RECT 30.505000 173.570000 31.015000 173.630000 ;
      RECT 31.400000  26.900000 31.930000  33.570000 ;
      RECT 31.400000  36.900000 31.930000  43.570000 ;
      RECT 31.400000  46.900000 31.930000  53.570000 ;
      RECT 31.400000  56.900000 31.930000  63.570000 ;
      RECT 31.400000  66.900000 31.930000  71.725000 ;
      RECT 31.400000 176.900000 31.930000 183.570000 ;
      RECT 31.400000 186.900000 31.930000 193.570000 ;
      RECT 31.410000  26.840000 31.920000  26.900000 ;
      RECT 31.410000  33.570000 31.920000  33.630000 ;
      RECT 31.410000  36.840000 31.920000  36.900000 ;
      RECT 31.410000  43.570000 31.920000  43.630000 ;
      RECT 31.410000  46.840000 31.920000  46.900000 ;
      RECT 31.410000  53.570000 31.920000  53.630000 ;
      RECT 31.410000  56.840000 31.920000  56.900000 ;
      RECT 31.410000  63.570000 31.920000  63.630000 ;
      RECT 31.410000  66.840000 31.920000  66.900000 ;
      RECT 31.410000 176.840000 31.920000 176.900000 ;
      RECT 31.410000 183.570000 31.920000 183.630000 ;
      RECT 31.410000 186.840000 31.920000 186.900000 ;
      RECT 31.410000 193.570000 31.920000 193.630000 ;
      RECT 32.585000 128.730000 33.115000 133.755000 ;
      RECT 32.585000 136.900000 33.115000 143.570000 ;
      RECT 32.585000 146.900000 33.115000 153.570000 ;
      RECT 32.585000 156.900000 33.115000 163.570000 ;
      RECT 32.585000 166.900000 33.115000 173.570000 ;
      RECT 32.785000  26.900000 33.315000  33.570000 ;
      RECT 32.785000  36.900000 33.315000  43.570000 ;
      RECT 32.785000  46.900000 33.315000  53.570000 ;
      RECT 32.785000  56.900000 33.315000  63.570000 ;
      RECT 32.785000  66.900000 33.315000  71.725000 ;
      RECT 32.785000 176.900000 33.315000 183.570000 ;
      RECT 32.785000 186.900000 33.315000 193.570000 ;
      RECT 33.590000  75.785000 33.760000  80.300000 ;
      RECT 33.590000  82.915000 33.760000  89.020000 ;
      RECT 33.590000  91.930000 33.760000  96.925000 ;
      RECT 33.590000 101.385000 33.760000 106.255000 ;
      RECT 33.590000 110.450000 33.760000 115.270000 ;
      RECT 33.595000 120.080000 33.765000 124.860000 ;
      RECT 34.170000  26.900000 34.700000  33.570000 ;
      RECT 34.170000  36.900000 34.700000  43.570000 ;
      RECT 34.170000  46.900000 34.700000  53.570000 ;
      RECT 34.170000  56.900000 34.700000  63.570000 ;
      RECT 34.170000  66.900000 34.700000  71.725000 ;
      RECT 34.170000 176.900000 34.700000 183.570000 ;
      RECT 34.170000 186.900000 34.700000 193.570000 ;
      RECT 34.180000  26.840000 34.690000  26.900000 ;
      RECT 34.180000  33.570000 34.690000  33.630000 ;
      RECT 34.180000  36.840000 34.690000  36.900000 ;
      RECT 34.180000  43.570000 34.690000  43.630000 ;
      RECT 34.180000  46.840000 34.690000  46.900000 ;
      RECT 34.180000  53.570000 34.690000  53.630000 ;
      RECT 34.180000  56.840000 34.690000  56.900000 ;
      RECT 34.180000  63.570000 34.690000  63.630000 ;
      RECT 34.180000  66.840000 34.690000  66.900000 ;
      RECT 34.180000 176.840000 34.690000 176.900000 ;
      RECT 34.180000 183.570000 34.690000 183.630000 ;
      RECT 34.180000 186.840000 34.690000 186.900000 ;
      RECT 34.180000 193.570000 34.690000 193.630000 ;
      RECT 34.675000 128.730000 35.205000 133.840000 ;
      RECT 34.675000 136.900000 35.205000 143.570000 ;
      RECT 34.675000 146.900000 35.205000 153.570000 ;
      RECT 34.675000 156.900000 35.205000 163.570000 ;
      RECT 34.675000 166.900000 35.205000 173.570000 ;
      RECT 34.685000 136.840000 35.195000 136.900000 ;
      RECT 34.685000 143.570000 35.195000 143.630000 ;
      RECT 34.685000 146.840000 35.195000 146.900000 ;
      RECT 34.685000 153.570000 35.195000 153.630000 ;
      RECT 34.685000 156.840000 35.195000 156.900000 ;
      RECT 34.685000 163.570000 35.195000 163.630000 ;
      RECT 34.685000 166.840000 35.195000 166.900000 ;
      RECT 34.685000 173.570000 35.195000 173.630000 ;
      RECT 35.555000  26.900000 36.085000  33.570000 ;
      RECT 35.555000  36.900000 36.085000  43.570000 ;
      RECT 35.555000  46.900000 36.085000  53.570000 ;
      RECT 35.555000  56.900000 36.085000  63.570000 ;
      RECT 35.555000  66.900000 36.085000  71.725000 ;
      RECT 35.555000 176.900000 36.085000 183.570000 ;
      RECT 35.555000 186.900000 36.085000 193.570000 ;
      RECT 36.765000 128.730000 37.295000 133.755000 ;
      RECT 36.765000 136.900000 37.295000 143.570000 ;
      RECT 36.765000 146.900000 37.295000 153.570000 ;
      RECT 36.765000 156.900000 37.295000 163.570000 ;
      RECT 36.765000 166.900000 37.295000 173.570000 ;
      RECT 36.940000  26.900000 37.470000  33.570000 ;
      RECT 36.940000  36.900000 37.470000  43.570000 ;
      RECT 36.940000  46.900000 37.470000  53.570000 ;
      RECT 36.940000  56.900000 37.470000  63.570000 ;
      RECT 36.940000  66.900000 37.470000  71.725000 ;
      RECT 36.940000 176.900000 37.470000 183.570000 ;
      RECT 36.940000 186.900000 37.470000 193.570000 ;
      RECT 36.950000  26.840000 37.460000  26.900000 ;
      RECT 36.950000  33.570000 37.460000  33.630000 ;
      RECT 36.950000  36.840000 37.460000  36.900000 ;
      RECT 36.950000  43.570000 37.460000  43.630000 ;
      RECT 36.950000  46.840000 37.460000  46.900000 ;
      RECT 36.950000  53.570000 37.460000  53.630000 ;
      RECT 36.950000  56.840000 37.460000  56.900000 ;
      RECT 36.950000  63.570000 37.460000  63.630000 ;
      RECT 36.950000  66.840000 37.460000  66.900000 ;
      RECT 36.950000 176.840000 37.460000 176.900000 ;
      RECT 36.950000 183.570000 37.460000 183.630000 ;
      RECT 36.950000 186.840000 37.460000 186.900000 ;
      RECT 36.950000 193.570000 37.460000 193.630000 ;
      RECT 38.325000  26.900000 38.855000  33.570000 ;
      RECT 38.325000  36.900000 38.855000  43.570000 ;
      RECT 38.325000  46.900000 38.855000  53.570000 ;
      RECT 38.325000  56.900000 38.855000  63.570000 ;
      RECT 38.325000  66.900000 38.855000  71.725000 ;
      RECT 38.325000 176.900000 38.855000 183.570000 ;
      RECT 38.325000 186.900000 38.855000 193.570000 ;
      RECT 38.855000 128.730000 39.385000 133.925000 ;
      RECT 38.855000 136.900000 39.385000 143.570000 ;
      RECT 38.855000 146.900000 39.385000 153.570000 ;
      RECT 38.855000 156.900000 39.385000 163.570000 ;
      RECT 38.855000 166.900000 39.385000 173.570000 ;
      RECT 38.865000 136.840000 39.375000 136.900000 ;
      RECT 38.865000 143.570000 39.375000 143.630000 ;
      RECT 38.865000 146.840000 39.375000 146.900000 ;
      RECT 38.865000 153.570000 39.375000 153.630000 ;
      RECT 38.865000 156.840000 39.375000 156.900000 ;
      RECT 38.865000 163.570000 39.375000 163.630000 ;
      RECT 38.865000 166.840000 39.375000 166.900000 ;
      RECT 38.865000 173.570000 39.375000 173.630000 ;
      RECT 39.710000  26.900000 40.240000  33.570000 ;
      RECT 39.710000  36.900000 40.240000  43.570000 ;
      RECT 39.710000  46.900000 40.240000  53.570000 ;
      RECT 39.710000  56.900000 40.240000  63.570000 ;
      RECT 39.710000  66.900000 40.240000  71.725000 ;
      RECT 39.710000 176.900000 40.240000 183.570000 ;
      RECT 39.710000 186.900000 40.240000 193.570000 ;
      RECT 39.720000  26.840000 40.230000  26.900000 ;
      RECT 39.720000  33.570000 40.230000  33.630000 ;
      RECT 39.720000  36.840000 40.230000  36.900000 ;
      RECT 39.720000  43.570000 40.230000  43.630000 ;
      RECT 39.720000  46.840000 40.230000  46.900000 ;
      RECT 39.720000  53.570000 40.230000  53.630000 ;
      RECT 39.720000  56.840000 40.230000  56.900000 ;
      RECT 39.720000  63.570000 40.230000  63.630000 ;
      RECT 39.720000  66.840000 40.230000  66.900000 ;
      RECT 39.720000 176.840000 40.230000 176.900000 ;
      RECT 39.720000 183.570000 40.230000 183.630000 ;
      RECT 39.720000 186.840000 40.230000 186.900000 ;
      RECT 39.720000 193.570000 40.230000 193.630000 ;
      RECT 40.945000 128.730000 41.475000 133.755000 ;
      RECT 40.945000 136.900000 41.475000 143.570000 ;
      RECT 40.945000 146.900000 41.475000 153.570000 ;
      RECT 40.945000 156.900000 41.475000 163.570000 ;
      RECT 40.945000 166.900000 41.475000 173.570000 ;
      RECT 41.095000  26.900000 41.625000  33.570000 ;
      RECT 41.095000  36.900000 41.625000  43.570000 ;
      RECT 41.095000  46.900000 41.625000  53.570000 ;
      RECT 41.095000  56.900000 41.625000  63.570000 ;
      RECT 41.095000  66.900000 41.625000  71.725000 ;
      RECT 41.095000 176.900000 41.625000 183.570000 ;
      RECT 41.095000 186.900000 41.625000 193.570000 ;
      RECT 41.870000  75.785000 42.040000  80.300000 ;
      RECT 41.870000  82.915000 42.040000  89.020000 ;
      RECT 41.870000  91.930000 42.040000  96.925000 ;
      RECT 41.870000 101.385000 42.040000 106.255000 ;
      RECT 41.870000 110.450000 42.040000 115.270000 ;
      RECT 41.870000 120.080000 42.040000 124.860000 ;
      RECT 42.480000  26.900000 43.010000  33.570000 ;
      RECT 42.480000  36.900000 43.010000  43.570000 ;
      RECT 42.480000  46.900000 43.010000  53.570000 ;
      RECT 42.480000  56.900000 43.010000  63.570000 ;
      RECT 42.480000  66.900000 43.010000  71.725000 ;
      RECT 42.480000 176.900000 43.010000 183.570000 ;
      RECT 42.480000 186.900000 43.010000 193.570000 ;
      RECT 42.490000  26.840000 43.000000  26.900000 ;
      RECT 42.490000  33.570000 43.000000  33.630000 ;
      RECT 42.490000  36.840000 43.000000  36.900000 ;
      RECT 42.490000  43.570000 43.000000  43.630000 ;
      RECT 42.490000  46.840000 43.000000  46.900000 ;
      RECT 42.490000  53.570000 43.000000  53.630000 ;
      RECT 42.490000  56.840000 43.000000  56.900000 ;
      RECT 42.490000  63.570000 43.000000  63.630000 ;
      RECT 42.490000  66.840000 43.000000  66.900000 ;
      RECT 42.490000 176.840000 43.000000 176.900000 ;
      RECT 42.490000 183.570000 43.000000 183.630000 ;
      RECT 42.490000 186.840000 43.000000 186.900000 ;
      RECT 42.490000 193.570000 43.000000 193.630000 ;
      RECT 43.035000 128.730000 43.565000 133.925000 ;
      RECT 43.035000 136.900000 43.565000 143.570000 ;
      RECT 43.035000 146.900000 43.565000 153.570000 ;
      RECT 43.035000 156.900000 43.565000 163.570000 ;
      RECT 43.035000 166.900000 43.565000 173.570000 ;
      RECT 43.045000 136.840000 43.555000 136.900000 ;
      RECT 43.045000 143.570000 43.555000 143.630000 ;
      RECT 43.045000 146.840000 43.555000 146.900000 ;
      RECT 43.045000 153.570000 43.555000 153.630000 ;
      RECT 43.045000 156.840000 43.555000 156.900000 ;
      RECT 43.045000 163.570000 43.555000 163.630000 ;
      RECT 43.045000 166.840000 43.555000 166.900000 ;
      RECT 43.045000 173.570000 43.555000 173.630000 ;
      RECT 43.865000  26.900000 44.395000  33.570000 ;
      RECT 43.865000  36.900000 44.395000  43.570000 ;
      RECT 43.865000  46.900000 44.395000  53.570000 ;
      RECT 43.865000  56.900000 44.395000  63.570000 ;
      RECT 43.865000  66.900000 44.395000  71.725000 ;
      RECT 43.865000 176.900000 44.395000 183.570000 ;
      RECT 43.865000 186.900000 44.395000 193.570000 ;
      RECT 45.125000 128.730000 45.655000 133.755000 ;
      RECT 45.125000 136.900000 45.655000 143.570000 ;
      RECT 45.125000 146.900000 45.655000 153.570000 ;
      RECT 45.125000 156.900000 45.655000 163.570000 ;
      RECT 45.125000 166.900000 45.655000 173.570000 ;
      RECT 45.250000  26.900000 45.780000  33.570000 ;
      RECT 45.250000  36.900000 45.780000  43.570000 ;
      RECT 45.250000  46.900000 45.780000  53.570000 ;
      RECT 45.250000  56.900000 45.780000  63.570000 ;
      RECT 45.250000  66.900000 45.780000  71.725000 ;
      RECT 45.250000 176.900000 45.780000 183.570000 ;
      RECT 45.250000 186.900000 45.780000 193.570000 ;
      RECT 45.260000  26.840000 45.770000  26.900000 ;
      RECT 45.260000  33.570000 45.770000  33.630000 ;
      RECT 45.260000  36.840000 45.770000  36.900000 ;
      RECT 45.260000  43.570000 45.770000  43.630000 ;
      RECT 45.260000  46.840000 45.770000  46.900000 ;
      RECT 45.260000  53.570000 45.770000  53.630000 ;
      RECT 45.260000  56.840000 45.770000  56.900000 ;
      RECT 45.260000  63.570000 45.770000  63.630000 ;
      RECT 45.260000  66.840000 45.770000  66.900000 ;
      RECT 45.260000 176.840000 45.770000 176.900000 ;
      RECT 45.260000 183.570000 45.770000 183.630000 ;
      RECT 45.260000 186.840000 45.770000 186.900000 ;
      RECT 45.260000 193.570000 45.770000 193.630000 ;
      RECT 46.635000  26.900000 47.165000  33.570000 ;
      RECT 46.635000  36.900000 47.165000  43.570000 ;
      RECT 46.635000  46.900000 47.165000  53.570000 ;
      RECT 46.635000  56.900000 47.165000  63.570000 ;
      RECT 46.635000  66.900000 47.165000  71.725000 ;
      RECT 46.635000 176.900000 47.165000 183.570000 ;
      RECT 46.635000 186.900000 47.165000 193.570000 ;
      RECT 47.215000 128.730000 47.745000 133.925000 ;
      RECT 47.215000 136.900000 47.745000 143.570000 ;
      RECT 47.215000 146.900000 47.745000 153.570000 ;
      RECT 47.215000 156.900000 47.745000 163.570000 ;
      RECT 47.215000 166.900000 47.745000 173.570000 ;
      RECT 47.225000 136.840000 47.735000 136.900000 ;
      RECT 47.225000 143.570000 47.735000 143.630000 ;
      RECT 47.225000 146.840000 47.735000 146.900000 ;
      RECT 47.225000 153.570000 47.735000 153.630000 ;
      RECT 47.225000 156.840000 47.735000 156.900000 ;
      RECT 47.225000 163.570000 47.735000 163.630000 ;
      RECT 47.225000 166.840000 47.735000 166.900000 ;
      RECT 47.225000 173.570000 47.735000 173.630000 ;
      RECT 48.020000  26.900000 48.550000  33.570000 ;
      RECT 48.020000  36.900000 48.550000  43.570000 ;
      RECT 48.020000  46.900000 48.550000  53.570000 ;
      RECT 48.020000  56.900000 48.550000  63.570000 ;
      RECT 48.020000  66.900000 48.550000  71.725000 ;
      RECT 48.020000 176.900000 48.550000 183.570000 ;
      RECT 48.020000 186.900000 48.550000 193.570000 ;
      RECT 48.030000  26.840000 48.540000  26.900000 ;
      RECT 48.030000  33.570000 48.540000  33.630000 ;
      RECT 48.030000  36.840000 48.540000  36.900000 ;
      RECT 48.030000  43.570000 48.540000  43.630000 ;
      RECT 48.030000  46.840000 48.540000  46.900000 ;
      RECT 48.030000  53.570000 48.540000  53.630000 ;
      RECT 48.030000  56.840000 48.540000  56.900000 ;
      RECT 48.030000  63.570000 48.540000  63.630000 ;
      RECT 48.030000  66.840000 48.540000  66.900000 ;
      RECT 48.030000 176.840000 48.540000 176.900000 ;
      RECT 48.030000 183.570000 48.540000 183.630000 ;
      RECT 48.030000 186.840000 48.540000 186.900000 ;
      RECT 48.030000 193.570000 48.540000 193.630000 ;
      RECT 49.305000 128.730000 49.835000 133.755000 ;
      RECT 49.305000 136.900000 49.835000 143.570000 ;
      RECT 49.305000 146.900000 49.835000 153.570000 ;
      RECT 49.305000 156.900000 49.835000 163.570000 ;
      RECT 49.305000 166.900000 49.835000 173.570000 ;
      RECT 49.405000  26.900000 49.935000  33.570000 ;
      RECT 49.405000  36.900000 49.935000  43.570000 ;
      RECT 49.405000  46.900000 49.935000  53.570000 ;
      RECT 49.405000  56.900000 49.935000  63.570000 ;
      RECT 49.405000  66.900000 49.935000  71.725000 ;
      RECT 49.405000 176.900000 49.935000 183.570000 ;
      RECT 49.405000 186.900000 49.935000 193.570000 ;
      RECT 50.150000  75.785000 50.320000  80.300000 ;
      RECT 50.150000  82.915000 50.320000  89.020000 ;
      RECT 50.150000  91.930000 50.320000  96.925000 ;
      RECT 50.150000 101.385000 50.320000 106.255000 ;
      RECT 50.150000 110.450000 50.320000 115.270000 ;
      RECT 50.150000 120.080000 50.320000 124.860000 ;
      RECT 50.790000  26.900000 51.320000  33.570000 ;
      RECT 50.790000  36.900000 51.320000  43.570000 ;
      RECT 50.790000  46.900000 51.320000  53.570000 ;
      RECT 50.790000  56.900000 51.320000  63.570000 ;
      RECT 50.790000  66.900000 51.320000  71.725000 ;
      RECT 50.790000 176.900000 51.320000 183.570000 ;
      RECT 50.790000 186.900000 51.320000 193.570000 ;
      RECT 50.800000  26.840000 51.310000  26.900000 ;
      RECT 50.800000  33.570000 51.310000  33.630000 ;
      RECT 50.800000  36.840000 51.310000  36.900000 ;
      RECT 50.800000  43.570000 51.310000  43.630000 ;
      RECT 50.800000  46.840000 51.310000  46.900000 ;
      RECT 50.800000  53.570000 51.310000  53.630000 ;
      RECT 50.800000  56.840000 51.310000  56.900000 ;
      RECT 50.800000  63.570000 51.310000  63.630000 ;
      RECT 50.800000  66.840000 51.310000  66.900000 ;
      RECT 50.800000 176.840000 51.310000 176.900000 ;
      RECT 50.800000 183.570000 51.310000 183.630000 ;
      RECT 50.800000 186.840000 51.310000 186.900000 ;
      RECT 50.800000 193.570000 51.310000 193.630000 ;
      RECT 51.395000 128.730000 51.925000 133.925000 ;
      RECT 51.395000 136.900000 51.925000 143.570000 ;
      RECT 51.395000 146.900000 51.925000 153.570000 ;
      RECT 51.395000 156.900000 51.925000 163.570000 ;
      RECT 51.395000 166.900000 51.925000 173.570000 ;
      RECT 51.405000 136.840000 51.915000 136.900000 ;
      RECT 51.405000 143.570000 51.915000 143.630000 ;
      RECT 51.405000 146.840000 51.915000 146.900000 ;
      RECT 51.405000 153.570000 51.915000 153.630000 ;
      RECT 51.405000 156.840000 51.915000 156.900000 ;
      RECT 51.405000 163.570000 51.915000 163.630000 ;
      RECT 51.405000 166.840000 51.915000 166.900000 ;
      RECT 51.405000 173.570000 51.915000 173.630000 ;
      RECT 52.175000  26.900000 52.705000  33.570000 ;
      RECT 52.175000  36.900000 52.705000  43.570000 ;
      RECT 52.175000  46.900000 52.705000  53.570000 ;
      RECT 52.175000  56.900000 52.705000  63.570000 ;
      RECT 52.175000  66.900000 52.705000  71.725000 ;
      RECT 52.175000 176.900000 52.705000 183.570000 ;
      RECT 52.175000 186.900000 52.705000 193.570000 ;
      RECT 53.485000 128.730000 54.015000 133.755000 ;
      RECT 53.485000 136.900000 54.015000 143.570000 ;
      RECT 53.485000 146.900000 54.015000 153.570000 ;
      RECT 53.485000 156.900000 54.015000 163.570000 ;
      RECT 53.485000 166.900000 54.015000 173.570000 ;
      RECT 53.560000  26.900000 54.090000  33.570000 ;
      RECT 53.560000  36.900000 54.090000  43.570000 ;
      RECT 53.560000  46.900000 54.090000  53.570000 ;
      RECT 53.560000  56.900000 54.090000  63.570000 ;
      RECT 53.560000  66.900000 54.090000  71.725000 ;
      RECT 53.560000 176.900000 54.090000 183.570000 ;
      RECT 53.560000 186.900000 54.090000 193.570000 ;
      RECT 53.570000  26.840000 54.080000  26.900000 ;
      RECT 53.570000  33.570000 54.080000  33.630000 ;
      RECT 53.570000  36.840000 54.080000  36.900000 ;
      RECT 53.570000  43.570000 54.080000  43.630000 ;
      RECT 53.570000  46.840000 54.080000  46.900000 ;
      RECT 53.570000  53.570000 54.080000  53.630000 ;
      RECT 53.570000  56.840000 54.080000  56.900000 ;
      RECT 53.570000  63.570000 54.080000  63.630000 ;
      RECT 53.570000  66.840000 54.080000  66.900000 ;
      RECT 53.570000 176.840000 54.080000 176.900000 ;
      RECT 53.570000 183.570000 54.080000 183.630000 ;
      RECT 53.570000 186.840000 54.080000 186.900000 ;
      RECT 53.570000 193.570000 54.080000 193.630000 ;
      RECT 54.945000  26.900000 55.475000  33.570000 ;
      RECT 54.945000  36.900000 55.475000  43.570000 ;
      RECT 54.945000  46.900000 55.475000  53.570000 ;
      RECT 54.945000  56.900000 55.475000  63.570000 ;
      RECT 54.945000  66.900000 55.475000  71.725000 ;
      RECT 54.945000 176.900000 55.475000 183.570000 ;
      RECT 54.945000 186.900000 55.475000 193.570000 ;
      RECT 55.575000 128.730000 56.105000 133.925000 ;
      RECT 55.575000 136.900000 56.105000 143.570000 ;
      RECT 55.575000 146.900000 56.105000 153.570000 ;
      RECT 55.575000 156.900000 56.105000 163.570000 ;
      RECT 55.575000 166.900000 56.105000 173.570000 ;
      RECT 55.585000 136.840000 56.095000 136.900000 ;
      RECT 55.585000 143.570000 56.095000 143.630000 ;
      RECT 55.585000 146.840000 56.095000 146.900000 ;
      RECT 55.585000 153.570000 56.095000 153.630000 ;
      RECT 55.585000 156.840000 56.095000 156.900000 ;
      RECT 55.585000 163.570000 56.095000 163.630000 ;
      RECT 55.585000 166.840000 56.095000 166.900000 ;
      RECT 55.585000 173.570000 56.095000 173.630000 ;
      RECT 56.330000  26.900000 56.860000  33.570000 ;
      RECT 56.330000  36.900000 56.860000  43.570000 ;
      RECT 56.330000  46.900000 56.860000  53.570000 ;
      RECT 56.330000  56.900000 56.860000  63.570000 ;
      RECT 56.330000  66.900000 56.860000  71.725000 ;
      RECT 56.330000 176.900000 56.860000 183.570000 ;
      RECT 56.330000 186.900000 56.860000 193.570000 ;
      RECT 56.340000  26.840000 56.850000  26.900000 ;
      RECT 56.340000  33.570000 56.850000  33.630000 ;
      RECT 56.340000  36.840000 56.850000  36.900000 ;
      RECT 56.340000  43.570000 56.850000  43.630000 ;
      RECT 56.340000  46.840000 56.850000  46.900000 ;
      RECT 56.340000  53.570000 56.850000  53.630000 ;
      RECT 56.340000  56.840000 56.850000  56.900000 ;
      RECT 56.340000  63.570000 56.850000  63.630000 ;
      RECT 56.340000  66.840000 56.850000  66.900000 ;
      RECT 56.340000 176.840000 56.850000 176.900000 ;
      RECT 56.340000 183.570000 56.850000 183.630000 ;
      RECT 56.340000 186.840000 56.850000 186.900000 ;
      RECT 56.340000 193.570000 56.850000 193.630000 ;
      RECT 56.980000  16.365000 57.510000  16.895000 ;
      RECT 57.665000 128.730000 58.195000 133.755000 ;
      RECT 57.665000 136.900000 58.195000 143.570000 ;
      RECT 57.665000 146.900000 58.195000 153.570000 ;
      RECT 57.665000 156.900000 58.195000 163.570000 ;
      RECT 57.665000 166.900000 58.195000 173.570000 ;
      RECT 57.715000  26.900000 58.245000  33.570000 ;
      RECT 57.715000  36.900000 58.245000  43.570000 ;
      RECT 57.715000  46.900000 58.245000  53.570000 ;
      RECT 57.715000  56.900000 58.245000  63.570000 ;
      RECT 57.715000  66.900000 58.245000  71.725000 ;
      RECT 57.715000 176.900000 58.245000 183.570000 ;
      RECT 57.715000 186.900000 58.245000 193.570000 ;
      RECT 58.430000  75.785000 58.600000  80.300000 ;
      RECT 58.430000  82.915000 58.600000  89.020000 ;
      RECT 58.430000  91.930000 58.600000  96.925000 ;
      RECT 58.430000 101.385000 58.600000 106.255000 ;
      RECT 58.430000 110.450000 58.600000 115.270000 ;
      RECT 58.430000 120.080000 58.600000 124.860000 ;
      RECT 59.100000  26.900000 59.630000  33.570000 ;
      RECT 59.100000  36.900000 59.630000  43.570000 ;
      RECT 59.100000  46.900000 59.630000  53.570000 ;
      RECT 59.100000  56.900000 59.630000  63.570000 ;
      RECT 59.100000  66.900000 59.630000  71.725000 ;
      RECT 59.100000 176.900000 59.630000 183.570000 ;
      RECT 59.100000 186.900000 59.630000 193.570000 ;
      RECT 59.110000  26.840000 59.620000  26.900000 ;
      RECT 59.110000  33.570000 59.620000  33.630000 ;
      RECT 59.110000  36.840000 59.620000  36.900000 ;
      RECT 59.110000  43.570000 59.620000  43.630000 ;
      RECT 59.110000  46.840000 59.620000  46.900000 ;
      RECT 59.110000  53.570000 59.620000  53.630000 ;
      RECT 59.110000  56.840000 59.620000  56.900000 ;
      RECT 59.110000  63.570000 59.620000  63.630000 ;
      RECT 59.110000  66.840000 59.620000  66.900000 ;
      RECT 59.110000 176.840000 59.620000 176.900000 ;
      RECT 59.110000 183.570000 59.620000 183.630000 ;
      RECT 59.110000 186.840000 59.620000 186.900000 ;
      RECT 59.110000 193.570000 59.620000 193.630000 ;
      RECT 59.755000 128.730000 60.285000 133.925000 ;
      RECT 59.755000 136.900000 60.285000 143.570000 ;
      RECT 59.755000 146.900000 60.285000 153.570000 ;
      RECT 59.755000 156.900000 60.285000 163.570000 ;
      RECT 59.755000 166.900000 60.285000 173.570000 ;
      RECT 59.765000 136.840000 60.275000 136.900000 ;
      RECT 59.765000 143.570000 60.275000 143.630000 ;
      RECT 59.765000 146.840000 60.275000 146.900000 ;
      RECT 59.765000 153.570000 60.275000 153.630000 ;
      RECT 59.765000 156.840000 60.275000 156.900000 ;
      RECT 59.765000 163.570000 60.275000 163.630000 ;
      RECT 59.765000 166.840000 60.275000 166.900000 ;
      RECT 59.765000 173.570000 60.275000 173.630000 ;
      RECT 60.485000  26.900000 61.015000  33.570000 ;
      RECT 60.485000  36.900000 61.015000  43.570000 ;
      RECT 60.485000  46.900000 61.015000  53.570000 ;
      RECT 60.485000  56.900000 61.015000  63.570000 ;
      RECT 60.485000  66.900000 61.015000  71.725000 ;
      RECT 60.485000 176.900000 61.015000 183.570000 ;
      RECT 60.485000 186.900000 61.015000 193.570000 ;
      RECT 61.845000 128.730000 62.375000 133.755000 ;
      RECT 61.845000 136.900000 62.375000 143.570000 ;
      RECT 61.845000 146.900000 62.375000 153.570000 ;
      RECT 61.845000 156.900000 62.375000 163.570000 ;
      RECT 61.845000 166.900000 62.375000 173.570000 ;
      RECT 61.870000  26.900000 62.400000  33.570000 ;
      RECT 61.870000  36.900000 62.400000  43.570000 ;
      RECT 61.870000  46.900000 62.400000  53.570000 ;
      RECT 61.870000  56.900000 62.400000  63.570000 ;
      RECT 61.870000  66.900000 62.400000  71.725000 ;
      RECT 61.870000 176.900000 62.400000 183.570000 ;
      RECT 61.870000 186.900000 62.400000 193.570000 ;
      RECT 61.880000  26.840000 62.390000  26.900000 ;
      RECT 61.880000  33.570000 62.390000  33.630000 ;
      RECT 61.880000  36.840000 62.390000  36.900000 ;
      RECT 61.880000  43.570000 62.390000  43.630000 ;
      RECT 61.880000  46.840000 62.390000  46.900000 ;
      RECT 61.880000  53.570000 62.390000  53.630000 ;
      RECT 61.880000  56.840000 62.390000  56.900000 ;
      RECT 61.880000  63.570000 62.390000  63.630000 ;
      RECT 61.880000  66.840000 62.390000  66.900000 ;
      RECT 61.880000 176.840000 62.390000 176.900000 ;
      RECT 61.880000 183.570000 62.390000 183.630000 ;
      RECT 61.880000 186.840000 62.390000 186.900000 ;
      RECT 61.880000 193.570000 62.390000 193.630000 ;
      RECT 63.255000  26.900000 63.785000  33.570000 ;
      RECT 63.255000  36.900000 63.785000  43.570000 ;
      RECT 63.255000  46.900000 63.785000  53.570000 ;
      RECT 63.255000  56.900000 63.785000  63.570000 ;
      RECT 63.255000  66.900000 63.785000  71.725000 ;
      RECT 63.255000 176.900000 63.785000 183.570000 ;
      RECT 63.255000 186.900000 63.785000 193.570000 ;
      RECT 63.935000 128.730000 64.465000 133.925000 ;
      RECT 63.935000 136.900000 64.465000 143.570000 ;
      RECT 63.935000 146.900000 64.465000 153.570000 ;
      RECT 63.935000 156.900000 64.465000 163.570000 ;
      RECT 63.935000 166.900000 64.465000 173.570000 ;
      RECT 63.945000 136.840000 64.455000 136.900000 ;
      RECT 63.945000 143.570000 64.455000 143.630000 ;
      RECT 63.945000 146.840000 64.455000 146.900000 ;
      RECT 63.945000 153.570000 64.455000 153.630000 ;
      RECT 63.945000 156.840000 64.455000 156.900000 ;
      RECT 63.945000 163.570000 64.455000 163.630000 ;
      RECT 63.945000 166.840000 64.455000 166.900000 ;
      RECT 63.945000 173.570000 64.455000 173.630000 ;
      RECT 64.640000  26.900000 65.170000  33.570000 ;
      RECT 64.640000  36.900000 65.170000  43.570000 ;
      RECT 64.640000  46.900000 65.170000  53.570000 ;
      RECT 64.640000  56.900000 65.170000  63.570000 ;
      RECT 64.640000  66.900000 65.170000  71.725000 ;
      RECT 64.640000 176.900000 65.170000 183.570000 ;
      RECT 64.640000 186.900000 65.170000 193.570000 ;
      RECT 64.650000  26.840000 65.160000  26.900000 ;
      RECT 64.650000  33.570000 65.160000  33.630000 ;
      RECT 64.650000  36.840000 65.160000  36.900000 ;
      RECT 64.650000  43.570000 65.160000  43.630000 ;
      RECT 64.650000  46.840000 65.160000  46.900000 ;
      RECT 64.650000  53.570000 65.160000  53.630000 ;
      RECT 64.650000  56.840000 65.160000  56.900000 ;
      RECT 64.650000  63.570000 65.160000  63.630000 ;
      RECT 64.650000  66.840000 65.160000  66.900000 ;
      RECT 64.650000 176.840000 65.160000 176.900000 ;
      RECT 64.650000 183.570000 65.160000 183.630000 ;
      RECT 64.650000 186.840000 65.160000 186.900000 ;
      RECT 64.650000 193.570000 65.160000 193.630000 ;
      RECT 66.025000  26.900000 66.555000  33.570000 ;
      RECT 66.025000  36.900000 66.555000  43.570000 ;
      RECT 66.025000  46.900000 66.555000  53.570000 ;
      RECT 66.025000  56.900000 66.555000  63.570000 ;
      RECT 66.025000  66.900000 66.555000  71.725000 ;
      RECT 66.025000 128.730000 66.555000 133.755000 ;
      RECT 66.025000 136.900000 66.555000 143.570000 ;
      RECT 66.025000 146.900000 66.555000 153.570000 ;
      RECT 66.025000 156.900000 66.555000 163.570000 ;
      RECT 66.025000 166.900000 66.555000 173.570000 ;
      RECT 66.025000 176.900000 66.555000 183.570000 ;
      RECT 66.025000 186.900000 66.555000 193.570000 ;
      RECT 66.700000   1.205000 67.230000   1.735000 ;
      RECT 66.710000  75.785000 66.880000  80.535000 ;
      RECT 66.710000  82.785000 66.880000  89.375000 ;
      RECT 66.710000  91.280000 66.880000  97.870000 ;
      RECT 66.710000 101.385000 66.880000 106.255000 ;
      RECT 66.710000 110.450000 66.880000 115.270000 ;
      RECT 66.710000 120.080000 66.880000 124.860000 ;
      RECT 67.290000  26.015000 68.140000  82.180000 ;
      RECT 67.290000  82.350000 68.140000  90.675000 ;
      RECT 67.290000  90.845000 68.140000  98.990000 ;
      RECT 67.575000 101.035000 68.495000 109.275000 ;
      RECT 67.575000 109.445000 68.495000 117.770000 ;
      RECT 67.575000 117.940000 68.495000 194.935000 ;
      RECT 67.610000   1.080000 73.375000   1.250000 ;
      RECT 67.615000   1.250000 67.785000  17.100000 ;
      RECT 67.615000  17.100000 73.375000  17.270000 ;
      RECT 68.110000   3.280000 68.280000   9.020000 ;
      RECT 68.110000   9.770000 68.280000  16.670000 ;
      RECT 68.335000   1.670000 72.655000   1.840000 ;
      RECT 68.335000   9.320000 72.655000   9.490000 ;
      RECT 68.570000   2.550000 68.740000   9.020000 ;
      RECT 68.570000  10.200000 68.740000  15.660000 ;
      RECT 69.030000   3.280000 69.200000   9.020000 ;
      RECT 69.030000   9.770000 69.200000  16.670000 ;
      RECT 69.190000  24.355000 69.720000  99.925000 ;
      RECT 69.190000 100.095000 69.720000 196.850000 ;
      RECT 69.490000   2.550000 69.660000   9.020000 ;
      RECT 69.490000  10.200000 69.660000  15.660000 ;
      RECT 69.530000  19.010000 70.265000  19.610000 ;
      RECT 69.950000   3.280000 70.120000   9.020000 ;
      RECT 69.950000   9.770000 70.120000  16.670000 ;
      RECT 70.410000   2.550000 70.580000   9.020000 ;
      RECT 70.410000  10.200000 70.580000  15.660000 ;
      RECT 70.495000  17.960000 71.095000  18.695000 ;
      RECT 70.870000   3.280000 71.040000   9.020000 ;
      RECT 70.870000   9.770000 71.040000  16.670000 ;
      RECT 71.330000   2.550000 71.500000   9.020000 ;
      RECT 71.330000  10.200000 71.500000  15.660000 ;
      RECT 71.790000   3.280000 71.960000   9.020000 ;
      RECT 71.790000   9.770000 71.960000  16.670000 ;
      RECT 72.250000   2.550000 72.420000   9.020000 ;
      RECT 72.250000  10.200000 72.420000  15.660000 ;
      RECT 72.710000   2.120000 72.880000   9.020000 ;
      RECT 72.710000   9.770000 72.880000  16.670000 ;
      RECT 73.205000   1.250000 73.375000  17.100000 ;
      RECT 73.875000 196.920000 74.755000 197.780000 ;
    LAYER met1 ;
      RECT  0.000000   0.000000 25.930000   0.295000 ;
      RECT  0.000000   0.000000 26.070000   0.310000 ;
      RECT  0.000000   0.295000 25.930000   0.310000 ;
      RECT  0.000000   0.310000 25.945000   0.325000 ;
      RECT  0.000000   0.310000 75.000000 198.000000 ;
      RECT  0.000000   0.325000 75.000000   3.330000 ;
      RECT  0.000000   3.330000  3.005000 194.995000 ;
      RECT  0.000000 194.995000 75.000000 198.000000 ;
      RECT  3.002000   3.002000 24.391000   3.070000 ;
      RECT  3.002000   3.002000 24.391000   3.070000 ;
      RECT  3.002000   3.070000 24.459000   3.140000 ;
      RECT  3.002000   3.070000 24.459000   3.140000 ;
      RECT  3.002000   3.140000 24.529000   3.210000 ;
      RECT  3.002000   3.140000 24.529000   3.210000 ;
      RECT  3.002000   3.210000 24.599000   3.280000 ;
      RECT  3.002000   3.210000 24.599000   3.280000 ;
      RECT  3.002000   3.280000 24.669000   3.325000 ;
      RECT  3.002000   3.280000 24.669000   3.325000 ;
      RECT  3.002000   3.327000 71.998000 194.998000 ;
      RECT 27.840000   0.000000 75.000000   0.310000 ;
      RECT 27.950000   0.320000 75.000000   0.325000 ;
      RECT 27.965000   0.305000 75.000000   0.320000 ;
      RECT 27.980000   0.000000 75.000000   0.290000 ;
      RECT 27.980000   0.290000 75.000000   0.305000 ;
      RECT 30.952000   3.002000 71.998000   6.332000 ;
      RECT 71.995000   3.330000 75.000000 194.995000 ;
    LAYER met2 ;
      RECT  0.000000   0.000000  0.220000 193.910000 ;
      RECT  0.000000   0.000000  0.220000 193.910000 ;
      RECT  0.000000 193.910000 75.000000 198.000000 ;
      RECT  0.000000 193.910000 75.000000 198.000000 ;
      RECT 10.700000   8.166000 11.735000   9.704000 ;
      RECT 10.700000   8.166000 11.735000   9.704000 ;
      RECT 10.700000   9.704000 11.735000   9.714000 ;
      RECT 10.705000   8.161000 11.735000   8.165000 ;
      RECT 10.705000   8.161000 11.735000   8.166000 ;
      RECT 10.706000   9.704000 11.735000   9.710000 ;
      RECT 10.710000   9.714000 11.514000   9.935000 ;
      RECT 10.711000   9.710000 11.735000   9.715000 ;
      RECT 10.721000   8.145000 11.719000   8.160000 ;
      RECT 10.781000   9.714000 11.664000   9.785000 ;
      RECT 10.791000   8.075000 11.649000   8.145000 ;
      RECT 10.851000   9.785000 11.594000   9.855000 ;
      RECT 10.861000   8.005000 11.579000   8.075000 ;
      RECT 10.921000   9.855000 11.524000   9.925000 ;
      RECT 10.931000   7.935000 11.509000   8.005000 ;
      RECT 10.931000   7.935000 11.735000   8.161000 ;
      RECT 10.931000   9.925000 11.514000   9.935000 ;
      RECT 14.030000  25.301000 65.465000  25.370000 ;
      RECT 14.030000  25.301000 65.465000  25.370000 ;
      RECT 14.030000  25.301000 65.860000  25.498000 ;
      RECT 14.030000  25.370000 65.534000  25.440000 ;
      RECT 14.030000  25.370000 65.534000  25.440000 ;
      RECT 14.030000  25.440000 65.604000  25.510000 ;
      RECT 14.030000  25.440000 65.604000  25.510000 ;
      RECT 14.030000  25.498000 65.860000  29.822000 ;
      RECT 14.030000  25.510000 65.674000  25.555000 ;
      RECT 14.030000  25.510000 65.674000  25.555000 ;
      RECT 14.030000  25.556000 65.720000  29.764000 ;
      RECT 14.030000  29.764000 65.649000  29.835000 ;
      RECT 14.030000  29.764000 65.649000  29.835000 ;
      RECT 14.030000  29.822000 64.812000  30.870000 ;
      RECT 14.030000  29.835000 65.579000  29.905000 ;
      RECT 14.030000  29.835000 65.579000  29.905000 ;
      RECT 14.030000  29.905000 65.509000  29.975000 ;
      RECT 14.030000  29.905000 65.509000  29.975000 ;
      RECT 14.030000  29.975000 65.439000  30.045000 ;
      RECT 14.030000  29.975000 65.439000  30.045000 ;
      RECT 14.030000  30.045000 65.369000  30.115000 ;
      RECT 14.030000  30.045000 65.369000  30.115000 ;
      RECT 14.030000  30.115000 65.299000  30.185000 ;
      RECT 14.030000  30.115000 65.299000  30.185000 ;
      RECT 14.030000  30.185000 65.229000  30.255000 ;
      RECT 14.030000  30.185000 65.229000  30.255000 ;
      RECT 14.030000  30.255000 65.159000  30.325000 ;
      RECT 14.030000  30.255000 65.159000  30.325000 ;
      RECT 14.030000  30.325000 65.089000  30.395000 ;
      RECT 14.030000  30.325000 65.089000  30.395000 ;
      RECT 14.030000  30.395000 65.019000  30.465000 ;
      RECT 14.030000  30.395000 65.019000  30.465000 ;
      RECT 14.030000  30.465000 64.949000  30.535000 ;
      RECT 14.030000  30.465000 64.949000  30.535000 ;
      RECT 14.030000  30.535000 64.879000  30.605000 ;
      RECT 14.030000  30.535000 64.879000  30.605000 ;
      RECT 14.030000  30.605000 64.809000  30.675000 ;
      RECT 14.030000  30.605000 64.809000  30.675000 ;
      RECT 14.030000  30.675000 64.754000  30.730000 ;
      RECT 14.030000  30.675000 64.754000  30.730000 ;
      RECT 14.030000  30.730000 15.855000  33.930000 ;
      RECT 14.030000  30.870000 15.995000  33.790000 ;
      RECT 14.030000  33.790000 65.860000  34.748000 ;
      RECT 14.030000  33.930000 64.844000  34.000000 ;
      RECT 14.030000  33.930000 64.844000  34.000000 ;
      RECT 14.030000  34.000000 64.914000  34.070000 ;
      RECT 14.030000  34.000000 64.914000  34.070000 ;
      RECT 14.030000  34.070000 64.984000  34.140000 ;
      RECT 14.030000  34.070000 64.984000  34.140000 ;
      RECT 14.030000  34.140000 65.054000  34.210000 ;
      RECT 14.030000  34.140000 65.054000  34.210000 ;
      RECT 14.030000  34.210000 65.124000  34.280000 ;
      RECT 14.030000  34.210000 65.124000  34.280000 ;
      RECT 14.030000  34.280000 65.194000  34.350000 ;
      RECT 14.030000  34.280000 65.194000  34.350000 ;
      RECT 14.030000  34.350000 65.264000  34.420000 ;
      RECT 14.030000  34.350000 65.264000  34.420000 ;
      RECT 14.030000  34.420000 65.334000  34.490000 ;
      RECT 14.030000  34.420000 65.334000  34.490000 ;
      RECT 14.030000  34.490000 65.404000  34.560000 ;
      RECT 14.030000  34.490000 65.404000  34.560000 ;
      RECT 14.030000  34.560000 65.474000  34.630000 ;
      RECT 14.030000  34.560000 65.474000  34.630000 ;
      RECT 14.030000  34.630000 65.544000  34.700000 ;
      RECT 14.030000  34.630000 65.544000  34.700000 ;
      RECT 14.030000  34.700000 65.614000  34.770000 ;
      RECT 14.030000  34.700000 65.614000  34.770000 ;
      RECT 14.030000  34.748000 65.860000  39.877000 ;
      RECT 14.030000  34.770000 65.684000  34.805000 ;
      RECT 14.030000  34.770000 65.684000  34.805000 ;
      RECT 14.030000  34.806000 65.720000  39.819000 ;
      RECT 14.030000  39.819000 65.649000  39.890000 ;
      RECT 14.030000  39.819000 65.649000  39.890000 ;
      RECT 14.030000  39.877000 64.887000  40.850000 ;
      RECT 14.030000  39.890000 65.579000  39.960000 ;
      RECT 14.030000  39.890000 65.579000  39.960000 ;
      RECT 14.030000  39.960000 65.509000  40.030000 ;
      RECT 14.030000  39.960000 65.509000  40.030000 ;
      RECT 14.030000  40.030000 65.439000  40.100000 ;
      RECT 14.030000  40.030000 65.439000  40.100000 ;
      RECT 14.030000  40.100000 65.369000  40.170000 ;
      RECT 14.030000  40.100000 65.369000  40.170000 ;
      RECT 14.030000  40.170000 65.299000  40.240000 ;
      RECT 14.030000  40.170000 65.299000  40.240000 ;
      RECT 14.030000  40.240000 65.229000  40.310000 ;
      RECT 14.030000  40.240000 65.229000  40.310000 ;
      RECT 14.030000  40.310000 65.159000  40.380000 ;
      RECT 14.030000  40.310000 65.159000  40.380000 ;
      RECT 14.030000  40.380000 65.089000  40.450000 ;
      RECT 14.030000  40.380000 65.089000  40.450000 ;
      RECT 14.030000  40.450000 65.019000  40.520000 ;
      RECT 14.030000  40.450000 65.019000  40.520000 ;
      RECT 14.030000  40.520000 64.949000  40.590000 ;
      RECT 14.030000  40.520000 64.949000  40.590000 ;
      RECT 14.030000  40.590000 64.879000  40.660000 ;
      RECT 14.030000  40.590000 64.879000  40.660000 ;
      RECT 14.030000  40.660000 64.829000  40.710000 ;
      RECT 14.030000  40.660000 64.829000  40.710000 ;
      RECT 14.030000  40.710000 15.855000  43.910000 ;
      RECT 14.030000  40.850000 15.995000  43.770000 ;
      RECT 14.030000  43.770000 65.860000  44.728000 ;
      RECT 14.030000  43.910000 64.844000  43.980000 ;
      RECT 14.030000  43.910000 64.844000  43.980000 ;
      RECT 14.030000  43.980000 64.914000  44.050000 ;
      RECT 14.030000  43.980000 64.914000  44.050000 ;
      RECT 14.030000  44.050000 64.984000  44.120000 ;
      RECT 14.030000  44.050000 64.984000  44.120000 ;
      RECT 14.030000  44.120000 65.054000  44.190000 ;
      RECT 14.030000  44.120000 65.054000  44.190000 ;
      RECT 14.030000  44.190000 65.124000  44.260000 ;
      RECT 14.030000  44.190000 65.124000  44.260000 ;
      RECT 14.030000  44.260000 65.194000  44.330000 ;
      RECT 14.030000  44.260000 65.194000  44.330000 ;
      RECT 14.030000  44.330000 65.264000  44.400000 ;
      RECT 14.030000  44.330000 65.264000  44.400000 ;
      RECT 14.030000  44.400000 65.334000  44.470000 ;
      RECT 14.030000  44.400000 65.334000  44.470000 ;
      RECT 14.030000  44.470000 65.404000  44.540000 ;
      RECT 14.030000  44.470000 65.404000  44.540000 ;
      RECT 14.030000  44.540000 65.474000  44.610000 ;
      RECT 14.030000  44.540000 65.474000  44.610000 ;
      RECT 14.030000  44.610000 65.544000  44.680000 ;
      RECT 14.030000  44.610000 65.544000  44.680000 ;
      RECT 14.030000  44.680000 65.614000  44.750000 ;
      RECT 14.030000  44.680000 65.614000  44.750000 ;
      RECT 14.030000  44.728000 65.860000  49.897000 ;
      RECT 14.030000  44.750000 65.684000  44.785000 ;
      RECT 14.030000  44.750000 65.684000  44.785000 ;
      RECT 14.030000  44.786000 65.720000  49.839000 ;
      RECT 14.030000  49.839000 65.649000  49.910000 ;
      RECT 14.030000  49.839000 65.649000  49.910000 ;
      RECT 14.030000  49.897000 64.887000  50.870000 ;
      RECT 14.030000  49.910000 65.579000  49.980000 ;
      RECT 14.030000  49.910000 65.579000  49.980000 ;
      RECT 14.030000  49.980000 65.509000  50.050000 ;
      RECT 14.030000  49.980000 65.509000  50.050000 ;
      RECT 14.030000  50.050000 65.439000  50.120000 ;
      RECT 14.030000  50.050000 65.439000  50.120000 ;
      RECT 14.030000  50.120000 65.369000  50.190000 ;
      RECT 14.030000  50.120000 65.369000  50.190000 ;
      RECT 14.030000  50.190000 65.299000  50.260000 ;
      RECT 14.030000  50.190000 65.299000  50.260000 ;
      RECT 14.030000  50.260000 65.229000  50.330000 ;
      RECT 14.030000  50.260000 65.229000  50.330000 ;
      RECT 14.030000  50.330000 65.159000  50.400000 ;
      RECT 14.030000  50.330000 65.159000  50.400000 ;
      RECT 14.030000  50.400000 65.089000  50.470000 ;
      RECT 14.030000  50.400000 65.089000  50.470000 ;
      RECT 14.030000  50.470000 65.019000  50.540000 ;
      RECT 14.030000  50.470000 65.019000  50.540000 ;
      RECT 14.030000  50.540000 64.949000  50.610000 ;
      RECT 14.030000  50.540000 64.949000  50.610000 ;
      RECT 14.030000  50.610000 64.879000  50.680000 ;
      RECT 14.030000  50.610000 64.879000  50.680000 ;
      RECT 14.030000  50.680000 64.829000  50.730000 ;
      RECT 14.030000  50.680000 64.829000  50.730000 ;
      RECT 14.030000  50.730000 15.855000  53.930000 ;
      RECT 14.030000  50.870000 15.995000  53.790000 ;
      RECT 14.030000  53.790000 65.855000  54.743000 ;
      RECT 14.030000  53.930000 64.844000  54.000000 ;
      RECT 14.030000  53.930000 64.844000  54.000000 ;
      RECT 14.030000  54.000000 64.914000  54.070000 ;
      RECT 14.030000  54.000000 64.914000  54.070000 ;
      RECT 14.030000  54.070000 64.984000  54.140000 ;
      RECT 14.030000  54.070000 64.984000  54.140000 ;
      RECT 14.030000  54.140000 65.054000  54.210000 ;
      RECT 14.030000  54.140000 65.054000  54.210000 ;
      RECT 14.030000  54.210000 65.124000  54.280000 ;
      RECT 14.030000  54.210000 65.124000  54.280000 ;
      RECT 14.030000  54.280000 65.194000  54.350000 ;
      RECT 14.030000  54.280000 65.194000  54.350000 ;
      RECT 14.030000  54.350000 65.264000  54.420000 ;
      RECT 14.030000  54.350000 65.264000  54.420000 ;
      RECT 14.030000  54.420000 65.334000  54.490000 ;
      RECT 14.030000  54.420000 65.334000  54.490000 ;
      RECT 14.030000  54.490000 65.404000  54.560000 ;
      RECT 14.030000  54.490000 65.404000  54.560000 ;
      RECT 14.030000  54.560000 65.474000  54.630000 ;
      RECT 14.030000  54.560000 65.474000  54.630000 ;
      RECT 14.030000  54.630000 65.544000  54.700000 ;
      RECT 14.030000  54.630000 65.544000  54.700000 ;
      RECT 14.030000  54.700000 65.614000  54.770000 ;
      RECT 14.030000  54.700000 65.614000  54.770000 ;
      RECT 14.030000  54.743000 65.855000  59.882000 ;
      RECT 14.030000  54.770000 65.684000  54.800000 ;
      RECT 14.030000  54.770000 65.684000  54.800000 ;
      RECT 14.030000  54.801000 65.715000  59.824000 ;
      RECT 14.030000  59.824000 65.644000  59.895000 ;
      RECT 14.030000  59.824000 65.644000  59.895000 ;
      RECT 14.030000  59.882000 64.887000  60.850000 ;
      RECT 14.030000  59.895000 65.574000  59.965000 ;
      RECT 14.030000  59.895000 65.574000  59.965000 ;
      RECT 14.030000  59.965000 65.504000  60.035000 ;
      RECT 14.030000  59.965000 65.504000  60.035000 ;
      RECT 14.030000  60.035000 65.434000  60.105000 ;
      RECT 14.030000  60.035000 65.434000  60.105000 ;
      RECT 14.030000  60.105000 65.364000  60.175000 ;
      RECT 14.030000  60.105000 65.364000  60.175000 ;
      RECT 14.030000  60.175000 65.294000  60.245000 ;
      RECT 14.030000  60.175000 65.294000  60.245000 ;
      RECT 14.030000  60.245000 65.224000  60.315000 ;
      RECT 14.030000  60.245000 65.224000  60.315000 ;
      RECT 14.030000  60.315000 65.154000  60.385000 ;
      RECT 14.030000  60.315000 65.154000  60.385000 ;
      RECT 14.030000  60.385000 65.084000  60.455000 ;
      RECT 14.030000  60.385000 65.084000  60.455000 ;
      RECT 14.030000  60.455000 65.014000  60.525000 ;
      RECT 14.030000  60.455000 65.014000  60.525000 ;
      RECT 14.030000  60.525000 64.944000  60.595000 ;
      RECT 14.030000  60.525000 64.944000  60.595000 ;
      RECT 14.030000  60.595000 64.874000  60.665000 ;
      RECT 14.030000  60.595000 64.874000  60.665000 ;
      RECT 14.030000  60.665000 64.829000  60.710000 ;
      RECT 14.030000  60.665000 64.829000  60.710000 ;
      RECT 14.030000  60.710000 15.855000  63.910000 ;
      RECT 14.030000  60.850000 15.995000  63.770000 ;
      RECT 14.030000  63.770000 65.855000  64.738000 ;
      RECT 14.030000  63.910000 64.829000  63.980000 ;
      RECT 14.030000  63.910000 64.829000  63.980000 ;
      RECT 14.030000  63.980000 64.899000  64.050000 ;
      RECT 14.030000  63.980000 64.899000  64.050000 ;
      RECT 14.030000  64.050000 64.969000  64.120000 ;
      RECT 14.030000  64.050000 64.969000  64.120000 ;
      RECT 14.030000  64.120000 65.039000  64.190000 ;
      RECT 14.030000  64.120000 65.039000  64.190000 ;
      RECT 14.030000  64.190000 65.109000  64.260000 ;
      RECT 14.030000  64.190000 65.109000  64.260000 ;
      RECT 14.030000  64.260000 65.179000  64.330000 ;
      RECT 14.030000  64.260000 65.179000  64.330000 ;
      RECT 14.030000  64.330000 65.249000  64.400000 ;
      RECT 14.030000  64.330000 65.249000  64.400000 ;
      RECT 14.030000  64.400000 65.319000  64.470000 ;
      RECT 14.030000  64.400000 65.319000  64.470000 ;
      RECT 14.030000  64.470000 65.389000  64.540000 ;
      RECT 14.030000  64.470000 65.389000  64.540000 ;
      RECT 14.030000  64.540000 65.459000  64.610000 ;
      RECT 14.030000  64.540000 65.459000  64.610000 ;
      RECT 14.030000  64.610000 65.529000  64.680000 ;
      RECT 14.030000  64.610000 65.529000  64.680000 ;
      RECT 14.030000  64.680000 65.599000  64.750000 ;
      RECT 14.030000  64.680000 65.599000  64.750000 ;
      RECT 14.030000  64.738000 65.855000  69.882000 ;
      RECT 14.030000  64.750000 65.669000  64.795000 ;
      RECT 14.030000  64.750000 65.669000  64.795000 ;
      RECT 14.030000  64.796000 65.715000  69.824000 ;
      RECT 14.030000  69.824000 65.644000  69.895000 ;
      RECT 14.030000  69.824000 65.644000  69.895000 ;
      RECT 14.030000  69.882000 64.887000  70.850000 ;
      RECT 14.030000  69.895000 65.574000  69.965000 ;
      RECT 14.030000  69.895000 65.574000  69.965000 ;
      RECT 14.030000  69.965000 65.504000  70.035000 ;
      RECT 14.030000  69.965000 65.504000  70.035000 ;
      RECT 14.030000  70.035000 65.434000  70.105000 ;
      RECT 14.030000  70.035000 65.434000  70.105000 ;
      RECT 14.030000  70.105000 65.364000  70.175000 ;
      RECT 14.030000  70.105000 65.364000  70.175000 ;
      RECT 14.030000  70.175000 65.294000  70.245000 ;
      RECT 14.030000  70.175000 65.294000  70.245000 ;
      RECT 14.030000  70.245000 65.224000  70.315000 ;
      RECT 14.030000  70.245000 65.224000  70.315000 ;
      RECT 14.030000  70.315000 65.154000  70.385000 ;
      RECT 14.030000  70.315000 65.154000  70.385000 ;
      RECT 14.030000  70.385000 65.084000  70.455000 ;
      RECT 14.030000  70.385000 65.084000  70.455000 ;
      RECT 14.030000  70.455000 65.014000  70.525000 ;
      RECT 14.030000  70.455000 65.014000  70.525000 ;
      RECT 14.030000  70.525000 64.944000  70.595000 ;
      RECT 14.030000  70.525000 64.944000  70.595000 ;
      RECT 14.030000  70.595000 64.874000  70.665000 ;
      RECT 14.030000  70.595000 64.874000  70.665000 ;
      RECT 14.030000  70.665000 64.829000  70.710000 ;
      RECT 14.030000  70.665000 64.829000  70.710000 ;
      RECT 14.030000  70.710000 15.855000  73.910000 ;
      RECT 14.030000  70.850000 15.995000  73.770000 ;
      RECT 14.030000  73.770000 65.551000  74.179000 ;
      RECT 14.030000  73.910000 65.084000  73.980000 ;
      RECT 14.030000  73.980000 65.154000  74.050000 ;
      RECT 14.030000  74.050000 65.224000  74.120000 ;
      RECT 14.030000  74.120000 65.294000  74.180000 ;
      RECT 14.030000  74.179000 65.761000  74.389000 ;
      RECT 14.066000  25.265000 65.429000  25.300000 ;
      RECT 14.066000  25.265000 65.429000  25.300000 ;
      RECT 14.101000  74.179000 65.353000  74.250000 ;
      RECT 14.136000  25.195000 65.359000  25.265000 ;
      RECT 14.136000  25.195000 65.359000  25.265000 ;
      RECT 14.171000  74.250000 65.424000  74.320000 ;
      RECT 14.206000  25.125000 65.289000  25.195000 ;
      RECT 14.206000  25.125000 65.289000  25.195000 ;
      RECT 14.240000  73.910000 65.084000  73.980000 ;
      RECT 14.240000  73.910000 65.084000  73.980000 ;
      RECT 14.240000  73.980000 65.154000  74.050000 ;
      RECT 14.240000  73.980000 65.154000  74.050000 ;
      RECT 14.240000  74.050000 65.224000  74.120000 ;
      RECT 14.240000  74.050000 65.224000  74.120000 ;
      RECT 14.240000  74.120000 65.294000  74.180000 ;
      RECT 14.240000  74.120000 65.294000  74.180000 ;
      RECT 14.240000  74.179000 65.353000  74.250000 ;
      RECT 14.240000  74.179000 65.353000  74.250000 ;
      RECT 14.240000  74.250000 65.424000  74.320000 ;
      RECT 14.240000  74.250000 65.424000  74.320000 ;
      RECT 14.240000  74.320000 65.494000  74.390000 ;
      RECT 14.240000  74.320000 65.494000  74.390000 ;
      RECT 14.240000  74.389000 65.563000  74.460000 ;
      RECT 14.240000  74.389000 65.563000  74.460000 ;
      RECT 14.240000  74.389000 65.860000  74.488000 ;
      RECT 14.240000  74.460000 65.634000  74.530000 ;
      RECT 14.240000  74.460000 65.634000  74.530000 ;
      RECT 14.240000  74.488000 65.860000  98.700000 ;
      RECT 14.240000  74.530000 65.704000  74.545000 ;
      RECT 14.240000  74.530000 65.704000  74.545000 ;
      RECT 14.240000  74.546000 65.720000  98.840000 ;
      RECT 14.240000  98.700000 75.000000 129.819000 ;
      RECT 14.240000  98.840000 75.000000 129.819000 ;
      RECT 14.240000 129.819000 75.000000 130.705000 ;
      RECT 14.240000 134.796000 75.000000 139.824000 ;
      RECT 14.240000 134.796000 75.000000 139.824000 ;
      RECT 14.240000 139.824000 75.000000 140.710000 ;
      RECT 14.240000 144.796000 75.000000 149.824000 ;
      RECT 14.240000 144.796000 75.000000 149.824000 ;
      RECT 14.240000 149.824000 75.000000 150.710000 ;
      RECT 14.240000 154.796000 75.000000 159.824000 ;
      RECT 14.240000 154.796000 75.000000 159.824000 ;
      RECT 14.240000 159.824000 75.000000 160.710000 ;
      RECT 14.240000 164.796000 75.000000 169.824000 ;
      RECT 14.240000 164.796000 75.000000 169.824000 ;
      RECT 14.240000 169.824000 75.000000 170.710000 ;
      RECT 14.240000 174.796000 75.000000 179.824000 ;
      RECT 14.240000 174.796000 75.000000 179.824000 ;
      RECT 14.240000 179.824000 75.000000 180.710000 ;
      RECT 14.240000 184.796000 75.000000 189.824000 ;
      RECT 14.240000 184.796000 75.000000 189.824000 ;
      RECT 14.240000 189.824000 75.000000 190.710000 ;
      RECT 14.241000  74.320000 65.494000  74.390000 ;
      RECT 14.276000  25.055000 65.219000  25.125000 ;
      RECT 14.276000  25.055000 65.219000  25.125000 ;
      RECT 14.286000 134.750000 75.000000 134.795000 ;
      RECT 14.286000 134.750000 75.000000 134.795000 ;
      RECT 14.286000 144.750000 75.000000 144.795000 ;
      RECT 14.286000 144.750000 75.000000 144.795000 ;
      RECT 14.286000 154.750000 75.000000 154.795000 ;
      RECT 14.286000 154.750000 75.000000 154.795000 ;
      RECT 14.286000 164.750000 75.000000 164.795000 ;
      RECT 14.286000 164.750000 75.000000 164.795000 ;
      RECT 14.286000 174.750000 75.000000 174.795000 ;
      RECT 14.286000 174.750000 75.000000 174.795000 ;
      RECT 14.286000 184.750000 75.000000 184.795000 ;
      RECT 14.286000 184.750000 75.000000 184.795000 ;
      RECT 14.311000 129.819000 75.000000 129.890000 ;
      RECT 14.311000 129.819000 75.000000 129.890000 ;
      RECT 14.311000 139.824000 75.000000 139.895000 ;
      RECT 14.311000 139.824000 75.000000 139.895000 ;
      RECT 14.311000 149.824000 75.000000 149.895000 ;
      RECT 14.311000 149.824000 75.000000 149.895000 ;
      RECT 14.311000 159.824000 75.000000 159.895000 ;
      RECT 14.311000 159.824000 75.000000 159.895000 ;
      RECT 14.311000 169.824000 75.000000 169.895000 ;
      RECT 14.311000 169.824000 75.000000 169.895000 ;
      RECT 14.311000 179.824000 75.000000 179.895000 ;
      RECT 14.311000 179.824000 75.000000 179.895000 ;
      RECT 14.311000 189.824000 75.000000 189.895000 ;
      RECT 14.311000 189.824000 75.000000 189.895000 ;
      RECT 14.346000  24.985000 65.149000  25.055000 ;
      RECT 14.346000  24.985000 65.149000  25.055000 ;
      RECT 14.356000 134.680000 75.000000 134.750000 ;
      RECT 14.356000 134.680000 75.000000 134.750000 ;
      RECT 14.356000 144.680000 75.000000 144.750000 ;
      RECT 14.356000 144.680000 75.000000 144.750000 ;
      RECT 14.356000 154.680000 75.000000 154.750000 ;
      RECT 14.356000 154.680000 75.000000 154.750000 ;
      RECT 14.356000 164.680000 75.000000 164.750000 ;
      RECT 14.356000 164.680000 75.000000 164.750000 ;
      RECT 14.356000 174.680000 75.000000 174.750000 ;
      RECT 14.356000 174.680000 75.000000 174.750000 ;
      RECT 14.356000 184.680000 75.000000 184.750000 ;
      RECT 14.356000 184.680000 75.000000 184.750000 ;
      RECT 14.381000 129.890000 75.000000 129.960000 ;
      RECT 14.381000 129.890000 75.000000 129.960000 ;
      RECT 14.381000 139.895000 75.000000 139.965000 ;
      RECT 14.381000 139.895000 75.000000 139.965000 ;
      RECT 14.381000 149.895000 75.000000 149.965000 ;
      RECT 14.381000 149.895000 75.000000 149.965000 ;
      RECT 14.381000 159.895000 75.000000 159.965000 ;
      RECT 14.381000 159.895000 75.000000 159.965000 ;
      RECT 14.381000 169.895000 75.000000 169.965000 ;
      RECT 14.381000 169.895000 75.000000 169.965000 ;
      RECT 14.381000 179.895000 75.000000 179.965000 ;
      RECT 14.381000 179.895000 75.000000 179.965000 ;
      RECT 14.381000 189.895000 75.000000 189.965000 ;
      RECT 14.381000 189.895000 75.000000 189.965000 ;
      RECT 14.416000  24.915000 65.079000  24.985000 ;
      RECT 14.416000  24.915000 65.079000  24.985000 ;
      RECT 14.426000 134.610000 75.000000 134.680000 ;
      RECT 14.426000 134.610000 75.000000 134.680000 ;
      RECT 14.426000 144.610000 75.000000 144.680000 ;
      RECT 14.426000 144.610000 75.000000 144.680000 ;
      RECT 14.426000 154.610000 75.000000 154.680000 ;
      RECT 14.426000 154.610000 75.000000 154.680000 ;
      RECT 14.426000 164.610000 75.000000 164.680000 ;
      RECT 14.426000 164.610000 75.000000 164.680000 ;
      RECT 14.426000 174.610000 75.000000 174.680000 ;
      RECT 14.426000 174.610000 75.000000 174.680000 ;
      RECT 14.426000 184.610000 75.000000 184.680000 ;
      RECT 14.426000 184.610000 75.000000 184.680000 ;
      RECT 14.451000 129.960000 75.000000 130.030000 ;
      RECT 14.451000 129.960000 75.000000 130.030000 ;
      RECT 14.451000 139.965000 75.000000 140.035000 ;
      RECT 14.451000 139.965000 75.000000 140.035000 ;
      RECT 14.451000 149.965000 75.000000 150.035000 ;
      RECT 14.451000 149.965000 75.000000 150.035000 ;
      RECT 14.451000 159.965000 75.000000 160.035000 ;
      RECT 14.451000 159.965000 75.000000 160.035000 ;
      RECT 14.451000 169.965000 75.000000 170.035000 ;
      RECT 14.451000 169.965000 75.000000 170.035000 ;
      RECT 14.451000 179.965000 75.000000 180.035000 ;
      RECT 14.451000 179.965000 75.000000 180.035000 ;
      RECT 14.451000 189.965000 75.000000 190.035000 ;
      RECT 14.451000 189.965000 75.000000 190.035000 ;
      RECT 14.486000  24.845000 65.009000  24.915000 ;
      RECT 14.486000  24.845000 65.009000  24.915000 ;
      RECT 14.496000 134.540000 75.000000 134.610000 ;
      RECT 14.496000 134.540000 75.000000 134.610000 ;
      RECT 14.496000 144.540000 75.000000 144.610000 ;
      RECT 14.496000 144.540000 75.000000 144.610000 ;
      RECT 14.496000 154.540000 75.000000 154.610000 ;
      RECT 14.496000 154.540000 75.000000 154.610000 ;
      RECT 14.496000 164.540000 75.000000 164.610000 ;
      RECT 14.496000 164.540000 75.000000 164.610000 ;
      RECT 14.496000 174.540000 75.000000 174.610000 ;
      RECT 14.496000 174.540000 75.000000 174.610000 ;
      RECT 14.496000 184.540000 75.000000 184.610000 ;
      RECT 14.496000 184.540000 75.000000 184.610000 ;
      RECT 14.521000 130.030000 75.000000 130.100000 ;
      RECT 14.521000 130.030000 75.000000 130.100000 ;
      RECT 14.521000 140.035000 75.000000 140.105000 ;
      RECT 14.521000 140.035000 75.000000 140.105000 ;
      RECT 14.521000 150.035000 75.000000 150.105000 ;
      RECT 14.521000 150.035000 75.000000 150.105000 ;
      RECT 14.521000 160.035000 75.000000 160.105000 ;
      RECT 14.521000 160.035000 75.000000 160.105000 ;
      RECT 14.521000 170.035000 75.000000 170.105000 ;
      RECT 14.521000 170.035000 75.000000 170.105000 ;
      RECT 14.521000 180.035000 75.000000 180.105000 ;
      RECT 14.521000 180.035000 75.000000 180.105000 ;
      RECT 14.521000 190.035000 75.000000 190.105000 ;
      RECT 14.521000 190.035000 75.000000 190.105000 ;
      RECT 14.556000  24.775000 64.939000  24.845000 ;
      RECT 14.556000  24.775000 64.939000  24.845000 ;
      RECT 14.566000 134.470000 75.000000 134.540000 ;
      RECT 14.566000 134.470000 75.000000 134.540000 ;
      RECT 14.566000 144.470000 75.000000 144.540000 ;
      RECT 14.566000 144.470000 75.000000 144.540000 ;
      RECT 14.566000 154.470000 75.000000 154.540000 ;
      RECT 14.566000 154.470000 75.000000 154.540000 ;
      RECT 14.566000 164.470000 75.000000 164.540000 ;
      RECT 14.566000 164.470000 75.000000 164.540000 ;
      RECT 14.566000 174.470000 75.000000 174.540000 ;
      RECT 14.566000 174.470000 75.000000 174.540000 ;
      RECT 14.566000 184.470000 75.000000 184.540000 ;
      RECT 14.566000 184.470000 75.000000 184.540000 ;
      RECT 14.591000 130.100000 75.000000 130.170000 ;
      RECT 14.591000 130.100000 75.000000 130.170000 ;
      RECT 14.591000 140.105000 75.000000 140.175000 ;
      RECT 14.591000 140.105000 75.000000 140.175000 ;
      RECT 14.591000 150.105000 75.000000 150.175000 ;
      RECT 14.591000 150.105000 75.000000 150.175000 ;
      RECT 14.591000 160.105000 75.000000 160.175000 ;
      RECT 14.591000 160.105000 75.000000 160.175000 ;
      RECT 14.591000 170.105000 75.000000 170.175000 ;
      RECT 14.591000 170.105000 75.000000 170.175000 ;
      RECT 14.591000 180.105000 75.000000 180.175000 ;
      RECT 14.591000 180.105000 75.000000 180.175000 ;
      RECT 14.591000 190.105000 75.000000 190.175000 ;
      RECT 14.591000 190.105000 75.000000 190.175000 ;
      RECT 14.626000  24.705000 64.869000  24.775000 ;
      RECT 14.626000  24.705000 64.869000  24.775000 ;
      RECT 14.636000 134.400000 75.000000 134.470000 ;
      RECT 14.636000 134.400000 75.000000 134.470000 ;
      RECT 14.636000 144.400000 75.000000 144.470000 ;
      RECT 14.636000 144.400000 75.000000 144.470000 ;
      RECT 14.636000 154.400000 75.000000 154.470000 ;
      RECT 14.636000 154.400000 75.000000 154.470000 ;
      RECT 14.636000 164.400000 75.000000 164.470000 ;
      RECT 14.636000 164.400000 75.000000 164.470000 ;
      RECT 14.636000 174.400000 75.000000 174.470000 ;
      RECT 14.636000 174.400000 75.000000 174.470000 ;
      RECT 14.636000 184.400000 75.000000 184.470000 ;
      RECT 14.636000 184.400000 75.000000 184.470000 ;
      RECT 14.661000 130.170000 75.000000 130.240000 ;
      RECT 14.661000 130.170000 75.000000 130.240000 ;
      RECT 14.661000 140.175000 75.000000 140.245000 ;
      RECT 14.661000 140.175000 75.000000 140.245000 ;
      RECT 14.661000 150.175000 75.000000 150.245000 ;
      RECT 14.661000 150.175000 75.000000 150.245000 ;
      RECT 14.661000 160.175000 75.000000 160.245000 ;
      RECT 14.661000 160.175000 75.000000 160.245000 ;
      RECT 14.661000 170.175000 75.000000 170.245000 ;
      RECT 14.661000 170.175000 75.000000 170.245000 ;
      RECT 14.661000 180.175000 75.000000 180.245000 ;
      RECT 14.661000 180.175000 75.000000 180.245000 ;
      RECT 14.661000 190.175000 75.000000 190.245000 ;
      RECT 14.661000 190.175000 75.000000 190.245000 ;
      RECT 14.696000  24.635000 64.799000  24.705000 ;
      RECT 14.696000  24.635000 64.799000  24.705000 ;
      RECT 14.706000 134.330000 75.000000 134.400000 ;
      RECT 14.706000 134.330000 75.000000 134.400000 ;
      RECT 14.706000 144.330000 75.000000 144.400000 ;
      RECT 14.706000 144.330000 75.000000 144.400000 ;
      RECT 14.706000 154.330000 75.000000 154.400000 ;
      RECT 14.706000 154.330000 75.000000 154.400000 ;
      RECT 14.706000 164.330000 75.000000 164.400000 ;
      RECT 14.706000 164.330000 75.000000 164.400000 ;
      RECT 14.706000 174.330000 75.000000 174.400000 ;
      RECT 14.706000 174.330000 75.000000 174.400000 ;
      RECT 14.706000 184.330000 75.000000 184.400000 ;
      RECT 14.706000 184.330000 75.000000 184.400000 ;
      RECT 14.731000 130.240000 75.000000 130.310000 ;
      RECT 14.731000 130.240000 75.000000 130.310000 ;
      RECT 14.731000 140.245000 75.000000 140.315000 ;
      RECT 14.731000 140.245000 75.000000 140.315000 ;
      RECT 14.731000 150.245000 75.000000 150.315000 ;
      RECT 14.731000 150.245000 75.000000 150.315000 ;
      RECT 14.731000 160.245000 75.000000 160.315000 ;
      RECT 14.731000 160.245000 75.000000 160.315000 ;
      RECT 14.731000 170.245000 75.000000 170.315000 ;
      RECT 14.731000 170.245000 75.000000 170.315000 ;
      RECT 14.731000 180.245000 75.000000 180.315000 ;
      RECT 14.731000 180.245000 75.000000 180.315000 ;
      RECT 14.731000 190.245000 75.000000 190.315000 ;
      RECT 14.731000 190.245000 75.000000 190.315000 ;
      RECT 14.766000  24.565000 64.729000  24.635000 ;
      RECT 14.766000  24.565000 64.729000  24.635000 ;
      RECT 14.776000 134.260000 75.000000 134.330000 ;
      RECT 14.776000 134.260000 75.000000 134.330000 ;
      RECT 14.776000 144.260000 75.000000 144.330000 ;
      RECT 14.776000 144.260000 75.000000 144.330000 ;
      RECT 14.776000 154.260000 75.000000 154.330000 ;
      RECT 14.776000 154.260000 75.000000 154.330000 ;
      RECT 14.776000 164.260000 75.000000 164.330000 ;
      RECT 14.776000 164.260000 75.000000 164.330000 ;
      RECT 14.776000 174.260000 75.000000 174.330000 ;
      RECT 14.776000 174.260000 75.000000 174.330000 ;
      RECT 14.776000 184.260000 75.000000 184.330000 ;
      RECT 14.776000 184.260000 75.000000 184.330000 ;
      RECT 14.801000 130.310000 75.000000 130.380000 ;
      RECT 14.801000 130.310000 75.000000 130.380000 ;
      RECT 14.801000 140.315000 75.000000 140.385000 ;
      RECT 14.801000 140.315000 75.000000 140.385000 ;
      RECT 14.801000 150.315000 75.000000 150.385000 ;
      RECT 14.801000 150.315000 75.000000 150.385000 ;
      RECT 14.801000 160.315000 75.000000 160.385000 ;
      RECT 14.801000 160.315000 75.000000 160.385000 ;
      RECT 14.801000 170.315000 75.000000 170.385000 ;
      RECT 14.801000 170.315000 75.000000 170.385000 ;
      RECT 14.801000 180.315000 75.000000 180.385000 ;
      RECT 14.801000 180.315000 75.000000 180.385000 ;
      RECT 14.801000 190.315000 75.000000 190.385000 ;
      RECT 14.801000 190.315000 75.000000 190.385000 ;
      RECT 14.836000  24.495000 64.659000  24.565000 ;
      RECT 14.836000  24.495000 64.659000  24.565000 ;
      RECT 14.846000 134.190000 75.000000 134.260000 ;
      RECT 14.846000 134.190000 75.000000 134.260000 ;
      RECT 14.846000 144.190000 75.000000 144.260000 ;
      RECT 14.846000 144.190000 75.000000 144.260000 ;
      RECT 14.846000 154.190000 75.000000 154.260000 ;
      RECT 14.846000 154.190000 75.000000 154.260000 ;
      RECT 14.846000 164.190000 75.000000 164.260000 ;
      RECT 14.846000 164.190000 75.000000 164.260000 ;
      RECT 14.846000 174.190000 75.000000 174.260000 ;
      RECT 14.846000 174.190000 75.000000 174.260000 ;
      RECT 14.846000 184.190000 75.000000 184.260000 ;
      RECT 14.846000 184.190000 75.000000 184.260000 ;
      RECT 14.871000 130.380000 75.000000 130.450000 ;
      RECT 14.871000 130.380000 75.000000 130.450000 ;
      RECT 14.871000 140.385000 75.000000 140.455000 ;
      RECT 14.871000 140.385000 75.000000 140.455000 ;
      RECT 14.871000 150.385000 75.000000 150.455000 ;
      RECT 14.871000 150.385000 75.000000 150.455000 ;
      RECT 14.871000 160.385000 75.000000 160.455000 ;
      RECT 14.871000 160.385000 75.000000 160.455000 ;
      RECT 14.871000 170.385000 75.000000 170.455000 ;
      RECT 14.871000 170.385000 75.000000 170.455000 ;
      RECT 14.871000 180.385000 75.000000 180.455000 ;
      RECT 14.871000 180.385000 75.000000 180.455000 ;
      RECT 14.871000 190.385000 75.000000 190.455000 ;
      RECT 14.871000 190.385000 75.000000 190.455000 ;
      RECT 14.906000  24.425000 64.589000  24.495000 ;
      RECT 14.906000  24.425000 64.589000  24.495000 ;
      RECT 14.916000 134.120000 75.000000 134.190000 ;
      RECT 14.916000 134.120000 75.000000 134.190000 ;
      RECT 14.916000 144.120000 75.000000 144.190000 ;
      RECT 14.916000 144.120000 75.000000 144.190000 ;
      RECT 14.916000 154.120000 75.000000 154.190000 ;
      RECT 14.916000 154.120000 75.000000 154.190000 ;
      RECT 14.916000 164.120000 75.000000 164.190000 ;
      RECT 14.916000 164.120000 75.000000 164.190000 ;
      RECT 14.916000 174.120000 75.000000 174.190000 ;
      RECT 14.916000 174.120000 75.000000 174.190000 ;
      RECT 14.916000 184.120000 75.000000 184.190000 ;
      RECT 14.916000 184.120000 75.000000 184.190000 ;
      RECT 14.941000 130.450000 75.000000 130.520000 ;
      RECT 14.941000 130.450000 75.000000 130.520000 ;
      RECT 14.941000 140.455000 75.000000 140.525000 ;
      RECT 14.941000 140.455000 75.000000 140.525000 ;
      RECT 14.941000 150.455000 75.000000 150.525000 ;
      RECT 14.941000 150.455000 75.000000 150.525000 ;
      RECT 14.941000 160.455000 75.000000 160.525000 ;
      RECT 14.941000 160.455000 75.000000 160.525000 ;
      RECT 14.941000 170.455000 75.000000 170.525000 ;
      RECT 14.941000 170.455000 75.000000 170.525000 ;
      RECT 14.941000 180.455000 75.000000 180.525000 ;
      RECT 14.941000 180.455000 75.000000 180.525000 ;
      RECT 14.941000 190.455000 75.000000 190.525000 ;
      RECT 14.941000 190.455000 75.000000 190.525000 ;
      RECT 14.976000  24.355000 64.519000  24.425000 ;
      RECT 14.976000  24.355000 64.519000  24.425000 ;
      RECT 14.986000 134.050000 75.000000 134.120000 ;
      RECT 14.986000 134.050000 75.000000 134.120000 ;
      RECT 14.986000 144.050000 75.000000 144.120000 ;
      RECT 14.986000 144.050000 75.000000 144.120000 ;
      RECT 14.986000 154.050000 75.000000 154.120000 ;
      RECT 14.986000 154.050000 75.000000 154.120000 ;
      RECT 14.986000 164.050000 75.000000 164.120000 ;
      RECT 14.986000 164.050000 75.000000 164.120000 ;
      RECT 14.986000 174.050000 75.000000 174.120000 ;
      RECT 14.986000 174.050000 75.000000 174.120000 ;
      RECT 14.986000 184.050000 75.000000 184.120000 ;
      RECT 14.986000 184.050000 75.000000 184.120000 ;
      RECT 15.011000 130.520000 75.000000 130.590000 ;
      RECT 15.011000 130.520000 75.000000 130.590000 ;
      RECT 15.011000 140.525000 75.000000 140.595000 ;
      RECT 15.011000 140.525000 75.000000 140.595000 ;
      RECT 15.011000 150.525000 75.000000 150.595000 ;
      RECT 15.011000 150.525000 75.000000 150.595000 ;
      RECT 15.011000 160.525000 75.000000 160.595000 ;
      RECT 15.011000 160.525000 75.000000 160.595000 ;
      RECT 15.011000 170.525000 75.000000 170.595000 ;
      RECT 15.011000 170.525000 75.000000 170.595000 ;
      RECT 15.011000 180.525000 75.000000 180.595000 ;
      RECT 15.011000 180.525000 75.000000 180.595000 ;
      RECT 15.011000 190.525000 75.000000 190.595000 ;
      RECT 15.011000 190.525000 75.000000 190.595000 ;
      RECT 15.046000  24.285000 64.449000  24.355000 ;
      RECT 15.046000  24.285000 64.449000  24.355000 ;
      RECT 15.056000 133.980000 75.000000 134.050000 ;
      RECT 15.056000 133.980000 75.000000 134.050000 ;
      RECT 15.056000 143.980000 75.000000 144.050000 ;
      RECT 15.056000 143.980000 75.000000 144.050000 ;
      RECT 15.056000 153.980000 75.000000 154.050000 ;
      RECT 15.056000 153.980000 75.000000 154.050000 ;
      RECT 15.056000 163.980000 75.000000 164.050000 ;
      RECT 15.056000 163.980000 75.000000 164.050000 ;
      RECT 15.056000 173.980000 75.000000 174.050000 ;
      RECT 15.056000 173.980000 75.000000 174.050000 ;
      RECT 15.056000 183.980000 75.000000 184.050000 ;
      RECT 15.056000 183.980000 75.000000 184.050000 ;
      RECT 15.081000 130.590000 75.000000 130.660000 ;
      RECT 15.081000 130.590000 75.000000 130.660000 ;
      RECT 15.081000 140.595000 75.000000 140.665000 ;
      RECT 15.081000 140.595000 75.000000 140.665000 ;
      RECT 15.081000 150.595000 75.000000 150.665000 ;
      RECT 15.081000 150.595000 75.000000 150.665000 ;
      RECT 15.081000 160.595000 75.000000 160.665000 ;
      RECT 15.081000 160.595000 75.000000 160.665000 ;
      RECT 15.081000 170.595000 75.000000 170.665000 ;
      RECT 15.081000 170.595000 75.000000 170.665000 ;
      RECT 15.081000 180.595000 75.000000 180.665000 ;
      RECT 15.081000 180.595000 75.000000 180.665000 ;
      RECT 15.081000 190.595000 75.000000 190.665000 ;
      RECT 15.081000 190.595000 75.000000 190.665000 ;
      RECT 15.116000  24.215000 64.379000  24.285000 ;
      RECT 15.116000  24.215000 64.379000  24.285000 ;
      RECT 15.126000 130.660000 75.000000 130.705000 ;
      RECT 15.126000 130.660000 75.000000 130.705000 ;
      RECT 15.126000 133.910000 75.000000 133.980000 ;
      RECT 15.126000 133.910000 75.000000 133.980000 ;
      RECT 15.126000 133.910000 75.000000 134.796000 ;
      RECT 15.126000 140.665000 75.000000 140.710000 ;
      RECT 15.126000 140.665000 75.000000 140.710000 ;
      RECT 15.126000 143.910000 75.000000 143.980000 ;
      RECT 15.126000 143.910000 75.000000 143.980000 ;
      RECT 15.126000 143.910000 75.000000 144.796000 ;
      RECT 15.126000 150.665000 75.000000 150.710000 ;
      RECT 15.126000 150.665000 75.000000 150.710000 ;
      RECT 15.126000 153.910000 75.000000 153.980000 ;
      RECT 15.126000 153.910000 75.000000 153.980000 ;
      RECT 15.126000 153.910000 75.000000 154.796000 ;
      RECT 15.126000 160.665000 75.000000 160.710000 ;
      RECT 15.126000 160.665000 75.000000 160.710000 ;
      RECT 15.126000 163.910000 75.000000 163.980000 ;
      RECT 15.126000 163.910000 75.000000 163.980000 ;
      RECT 15.126000 163.910000 75.000000 164.796000 ;
      RECT 15.126000 170.665000 75.000000 170.710000 ;
      RECT 15.126000 170.665000 75.000000 170.710000 ;
      RECT 15.126000 173.910000 75.000000 173.980000 ;
      RECT 15.126000 173.910000 75.000000 173.980000 ;
      RECT 15.126000 173.910000 75.000000 174.796000 ;
      RECT 15.126000 180.665000 75.000000 180.710000 ;
      RECT 15.126000 180.665000 75.000000 180.710000 ;
      RECT 15.126000 183.910000 75.000000 183.980000 ;
      RECT 15.126000 183.910000 75.000000 183.980000 ;
      RECT 15.126000 183.910000 75.000000 184.796000 ;
      RECT 15.126000 190.665000 75.000000 190.710000 ;
      RECT 15.126000 190.665000 75.000000 190.710000 ;
      RECT 15.186000  24.145000 64.309000  24.215000 ;
      RECT 15.186000  24.145000 64.309000  24.215000 ;
      RECT 15.256000  24.075000 64.239000  24.145000 ;
      RECT 15.256000  24.075000 64.239000  24.145000 ;
      RECT 15.326000  24.005000 64.169000  24.075000 ;
      RECT 15.326000  24.005000 64.169000  24.075000 ;
      RECT 15.396000  23.935000 64.099000  24.005000 ;
      RECT 15.396000  23.935000 64.099000  24.005000 ;
      RECT 15.466000  23.865000 64.029000  23.935000 ;
      RECT 15.466000  23.865000 64.029000  23.935000 ;
      RECT 15.522000 130.705000 75.000000 130.845000 ;
      RECT 15.522000 140.710000 75.000000 140.850000 ;
      RECT 15.522000 150.710000 75.000000 150.850000 ;
      RECT 15.522000 160.710000 75.000000 160.850000 ;
      RECT 15.522000 170.710000 75.000000 170.850000 ;
      RECT 15.522000 180.710000 75.000000 180.850000 ;
      RECT 15.522000 190.710000 75.000000 190.850000 ;
      RECT 15.536000  23.795000 63.959000  23.865000 ;
      RECT 15.536000  23.795000 63.959000  23.865000 ;
      RECT 15.606000  23.725000 63.889000  23.795000 ;
      RECT 15.606000  23.725000 63.889000  23.795000 ;
      RECT 15.662000 133.770000 75.000000 133.910000 ;
      RECT 15.662000 143.770000 75.000000 143.910000 ;
      RECT 15.662000 153.770000 75.000000 153.910000 ;
      RECT 15.662000 163.770000 75.000000 163.910000 ;
      RECT 15.662000 173.770000 75.000000 173.910000 ;
      RECT 15.662000 183.770000 75.000000 183.910000 ;
      RECT 15.676000  23.655000 63.819000  23.725000 ;
      RECT 15.676000  23.655000 63.819000  23.725000 ;
      RECT 15.746000  23.585000 63.749000  23.655000 ;
      RECT 15.746000  23.585000 63.749000  23.655000 ;
      RECT 15.816000  23.515000 63.679000  23.585000 ;
      RECT 15.816000  23.515000 63.679000  23.585000 ;
      RECT 15.886000  23.445000 63.609000  23.515000 ;
      RECT 15.886000  23.445000 63.609000  23.515000 ;
      RECT 15.956000  23.375000 63.539000  23.445000 ;
      RECT 15.956000  23.375000 63.539000  23.445000 ;
      RECT 16.026000  23.305000 63.469000  23.375000 ;
      RECT 16.026000  23.305000 63.469000  23.375000 ;
      RECT 16.096000  23.235000 63.399000  23.305000 ;
      RECT 16.096000  23.235000 63.399000  23.305000 ;
      RECT 16.166000  23.165000 63.329000  23.235000 ;
      RECT 16.166000  23.165000 63.329000  23.235000 ;
      RECT 16.236000  23.095000 63.259000  23.165000 ;
      RECT 16.236000  23.095000 63.259000  23.165000 ;
      RECT 16.306000  23.025000 63.189000  23.095000 ;
      RECT 16.306000  23.025000 63.189000  23.095000 ;
      RECT 16.376000  22.955000 63.119000  23.025000 ;
      RECT 16.376000  22.955000 63.119000  23.025000 ;
      RECT 16.446000  22.885000 63.049000  22.955000 ;
      RECT 16.446000  22.885000 63.049000  22.955000 ;
      RECT 16.516000  22.815000 62.979000  22.885000 ;
      RECT 16.516000  22.815000 62.979000  22.885000 ;
      RECT 16.586000  22.745000 62.909000  22.815000 ;
      RECT 16.586000  22.745000 62.909000  22.815000 ;
      RECT 16.656000  22.675000 62.839000  22.745000 ;
      RECT 16.656000  22.675000 62.839000  22.745000 ;
      RECT 16.726000  22.605000 62.769000  22.675000 ;
      RECT 16.726000  22.605000 62.769000  22.675000 ;
      RECT 16.796000  22.535000 62.699000  22.605000 ;
      RECT 16.796000  22.535000 62.699000  22.605000 ;
      RECT 16.866000  22.465000 62.629000  22.535000 ;
      RECT 16.866000  22.465000 62.629000  22.535000 ;
      RECT 16.936000  22.395000 62.559000  22.465000 ;
      RECT 16.936000  22.395000 62.559000  22.465000 ;
      RECT 17.006000  22.325000 62.489000  22.395000 ;
      RECT 17.006000  22.325000 62.489000  22.395000 ;
      RECT 17.076000  22.255000 62.419000  22.325000 ;
      RECT 17.076000  22.255000 62.419000  22.325000 ;
      RECT 17.140000   5.236000 17.350000   9.249000 ;
      RECT 17.140000   5.236000 17.490000   9.249000 ;
      RECT 17.140000   9.249000 17.490000   9.599000 ;
      RECT 17.146000  22.185000 62.349000  22.255000 ;
      RECT 17.146000  22.185000 62.349000  22.255000 ;
      RECT 17.211000   5.165000 17.350000   5.235000 ;
      RECT 17.211000   9.249000 17.350000   9.320000 ;
      RECT 17.216000  22.115000 62.279000  22.185000 ;
      RECT 17.216000  22.115000 62.279000  22.185000 ;
      RECT 17.281000   5.095000 17.350000   5.165000 ;
      RECT 17.281000   9.320000 17.350000   9.390000 ;
      RECT 17.286000  22.045000 62.209000  22.115000 ;
      RECT 17.286000  22.045000 62.209000  22.115000 ;
      RECT 17.319000   5.057000 17.490000   5.236000 ;
      RECT 17.356000  21.975000 62.139000  22.045000 ;
      RECT 17.356000  21.975000 62.139000  22.045000 ;
      RECT 17.426000  21.905000 53.815000  21.975000 ;
      RECT 17.426000  21.905000 53.815000  21.975000 ;
      RECT 17.496000  21.835000 53.815000  21.905000 ;
      RECT 17.496000  21.835000 53.815000  21.905000 ;
      RECT 17.496000  21.835000 65.663000  25.301000 ;
      RECT 17.566000  21.765000 53.815000  21.835000 ;
      RECT 17.566000  21.765000 53.815000  21.835000 ;
      RECT 17.571000   9.680000 55.882000   9.800000 ;
      RECT 17.636000  21.695000 53.815000  21.765000 ;
      RECT 17.636000  21.695000 53.815000  21.765000 ;
      RECT 17.706000  21.625000 53.815000  21.695000 ;
      RECT 17.706000  21.625000 53.815000  21.695000 ;
      RECT 17.776000  21.555000 53.815000  21.625000 ;
      RECT 17.776000  21.555000 53.815000  21.625000 ;
      RECT 17.846000  21.485000 53.815000  21.555000 ;
      RECT 17.846000  21.485000 53.815000  21.555000 ;
      RECT 17.916000  21.415000 53.815000  21.485000 ;
      RECT 17.916000  21.415000 53.815000  21.485000 ;
      RECT 17.986000  21.345000 53.815000  21.415000 ;
      RECT 17.986000  21.345000 53.815000  21.415000 ;
      RECT 18.056000  21.275000 53.815000  21.345000 ;
      RECT 18.056000  21.275000 53.815000  21.345000 ;
      RECT 18.126000  21.205000 53.815000  21.275000 ;
      RECT 18.126000  21.205000 53.815000  21.275000 ;
      RECT 18.196000  21.135000 53.815000  21.205000 ;
      RECT 18.196000  21.135000 53.815000  21.205000 ;
      RECT 18.266000  21.065000 53.815000  21.135000 ;
      RECT 18.266000  21.065000 53.815000  21.135000 ;
      RECT 18.336000  20.995000 53.815000  21.065000 ;
      RECT 18.336000  20.995000 53.815000  21.065000 ;
      RECT 18.406000  20.925000 53.815000  20.995000 ;
      RECT 18.406000  20.925000 53.815000  20.995000 ;
      RECT 18.476000  20.855000 53.815000  20.925000 ;
      RECT 18.476000  20.855000 53.815000  20.925000 ;
      RECT 18.546000  20.785000 53.815000  20.855000 ;
      RECT 18.546000  20.785000 53.815000  20.855000 ;
      RECT 18.582000 193.770000 75.000000 193.910000 ;
      RECT 18.616000  20.715000 53.815000  20.785000 ;
      RECT 18.616000  20.715000 53.815000  20.785000 ;
      RECT 18.686000  20.645000 53.815000  20.715000 ;
      RECT 18.686000  20.645000 53.815000  20.715000 ;
      RECT 18.756000  20.575000 53.815000  20.645000 ;
      RECT 18.756000  20.575000 53.815000  20.645000 ;
      RECT 18.826000  20.505000 53.815000  20.575000 ;
      RECT 18.826000  20.505000 53.815000  20.575000 ;
      RECT 18.896000  20.435000 53.815000  20.505000 ;
      RECT 18.896000  20.435000 53.815000  20.505000 ;
      RECT 18.966000  20.365000 53.815000  20.435000 ;
      RECT 18.966000  20.365000 53.815000  20.435000 ;
      RECT 19.036000  20.295000 53.815000  20.365000 ;
      RECT 19.036000  20.295000 53.815000  20.365000 ;
      RECT 19.106000  20.225000 53.815000  20.295000 ;
      RECT 19.106000  20.225000 53.815000  20.295000 ;
      RECT 19.176000  20.155000 53.815000  20.225000 ;
      RECT 19.176000  20.155000 53.815000  20.225000 ;
      RECT 19.246000  20.085000 53.815000  20.155000 ;
      RECT 19.246000  20.085000 53.815000  20.155000 ;
      RECT 19.316000  20.015000 53.815000  20.085000 ;
      RECT 19.316000  20.015000 53.815000  20.085000 ;
      RECT 19.386000  19.945000 53.815000  20.015000 ;
      RECT 19.386000  19.945000 53.815000  20.015000 ;
      RECT 19.399000  19.932000 53.955000  21.835000 ;
      RECT 19.457000  19.874000 53.815000  19.945000 ;
      RECT 19.457000  19.874000 53.815000  19.945000 ;
      RECT 19.511000  19.820000 53.814000  19.875000 ;
      RECT 19.511000  19.820000 53.814000  19.875000 ;
      RECT 19.581000  19.750000 53.869000  19.820000 ;
      RECT 19.581000  19.750000 53.869000  19.820000 ;
      RECT 19.651000  19.680000 53.939000  19.750000 ;
      RECT 19.651000  19.680000 53.939000  19.750000 ;
      RECT 19.721000  19.610000 54.009000  19.680000 ;
      RECT 19.721000  19.610000 54.009000  19.680000 ;
      RECT 19.791000  19.540000 54.079000  19.610000 ;
      RECT 19.791000  19.540000 54.079000  19.610000 ;
      RECT 19.861000  19.470000 54.149000  19.540000 ;
      RECT 19.861000  19.470000 54.149000  19.540000 ;
      RECT 19.931000  19.400000 54.219000  19.470000 ;
      RECT 19.931000  19.400000 54.219000  19.470000 ;
      RECT 20.001000  19.330000 54.289000  19.400000 ;
      RECT 20.001000  19.330000 54.289000  19.400000 ;
      RECT 20.071000  19.260000 54.359000  19.330000 ;
      RECT 20.071000  19.260000 54.359000  19.330000 ;
      RECT 20.141000  19.190000 54.429000  19.260000 ;
      RECT 20.141000  19.190000 54.429000  19.260000 ;
      RECT 20.211000  19.120000 54.499000  19.190000 ;
      RECT 20.211000  19.120000 54.499000  19.190000 ;
      RECT 20.281000  19.050000 54.569000  19.120000 ;
      RECT 20.281000  19.050000 54.569000  19.120000 ;
      RECT 20.351000  18.980000 54.639000  19.050000 ;
      RECT 20.351000  18.980000 54.639000  19.050000 ;
      RECT 20.421000  18.910000 54.709000  18.980000 ;
      RECT 20.421000  18.910000 54.709000  18.980000 ;
      RECT 20.491000  18.840000 54.779000  18.910000 ;
      RECT 20.491000  18.840000 54.779000  18.910000 ;
      RECT 20.561000  18.770000 54.849000  18.840000 ;
      RECT 20.561000  18.770000 54.849000  18.840000 ;
      RECT 20.631000  18.700000 54.919000  18.770000 ;
      RECT 20.631000  18.700000 54.919000  18.770000 ;
      RECT 20.701000  18.630000 54.989000  18.700000 ;
      RECT 20.701000  18.630000 54.989000  18.700000 ;
      RECT 20.771000  18.560000 55.059000  18.630000 ;
      RECT 20.771000  18.560000 55.059000  18.630000 ;
      RECT 20.775000   0.000000 20.785000   1.601000 ;
      RECT 20.775000   1.601000 20.785000   1.762000 ;
      RECT 20.841000  18.490000 55.129000  18.560000 ;
      RECT 20.841000  18.490000 55.129000  18.560000 ;
      RECT 20.911000  18.420000 55.199000  18.490000 ;
      RECT 20.911000  18.420000 55.199000  18.490000 ;
      RECT 20.981000  18.350000 55.269000  18.420000 ;
      RECT 20.981000  18.350000 55.269000  18.420000 ;
      RECT 21.051000  18.280000 55.339000  18.350000 ;
      RECT 21.051000  18.280000 55.339000  18.350000 ;
      RECT 21.121000  18.210000 55.409000  18.280000 ;
      RECT 21.121000  18.210000 55.409000  18.280000 ;
      RECT 21.191000  18.140000 55.479000  18.210000 ;
      RECT 21.191000  18.140000 55.479000  18.210000 ;
      RECT 21.261000  18.070000 55.549000  18.140000 ;
      RECT 21.261000  18.070000 55.549000  18.140000 ;
      RECT 21.331000  18.000000 55.619000  18.070000 ;
      RECT 21.331000  18.000000 55.619000  18.070000 ;
      RECT 21.401000  17.930000 55.689000  18.000000 ;
      RECT 21.401000  17.930000 55.689000  18.000000 ;
      RECT 21.471000  17.860000 55.759000  17.930000 ;
      RECT 21.471000  17.860000 55.759000  17.930000 ;
      RECT 21.541000  17.790000 55.829000  17.860000 ;
      RECT 21.541000  17.790000 55.829000  17.860000 ;
      RECT 21.554000  17.777000 53.955000  19.932000 ;
      RECT 21.612000  17.719000 55.899000  17.790000 ;
      RECT 21.612000  17.719000 55.899000  17.790000 ;
      RECT 21.621000  17.710000 55.970000  17.720000 ;
      RECT 21.621000  17.710000 55.970000  17.720000 ;
      RECT 21.691000  17.640000 55.970000  17.710000 ;
      RECT 21.691000  17.640000 55.970000  17.710000 ;
      RECT 21.761000  17.570000 55.970000  17.640000 ;
      RECT 21.761000  17.570000 55.970000  17.640000 ;
      RECT 21.831000  17.500000 55.970000  17.570000 ;
      RECT 21.831000  17.500000 55.970000  17.570000 ;
      RECT 21.901000  17.430000 55.970000  17.500000 ;
      RECT 21.901000  17.430000 55.970000  17.500000 ;
      RECT 21.971000  17.360000 55.970000  17.430000 ;
      RECT 21.971000  17.360000 55.970000  17.430000 ;
      RECT 21.971000  17.360000 56.110000  17.777000 ;
      RECT 53.675000   0.000000 53.955000   7.873000 ;
      RECT 53.675000   7.873000 55.762000   9.680000 ;
      RECT 53.815000   8.000000 53.884000   8.070000 ;
      RECT 53.815000   8.070000 53.954000   8.140000 ;
      RECT 53.815000   8.140000 54.024000   8.210000 ;
      RECT 53.815000   8.210000 54.094000   8.280000 ;
      RECT 53.815000   8.280000 54.164000   8.350000 ;
      RECT 53.815000   8.350000 54.234000   8.420000 ;
      RECT 53.815000   8.420000 54.304000   8.490000 ;
      RECT 53.815000   8.490000 54.374000   8.560000 ;
      RECT 53.815000   8.560000 54.444000   8.630000 ;
      RECT 53.815000   8.630000 54.514000   8.700000 ;
      RECT 53.815000   8.700000 54.584000   8.770000 ;
      RECT 53.815000   8.770000 54.654000   8.840000 ;
      RECT 53.815000   8.840000 54.724000   8.910000 ;
      RECT 53.815000   8.910000 54.794000   8.980000 ;
      RECT 53.815000   8.980000 54.864000   9.050000 ;
      RECT 53.815000   9.050000 54.934000   9.120000 ;
      RECT 53.815000   9.120000 55.004000   9.190000 ;
      RECT 53.815000   9.190000 55.074000   9.260000 ;
      RECT 53.815000   9.260000 55.144000   9.330000 ;
      RECT 53.815000   9.330000 55.214000   9.400000 ;
      RECT 53.815000   9.400000 55.284000   9.470000 ;
      RECT 53.815000   9.470000 55.354000   9.540000 ;
      RECT 53.815000   9.540000 55.424000   9.610000 ;
      RECT 53.815000   9.610000 55.494000   9.680000 ;
      RECT 53.815000   9.680000 55.564000   9.750000 ;
      RECT 53.815000   9.750000 55.634000   9.800000 ;
      RECT 55.875000   9.800000 56.110000  10.028000 ;
      RECT 55.875000  10.028000 56.110000  17.360000 ;
      RECT 68.150000  74.488000 75.000000  98.700000 ;
      RECT 68.150000 130.845000 75.000000 133.770000 ;
      RECT 68.150000 140.850000 75.000000 143.770000 ;
      RECT 68.150000 150.850000 75.000000 153.770000 ;
      RECT 68.150000 160.850000 75.000000 163.770000 ;
      RECT 68.150000 170.850000 75.000000 173.770000 ;
      RECT 68.150000 180.850000 75.000000 183.770000 ;
      RECT 68.150000 190.850000 75.000000 193.770000 ;
      RECT 68.290000  74.546000 75.000000  98.840000 ;
      RECT 68.290000 130.705000 75.000000 133.910000 ;
      RECT 68.290000 140.710000 75.000000 143.910000 ;
      RECT 68.290000 150.710000 75.000000 153.910000 ;
      RECT 68.290000 160.710000 75.000000 163.910000 ;
      RECT 68.290000 170.710000 75.000000 173.910000 ;
      RECT 68.290000 180.710000 75.000000 183.910000 ;
      RECT 68.290000 190.710000 75.000000 193.910000 ;
      RECT 68.296000  74.540000 75.000000  74.545000 ;
      RECT 68.296000  74.540000 75.000000  74.545000 ;
      RECT 68.366000  74.470000 75.000000  74.540000 ;
      RECT 68.366000  74.470000 75.000000  74.540000 ;
      RECT 68.436000  74.400000 75.000000  74.470000 ;
      RECT 68.436000  74.400000 75.000000  74.470000 ;
      RECT 68.506000  74.330000 75.000000  74.400000 ;
      RECT 68.506000  74.330000 75.000000  74.400000 ;
      RECT 68.576000  74.260000 75.000000  74.330000 ;
      RECT 68.576000  74.260000 75.000000  74.330000 ;
      RECT 68.646000  74.190000 75.000000  74.260000 ;
      RECT 68.646000  74.190000 75.000000  74.260000 ;
      RECT 68.716000  74.120000 75.000000  74.190000 ;
      RECT 68.716000  74.120000 75.000000  74.190000 ;
      RECT 68.786000  74.050000 75.000000  74.120000 ;
      RECT 68.786000  74.050000 75.000000  74.120000 ;
      RECT 68.856000  73.980000 75.000000  74.050000 ;
      RECT 68.856000  73.980000 75.000000  74.050000 ;
      RECT 68.868000  73.770000 75.000000  74.488000 ;
      RECT 68.926000  73.910000 75.000000  73.980000 ;
      RECT 68.926000  73.910000 75.000000  73.980000 ;
      RECT 74.840000   0.000000 75.000000  73.770000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000  0.200000 171.495000 ;
      RECT  0.000000 171.495000 15.205000 189.915000 ;
      RECT  0.000000 171.595000 15.205000 189.915000 ;
      RECT  0.000000 171.595000 15.205000 198.000000 ;
      RECT  0.000000 189.915000 75.000000 198.000000 ;
      RECT  0.000000 189.915000 75.000000 198.000000 ;
      RECT 13.200000  94.384000 15.205000 171.495000 ;
      RECT 13.300000  94.426000 15.205000 171.595000 ;
      RECT 13.440000  94.144000 15.205000  94.384000 ;
      RECT 13.441000  94.285000 15.205000  94.425000 ;
      RECT 13.582000  94.144000 15.205000  94.285000 ;
      RECT 13.726000  94.000000 15.204000  94.145000 ;
      RECT 13.876000  93.850000 15.349000  94.000000 ;
      RECT 14.026000  93.700000 15.499000  93.850000 ;
      RECT 14.176000  93.550000 15.649000  93.700000 ;
      RECT 14.326000  93.400000 15.799000  93.550000 ;
      RECT 14.476000  93.250000 15.949000  93.400000 ;
      RECT 14.626000  93.100000 16.099000  93.250000 ;
      RECT 14.776000  92.950000 16.249000  93.100000 ;
      RECT 14.926000  92.800000 16.399000  92.950000 ;
      RECT 15.076000  92.650000 16.549000  92.800000 ;
      RECT 15.226000  92.500000 16.699000  92.650000 ;
      RECT 15.376000  92.350000 16.849000  92.500000 ;
      RECT 15.526000  92.200000 16.999000  92.350000 ;
      RECT 15.676000  92.050000 17.149000  92.200000 ;
      RECT 15.826000  91.900000 17.299000  92.050000 ;
      RECT 15.976000  91.750000 17.449000  91.900000 ;
      RECT 16.126000  91.600000 17.599000  91.750000 ;
      RECT 16.276000  91.450000 17.749000  91.600000 ;
      RECT 16.426000  91.300000 17.899000  91.450000 ;
      RECT 16.576000  91.150000 18.049000  91.300000 ;
      RECT 16.726000  91.000000 18.199000  91.150000 ;
      RECT 16.876000  90.850000 18.349000  91.000000 ;
      RECT 17.026000  90.700000 18.499000  90.850000 ;
      RECT 17.176000  90.550000 18.649000  90.700000 ;
      RECT 17.326000  90.400000 18.799000  90.550000 ;
      RECT 17.476000  90.250000 18.949000  90.400000 ;
      RECT 17.626000  90.100000 19.099000  90.250000 ;
      RECT 17.776000  89.950000 19.249000  90.100000 ;
      RECT 17.926000  89.800000 19.399000  89.950000 ;
      RECT 18.076000  89.650000 19.549000  89.800000 ;
      RECT 18.226000  89.500000 19.699000  89.650000 ;
      RECT 18.376000  89.350000 19.849000  89.500000 ;
      RECT 18.526000  89.200000 19.999000  89.350000 ;
      RECT 18.676000  89.050000 20.149000  89.200000 ;
      RECT 18.826000  88.900000 20.299000  89.050000 ;
      RECT 18.976000  88.750000 20.449000  88.900000 ;
      RECT 19.126000  88.600000 20.599000  88.750000 ;
      RECT 19.276000  88.450000 20.749000  88.600000 ;
      RECT 19.426000  88.300000 20.899000  88.450000 ;
      RECT 19.576000  88.150000 21.049000  88.300000 ;
      RECT 19.726000  88.000000 21.199000  88.150000 ;
      RECT 19.876000  87.850000 21.349000  88.000000 ;
      RECT 20.026000  87.700000 21.499000  87.850000 ;
      RECT 20.176000  87.550000 21.649000  87.700000 ;
      RECT 20.326000  87.400000 21.799000  87.550000 ;
      RECT 20.476000  87.250000 21.949000  87.400000 ;
      RECT 20.626000  87.100000 22.099000  87.250000 ;
      RECT 20.776000  86.950000 22.249000  87.100000 ;
      RECT 20.926000  86.800000 22.399000  86.950000 ;
      RECT 21.076000  86.650000 22.549000  86.800000 ;
      RECT 21.226000  86.500000 22.699000  86.650000 ;
      RECT 21.376000  86.350000 22.849000  86.500000 ;
      RECT 21.526000  86.200000 22.999000  86.350000 ;
      RECT 21.676000  86.050000 23.149000  86.200000 ;
      RECT 21.827000  85.899000 23.299000  86.050000 ;
      RECT 21.951000  85.775000 23.450000  85.900000 ;
      RECT 22.005000  96.956000 25.635000 166.934000 ;
      RECT 22.005000  96.956000 25.635000 166.934000 ;
      RECT 22.005000 166.934000 25.635000 170.444000 ;
      RECT 22.076000  96.885000 25.635000  96.955000 ;
      RECT 22.101000  85.625000 23.450000  85.775000 ;
      RECT 22.156000 166.934000 25.635000 167.085000 ;
      RECT 22.226000  96.735000 25.635000  96.885000 ;
      RECT 22.251000  85.475000 23.450000  85.625000 ;
      RECT 22.306000 167.085000 25.635000 167.235000 ;
      RECT 22.376000  96.585000 25.635000  96.735000 ;
      RECT 22.401000  85.325000 23.450000  85.475000 ;
      RECT 22.456000 167.235000 25.635000 167.385000 ;
      RECT 22.526000  96.435000 25.635000  96.585000 ;
      RECT 22.551000  85.175000 23.450000  85.325000 ;
      RECT 22.606000 167.385000 25.635000 167.535000 ;
      RECT 22.676000  96.285000 25.635000  96.435000 ;
      RECT 22.701000  85.025000 23.450000  85.175000 ;
      RECT 22.756000 167.535000 25.635000 167.685000 ;
      RECT 22.826000  96.135000 25.635000  96.285000 ;
      RECT 22.851000  84.875000 23.450000  85.025000 ;
      RECT 22.906000 167.685000 25.635000 167.835000 ;
      RECT 22.976000  95.985000 25.635000  96.135000 ;
      RECT 23.001000  84.725000 23.450000  84.875000 ;
      RECT 23.056000 167.835000 25.635000 167.985000 ;
      RECT 23.100000  84.484000 23.450000  85.899000 ;
      RECT 23.126000  95.835000 25.635000  95.985000 ;
      RECT 23.151000  84.575000 23.450000  84.725000 ;
      RECT 23.206000 167.985000 25.635000 168.135000 ;
      RECT 23.276000  95.685000 25.635000  95.835000 ;
      RECT 23.301000  84.425000 23.450000  84.575000 ;
      RECT 23.356000 168.135000 25.635000 168.285000 ;
      RECT 23.426000  95.535000 25.635000  95.685000 ;
      RECT 23.506000 168.285000 25.635000 168.435000 ;
      RECT 23.576000  95.385000 25.635000  95.535000 ;
      RECT 23.656000 168.435000 25.635000 168.585000 ;
      RECT 23.726000  95.235000 25.635000  95.385000 ;
      RECT 23.806000 168.585000 25.635000 168.735000 ;
      RECT 23.876000  95.085000 25.635000  95.235000 ;
      RECT 23.956000 168.735000 25.635000 168.885000 ;
      RECT 24.026000  94.935000 25.635000  95.085000 ;
      RECT 24.106000 168.885000 25.635000 169.035000 ;
      RECT 24.176000  94.785000 25.635000  94.935000 ;
      RECT 24.256000 169.035000 25.635000 169.185000 ;
      RECT 24.326000  94.635000 25.635000  94.785000 ;
      RECT 24.406000 169.185000 25.635000 169.335000 ;
      RECT 24.476000  94.485000 25.635000  94.635000 ;
      RECT 24.556000 169.335000 25.635000 169.485000 ;
      RECT 24.627000  94.334000 25.635000  94.485000 ;
      RECT 24.627000  94.334000 25.635000  96.956000 ;
      RECT 24.706000 169.485000 25.635000 169.635000 ;
      RECT 24.746000  94.215000 25.634000  94.335000 ;
      RECT 24.800000   0.000000 25.600000  82.334000 ;
      RECT 24.800000  82.334000 25.150000  82.784000 ;
      RECT 24.856000 169.635000 25.635000 169.785000 ;
      RECT 24.896000  94.065000 25.754000  94.215000 ;
      RECT 24.900000   0.000000 25.600000  82.334000 ;
      RECT 24.900000  82.334000 25.449000  82.485000 ;
      RECT 24.900000  82.485000 25.299000  82.635000 ;
      RECT 24.900000  82.635000 25.149000  82.785000 ;
      RECT 24.900000  82.785000 24.999000  82.935000 ;
      RECT 25.006000 169.785000 25.635000 169.935000 ;
      RECT 25.046000  93.915000 25.904000  94.065000 ;
      RECT 25.156000 169.935000 25.635000 170.085000 ;
      RECT 25.196000  93.765000 26.054000  93.915000 ;
      RECT 25.306000 170.085000 25.635000 170.235000 ;
      RECT 25.346000  93.615000 26.204000  93.765000 ;
      RECT 25.456000 170.235000 25.635000 170.385000 ;
      RECT 25.496000  93.465000 26.354000  93.615000 ;
      RECT 25.515000 170.444000 25.635000 189.915000 ;
      RECT 25.606000 170.385000 25.635000 170.535000 ;
      RECT 25.646000  93.315000 26.504000  93.465000 ;
      RECT 25.796000  93.165000 26.654000  93.315000 ;
      RECT 25.946000  93.015000 26.804000  93.165000 ;
      RECT 26.096000  92.865000 26.954000  93.015000 ;
      RECT 26.246000  92.715000 27.104000  92.865000 ;
      RECT 26.396000  92.565000 27.254000  92.715000 ;
      RECT 26.546000  92.415000 27.404000  92.565000 ;
      RECT 26.696000  92.265000 27.554000  92.415000 ;
      RECT 26.846000  92.115000 27.704000  92.265000 ;
      RECT 26.996000  91.965000 27.854000  92.115000 ;
      RECT 27.146000  91.815000 28.004000  91.965000 ;
      RECT 27.296000  91.665000 28.154000  91.815000 ;
      RECT 27.446000  91.515000 28.304000  91.665000 ;
      RECT 27.596000  91.365000 28.454000  91.515000 ;
      RECT 27.746000  91.215000 28.604000  91.365000 ;
      RECT 27.896000  91.065000 28.754000  91.215000 ;
      RECT 28.046000  90.915000 28.904000  91.065000 ;
      RECT 28.196000  90.765000 29.054000  90.915000 ;
      RECT 28.346000  90.615000 29.204000  90.765000 ;
      RECT 28.496000  90.465000 29.354000  90.615000 ;
      RECT 28.646000  90.315000 29.504000  90.465000 ;
      RECT 28.796000  90.165000 29.654000  90.315000 ;
      RECT 28.946000  90.015000 29.804000  90.165000 ;
      RECT 29.096000  89.865000 29.954000  90.015000 ;
      RECT 29.246000  89.715000 30.104000  89.865000 ;
      RECT 29.396000  89.565000 30.254000  89.715000 ;
      RECT 29.546000  89.415000 30.404000  89.565000 ;
      RECT 29.696000  89.265000 30.554000  89.415000 ;
      RECT 29.846000  89.115000 30.704000  89.265000 ;
      RECT 29.996000  88.965000 30.854000  89.115000 ;
      RECT 30.146000  88.815000 31.004000  88.965000 ;
      RECT 30.296000  88.665000 31.154000  88.815000 ;
      RECT 30.446000  88.515000 31.304000  88.665000 ;
      RECT 30.596000  88.365000 31.454000  88.515000 ;
      RECT 30.746000  88.215000 31.604000  88.365000 ;
      RECT 30.896000  88.065000 31.754000  88.215000 ;
      RECT 31.046000  87.915000 31.904000  88.065000 ;
      RECT 31.196000  87.765000 32.054000  87.915000 ;
      RECT 31.346000  87.615000 32.204000  87.765000 ;
      RECT 31.496000  87.465000 32.354000  87.615000 ;
      RECT 31.646000  87.315000 32.504000  87.465000 ;
      RECT 31.796000  87.165000 32.654000  87.315000 ;
      RECT 31.946000  87.015000 32.804000  87.165000 ;
      RECT 32.096000  86.865000 32.954000  87.015000 ;
      RECT 32.246000  86.715000 33.104000  86.865000 ;
      RECT 32.396000  86.565000 33.254000  86.715000 ;
      RECT 32.435000  93.556000 40.410000  93.705000 ;
      RECT 32.435000  93.556000 42.435000  95.581000 ;
      RECT 32.435000  93.705000 40.559000  93.855000 ;
      RECT 32.435000  93.855000 40.709000  94.005000 ;
      RECT 32.435000  94.005000 40.859000  94.155000 ;
      RECT 32.435000  94.155000 41.009000  94.305000 ;
      RECT 32.435000  94.305000 41.159000  94.455000 ;
      RECT 32.435000  94.455000 41.309000  94.605000 ;
      RECT 32.435000  94.605000 41.459000  94.755000 ;
      RECT 32.435000  94.755000 41.609000  94.905000 ;
      RECT 32.435000  94.905000 41.759000  95.055000 ;
      RECT 32.435000  95.055000 41.909000  95.205000 ;
      RECT 32.435000  95.205000 42.059000  95.355000 ;
      RECT 32.435000  95.355000 42.209000  95.505000 ;
      RECT 32.435000  95.505000 42.359000  95.580000 ;
      RECT 32.435000  95.581000 35.440000 159.399000 ;
      RECT 32.435000  95.581000 42.435000 162.404000 ;
      RECT 32.435000 159.399000 36.681000 162.404000 ;
      RECT 32.435000 162.404000 42.435000 163.969000 ;
      RECT 32.516000  93.475000 40.329000  93.555000 ;
      RECT 32.545000  84.856000 34.105000  85.864000 ;
      RECT 32.545000  84.856000 34.105000  85.864000 ;
      RECT 32.545000  85.864000 33.553000  86.416000 ;
      RECT 32.545000  85.864000 33.954000  86.015000 ;
      RECT 32.545000  86.015000 33.804000  86.165000 ;
      RECT 32.545000  86.165000 33.654000  86.315000 ;
      RECT 32.545000  86.315000 33.554000  86.415000 ;
      RECT 32.545000  86.416000 33.404000  86.565000 ;
      RECT 32.571000  84.830000 34.079000  84.855000 ;
      RECT 32.586000 162.404000 42.435000 162.555000 ;
      RECT 32.666000  93.325000 40.179000  93.475000 ;
      RECT 32.721000  84.680000 33.929000  84.830000 ;
      RECT 32.736000 162.555000 42.435000 162.705000 ;
      RECT 32.816000  93.175000 40.029000  93.325000 ;
      RECT 32.871000  84.530000 33.779000  84.680000 ;
      RECT 32.886000 162.705000 42.435000 162.855000 ;
      RECT 32.966000  93.025000 39.879000  93.175000 ;
      RECT 33.021000  84.380000 33.629000  84.530000 ;
      RECT 33.021000  84.380000 34.105000  84.856000 ;
      RECT 33.036000 162.855000 42.435000 163.005000 ;
      RECT 33.116000  92.875000 39.729000  93.025000 ;
      RECT 33.186000 163.005000 42.435000 163.155000 ;
      RECT 33.266000  92.725000 39.579000  92.875000 ;
      RECT 33.336000 163.155000 42.435000 163.305000 ;
      RECT 33.416000  92.575000 39.429000  92.725000 ;
      RECT 33.486000 163.305000 42.435000 163.455000 ;
      RECT 33.566000  92.425000 39.279000  92.575000 ;
      RECT 33.636000 163.455000 42.435000 163.605000 ;
      RECT 33.716000  92.275000 39.129000  92.425000 ;
      RECT 33.786000 163.605000 42.435000 163.755000 ;
      RECT 33.866000  92.125000 38.979000  92.275000 ;
      RECT 33.936000 163.755000 42.435000 163.905000 ;
      RECT 34.000000 163.969000 39.110000 167.294000 ;
      RECT 34.001000 163.905000 42.435000 163.970000 ;
      RECT 34.016000  91.975000 38.829000  92.125000 ;
      RECT 34.151000 163.969000 42.284000 164.120000 ;
      RECT 34.166000  91.825000 38.679000  91.975000 ;
      RECT 34.301000 164.120000 42.134000 164.270000 ;
      RECT 34.316000  91.675000 38.529000  91.825000 ;
      RECT 34.451000 164.270000 41.984000 164.420000 ;
      RECT 34.466000  91.525000 38.379000  91.675000 ;
      RECT 34.601000 164.420000 41.834000 164.570000 ;
      RECT 34.616000  91.375000 38.229000  91.525000 ;
      RECT 34.751000 164.570000 41.684000 164.720000 ;
      RECT 34.766000  91.225000 38.079000  91.375000 ;
      RECT 34.901000 164.720000 41.534000 164.870000 ;
      RECT 34.916000  91.075000 37.929000  91.225000 ;
      RECT 35.051000 164.870000 41.384000 165.020000 ;
      RECT 35.066000  90.925000 37.779000  91.075000 ;
      RECT 35.201000 165.020000 41.234000 165.170000 ;
      RECT 35.216000  90.775000 37.629000  90.925000 ;
      RECT 35.216000  90.775000 40.410000  93.556000 ;
      RECT 35.351000 165.170000 41.084000 165.320000 ;
      RECT 35.437000  94.800000 37.408000  94.950000 ;
      RECT 35.437000  94.800000 37.408000  94.950000 ;
      RECT 35.437000  94.950000 37.558000  95.100000 ;
      RECT 35.437000  94.950000 37.558000  95.100000 ;
      RECT 35.437000  95.100000 37.708000  95.250000 ;
      RECT 35.437000  95.100000 37.708000  95.250000 ;
      RECT 35.437000  95.250000 37.858000  95.400000 ;
      RECT 35.437000  95.250000 37.858000  95.400000 ;
      RECT 35.437000  95.400000 38.008000  95.550000 ;
      RECT 35.437000  95.400000 38.008000  95.550000 ;
      RECT 35.437000  95.550000 38.158000  95.700000 ;
      RECT 35.437000  95.550000 38.158000  95.700000 ;
      RECT 35.437000  95.700000 38.308000  95.850000 ;
      RECT 35.437000  95.700000 38.308000  95.850000 ;
      RECT 35.437000  95.850000 38.458000  96.000000 ;
      RECT 35.437000  95.850000 38.458000  96.000000 ;
      RECT 35.437000  96.000000 38.608000  96.150000 ;
      RECT 35.437000  96.000000 38.608000  96.150000 ;
      RECT 35.437000  96.150000 38.758000  96.300000 ;
      RECT 35.437000  96.150000 38.758000  96.300000 ;
      RECT 35.437000  96.300000 38.908000  96.450000 ;
      RECT 35.437000  96.300000 38.908000  96.450000 ;
      RECT 35.437000  96.450000 39.058000  96.600000 ;
      RECT 35.437000  96.450000 39.058000  96.600000 ;
      RECT 35.437000  96.600000 39.208000  96.750000 ;
      RECT 35.437000  96.600000 39.208000  96.750000 ;
      RECT 35.437000  96.750000 39.358000  96.825000 ;
      RECT 35.437000  96.750000 39.358000  96.825000 ;
      RECT 35.437000  96.825000 39.433000 161.160000 ;
      RECT 35.501000 165.320000 40.934000 165.470000 ;
      RECT 35.522000  94.715000 37.323000  94.800000 ;
      RECT 35.522000  94.715000 37.323000  94.800000 ;
      RECT 35.587000 161.160000 39.433000 161.310000 ;
      RECT 35.587000 161.160000 39.433000 161.310000 ;
      RECT 35.651000 165.470000 40.784000 165.620000 ;
      RECT 35.672000  94.565000 37.173000  94.715000 ;
      RECT 35.672000  94.565000 37.173000  94.715000 ;
      RECT 35.737000 161.310000 39.433000 161.460000 ;
      RECT 35.737000 161.310000 39.433000 161.460000 ;
      RECT 35.801000 165.620000 40.634000 165.770000 ;
      RECT 35.822000  94.415000 37.023000  94.565000 ;
      RECT 35.822000  94.415000 37.023000  94.565000 ;
      RECT 35.887000 161.460000 39.433000 161.610000 ;
      RECT 35.887000 161.460000 39.433000 161.610000 ;
      RECT 35.951000 165.770000 40.484000 165.920000 ;
      RECT 35.973000  94.265000 36.873000  94.415000 ;
      RECT 35.973000  94.265000 36.873000  94.415000 ;
      RECT 36.037000 161.610000 39.433000 161.760000 ;
      RECT 36.037000 161.610000 39.433000 161.760000 ;
      RECT 36.101000 165.920000 40.334000 166.070000 ;
      RECT 36.123000  94.115000 36.723000  94.265000 ;
      RECT 36.123000  94.115000 36.723000  94.265000 ;
      RECT 36.187000 161.760000 39.433000 161.910000 ;
      RECT 36.187000 161.760000 39.433000 161.910000 ;
      RECT 36.251000 166.070000 40.184000 166.220000 ;
      RECT 36.273000  93.965000 36.573000  94.115000 ;
      RECT 36.273000  93.965000 36.573000  94.115000 ;
      RECT 36.337000 161.910000 39.433000 162.060000 ;
      RECT 36.337000 161.910000 39.433000 162.060000 ;
      RECT 36.401000 166.220000 40.034000 166.370000 ;
      RECT 36.487000 162.060000 39.433000 162.210000 ;
      RECT 36.487000 162.060000 39.433000 162.210000 ;
      RECT 36.551000 166.370000 39.884000 166.520000 ;
      RECT 36.637000 162.210000 39.433000 162.360000 ;
      RECT 36.637000 162.210000 39.433000 162.360000 ;
      RECT 36.701000 166.520000 39.734000 166.670000 ;
      RECT 36.787000 162.360000 39.433000 162.510000 ;
      RECT 36.787000 162.360000 39.433000 162.510000 ;
      RECT 36.851000 166.670000 39.584000 166.820000 ;
      RECT 36.937000 162.510000 39.433000 162.660000 ;
      RECT 36.937000 162.510000 39.433000 162.660000 ;
      RECT 37.001000 166.820000 39.434000 166.970000 ;
      RECT 37.002000 162.660000 39.433000 162.725000 ;
      RECT 37.002000 162.660000 39.433000 162.725000 ;
      RECT 37.151000 166.970000 39.284000 167.120000 ;
      RECT 37.152000 162.725000 39.283000 162.875000 ;
      RECT 37.152000 162.725000 39.283000 162.875000 ;
      RECT 37.280000   0.000000 37.980000  69.890000 ;
      RECT 37.280000   0.000000 37.980000  69.890000 ;
      RECT 37.280000  69.890000 50.355000  70.939000 ;
      RECT 37.280000  69.890000 50.355000  74.340000 ;
      RECT 37.280000  69.890000 50.455000  70.939000 ;
      RECT 37.280000  70.939000 50.455000  74.340000 ;
      RECT 37.301000 167.120000 39.134000 167.270000 ;
      RECT 37.302000 162.875000 39.133000 163.025000 ;
      RECT 37.302000 162.875000 39.133000 163.025000 ;
      RECT 37.325000 167.294000 37.545000 168.859000 ;
      RECT 37.325000 167.294000 38.959000 167.445000 ;
      RECT 37.325000 167.445000 38.809000 167.595000 ;
      RECT 37.325000 167.595000 38.659000 167.745000 ;
      RECT 37.325000 167.745000 38.509000 167.895000 ;
      RECT 37.325000 167.895000 38.359000 168.045000 ;
      RECT 37.325000 168.045000 38.209000 168.195000 ;
      RECT 37.325000 168.195000 38.059000 168.345000 ;
      RECT 37.325000 168.345000 37.909000 168.495000 ;
      RECT 37.325000 168.495000 37.759000 168.645000 ;
      RECT 37.325000 168.645000 37.609000 168.795000 ;
      RECT 37.325000 168.795000 37.459000 168.945000 ;
      RECT 37.325000 168.859000 37.545000 189.915000 ;
      RECT 37.326000 167.270000 39.109000 167.295000 ;
      RECT 37.431000  70.939000 50.355000  71.090000 ;
      RECT 37.431000  70.939000 50.355000  71.090000 ;
      RECT 37.452000 163.025000 38.983000 163.175000 ;
      RECT 37.452000 163.025000 38.983000 163.175000 ;
      RECT 37.581000  71.090000 50.355000  71.240000 ;
      RECT 37.581000  71.090000 50.355000  71.240000 ;
      RECT 37.602000 163.175000 38.833000 163.325000 ;
      RECT 37.602000 163.175000 38.833000 163.325000 ;
      RECT 37.731000  71.240000 50.355000  71.390000 ;
      RECT 37.731000  71.240000 50.355000  71.390000 ;
      RECT 37.752000 163.325000 38.684000 163.475000 ;
      RECT 37.752000 163.325000 38.684000 163.475000 ;
      RECT 37.881000  71.390000 50.355000  71.540000 ;
      RECT 37.881000  71.390000 50.355000  71.540000 ;
      RECT 37.902000 163.475000 38.534000 163.625000 ;
      RECT 37.902000 163.475000 38.534000 163.625000 ;
      RECT 38.031000  71.540000 50.355000  71.690000 ;
      RECT 38.031000  71.540000 50.355000  71.690000 ;
      RECT 38.052000 163.625000 38.384000 163.775000 ;
      RECT 38.052000 163.625000 38.384000 163.775000 ;
      RECT 38.181000  71.690000 50.355000  71.840000 ;
      RECT 38.181000  71.690000 50.355000  71.840000 ;
      RECT 38.189000  95.581000 42.435000  98.586000 ;
      RECT 38.202000 163.775000 38.234000 163.925000 ;
      RECT 38.202000 163.775000 38.234000 163.925000 ;
      RECT 38.217000 163.925000 38.218000 163.940000 ;
      RECT 38.217000 163.925000 38.218000 163.940000 ;
      RECT 38.331000  71.840000 50.355000  71.990000 ;
      RECT 38.331000  71.840000 50.355000  71.990000 ;
      RECT 38.481000  71.990000 50.355000  72.140000 ;
      RECT 38.481000  71.990000 50.355000  72.140000 ;
      RECT 38.631000  72.140000 50.355000  72.290000 ;
      RECT 38.631000  72.140000 50.355000  72.290000 ;
      RECT 38.781000  72.290000 50.355000  72.440000 ;
      RECT 38.781000  72.290000 50.355000  72.440000 ;
      RECT 38.931000  72.440000 50.355000  72.590000 ;
      RECT 38.931000  72.440000 50.355000  72.590000 ;
      RECT 39.081000  72.590000 50.355000  72.740000 ;
      RECT 39.081000  72.590000 50.355000  72.740000 ;
      RECT 39.231000  72.740000 50.355000  72.890000 ;
      RECT 39.231000  72.740000 50.355000  72.890000 ;
      RECT 39.381000  72.890000 50.355000  73.040000 ;
      RECT 39.381000  72.890000 50.355000  73.040000 ;
      RECT 39.430000  98.586000 42.435000 162.404000 ;
      RECT 39.531000  73.040000 50.355000  73.190000 ;
      RECT 39.531000  73.040000 50.355000  73.190000 ;
      RECT 39.681000  73.190000 50.355000  73.340000 ;
      RECT 39.681000  73.190000 50.355000  73.340000 ;
      RECT 39.785000  84.856000 41.210000  87.194000 ;
      RECT 39.785000  84.856000 41.210000  87.194000 ;
      RECT 39.785000  87.194000 41.210000  87.611000 ;
      RECT 39.811000  84.830000 41.184000  84.855000 ;
      RECT 39.831000  73.340000 50.355000  73.490000 ;
      RECT 39.831000  73.340000 50.355000  73.490000 ;
      RECT 39.936000  87.194000 41.210000  87.345000 ;
      RECT 39.961000  84.680000 41.034000  84.830000 ;
      RECT 39.981000  73.490000 50.355000  73.640000 ;
      RECT 39.981000  73.490000 50.355000  73.640000 ;
      RECT 40.086000  87.345000 41.210000  87.495000 ;
      RECT 40.111000  84.530000 40.884000  84.680000 ;
      RECT 40.131000  73.640000 50.355000  73.790000 ;
      RECT 40.131000  73.640000 50.355000  73.790000 ;
      RECT 40.201000  87.495000 41.210000  87.610000 ;
      RECT 40.202000  87.611000 50.243000  96.644000 ;
      RECT 40.261000  84.380000 40.734000  84.530000 ;
      RECT 40.261000  84.380000 41.210000  84.856000 ;
      RECT 40.281000  73.790000 50.355000  73.940000 ;
      RECT 40.281000  73.790000 50.355000  73.940000 ;
      RECT 40.351000  87.611000 41.210000  87.760000 ;
      RECT 40.431000  73.940000 50.355000  74.090000 ;
      RECT 40.431000  73.940000 50.355000  74.090000 ;
      RECT 40.501000  87.760000 41.359000  87.910000 ;
      RECT 40.581000  74.090000 50.355000  74.240000 ;
      RECT 40.581000  74.090000 50.355000  74.240000 ;
      RECT 40.651000  87.910000 41.509000  88.060000 ;
      RECT 40.681000  74.240000 50.355000  74.340000 ;
      RECT 40.681000  74.240000 50.355000  74.340000 ;
      RECT 40.801000  88.060000 41.659000  88.210000 ;
      RECT 40.951000  88.210000 41.809000  88.360000 ;
      RECT 41.101000  88.360000 41.959000  88.510000 ;
      RECT 41.251000  88.510000 42.109000  88.660000 ;
      RECT 41.401000  88.660000 42.259000  88.810000 ;
      RECT 41.551000  88.810000 42.409000  88.960000 ;
      RECT 41.701000  88.960000 42.559000  89.110000 ;
      RECT 41.851000  89.110000 42.709000  89.260000 ;
      RECT 42.001000  89.260000 42.859000  89.410000 ;
      RECT 42.151000  89.410000 43.009000  89.560000 ;
      RECT 42.301000  89.560000 43.159000  89.710000 ;
      RECT 42.451000  89.710000 43.309000  89.860000 ;
      RECT 42.601000  89.860000 43.459000  90.010000 ;
      RECT 42.751000  90.010000 43.609000  90.160000 ;
      RECT 42.901000  90.160000 43.759000  90.310000 ;
      RECT 43.051000  90.310000 43.909000  90.460000 ;
      RECT 43.201000  90.460000 44.059000  90.610000 ;
      RECT 43.351000  90.610000 44.209000  90.760000 ;
      RECT 43.501000  90.760000 44.359000  90.910000 ;
      RECT 43.651000  90.910000 44.509000  91.060000 ;
      RECT 43.801000  91.060000 44.659000  91.210000 ;
      RECT 43.951000  91.210000 44.809000  91.360000 ;
      RECT 44.101000  91.360000 44.959000  91.510000 ;
      RECT 44.251000  91.510000 45.109000  91.660000 ;
      RECT 44.401000  91.660000 45.259000  91.810000 ;
      RECT 44.551000  91.810000 45.409000  91.960000 ;
      RECT 44.701000  91.960000 45.559000  92.110000 ;
      RECT 44.851000  92.110000 45.709000  92.260000 ;
      RECT 45.001000  92.260000 45.859000  92.410000 ;
      RECT 45.151000  92.410000 46.009000  92.560000 ;
      RECT 45.301000  92.560000 46.159000  92.710000 ;
      RECT 45.451000  92.710000 46.309000  92.860000 ;
      RECT 45.601000  92.860000 46.459000  93.010000 ;
      RECT 45.751000  93.010000 46.609000  93.160000 ;
      RECT 45.901000  93.160000 46.759000  93.310000 ;
      RECT 46.051000  93.310000 46.909000  93.460000 ;
      RECT 46.201000  93.460000 47.059000  93.610000 ;
      RECT 46.351000  93.610000 47.209000  93.760000 ;
      RECT 46.501000  93.760000 47.359000  93.910000 ;
      RECT 46.651000  93.910000 47.509000  94.060000 ;
      RECT 46.801000  94.060000 47.659000  94.210000 ;
      RECT 46.951000  94.210000 47.809000  94.360000 ;
      RECT 46.961000  74.340000 50.455000  76.649000 ;
      RECT 47.101000  94.360000 47.959000  94.510000 ;
      RECT 47.111000  74.340000 50.355000  74.490000 ;
      RECT 47.111000  74.340000 50.355000  74.490000 ;
      RECT 47.251000  94.510000 48.109000  94.660000 ;
      RECT 47.261000  74.490000 50.355000  74.640000 ;
      RECT 47.261000  74.490000 50.355000  74.640000 ;
      RECT 47.401000  94.660000 48.259000  94.810000 ;
      RECT 47.411000  74.640000 50.355000  74.790000 ;
      RECT 47.411000  74.640000 50.355000  74.790000 ;
      RECT 47.551000  94.810000 48.409000  94.960000 ;
      RECT 47.561000  74.790000 50.355000  74.940000 ;
      RECT 47.561000  74.790000 50.355000  74.940000 ;
      RECT 47.701000  94.960000 48.559000  95.110000 ;
      RECT 47.711000  74.940000 50.355000  75.090000 ;
      RECT 47.711000  74.940000 50.355000  75.090000 ;
      RECT 47.851000  95.110000 48.709000  95.260000 ;
      RECT 47.861000  75.090000 50.355000  75.240000 ;
      RECT 47.861000  75.090000 50.355000  75.240000 ;
      RECT 48.001000  95.260000 48.859000  95.410000 ;
      RECT 48.011000  75.240000 50.355000  75.390000 ;
      RECT 48.011000  75.240000 50.355000  75.390000 ;
      RECT 48.151000  95.410000 49.009000  95.560000 ;
      RECT 48.161000  75.390000 50.355000  75.540000 ;
      RECT 48.161000  75.390000 50.355000  75.540000 ;
      RECT 48.301000  95.560000 49.159000  95.710000 ;
      RECT 48.311000  75.540000 50.355000  75.690000 ;
      RECT 48.311000  75.540000 50.355000  75.690000 ;
      RECT 48.451000  95.710000 49.309000  95.860000 ;
      RECT 48.461000  75.690000 50.355000  75.840000 ;
      RECT 48.461000  75.690000 50.355000  75.840000 ;
      RECT 48.601000  95.860000 49.459000  96.010000 ;
      RECT 48.611000  75.840000 50.355000  75.990000 ;
      RECT 48.611000  75.840000 50.355000  75.990000 ;
      RECT 48.751000  96.010000 49.609000  96.160000 ;
      RECT 48.761000  75.990000 50.355000  76.140000 ;
      RECT 48.761000  75.990000 50.355000  76.140000 ;
      RECT 48.901000  96.160000 49.759000  96.310000 ;
      RECT 48.911000  76.140000 50.355000  76.290000 ;
      RECT 48.911000  76.140000 50.355000  76.290000 ;
      RECT 49.051000  96.310000 49.909000  96.460000 ;
      RECT 49.061000  76.290000 50.355000  76.440000 ;
      RECT 49.061000  76.290000 50.355000  76.440000 ;
      RECT 49.201000  96.460000 50.059000  96.610000 ;
      RECT 49.211000  76.440000 50.355000  76.590000 ;
      RECT 49.211000  76.440000 50.355000  76.590000 ;
      RECT 49.235000  96.644000 50.243000  96.795000 ;
      RECT 49.235000  96.644000 53.930000 100.331000 ;
      RECT 49.235000  96.795000 50.394000  96.945000 ;
      RECT 49.235000  96.945000 50.544000  97.095000 ;
      RECT 49.235000  97.095000 50.694000  97.245000 ;
      RECT 49.235000  97.245000 50.844000  97.395000 ;
      RECT 49.235000  97.395000 50.994000  97.545000 ;
      RECT 49.235000  97.545000 51.144000  97.695000 ;
      RECT 49.235000  97.695000 51.294000  97.845000 ;
      RECT 49.235000  97.845000 51.444000  97.995000 ;
      RECT 49.235000  97.995000 51.594000  98.145000 ;
      RECT 49.235000  98.145000 51.744000  98.295000 ;
      RECT 49.235000  98.295000 51.894000  98.445000 ;
      RECT 49.235000  98.445000 52.044000  98.595000 ;
      RECT 49.235000  98.595000 52.194000  98.745000 ;
      RECT 49.235000  98.745000 52.344000  98.895000 ;
      RECT 49.235000  98.895000 52.494000  99.045000 ;
      RECT 49.235000  99.045000 52.644000  99.195000 ;
      RECT 49.235000  99.195000 52.794000  99.345000 ;
      RECT 49.235000  99.345000 52.944000  99.495000 ;
      RECT 49.235000  99.495000 53.094000  99.645000 ;
      RECT 49.235000  99.645000 53.244000  99.795000 ;
      RECT 49.235000  99.795000 53.394000  99.945000 ;
      RECT 49.235000  99.945000 53.544000 100.095000 ;
      RECT 49.235000 100.095000 53.694000 100.245000 ;
      RECT 49.235000 100.245000 53.844000 100.330000 ;
      RECT 49.235000 100.331000 53.930000 164.294000 ;
      RECT 49.235000 100.331000 53.930000 164.294000 ;
      RECT 49.235000 164.294000 49.470000 168.754000 ;
      RECT 49.235000 164.294000 53.779000 164.445000 ;
      RECT 49.235000 164.445000 53.629000 164.595000 ;
      RECT 49.235000 164.595000 53.479000 164.745000 ;
      RECT 49.235000 164.745000 53.329000 164.895000 ;
      RECT 49.235000 164.895000 53.179000 165.045000 ;
      RECT 49.235000 165.045000 53.029000 165.195000 ;
      RECT 49.235000 165.195000 52.879000 165.345000 ;
      RECT 49.235000 165.345000 52.729000 165.495000 ;
      RECT 49.235000 165.495000 52.579000 165.645000 ;
      RECT 49.235000 165.645000 52.429000 165.795000 ;
      RECT 49.235000 165.795000 52.279000 165.945000 ;
      RECT 49.235000 165.945000 52.129000 166.095000 ;
      RECT 49.235000 166.095000 51.979000 166.245000 ;
      RECT 49.235000 166.245000 51.829000 166.395000 ;
      RECT 49.235000 166.395000 51.679000 166.545000 ;
      RECT 49.235000 166.545000 51.529000 166.695000 ;
      RECT 49.235000 166.695000 51.379000 166.845000 ;
      RECT 49.235000 166.845000 51.229000 166.995000 ;
      RECT 49.235000 166.995000 51.079000 167.145000 ;
      RECT 49.235000 167.145000 50.929000 167.295000 ;
      RECT 49.235000 167.295000 50.779000 167.445000 ;
      RECT 49.235000 167.445000 50.629000 167.595000 ;
      RECT 49.235000 167.595000 50.479000 167.745000 ;
      RECT 49.235000 167.745000 50.329000 167.895000 ;
      RECT 49.235000 167.895000 50.179000 168.045000 ;
      RECT 49.235000 168.045000 50.029000 168.195000 ;
      RECT 49.235000 168.195000 49.879000 168.345000 ;
      RECT 49.235000 168.345000 49.729000 168.495000 ;
      RECT 49.235000 168.495000 49.579000 168.645000 ;
      RECT 49.235000 168.645000 49.429000 168.795000 ;
      RECT 49.235000 168.754000 49.470000 189.915000 ;
      RECT 49.235000 168.795000 49.279000 168.945000 ;
      RECT 49.236000  96.610000 50.209000  96.645000 ;
      RECT 49.270000  76.649000 50.455000  84.589000 ;
      RECT 49.270000  77.734000 50.355000  84.631000 ;
      RECT 49.270000  84.589000 50.510000  84.644000 ;
      RECT 49.270000  84.631000 50.355000  84.635000 ;
      RECT 49.270000  84.635000 50.359000  84.640000 ;
      RECT 49.270000  84.640000 50.364000  84.645000 ;
      RECT 49.270000  84.644000 52.660000  86.794000 ;
      RECT 49.271000  76.590000 50.355000  76.650000 ;
      RECT 49.271000  76.590000 50.355000  76.650000 ;
      RECT 49.421000  76.649000 50.355000  76.800000 ;
      RECT 49.421000  76.649000 50.355000  76.800000 ;
      RECT 49.421000  84.644000 50.368000  84.795000 ;
      RECT 49.571000  76.800000 50.355000  76.950000 ;
      RECT 49.571000  76.800000 50.355000  76.950000 ;
      RECT 49.571000  84.795000 50.519000  84.945000 ;
      RECT 49.655000   0.000000 50.355000  69.890000 ;
      RECT 49.655000   0.000000 50.455000  69.890000 ;
      RECT 49.721000  76.950000 50.355000  77.100000 ;
      RECT 49.721000  76.950000 50.355000  77.100000 ;
      RECT 49.721000  84.945000 50.669000  85.095000 ;
      RECT 49.871000  77.100000 50.355000  77.250000 ;
      RECT 49.871000  77.100000 50.355000  77.250000 ;
      RECT 49.871000  85.095000 50.819000  85.245000 ;
      RECT 50.021000  77.250000 50.355000  77.400000 ;
      RECT 50.021000  77.250000 50.355000  77.400000 ;
      RECT 50.021000  85.245000 50.969000  85.395000 ;
      RECT 50.171000  77.400000 50.355000  77.550000 ;
      RECT 50.171000  77.400000 50.355000  77.550000 ;
      RECT 50.171000  85.395000 51.119000  85.545000 ;
      RECT 50.321000  77.550000 50.355000  77.700000 ;
      RECT 50.321000  77.550000 50.355000  77.700000 ;
      RECT 50.321000  85.545000 51.269000  85.695000 ;
      RECT 50.471000  85.695000 51.419000  85.845000 ;
      RECT 50.621000  85.845000 51.569000  85.995000 ;
      RECT 50.771000  85.995000 51.719000  86.145000 ;
      RECT 50.921000  86.145000 51.869000  86.295000 ;
      RECT 51.071000  86.295000 52.019000  86.445000 ;
      RECT 51.221000  86.445000 52.169000  86.595000 ;
      RECT 51.371000  86.595000 52.319000  86.745000 ;
      RECT 51.420000  86.794000 52.518000  86.945000 ;
      RECT 51.420000  86.794000 54.075000  88.209000 ;
      RECT 51.420000  86.945000 52.669000  87.095000 ;
      RECT 51.420000  87.095000 52.819000  87.245000 ;
      RECT 51.420000  87.245000 52.969000  87.395000 ;
      RECT 51.420000  87.395000 53.119000  87.545000 ;
      RECT 51.420000  87.545000 53.269000  87.695000 ;
      RECT 51.420000  87.695000 53.419000  87.845000 ;
      RECT 51.420000  87.845000 53.569000  87.995000 ;
      RECT 51.420000  87.995000 53.719000  88.145000 ;
      RECT 51.420000  88.145000 53.869000  88.210000 ;
      RECT 51.420000  88.209000 61.745000  95.879000 ;
      RECT 51.421000  86.745000 52.469000  86.795000 ;
      RECT 51.571000  88.209000 53.933000  88.360000 ;
      RECT 51.721000  88.360000 54.084000  88.510000 ;
      RECT 51.871000  88.510000 54.234000  88.660000 ;
      RECT 52.021000  88.660000 54.384000  88.810000 ;
      RECT 52.171000  88.810000 54.534000  88.960000 ;
      RECT 52.321000  88.960000 54.684000  89.110000 ;
      RECT 52.471000  89.110000 54.834000  89.260000 ;
      RECT 52.621000  89.260000 54.984000  89.410000 ;
      RECT 52.771000  89.410000 55.134000  89.560000 ;
      RECT 52.921000  89.560000 55.284000  89.710000 ;
      RECT 53.071000  89.710000 55.434000  89.860000 ;
      RECT 53.221000  89.860000 55.584000  90.010000 ;
      RECT 53.371000  90.010000 55.734000  90.160000 ;
      RECT 53.521000  90.160000 55.884000  90.310000 ;
      RECT 53.671000  90.310000 56.034000  90.460000 ;
      RECT 53.821000  90.460000 56.184000  90.610000 ;
      RECT 53.971000  90.610000 56.334000  90.760000 ;
      RECT 54.121000  90.760000 56.484000  90.910000 ;
      RECT 54.271000  90.910000 56.634000  91.060000 ;
      RECT 54.421000  91.060000 56.784000  91.210000 ;
      RECT 54.571000  91.210000 56.934000  91.360000 ;
      RECT 54.721000  91.360000 57.084000  91.510000 ;
      RECT 54.871000  91.510000 57.234000  91.660000 ;
      RECT 55.021000  91.660000 57.384000  91.810000 ;
      RECT 55.171000  91.810000 57.534000  91.960000 ;
      RECT 55.321000  91.960000 57.684000  92.110000 ;
      RECT 55.471000  92.110000 57.834000  92.260000 ;
      RECT 55.621000  92.260000 57.984000  92.410000 ;
      RECT 55.771000  92.410000 58.134000  92.560000 ;
      RECT 55.921000  92.560000 58.284000  92.710000 ;
      RECT 56.071000  92.710000 58.434000  92.860000 ;
      RECT 56.221000  92.860000 58.584000  93.010000 ;
      RECT 56.371000  93.010000 58.734000  93.160000 ;
      RECT 56.521000  93.160000 58.884000  93.310000 ;
      RECT 56.671000  93.310000 59.034000  93.460000 ;
      RECT 56.821000  93.460000 59.184000  93.610000 ;
      RECT 56.971000  93.610000 59.334000  93.760000 ;
      RECT 57.121000  93.760000 59.484000  93.910000 ;
      RECT 57.271000  93.910000 59.634000  94.060000 ;
      RECT 57.421000  94.060000 59.784000  94.210000 ;
      RECT 57.571000  94.210000 59.934000  94.360000 ;
      RECT 57.721000  94.360000 60.084000  94.510000 ;
      RECT 57.871000  94.510000 60.234000  94.660000 ;
      RECT 58.021000  94.660000 60.384000  94.810000 ;
      RECT 58.171000  94.810000 60.534000  94.960000 ;
      RECT 58.321000  94.960000 60.684000  95.110000 ;
      RECT 58.471000  95.110000 60.834000  95.260000 ;
      RECT 58.621000  95.260000 60.984000  95.410000 ;
      RECT 58.771000  95.410000 61.134000  95.560000 ;
      RECT 58.921000  95.560000 61.284000  95.710000 ;
      RECT 59.071000  95.710000 61.434000  95.860000 ;
      RECT 59.090000  95.879000 61.745000  97.519000 ;
      RECT 59.131000  95.860000 61.584000  95.920000 ;
      RECT 59.281000  95.921000 61.645000  96.070000 ;
      RECT 59.431000  96.070000 61.645000  96.220000 ;
      RECT 59.581000  96.220000 61.645000  96.370000 ;
      RECT 59.731000  96.370000 61.645000  96.520000 ;
      RECT 59.881000  96.520000 61.645000  96.670000 ;
      RECT 60.031000  96.670000 61.645000  96.820000 ;
      RECT 60.181000  96.820000 61.645000  96.970000 ;
      RECT 60.331000  96.970000 61.645000  97.120000 ;
      RECT 60.481000  97.120000 61.645000  97.270000 ;
      RECT 60.631000  97.270000 61.645000  97.420000 ;
      RECT 60.730000  97.519000 61.645000 172.635000 ;
      RECT 60.730000  97.519000 61.745000 172.535000 ;
      RECT 60.730000 172.535000 75.000000 189.915000 ;
      RECT 60.730000 172.635000 75.000000 189.915000 ;
      RECT 60.730000 172.635000 75.000000 198.000000 ;
      RECT 60.731000  97.420000 61.645000  97.520000 ;
    LAYER met4 ;
      RECT  4.820000 102.300000  7.470000 164.545000 ;
      RECT  5.440000 101.650000  5.945000 102.180000 ;
      RECT  5.440000 164.605000  5.945000 165.135000 ;
      RECT  6.070000 101.090000  8.445000 102.160000 ;
      RECT  6.070000 164.625000  8.445000 165.695000 ;
      RECT  6.555000 100.535000  7.060000 101.065000 ;
      RECT  6.555000 165.720000  7.060000 166.250000 ;
      RECT  7.350000  99.950000  9.725000 101.020000 ;
      RECT  7.350000 165.765000  9.725000 166.835000 ;
      RECT  7.535000 102.245000  8.040000 102.775000 ;
      RECT  7.535000 164.010000  8.040000 164.540000 ;
      RECT  7.750000  99.340000  8.255000  99.870000 ;
      RECT  7.750000 166.915000  8.255000 167.445000 ;
      RECT  8.340000  98.810000 10.715000  99.880000 ;
      RECT  8.415000 166.915000 10.700000 167.865000 ;
      RECT  8.650000 101.130000  9.155000 101.660000 ;
      RECT  8.650000 165.125000  9.155000 165.655000 ;
      RECT  8.825000  98.265000  9.330000  98.795000 ;
      RECT  8.825000 167.990000  9.330000 168.520000 ;
      RECT  9.460000  97.645000 11.835000  98.715000 ;
      RECT  9.460000 168.025000 11.835000 169.095000 ;
      RECT  9.845000  99.935000 10.350000 100.465000 ;
      RECT  9.845000 166.320000 10.350000 166.850000 ;
      RECT  9.985000  97.070000 10.490000  97.600000 ;
      RECT  9.985000 169.150000 10.490000 169.680000 ;
      RECT 10.595000  96.475000 11.850000  96.480000 ;
      RECT 10.595000  96.480000 11.835000  97.545000 ;
      RECT 10.610000 169.340000 11.745000 170.260000 ;
      RECT 10.920000  98.860000 11.425000  99.390000 ;
      RECT 10.920000 167.395000 11.425000 167.925000 ;
      RECT 11.095000  95.950000 11.850000  96.475000 ;
      RECT 11.095000 170.260000 11.850000 170.790000 ;
      RECT 11.965000  95.795000 12.835000  98.295000 ;
      RECT 11.965000 168.490000 12.835000 170.990000 ;
      RECT 25.035000  17.815000 25.465000  22.250000 ;
      RECT 25.035000  39.785000 25.365000  41.435000 ;
      RECT 62.225000  95.795000 63.095000  98.295000 ;
      RECT 62.225000 168.490000 63.095000 170.990000 ;
      RECT 63.225000  96.475000 64.465000  97.545000 ;
      RECT 63.225000  97.645000 65.600000  98.715000 ;
      RECT 63.225000 169.160000 64.465000 170.230000 ;
      RECT 63.235000 168.165000 65.495000 169.005000 ;
      RECT 63.635000  98.860000 64.140000  99.390000 ;
      RECT 63.635000 167.395000 64.140000 167.925000 ;
      RECT 64.345000  98.810000 66.720000  99.880000 ;
      RECT 64.345000 166.905000 66.720000 167.975000 ;
      RECT 64.570000  97.070000 65.075000  97.600000 ;
      RECT 64.570000 169.150000 65.075000 169.680000 ;
      RECT 64.710000  99.935000 65.215000 100.465000 ;
      RECT 64.710000 166.320000 65.215000 166.850000 ;
      RECT 65.335000  99.950000 67.710000 101.020000 ;
      RECT 65.335000 165.765000 67.710000 166.835000 ;
      RECT 65.730000  98.265000 66.235000  98.795000 ;
      RECT 65.730000 167.990000 66.235000 168.520000 ;
      RECT 65.905000 101.130000 66.410000 101.660000 ;
      RECT 65.905000 165.125000 66.410000 165.655000 ;
      RECT 66.615000 101.090000 68.990000 102.160000 ;
      RECT 66.615000 164.625000 68.990000 165.695000 ;
      RECT 66.805000  99.340000 67.310000  99.870000 ;
      RECT 66.805000 166.915000 67.310000 167.445000 ;
      RECT 67.020000 102.245000 70.110000 102.775000 ;
      RECT 67.020000 164.010000 70.165000 164.350000 ;
      RECT 67.020000 164.350000 67.525000 164.540000 ;
      RECT 67.515000 103.000000 70.165000 164.010000 ;
      RECT 68.000000 100.535000 68.505000 101.065000 ;
      RECT 68.000000 165.720000 68.505000 166.250000 ;
      RECT 69.115000 101.650000 69.620000 102.180000 ;
      RECT 69.115000 164.605000 69.620000 165.135000 ;
  END
END sky130_fd_io__top_ground_lvc_wpad
END LIBRARY
