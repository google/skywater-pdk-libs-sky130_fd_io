# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__corner_bus_overlay
  CLASS BLOCK ;
  FOREIGN sky130_fd_io__corner_bus_overlay ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  200.0000 BY  203.6650 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 56.790000 22.910000 59.770000 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.125000 0.000000 56.105000 18.475000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 52.030000 20.935000 55.010000 ;
    END
    PORT
      LAYER met4 ;
        RECT 48.365000 0.000000 51.345000 20.875000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 12.550000 3.785000 17.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.885000 0.000000 13.535000 1.270000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 12.650000 3.785000 17.100000 ;
    END
    PORT
      LAYER met5 ;
        RECT 8.985000 0.000000 13.435000 1.270000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 5.700000 2.350000 11.150000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.035000 0.000000 7.485000 1.270000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 5.800000 2.350000 11.050000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2.135000 0.000000 7.385000 1.270000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 18.600000 1.470000 22.050000 ;
    END
    PORT
      LAYER met4 ;
        RECT 14.935000 0.000000 18.385000 1.255000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 18.700000 1.470000 21.950000 ;
    END
    PORT
      LAYER met5 ;
        RECT 15.035000 0.000000 18.285000 1.255000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 23.450000 1.525000 28.100000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 73.700000 2.645000 98.665000 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.785000 0.000000 24.435000 1.270000 ;
    END
    PORT
      LAYER met4 ;
        RECT 70.035000 0.000000 95.000000 1.520000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 23.550000 1.525000 28.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 73.700000 2.645000 98.650000 ;
    END
    PORT
      LAYER met5 ;
        RECT 19.885000 0.000000 24.335000 1.270000 ;
    END
    PORT
      LAYER met5 ;
        RECT 70.035000 0.000000 94.985000 1.520000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 67.750000 1.480000 72.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.085000 0.000000 68.535000 1.270000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 67.850000 1.480000 72.100000 ;
    END
    PORT
      LAYER met5 ;
        RECT 64.185000 0.000000 68.435000 1.270000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 40.400000 1.335000 43.850000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.400000 19.575000 51.730000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 55.310000 21.550000 56.490000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 60.070000 23.175000 60.400000 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.735000 0.000000 40.185000 1.270000 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.735000 0.000000 48.065000 23.240000 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.645000 0.000000 52.825000 21.555000 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.405000 0.000000 56.735000 26.840000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 40.500000 1.335000 43.750000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 51.400000 23.155000 60.400000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.630000 54.950000 0.640000 54.960000 ;
    END
    PORT
      LAYER met5 ;
        RECT 36.840000 0.000000 40.085000 1.270000 ;
    END
    PORT
      LAYER met5 ;
        RECT 47.735000 0.000000 56.735000 26.820000 ;
    END
    PORT
      LAYER met5 ;
        RECT 52.020000 0.630000 52.030000 0.640000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 45.250000 1.475000 49.900000 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.585000 0.000000 46.235000 1.270000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 45.350000 1.475000 49.800000 ;
    END
    PORT
      LAYER met5 ;
        RECT 41.685000 0.000000 46.135000 1.270000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 179.450000 1.435000 203.665000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 29.500000 1.600000 34.150000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.630000 194.530000 0.640000 194.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 175.785000 0.000000 200.000000 1.270000 ;
    END
    PORT
      LAYER met4 ;
        RECT 190.865000 0.630000 190.875000 0.640000 ;
    END
    PORT
      LAYER met4 ;
        RECT 25.835000 0.000000 30.485000 1.270000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 179.450000 1.435000 203.665000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 29.600000 1.600000 34.050000 ;
    END
    PORT
      LAYER met5 ;
        RECT 175.785000 0.000000 200.000000 1.270000 ;
    END
    PORT
      LAYER met5 ;
        RECT 25.935000 0.000000 30.385000 1.270000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 61.900000 1.625000 66.350000 ;
    END
    PORT
      LAYER met4 ;
        RECT 58.235000 0.000000 62.685000 1.270000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 62.000000 1.625000 66.250000 ;
    END
    PORT
      LAYER met5 ;
        RECT 58.335000 0.000000 62.585000 1.270000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 35.550000 1.385000 39.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 31.885000 0.000000 35.335000 1.270000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 35.650000 1.385000 38.900000 ;
    END
    PORT
      LAYER met5 ;
        RECT 31.985000 0.000000 35.235000 1.270000 ;
    END
  END VSWITCH
  OBS
    LAYER met4 ;
      RECT  0.000000   1.255000   1.635000   1.670000 ;
      RECT  0.000000   1.670000  47.335000   5.300000 ;
      RECT  0.000000  11.550000  47.335000  12.150000 ;
      RECT  0.000000  17.600000  47.335000  18.200000 ;
      RECT  0.000000  22.450000  47.335000  23.050000 ;
      RECT  0.000000  28.500000 200.000000  29.100000 ;
      RECT  0.000000  34.550000 200.000000  35.150000 ;
      RECT  0.000000  39.400000 200.000000  40.000000 ;
      RECT  0.000000  44.250000 200.000000  44.850000 ;
      RECT  0.000000  50.300000 200.000000  51.000000 ;
      RECT  0.000000  60.800000 200.000000  61.500000 ;
      RECT  0.000000  66.750000 200.000000  67.350000 ;
      RECT  0.000000  72.600000 200.000000  73.300000 ;
      RECT  0.000000  99.065000 200.000000 179.050000 ;
      RECT  1.735000  40.000000 200.000000  44.250000 ;
      RECT  1.785000  35.150000 200.000000  39.400000 ;
      RECT  1.835000 179.050000 200.000000 203.665000 ;
      RECT  1.870000  18.200000  47.335000  22.450000 ;
      RECT  1.875000  44.850000 200.000000  50.300000 ;
      RECT  1.880000  67.350000 200.000000  72.600000 ;
      RECT  1.925000  23.050000  47.335000  23.640000 ;
      RECT  1.925000  23.640000  56.005000  27.240000 ;
      RECT  1.925000  27.240000 200.000000  28.500000 ;
      RECT  2.000000  29.100000 200.000000  34.550000 ;
      RECT  2.025000  61.500000 200.000000  66.750000 ;
      RECT  2.750000   5.300000  47.335000  11.550000 ;
      RECT  3.045000  73.300000 200.000000  99.065000 ;
      RECT  4.185000  12.150000  47.335000  17.600000 ;
      RECT  7.885000   1.255000   8.485000   1.670000 ;
      RECT 13.935000   1.255000  14.535000   1.655000 ;
      RECT 13.935000   1.655000  19.385000   1.670000 ;
      RECT 18.785000   1.255000  19.385000   1.655000 ;
      RECT 19.975000  51.000000 200.000000  51.630000 ;
      RECT 21.335000  51.630000 200.000000  54.910000 ;
      RECT 21.950000  54.910000 200.000000  56.390000 ;
      RECT 23.310000  56.390000 200.000000  59.670000 ;
      RECT 23.575000  59.670000 200.000000  60.800000 ;
      RECT 24.835000   1.255000  25.435000   1.670000 ;
      RECT 30.885000   1.255000  31.485000   1.670000 ;
      RECT 35.735000   1.255000  36.335000   1.670000 ;
      RECT 40.585000   1.255000  41.185000   1.670000 ;
      RECT 46.635000   1.255000  47.335000   1.670000 ;
      RECT 48.465000  21.275000  51.245000  21.955000 ;
      RECT 48.465000  21.955000  56.005000  23.640000 ;
      RECT 53.225000  18.875000  56.005000  21.955000 ;
      RECT 57.135000   1.255000  57.835000   1.670000 ;
      RECT 57.135000   1.670000  69.635000   1.920000 ;
      RECT 57.135000   1.920000 200.000000  27.240000 ;
      RECT 63.085000   1.255000  63.685000   1.670000 ;
      RECT 68.935000   1.255000  69.635000   1.670000 ;
      RECT 95.400000   1.255000 175.385000   1.670000 ;
      RECT 95.400000   1.670000 200.000000   1.920000 ;
    LAYER met5 ;
      RECT  0.000000   0.000000   0.535000   2.870000 ;
      RECT  0.000000   2.870000  46.135000   4.200000 ;
      RECT  0.000000 100.250000 200.000000 177.850000 ;
      RECT  2.935000  40.500000 200.000000  43.750000 ;
      RECT  2.985000  35.650000 200.000000  40.500000 ;
      RECT  3.035000 177.850000 200.000000 203.665000 ;
      RECT  3.070000  18.700000  46.135000  21.950000 ;
      RECT  3.075000  43.750000 200.000000  49.800000 ;
      RECT  3.080000  67.850000 200.000000  72.100000 ;
      RECT  3.125000  21.950000  46.135000  28.000000 ;
      RECT  3.200000  28.000000  46.135000  28.420000 ;
      RECT  3.200000  28.420000 200.000000  35.650000 ;
      RECT  3.225000  62.000000 200.000000  67.850000 ;
      RECT  3.950000   4.200000  46.135000  11.050000 ;
      RECT  4.245000  72.100000 200.000000 100.250000 ;
      RECT  5.385000  11.050000  46.135000  18.700000 ;
      RECT 15.035000   2.855000  18.285000   2.870000 ;
      RECT 24.755000  49.800000 200.000000  62.000000 ;
      RECT 58.335000   2.870000  68.435000   3.120000 ;
      RECT 58.335000   3.120000 200.000000  28.420000 ;
      RECT 96.585000   0.000000 174.185000   2.870000 ;
      RECT 96.585000   2.870000 200.000000   3.120000 ;
  END
END sky130_fd_io__corner_bus_overlay
END LIBRARY
