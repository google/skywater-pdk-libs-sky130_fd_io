# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_io__overlay_vddio_lvc
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 198 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 1.270000 54.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 1.270000 49.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 6.885000 1.270000 11.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 6.885000 75.000000 11.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 6.985000 1.270000 11.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 0.035000 1.270000 5.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 0.035000 75.000000 5.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 0.135000 1.270000 5.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 12.935000 0.965000 16.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 12.935000 75.000000 16.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 13.035000 0.965000 16.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.595000 68.035000 24.495000 82.665000 ;
        RECT 0.595000 82.665000 24.345000 82.815000 ;
        RECT 0.595000 82.815000 24.195000 82.965000 ;
        RECT 0.595000 82.965000 24.045000 83.115000 ;
        RECT 0.595000 83.115000 23.895000 83.265000 ;
        RECT 0.595000 83.265000 23.745000 83.415000 ;
        RECT 0.595000 83.415000 23.595000 83.565000 ;
        RECT 0.595000 83.565000 23.445000 83.715000 ;
        RECT 0.595000 83.715000 23.295000 83.865000 ;
        RECT 0.595000 83.865000 23.145000 84.015000 ;
        RECT 0.595000 84.015000 22.995000 84.165000 ;
        RECT 0.595000 84.165000 22.845000 84.315000 ;
        RECT 0.595000 84.315000 22.695000 84.465000 ;
        RECT 0.595000 84.465000 22.545000 84.615000 ;
        RECT 0.595000 84.615000 22.395000 84.765000 ;
        RECT 0.595000 84.765000 22.245000 84.915000 ;
        RECT 0.595000 84.915000 22.095000 85.065000 ;
        RECT 0.595000 85.065000 21.945000 85.215000 ;
        RECT 0.595000 85.215000 21.795000 85.365000 ;
        RECT 0.595000 85.365000 21.645000 85.515000 ;
        RECT 0.595000 85.515000 21.495000 85.665000 ;
        RECT 0.595000 85.665000 21.345000 85.815000 ;
        RECT 0.595000 85.815000 21.195000 85.965000 ;
        RECT 0.595000 85.965000 21.045000 86.115000 ;
        RECT 0.595000 86.115000 20.895000 86.265000 ;
        RECT 0.595000 86.265000 20.745000 86.415000 ;
        RECT 0.595000 86.415000 20.595000 86.565000 ;
        RECT 0.595000 86.565000 20.445000 86.715000 ;
        RECT 0.595000 86.715000 20.295000 86.865000 ;
        RECT 0.595000 86.865000 20.145000 87.015000 ;
        RECT 0.595000 87.015000 19.995000 87.165000 ;
        RECT 0.595000 87.165000 19.845000 87.315000 ;
        RECT 0.595000 87.315000 19.695000 87.465000 ;
        RECT 0.595000 87.465000 19.545000 87.615000 ;
        RECT 0.595000 87.615000 19.395000 87.765000 ;
        RECT 0.595000 87.765000 19.245000 87.915000 ;
        RECT 0.595000 87.915000 19.095000 88.065000 ;
        RECT 0.595000 88.065000 18.945000 88.215000 ;
        RECT 0.595000 88.215000 18.795000 88.365000 ;
        RECT 0.595000 88.365000 18.645000 88.515000 ;
        RECT 0.595000 88.515000 18.495000 88.665000 ;
        RECT 0.595000 88.665000 18.345000 88.815000 ;
        RECT 0.595000 88.815000 18.195000 88.965000 ;
        RECT 0.595000 88.965000 18.045000 89.115000 ;
        RECT 0.595000 89.115000 17.895000 89.265000 ;
        RECT 0.595000 89.265000 17.745000 89.415000 ;
        RECT 0.595000 89.415000 17.595000 89.565000 ;
        RECT 0.595000 89.565000 17.445000 89.715000 ;
        RECT 0.595000 89.715000 17.295000 89.865000 ;
        RECT 0.595000 89.865000 17.145000 90.015000 ;
        RECT 0.595000 90.015000 16.995000 90.165000 ;
        RECT 0.595000 90.165000 16.845000 90.315000 ;
        RECT 0.595000 90.315000 16.695000 90.465000 ;
        RECT 0.595000 90.465000 16.545000 90.615000 ;
        RECT 0.595000 90.615000 16.395000 90.765000 ;
        RECT 0.595000 90.765000 16.245000 90.915000 ;
        RECT 0.595000 90.915000 16.095000 91.065000 ;
        RECT 0.595000 91.065000 15.945000 91.215000 ;
        RECT 0.595000 91.215000 15.795000 91.365000 ;
        RECT 0.595000 91.365000 15.645000 91.515000 ;
        RECT 0.595000 91.515000 15.495000 91.665000 ;
        RECT 0.595000 91.665000 15.345000 91.815000 ;
        RECT 0.595000 91.815000 15.195000 91.965000 ;
        RECT 0.595000 91.965000 15.045000 92.115000 ;
        RECT 0.595000 92.115000 14.895000 92.265000 ;
        RECT 0.595000 92.265000 14.745000 92.415000 ;
        RECT 0.595000 92.415000 14.595000 92.565000 ;
        RECT 0.595000 92.565000 14.445000 92.715000 ;
        RECT 0.595000 92.715000 14.295000 92.865000 ;
        RECT 0.595000 92.865000 14.205000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.600000 17.790000 24.500000 22.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000 17.790000 74.655000 22.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.760000 68.035000 74.660000 82.665000 ;
        RECT 50.910000 82.665000 74.660000 82.815000 ;
        RECT 51.060000 82.815000 74.660000 82.965000 ;
        RECT 51.210000 82.965000 74.660000 83.115000 ;
        RECT 51.360000 83.115000 74.660000 83.265000 ;
        RECT 51.510000 83.265000 74.660000 83.415000 ;
        RECT 51.660000 83.415000 74.660000 83.565000 ;
        RECT 51.810000 83.565000 74.660000 83.715000 ;
        RECT 51.960000 83.715000 74.660000 83.865000 ;
        RECT 52.110000 83.865000 74.660000 84.015000 ;
        RECT 52.260000 84.015000 74.660000 84.165000 ;
        RECT 52.410000 84.165000 74.660000 84.315000 ;
        RECT 52.560000 84.315000 74.660000 84.465000 ;
        RECT 52.710000 84.465000 74.660000 84.615000 ;
        RECT 52.860000 84.615000 74.660000 84.765000 ;
        RECT 53.010000 84.765000 74.660000 84.915000 ;
        RECT 53.160000 84.915000 74.660000 85.065000 ;
        RECT 53.310000 85.065000 74.660000 85.215000 ;
        RECT 53.460000 85.215000 74.660000 85.365000 ;
        RECT 53.610000 85.365000 74.660000 85.515000 ;
        RECT 53.760000 85.515000 74.660000 85.665000 ;
        RECT 53.910000 85.665000 74.660000 85.815000 ;
        RECT 54.060000 85.815000 74.660000 85.965000 ;
        RECT 54.210000 85.965000 74.660000 86.115000 ;
        RECT 54.360000 86.115000 74.660000 86.265000 ;
        RECT 54.510000 86.265000 74.660000 86.415000 ;
        RECT 54.660000 86.415000 74.660000 86.565000 ;
        RECT 54.810000 86.565000 74.660000 86.715000 ;
        RECT 54.960000 86.715000 74.660000 86.865000 ;
        RECT 55.110000 86.865000 74.660000 87.015000 ;
        RECT 55.260000 87.015000 74.660000 87.165000 ;
        RECT 55.410000 87.165000 74.660000 87.315000 ;
        RECT 55.560000 87.315000 74.660000 87.465000 ;
        RECT 55.710000 87.465000 74.660000 87.615000 ;
        RECT 55.860000 87.615000 74.660000 87.765000 ;
        RECT 56.010000 87.765000 74.660000 87.915000 ;
        RECT 56.160000 87.915000 74.660000 88.065000 ;
        RECT 56.310000 88.065000 74.660000 88.215000 ;
        RECT 56.460000 88.215000 74.660000 88.365000 ;
        RECT 56.610000 88.365000 74.660000 88.515000 ;
        RECT 56.760000 88.515000 74.660000 88.665000 ;
        RECT 56.910000 88.665000 74.660000 88.815000 ;
        RECT 57.060000 88.815000 74.660000 88.965000 ;
        RECT 57.210000 88.965000 74.660000 89.115000 ;
        RECT 57.360000 89.115000 74.660000 89.265000 ;
        RECT 57.510000 89.265000 74.660000 89.415000 ;
        RECT 57.660000 89.415000 74.660000 89.565000 ;
        RECT 57.810000 89.565000 74.660000 89.715000 ;
        RECT 57.960000 89.715000 74.660000 89.865000 ;
        RECT 58.110000 89.865000 74.660000 90.015000 ;
        RECT 58.260000 90.015000 74.660000 90.165000 ;
        RECT 58.410000 90.165000 74.660000 90.315000 ;
        RECT 58.560000 90.315000 74.660000 90.465000 ;
        RECT 58.710000 90.465000 74.660000 90.615000 ;
        RECT 58.860000 90.615000 74.660000 90.765000 ;
        RECT 59.010000 90.765000 74.660000 90.915000 ;
        RECT 59.160000 90.915000 74.660000 91.065000 ;
        RECT 59.310000 91.065000 74.660000 91.215000 ;
        RECT 59.460000 91.215000 74.660000 91.365000 ;
        RECT 59.610000 91.365000 74.660000 91.515000 ;
        RECT 59.760000 91.515000 74.660000 91.665000 ;
        RECT 59.910000 91.665000 74.660000 91.815000 ;
        RECT 60.060000 91.815000 74.660000 91.965000 ;
        RECT 60.210000 91.965000 74.660000 92.115000 ;
        RECT 60.360000 92.115000 74.660000 92.265000 ;
        RECT 60.510000 92.265000 74.660000 92.415000 ;
        RECT 60.660000 92.415000 74.660000 92.565000 ;
        RECT 60.810000 92.565000 74.660000 92.715000 ;
        RECT 60.960000 92.715000 74.660000 92.865000 ;
        RECT 61.055000 92.865000 74.660000 92.960000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 17.785000 24.475000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 68.035000  1.270000 68.060000 ;
        RECT 0.000000 68.060000 24.500000 82.625000 ;
        RECT 0.000000 82.625000  1.270000 82.790000 ;
        RECT 0.000000 82.790000 14.105000 92.960000 ;
        RECT 0.000000 92.960000  1.270000 93.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 14.255000 90.950000 15.365000 91.710000 ;
    END
    PORT
      LAYER met4 ;
        RECT 14.270000 88.345000 16.250000 90.820000 ;
    END
    PORT
      LAYER met4 ;
        RECT 14.375000 82.990000 18.855000 88.140000 ;
    END
    PORT
      LAYER met4 ;
        RECT 16.415000 88.365000 17.525000 89.530000 ;
    END
    PORT
      LAYER met4 ;
        RECT 18.995000 85.810000 20.065000 87.015000 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.170000 82.945000 21.450000 85.590000 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.650000 82.855000 22.770000 84.285000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.755000 68.060000 75.000000 82.625000 ;
        RECT 61.150000 82.785000 75.000000 92.965000 ;
        RECT 73.730000 68.035000 75.000000 68.060000 ;
        RECT 73.730000 82.625000 75.000000 82.785000 ;
        RECT 73.730000 92.965000 75.000000 93.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.780000 17.785000 75.000000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 52.485000 82.855000 53.605000 84.285000 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.805000 82.945000 56.085000 85.590000 ;
    END
    PORT
      LAYER met4 ;
        RECT 55.190000 85.810000 56.260000 87.015000 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.400000 82.990000 60.880000 88.140000 ;
    END
    PORT
      LAYER met4 ;
        RECT 57.730000 88.365000 58.840000 89.530000 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.005000 88.345000 60.985000 90.820000 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.890000 90.950000 61.000000 91.710000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 17.885000 1.270000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 68.035000 1.270000 92.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 17.885000 75.000000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.690000 17.860000  0.890000 18.060000 ;
        RECT  0.690000 18.290000  0.890000 18.490000 ;
        RECT  0.690000 18.720000  0.890000 18.920000 ;
        RECT  0.690000 19.150000  0.890000 19.350000 ;
        RECT  0.690000 19.580000  0.890000 19.780000 ;
        RECT  0.690000 20.010000  0.890000 20.210000 ;
        RECT  0.690000 20.440000  0.890000 20.640000 ;
        RECT  0.690000 20.870000  0.890000 21.070000 ;
        RECT  0.690000 21.300000  0.890000 21.500000 ;
        RECT  0.690000 21.730000  0.890000 21.930000 ;
        RECT  0.690000 22.160000  0.890000 22.360000 ;
        RECT  0.735000 82.855000  0.935000 83.055000 ;
        RECT  0.735000 83.265000  0.935000 83.465000 ;
        RECT  0.735000 83.675000  0.935000 83.875000 ;
        RECT  0.735000 84.085000  0.935000 84.285000 ;
        RECT  0.735000 84.495000  0.935000 84.695000 ;
        RECT  0.735000 84.905000  0.935000 85.105000 ;
        RECT  0.735000 85.315000  0.935000 85.515000 ;
        RECT  0.735000 85.725000  0.935000 85.925000 ;
        RECT  0.735000 86.135000  0.935000 86.335000 ;
        RECT  0.735000 86.545000  0.935000 86.745000 ;
        RECT  0.735000 86.955000  0.935000 87.155000 ;
        RECT  0.735000 87.365000  0.935000 87.565000 ;
        RECT  0.735000 87.775000  0.935000 87.975000 ;
        RECT  0.735000 88.185000  0.935000 88.385000 ;
        RECT  0.735000 88.595000  0.935000 88.795000 ;
        RECT  0.735000 89.005000  0.935000 89.205000 ;
        RECT  0.735000 89.415000  0.935000 89.615000 ;
        RECT  0.735000 89.825000  0.935000 90.025000 ;
        RECT  0.735000 90.235000  0.935000 90.435000 ;
        RECT  0.735000 90.645000  0.935000 90.845000 ;
        RECT  0.735000 91.055000  0.935000 91.255000 ;
        RECT  0.735000 91.465000  0.935000 91.665000 ;
        RECT  0.735000 91.875000  0.935000 92.075000 ;
        RECT  0.735000 92.285000  0.935000 92.485000 ;
        RECT  0.735000 92.695000  0.935000 92.895000 ;
        RECT  0.845000 68.125000  1.045000 68.325000 ;
        RECT  0.845000 68.535000  1.045000 68.735000 ;
        RECT  0.845000 68.945000  1.045000 69.145000 ;
        RECT  0.845000 69.355000  1.045000 69.555000 ;
        RECT  0.845000 69.765000  1.045000 69.965000 ;
        RECT  0.845000 70.175000  1.045000 70.375000 ;
        RECT  0.845000 70.585000  1.045000 70.785000 ;
        RECT  0.845000 70.995000  1.045000 71.195000 ;
        RECT  0.845000 71.405000  1.045000 71.605000 ;
        RECT  0.845000 71.815000  1.045000 72.015000 ;
        RECT  0.845000 72.225000  1.045000 72.425000 ;
        RECT  0.845000 72.635000  1.045000 72.835000 ;
        RECT  0.845000 73.045000  1.045000 73.245000 ;
        RECT  0.845000 73.450000  1.045000 73.650000 ;
        RECT  0.845000 73.855000  1.045000 74.055000 ;
        RECT  0.845000 74.260000  1.045000 74.460000 ;
        RECT  0.845000 74.665000  1.045000 74.865000 ;
        RECT  0.845000 75.070000  1.045000 75.270000 ;
        RECT  0.845000 75.475000  1.045000 75.675000 ;
        RECT  0.845000 75.880000  1.045000 76.080000 ;
        RECT  0.845000 76.285000  1.045000 76.485000 ;
        RECT  0.845000 76.690000  1.045000 76.890000 ;
        RECT  0.845000 77.095000  1.045000 77.295000 ;
        RECT  0.845000 77.500000  1.045000 77.700000 ;
        RECT  0.845000 77.905000  1.045000 78.105000 ;
        RECT  0.845000 78.310000  1.045000 78.510000 ;
        RECT  0.845000 78.715000  1.045000 78.915000 ;
        RECT  0.845000 79.120000  1.045000 79.320000 ;
        RECT  0.845000 79.525000  1.045000 79.725000 ;
        RECT  0.845000 79.930000  1.045000 80.130000 ;
        RECT  0.845000 80.335000  1.045000 80.535000 ;
        RECT  0.845000 80.740000  1.045000 80.940000 ;
        RECT  0.845000 81.145000  1.045000 81.345000 ;
        RECT  0.845000 81.550000  1.045000 81.750000 ;
        RECT  0.845000 81.955000  1.045000 82.155000 ;
        RECT  0.845000 82.360000  1.045000 82.560000 ;
        RECT  1.095000 17.860000  1.295000 18.060000 ;
        RECT  1.095000 18.290000  1.295000 18.490000 ;
        RECT  1.095000 18.720000  1.295000 18.920000 ;
        RECT  1.095000 19.150000  1.295000 19.350000 ;
        RECT  1.095000 19.580000  1.295000 19.780000 ;
        RECT  1.095000 20.010000  1.295000 20.210000 ;
        RECT  1.095000 20.440000  1.295000 20.640000 ;
        RECT  1.095000 20.870000  1.295000 21.070000 ;
        RECT  1.095000 21.300000  1.295000 21.500000 ;
        RECT  1.095000 21.730000  1.295000 21.930000 ;
        RECT  1.095000 22.160000  1.295000 22.360000 ;
        RECT  1.145000 82.855000  1.345000 83.055000 ;
        RECT  1.145000 83.265000  1.345000 83.465000 ;
        RECT  1.145000 83.675000  1.345000 83.875000 ;
        RECT  1.145000 84.085000  1.345000 84.285000 ;
        RECT  1.145000 84.495000  1.345000 84.695000 ;
        RECT  1.145000 84.905000  1.345000 85.105000 ;
        RECT  1.145000 85.315000  1.345000 85.515000 ;
        RECT  1.145000 85.725000  1.345000 85.925000 ;
        RECT  1.145000 86.135000  1.345000 86.335000 ;
        RECT  1.145000 86.545000  1.345000 86.745000 ;
        RECT  1.145000 86.955000  1.345000 87.155000 ;
        RECT  1.145000 87.365000  1.345000 87.565000 ;
        RECT  1.145000 87.775000  1.345000 87.975000 ;
        RECT  1.145000 88.185000  1.345000 88.385000 ;
        RECT  1.145000 88.595000  1.345000 88.795000 ;
        RECT  1.145000 89.005000  1.345000 89.205000 ;
        RECT  1.145000 89.415000  1.345000 89.615000 ;
        RECT  1.145000 89.825000  1.345000 90.025000 ;
        RECT  1.145000 90.235000  1.345000 90.435000 ;
        RECT  1.145000 90.645000  1.345000 90.845000 ;
        RECT  1.145000 91.055000  1.345000 91.255000 ;
        RECT  1.145000 91.465000  1.345000 91.665000 ;
        RECT  1.145000 91.875000  1.345000 92.075000 ;
        RECT  1.145000 92.285000  1.345000 92.485000 ;
        RECT  1.145000 92.695000  1.345000 92.895000 ;
        RECT  1.245000 68.125000  1.445000 68.325000 ;
        RECT  1.245000 68.535000  1.445000 68.735000 ;
        RECT  1.245000 68.945000  1.445000 69.145000 ;
        RECT  1.245000 69.355000  1.445000 69.555000 ;
        RECT  1.245000 69.765000  1.445000 69.965000 ;
        RECT  1.245000 70.175000  1.445000 70.375000 ;
        RECT  1.245000 70.585000  1.445000 70.785000 ;
        RECT  1.245000 70.995000  1.445000 71.195000 ;
        RECT  1.245000 71.405000  1.445000 71.605000 ;
        RECT  1.245000 71.815000  1.445000 72.015000 ;
        RECT  1.245000 72.225000  1.445000 72.425000 ;
        RECT  1.245000 72.635000  1.445000 72.835000 ;
        RECT  1.245000 73.045000  1.445000 73.245000 ;
        RECT  1.245000 73.450000  1.445000 73.650000 ;
        RECT  1.245000 73.855000  1.445000 74.055000 ;
        RECT  1.245000 74.260000  1.445000 74.460000 ;
        RECT  1.245000 74.665000  1.445000 74.865000 ;
        RECT  1.245000 75.070000  1.445000 75.270000 ;
        RECT  1.245000 75.475000  1.445000 75.675000 ;
        RECT  1.245000 75.880000  1.445000 76.080000 ;
        RECT  1.245000 76.285000  1.445000 76.485000 ;
        RECT  1.245000 76.690000  1.445000 76.890000 ;
        RECT  1.245000 77.095000  1.445000 77.295000 ;
        RECT  1.245000 77.500000  1.445000 77.700000 ;
        RECT  1.245000 77.905000  1.445000 78.105000 ;
        RECT  1.245000 78.310000  1.445000 78.510000 ;
        RECT  1.245000 78.715000  1.445000 78.915000 ;
        RECT  1.245000 79.120000  1.445000 79.320000 ;
        RECT  1.245000 79.525000  1.445000 79.725000 ;
        RECT  1.245000 79.930000  1.445000 80.130000 ;
        RECT  1.245000 80.335000  1.445000 80.535000 ;
        RECT  1.245000 80.740000  1.445000 80.940000 ;
        RECT  1.245000 81.145000  1.445000 81.345000 ;
        RECT  1.245000 81.550000  1.445000 81.750000 ;
        RECT  1.245000 81.955000  1.445000 82.155000 ;
        RECT  1.245000 82.360000  1.445000 82.560000 ;
        RECT  1.500000 17.860000  1.700000 18.060000 ;
        RECT  1.500000 18.290000  1.700000 18.490000 ;
        RECT  1.500000 18.720000  1.700000 18.920000 ;
        RECT  1.500000 19.150000  1.700000 19.350000 ;
        RECT  1.500000 19.580000  1.700000 19.780000 ;
        RECT  1.500000 20.010000  1.700000 20.210000 ;
        RECT  1.500000 20.440000  1.700000 20.640000 ;
        RECT  1.500000 20.870000  1.700000 21.070000 ;
        RECT  1.500000 21.300000  1.700000 21.500000 ;
        RECT  1.500000 21.730000  1.700000 21.930000 ;
        RECT  1.500000 22.160000  1.700000 22.360000 ;
        RECT  1.555000 82.855000  1.755000 83.055000 ;
        RECT  1.555000 83.265000  1.755000 83.465000 ;
        RECT  1.555000 83.675000  1.755000 83.875000 ;
        RECT  1.555000 84.085000  1.755000 84.285000 ;
        RECT  1.555000 84.495000  1.755000 84.695000 ;
        RECT  1.555000 84.905000  1.755000 85.105000 ;
        RECT  1.555000 85.315000  1.755000 85.515000 ;
        RECT  1.555000 85.725000  1.755000 85.925000 ;
        RECT  1.555000 86.135000  1.755000 86.335000 ;
        RECT  1.555000 86.545000  1.755000 86.745000 ;
        RECT  1.555000 86.955000  1.755000 87.155000 ;
        RECT  1.555000 87.365000  1.755000 87.565000 ;
        RECT  1.555000 87.775000  1.755000 87.975000 ;
        RECT  1.555000 88.185000  1.755000 88.385000 ;
        RECT  1.555000 88.595000  1.755000 88.795000 ;
        RECT  1.555000 89.005000  1.755000 89.205000 ;
        RECT  1.555000 89.415000  1.755000 89.615000 ;
        RECT  1.555000 89.825000  1.755000 90.025000 ;
        RECT  1.555000 90.235000  1.755000 90.435000 ;
        RECT  1.555000 90.645000  1.755000 90.845000 ;
        RECT  1.555000 91.055000  1.755000 91.255000 ;
        RECT  1.555000 91.465000  1.755000 91.665000 ;
        RECT  1.555000 91.875000  1.755000 92.075000 ;
        RECT  1.555000 92.285000  1.755000 92.485000 ;
        RECT  1.555000 92.695000  1.755000 92.895000 ;
        RECT  1.645000 68.125000  1.845000 68.325000 ;
        RECT  1.645000 68.535000  1.845000 68.735000 ;
        RECT  1.645000 68.945000  1.845000 69.145000 ;
        RECT  1.645000 69.355000  1.845000 69.555000 ;
        RECT  1.645000 69.765000  1.845000 69.965000 ;
        RECT  1.645000 70.175000  1.845000 70.375000 ;
        RECT  1.645000 70.585000  1.845000 70.785000 ;
        RECT  1.645000 70.995000  1.845000 71.195000 ;
        RECT  1.645000 71.405000  1.845000 71.605000 ;
        RECT  1.645000 71.815000  1.845000 72.015000 ;
        RECT  1.645000 72.225000  1.845000 72.425000 ;
        RECT  1.645000 72.635000  1.845000 72.835000 ;
        RECT  1.645000 73.045000  1.845000 73.245000 ;
        RECT  1.645000 73.450000  1.845000 73.650000 ;
        RECT  1.645000 73.855000  1.845000 74.055000 ;
        RECT  1.645000 74.260000  1.845000 74.460000 ;
        RECT  1.645000 74.665000  1.845000 74.865000 ;
        RECT  1.645000 75.070000  1.845000 75.270000 ;
        RECT  1.645000 75.475000  1.845000 75.675000 ;
        RECT  1.645000 75.880000  1.845000 76.080000 ;
        RECT  1.645000 76.285000  1.845000 76.485000 ;
        RECT  1.645000 76.690000  1.845000 76.890000 ;
        RECT  1.645000 77.095000  1.845000 77.295000 ;
        RECT  1.645000 77.500000  1.845000 77.700000 ;
        RECT  1.645000 77.905000  1.845000 78.105000 ;
        RECT  1.645000 78.310000  1.845000 78.510000 ;
        RECT  1.645000 78.715000  1.845000 78.915000 ;
        RECT  1.645000 79.120000  1.845000 79.320000 ;
        RECT  1.645000 79.525000  1.845000 79.725000 ;
        RECT  1.645000 79.930000  1.845000 80.130000 ;
        RECT  1.645000 80.335000  1.845000 80.535000 ;
        RECT  1.645000 80.740000  1.845000 80.940000 ;
        RECT  1.645000 81.145000  1.845000 81.345000 ;
        RECT  1.645000 81.550000  1.845000 81.750000 ;
        RECT  1.645000 81.955000  1.845000 82.155000 ;
        RECT  1.645000 82.360000  1.845000 82.560000 ;
        RECT  1.905000 17.860000  2.105000 18.060000 ;
        RECT  1.905000 18.290000  2.105000 18.490000 ;
        RECT  1.905000 18.720000  2.105000 18.920000 ;
        RECT  1.905000 19.150000  2.105000 19.350000 ;
        RECT  1.905000 19.580000  2.105000 19.780000 ;
        RECT  1.905000 20.010000  2.105000 20.210000 ;
        RECT  1.905000 20.440000  2.105000 20.640000 ;
        RECT  1.905000 20.870000  2.105000 21.070000 ;
        RECT  1.905000 21.300000  2.105000 21.500000 ;
        RECT  1.905000 21.730000  2.105000 21.930000 ;
        RECT  1.905000 22.160000  2.105000 22.360000 ;
        RECT  1.965000 82.855000  2.165000 83.055000 ;
        RECT  1.965000 83.265000  2.165000 83.465000 ;
        RECT  1.965000 83.675000  2.165000 83.875000 ;
        RECT  1.965000 84.085000  2.165000 84.285000 ;
        RECT  1.965000 84.495000  2.165000 84.695000 ;
        RECT  1.965000 84.905000  2.165000 85.105000 ;
        RECT  1.965000 85.315000  2.165000 85.515000 ;
        RECT  1.965000 85.725000  2.165000 85.925000 ;
        RECT  1.965000 86.135000  2.165000 86.335000 ;
        RECT  1.965000 86.545000  2.165000 86.745000 ;
        RECT  1.965000 86.955000  2.165000 87.155000 ;
        RECT  1.965000 87.365000  2.165000 87.565000 ;
        RECT  1.965000 87.775000  2.165000 87.975000 ;
        RECT  1.965000 88.185000  2.165000 88.385000 ;
        RECT  1.965000 88.595000  2.165000 88.795000 ;
        RECT  1.965000 89.005000  2.165000 89.205000 ;
        RECT  1.965000 89.415000  2.165000 89.615000 ;
        RECT  1.965000 89.825000  2.165000 90.025000 ;
        RECT  1.965000 90.235000  2.165000 90.435000 ;
        RECT  1.965000 90.645000  2.165000 90.845000 ;
        RECT  1.965000 91.055000  2.165000 91.255000 ;
        RECT  1.965000 91.465000  2.165000 91.665000 ;
        RECT  1.965000 91.875000  2.165000 92.075000 ;
        RECT  1.965000 92.285000  2.165000 92.485000 ;
        RECT  1.965000 92.695000  2.165000 92.895000 ;
        RECT  2.045000 68.125000  2.245000 68.325000 ;
        RECT  2.045000 68.535000  2.245000 68.735000 ;
        RECT  2.045000 68.945000  2.245000 69.145000 ;
        RECT  2.045000 69.355000  2.245000 69.555000 ;
        RECT  2.045000 69.765000  2.245000 69.965000 ;
        RECT  2.045000 70.175000  2.245000 70.375000 ;
        RECT  2.045000 70.585000  2.245000 70.785000 ;
        RECT  2.045000 70.995000  2.245000 71.195000 ;
        RECT  2.045000 71.405000  2.245000 71.605000 ;
        RECT  2.045000 71.815000  2.245000 72.015000 ;
        RECT  2.045000 72.225000  2.245000 72.425000 ;
        RECT  2.045000 72.635000  2.245000 72.835000 ;
        RECT  2.045000 73.045000  2.245000 73.245000 ;
        RECT  2.045000 73.450000  2.245000 73.650000 ;
        RECT  2.045000 73.855000  2.245000 74.055000 ;
        RECT  2.045000 74.260000  2.245000 74.460000 ;
        RECT  2.045000 74.665000  2.245000 74.865000 ;
        RECT  2.045000 75.070000  2.245000 75.270000 ;
        RECT  2.045000 75.475000  2.245000 75.675000 ;
        RECT  2.045000 75.880000  2.245000 76.080000 ;
        RECT  2.045000 76.285000  2.245000 76.485000 ;
        RECT  2.045000 76.690000  2.245000 76.890000 ;
        RECT  2.045000 77.095000  2.245000 77.295000 ;
        RECT  2.045000 77.500000  2.245000 77.700000 ;
        RECT  2.045000 77.905000  2.245000 78.105000 ;
        RECT  2.045000 78.310000  2.245000 78.510000 ;
        RECT  2.045000 78.715000  2.245000 78.915000 ;
        RECT  2.045000 79.120000  2.245000 79.320000 ;
        RECT  2.045000 79.525000  2.245000 79.725000 ;
        RECT  2.045000 79.930000  2.245000 80.130000 ;
        RECT  2.045000 80.335000  2.245000 80.535000 ;
        RECT  2.045000 80.740000  2.245000 80.940000 ;
        RECT  2.045000 81.145000  2.245000 81.345000 ;
        RECT  2.045000 81.550000  2.245000 81.750000 ;
        RECT  2.045000 81.955000  2.245000 82.155000 ;
        RECT  2.045000 82.360000  2.245000 82.560000 ;
        RECT  2.310000 17.860000  2.510000 18.060000 ;
        RECT  2.310000 18.290000  2.510000 18.490000 ;
        RECT  2.310000 18.720000  2.510000 18.920000 ;
        RECT  2.310000 19.150000  2.510000 19.350000 ;
        RECT  2.310000 19.580000  2.510000 19.780000 ;
        RECT  2.310000 20.010000  2.510000 20.210000 ;
        RECT  2.310000 20.440000  2.510000 20.640000 ;
        RECT  2.310000 20.870000  2.510000 21.070000 ;
        RECT  2.310000 21.300000  2.510000 21.500000 ;
        RECT  2.310000 21.730000  2.510000 21.930000 ;
        RECT  2.310000 22.160000  2.510000 22.360000 ;
        RECT  2.375000 82.855000  2.575000 83.055000 ;
        RECT  2.375000 83.265000  2.575000 83.465000 ;
        RECT  2.375000 83.675000  2.575000 83.875000 ;
        RECT  2.375000 84.085000  2.575000 84.285000 ;
        RECT  2.375000 84.495000  2.575000 84.695000 ;
        RECT  2.375000 84.905000  2.575000 85.105000 ;
        RECT  2.375000 85.315000  2.575000 85.515000 ;
        RECT  2.375000 85.725000  2.575000 85.925000 ;
        RECT  2.375000 86.135000  2.575000 86.335000 ;
        RECT  2.375000 86.545000  2.575000 86.745000 ;
        RECT  2.375000 86.955000  2.575000 87.155000 ;
        RECT  2.375000 87.365000  2.575000 87.565000 ;
        RECT  2.375000 87.775000  2.575000 87.975000 ;
        RECT  2.375000 88.185000  2.575000 88.385000 ;
        RECT  2.375000 88.595000  2.575000 88.795000 ;
        RECT  2.375000 89.005000  2.575000 89.205000 ;
        RECT  2.375000 89.415000  2.575000 89.615000 ;
        RECT  2.375000 89.825000  2.575000 90.025000 ;
        RECT  2.375000 90.235000  2.575000 90.435000 ;
        RECT  2.375000 90.645000  2.575000 90.845000 ;
        RECT  2.375000 91.055000  2.575000 91.255000 ;
        RECT  2.375000 91.465000  2.575000 91.665000 ;
        RECT  2.375000 91.875000  2.575000 92.075000 ;
        RECT  2.375000 92.285000  2.575000 92.485000 ;
        RECT  2.375000 92.695000  2.575000 92.895000 ;
        RECT  2.445000 68.125000  2.645000 68.325000 ;
        RECT  2.445000 68.535000  2.645000 68.735000 ;
        RECT  2.445000 68.945000  2.645000 69.145000 ;
        RECT  2.445000 69.355000  2.645000 69.555000 ;
        RECT  2.445000 69.765000  2.645000 69.965000 ;
        RECT  2.445000 70.175000  2.645000 70.375000 ;
        RECT  2.445000 70.585000  2.645000 70.785000 ;
        RECT  2.445000 70.995000  2.645000 71.195000 ;
        RECT  2.445000 71.405000  2.645000 71.605000 ;
        RECT  2.445000 71.815000  2.645000 72.015000 ;
        RECT  2.445000 72.225000  2.645000 72.425000 ;
        RECT  2.445000 72.635000  2.645000 72.835000 ;
        RECT  2.445000 73.045000  2.645000 73.245000 ;
        RECT  2.445000 73.450000  2.645000 73.650000 ;
        RECT  2.445000 73.855000  2.645000 74.055000 ;
        RECT  2.445000 74.260000  2.645000 74.460000 ;
        RECT  2.445000 74.665000  2.645000 74.865000 ;
        RECT  2.445000 75.070000  2.645000 75.270000 ;
        RECT  2.445000 75.475000  2.645000 75.675000 ;
        RECT  2.445000 75.880000  2.645000 76.080000 ;
        RECT  2.445000 76.285000  2.645000 76.485000 ;
        RECT  2.445000 76.690000  2.645000 76.890000 ;
        RECT  2.445000 77.095000  2.645000 77.295000 ;
        RECT  2.445000 77.500000  2.645000 77.700000 ;
        RECT  2.445000 77.905000  2.645000 78.105000 ;
        RECT  2.445000 78.310000  2.645000 78.510000 ;
        RECT  2.445000 78.715000  2.645000 78.915000 ;
        RECT  2.445000 79.120000  2.645000 79.320000 ;
        RECT  2.445000 79.525000  2.645000 79.725000 ;
        RECT  2.445000 79.930000  2.645000 80.130000 ;
        RECT  2.445000 80.335000  2.645000 80.535000 ;
        RECT  2.445000 80.740000  2.645000 80.940000 ;
        RECT  2.445000 81.145000  2.645000 81.345000 ;
        RECT  2.445000 81.550000  2.645000 81.750000 ;
        RECT  2.445000 81.955000  2.645000 82.155000 ;
        RECT  2.445000 82.360000  2.645000 82.560000 ;
        RECT  2.715000 17.860000  2.915000 18.060000 ;
        RECT  2.715000 18.290000  2.915000 18.490000 ;
        RECT  2.715000 18.720000  2.915000 18.920000 ;
        RECT  2.715000 19.150000  2.915000 19.350000 ;
        RECT  2.715000 19.580000  2.915000 19.780000 ;
        RECT  2.715000 20.010000  2.915000 20.210000 ;
        RECT  2.715000 20.440000  2.915000 20.640000 ;
        RECT  2.715000 20.870000  2.915000 21.070000 ;
        RECT  2.715000 21.300000  2.915000 21.500000 ;
        RECT  2.715000 21.730000  2.915000 21.930000 ;
        RECT  2.715000 22.160000  2.915000 22.360000 ;
        RECT  2.785000 82.855000  2.985000 83.055000 ;
        RECT  2.785000 83.265000  2.985000 83.465000 ;
        RECT  2.785000 83.675000  2.985000 83.875000 ;
        RECT  2.785000 84.085000  2.985000 84.285000 ;
        RECT  2.785000 84.495000  2.985000 84.695000 ;
        RECT  2.785000 84.905000  2.985000 85.105000 ;
        RECT  2.785000 85.315000  2.985000 85.515000 ;
        RECT  2.785000 85.725000  2.985000 85.925000 ;
        RECT  2.785000 86.135000  2.985000 86.335000 ;
        RECT  2.785000 86.545000  2.985000 86.745000 ;
        RECT  2.785000 86.955000  2.985000 87.155000 ;
        RECT  2.785000 87.365000  2.985000 87.565000 ;
        RECT  2.785000 87.775000  2.985000 87.975000 ;
        RECT  2.785000 88.185000  2.985000 88.385000 ;
        RECT  2.785000 88.595000  2.985000 88.795000 ;
        RECT  2.785000 89.005000  2.985000 89.205000 ;
        RECT  2.785000 89.415000  2.985000 89.615000 ;
        RECT  2.785000 89.825000  2.985000 90.025000 ;
        RECT  2.785000 90.235000  2.985000 90.435000 ;
        RECT  2.785000 90.645000  2.985000 90.845000 ;
        RECT  2.785000 91.055000  2.985000 91.255000 ;
        RECT  2.785000 91.465000  2.985000 91.665000 ;
        RECT  2.785000 91.875000  2.985000 92.075000 ;
        RECT  2.785000 92.285000  2.985000 92.485000 ;
        RECT  2.785000 92.695000  2.985000 92.895000 ;
        RECT  2.845000 68.125000  3.045000 68.325000 ;
        RECT  2.845000 68.535000  3.045000 68.735000 ;
        RECT  2.845000 68.945000  3.045000 69.145000 ;
        RECT  2.845000 69.355000  3.045000 69.555000 ;
        RECT  2.845000 69.765000  3.045000 69.965000 ;
        RECT  2.845000 70.175000  3.045000 70.375000 ;
        RECT  2.845000 70.585000  3.045000 70.785000 ;
        RECT  2.845000 70.995000  3.045000 71.195000 ;
        RECT  2.845000 71.405000  3.045000 71.605000 ;
        RECT  2.845000 71.815000  3.045000 72.015000 ;
        RECT  2.845000 72.225000  3.045000 72.425000 ;
        RECT  2.845000 72.635000  3.045000 72.835000 ;
        RECT  2.845000 73.045000  3.045000 73.245000 ;
        RECT  2.845000 73.450000  3.045000 73.650000 ;
        RECT  2.845000 73.855000  3.045000 74.055000 ;
        RECT  2.845000 74.260000  3.045000 74.460000 ;
        RECT  2.845000 74.665000  3.045000 74.865000 ;
        RECT  2.845000 75.070000  3.045000 75.270000 ;
        RECT  2.845000 75.475000  3.045000 75.675000 ;
        RECT  2.845000 75.880000  3.045000 76.080000 ;
        RECT  2.845000 76.285000  3.045000 76.485000 ;
        RECT  2.845000 76.690000  3.045000 76.890000 ;
        RECT  2.845000 77.095000  3.045000 77.295000 ;
        RECT  2.845000 77.500000  3.045000 77.700000 ;
        RECT  2.845000 77.905000  3.045000 78.105000 ;
        RECT  2.845000 78.310000  3.045000 78.510000 ;
        RECT  2.845000 78.715000  3.045000 78.915000 ;
        RECT  2.845000 79.120000  3.045000 79.320000 ;
        RECT  2.845000 79.525000  3.045000 79.725000 ;
        RECT  2.845000 79.930000  3.045000 80.130000 ;
        RECT  2.845000 80.335000  3.045000 80.535000 ;
        RECT  2.845000 80.740000  3.045000 80.940000 ;
        RECT  2.845000 81.145000  3.045000 81.345000 ;
        RECT  2.845000 81.550000  3.045000 81.750000 ;
        RECT  2.845000 81.955000  3.045000 82.155000 ;
        RECT  2.845000 82.360000  3.045000 82.560000 ;
        RECT  3.120000 17.860000  3.320000 18.060000 ;
        RECT  3.120000 18.290000  3.320000 18.490000 ;
        RECT  3.120000 18.720000  3.320000 18.920000 ;
        RECT  3.120000 19.150000  3.320000 19.350000 ;
        RECT  3.120000 19.580000  3.320000 19.780000 ;
        RECT  3.120000 20.010000  3.320000 20.210000 ;
        RECT  3.120000 20.440000  3.320000 20.640000 ;
        RECT  3.120000 20.870000  3.320000 21.070000 ;
        RECT  3.120000 21.300000  3.320000 21.500000 ;
        RECT  3.120000 21.730000  3.320000 21.930000 ;
        RECT  3.120000 22.160000  3.320000 22.360000 ;
        RECT  3.195000 82.855000  3.395000 83.055000 ;
        RECT  3.195000 83.265000  3.395000 83.465000 ;
        RECT  3.195000 83.675000  3.395000 83.875000 ;
        RECT  3.195000 84.085000  3.395000 84.285000 ;
        RECT  3.195000 84.495000  3.395000 84.695000 ;
        RECT  3.195000 84.905000  3.395000 85.105000 ;
        RECT  3.195000 85.315000  3.395000 85.515000 ;
        RECT  3.195000 85.725000  3.395000 85.925000 ;
        RECT  3.195000 86.135000  3.395000 86.335000 ;
        RECT  3.195000 86.545000  3.395000 86.745000 ;
        RECT  3.195000 86.955000  3.395000 87.155000 ;
        RECT  3.195000 87.365000  3.395000 87.565000 ;
        RECT  3.195000 87.775000  3.395000 87.975000 ;
        RECT  3.195000 88.185000  3.395000 88.385000 ;
        RECT  3.195000 88.595000  3.395000 88.795000 ;
        RECT  3.195000 89.005000  3.395000 89.205000 ;
        RECT  3.195000 89.415000  3.395000 89.615000 ;
        RECT  3.195000 89.825000  3.395000 90.025000 ;
        RECT  3.195000 90.235000  3.395000 90.435000 ;
        RECT  3.195000 90.645000  3.395000 90.845000 ;
        RECT  3.195000 91.055000  3.395000 91.255000 ;
        RECT  3.195000 91.465000  3.395000 91.665000 ;
        RECT  3.195000 91.875000  3.395000 92.075000 ;
        RECT  3.195000 92.285000  3.395000 92.485000 ;
        RECT  3.195000 92.695000  3.395000 92.895000 ;
        RECT  3.245000 68.125000  3.445000 68.325000 ;
        RECT  3.245000 68.535000  3.445000 68.735000 ;
        RECT  3.245000 68.945000  3.445000 69.145000 ;
        RECT  3.245000 69.355000  3.445000 69.555000 ;
        RECT  3.245000 69.765000  3.445000 69.965000 ;
        RECT  3.245000 70.175000  3.445000 70.375000 ;
        RECT  3.245000 70.585000  3.445000 70.785000 ;
        RECT  3.245000 70.995000  3.445000 71.195000 ;
        RECT  3.245000 71.405000  3.445000 71.605000 ;
        RECT  3.245000 71.815000  3.445000 72.015000 ;
        RECT  3.245000 72.225000  3.445000 72.425000 ;
        RECT  3.245000 72.635000  3.445000 72.835000 ;
        RECT  3.245000 73.045000  3.445000 73.245000 ;
        RECT  3.245000 73.450000  3.445000 73.650000 ;
        RECT  3.245000 73.855000  3.445000 74.055000 ;
        RECT  3.245000 74.260000  3.445000 74.460000 ;
        RECT  3.245000 74.665000  3.445000 74.865000 ;
        RECT  3.245000 75.070000  3.445000 75.270000 ;
        RECT  3.245000 75.475000  3.445000 75.675000 ;
        RECT  3.245000 75.880000  3.445000 76.080000 ;
        RECT  3.245000 76.285000  3.445000 76.485000 ;
        RECT  3.245000 76.690000  3.445000 76.890000 ;
        RECT  3.245000 77.095000  3.445000 77.295000 ;
        RECT  3.245000 77.500000  3.445000 77.700000 ;
        RECT  3.245000 77.905000  3.445000 78.105000 ;
        RECT  3.245000 78.310000  3.445000 78.510000 ;
        RECT  3.245000 78.715000  3.445000 78.915000 ;
        RECT  3.245000 79.120000  3.445000 79.320000 ;
        RECT  3.245000 79.525000  3.445000 79.725000 ;
        RECT  3.245000 79.930000  3.445000 80.130000 ;
        RECT  3.245000 80.335000  3.445000 80.535000 ;
        RECT  3.245000 80.740000  3.445000 80.940000 ;
        RECT  3.245000 81.145000  3.445000 81.345000 ;
        RECT  3.245000 81.550000  3.445000 81.750000 ;
        RECT  3.245000 81.955000  3.445000 82.155000 ;
        RECT  3.245000 82.360000  3.445000 82.560000 ;
        RECT  3.525000 17.860000  3.725000 18.060000 ;
        RECT  3.525000 18.290000  3.725000 18.490000 ;
        RECT  3.525000 18.720000  3.725000 18.920000 ;
        RECT  3.525000 19.150000  3.725000 19.350000 ;
        RECT  3.525000 19.580000  3.725000 19.780000 ;
        RECT  3.525000 20.010000  3.725000 20.210000 ;
        RECT  3.525000 20.440000  3.725000 20.640000 ;
        RECT  3.525000 20.870000  3.725000 21.070000 ;
        RECT  3.525000 21.300000  3.725000 21.500000 ;
        RECT  3.525000 21.730000  3.725000 21.930000 ;
        RECT  3.525000 22.160000  3.725000 22.360000 ;
        RECT  3.605000 82.855000  3.805000 83.055000 ;
        RECT  3.605000 83.265000  3.805000 83.465000 ;
        RECT  3.605000 83.675000  3.805000 83.875000 ;
        RECT  3.605000 84.085000  3.805000 84.285000 ;
        RECT  3.605000 84.495000  3.805000 84.695000 ;
        RECT  3.605000 84.905000  3.805000 85.105000 ;
        RECT  3.605000 85.315000  3.805000 85.515000 ;
        RECT  3.605000 85.725000  3.805000 85.925000 ;
        RECT  3.605000 86.135000  3.805000 86.335000 ;
        RECT  3.605000 86.545000  3.805000 86.745000 ;
        RECT  3.605000 86.955000  3.805000 87.155000 ;
        RECT  3.605000 87.365000  3.805000 87.565000 ;
        RECT  3.605000 87.775000  3.805000 87.975000 ;
        RECT  3.605000 88.185000  3.805000 88.385000 ;
        RECT  3.605000 88.595000  3.805000 88.795000 ;
        RECT  3.605000 89.005000  3.805000 89.205000 ;
        RECT  3.605000 89.415000  3.805000 89.615000 ;
        RECT  3.605000 89.825000  3.805000 90.025000 ;
        RECT  3.605000 90.235000  3.805000 90.435000 ;
        RECT  3.605000 90.645000  3.805000 90.845000 ;
        RECT  3.605000 91.055000  3.805000 91.255000 ;
        RECT  3.605000 91.465000  3.805000 91.665000 ;
        RECT  3.605000 91.875000  3.805000 92.075000 ;
        RECT  3.605000 92.285000  3.805000 92.485000 ;
        RECT  3.605000 92.695000  3.805000 92.895000 ;
        RECT  3.645000 68.125000  3.845000 68.325000 ;
        RECT  3.645000 68.535000  3.845000 68.735000 ;
        RECT  3.645000 68.945000  3.845000 69.145000 ;
        RECT  3.645000 69.355000  3.845000 69.555000 ;
        RECT  3.645000 69.765000  3.845000 69.965000 ;
        RECT  3.645000 70.175000  3.845000 70.375000 ;
        RECT  3.645000 70.585000  3.845000 70.785000 ;
        RECT  3.645000 70.995000  3.845000 71.195000 ;
        RECT  3.645000 71.405000  3.845000 71.605000 ;
        RECT  3.645000 71.815000  3.845000 72.015000 ;
        RECT  3.645000 72.225000  3.845000 72.425000 ;
        RECT  3.645000 72.635000  3.845000 72.835000 ;
        RECT  3.645000 73.045000  3.845000 73.245000 ;
        RECT  3.645000 73.450000  3.845000 73.650000 ;
        RECT  3.645000 73.855000  3.845000 74.055000 ;
        RECT  3.645000 74.260000  3.845000 74.460000 ;
        RECT  3.645000 74.665000  3.845000 74.865000 ;
        RECT  3.645000 75.070000  3.845000 75.270000 ;
        RECT  3.645000 75.475000  3.845000 75.675000 ;
        RECT  3.645000 75.880000  3.845000 76.080000 ;
        RECT  3.645000 76.285000  3.845000 76.485000 ;
        RECT  3.645000 76.690000  3.845000 76.890000 ;
        RECT  3.645000 77.095000  3.845000 77.295000 ;
        RECT  3.645000 77.500000  3.845000 77.700000 ;
        RECT  3.645000 77.905000  3.845000 78.105000 ;
        RECT  3.645000 78.310000  3.845000 78.510000 ;
        RECT  3.645000 78.715000  3.845000 78.915000 ;
        RECT  3.645000 79.120000  3.845000 79.320000 ;
        RECT  3.645000 79.525000  3.845000 79.725000 ;
        RECT  3.645000 79.930000  3.845000 80.130000 ;
        RECT  3.645000 80.335000  3.845000 80.535000 ;
        RECT  3.645000 80.740000  3.845000 80.940000 ;
        RECT  3.645000 81.145000  3.845000 81.345000 ;
        RECT  3.645000 81.550000  3.845000 81.750000 ;
        RECT  3.645000 81.955000  3.845000 82.155000 ;
        RECT  3.645000 82.360000  3.845000 82.560000 ;
        RECT  3.930000 17.860000  4.130000 18.060000 ;
        RECT  3.930000 18.290000  4.130000 18.490000 ;
        RECT  3.930000 18.720000  4.130000 18.920000 ;
        RECT  3.930000 19.150000  4.130000 19.350000 ;
        RECT  3.930000 19.580000  4.130000 19.780000 ;
        RECT  3.930000 20.010000  4.130000 20.210000 ;
        RECT  3.930000 20.440000  4.130000 20.640000 ;
        RECT  3.930000 20.870000  4.130000 21.070000 ;
        RECT  3.930000 21.300000  4.130000 21.500000 ;
        RECT  3.930000 21.730000  4.130000 21.930000 ;
        RECT  3.930000 22.160000  4.130000 22.360000 ;
        RECT  4.015000 82.855000  4.215000 83.055000 ;
        RECT  4.015000 83.265000  4.215000 83.465000 ;
        RECT  4.015000 83.675000  4.215000 83.875000 ;
        RECT  4.015000 84.085000  4.215000 84.285000 ;
        RECT  4.015000 84.495000  4.215000 84.695000 ;
        RECT  4.015000 84.905000  4.215000 85.105000 ;
        RECT  4.015000 85.315000  4.215000 85.515000 ;
        RECT  4.015000 85.725000  4.215000 85.925000 ;
        RECT  4.015000 86.135000  4.215000 86.335000 ;
        RECT  4.015000 86.545000  4.215000 86.745000 ;
        RECT  4.015000 86.955000  4.215000 87.155000 ;
        RECT  4.015000 87.365000  4.215000 87.565000 ;
        RECT  4.015000 87.775000  4.215000 87.975000 ;
        RECT  4.015000 88.185000  4.215000 88.385000 ;
        RECT  4.015000 88.595000  4.215000 88.795000 ;
        RECT  4.015000 89.005000  4.215000 89.205000 ;
        RECT  4.015000 89.415000  4.215000 89.615000 ;
        RECT  4.015000 89.825000  4.215000 90.025000 ;
        RECT  4.015000 90.235000  4.215000 90.435000 ;
        RECT  4.015000 90.645000  4.215000 90.845000 ;
        RECT  4.015000 91.055000  4.215000 91.255000 ;
        RECT  4.015000 91.465000  4.215000 91.665000 ;
        RECT  4.015000 91.875000  4.215000 92.075000 ;
        RECT  4.015000 92.285000  4.215000 92.485000 ;
        RECT  4.015000 92.695000  4.215000 92.895000 ;
        RECT  4.045000 68.125000  4.245000 68.325000 ;
        RECT  4.045000 68.535000  4.245000 68.735000 ;
        RECT  4.045000 68.945000  4.245000 69.145000 ;
        RECT  4.045000 69.355000  4.245000 69.555000 ;
        RECT  4.045000 69.765000  4.245000 69.965000 ;
        RECT  4.045000 70.175000  4.245000 70.375000 ;
        RECT  4.045000 70.585000  4.245000 70.785000 ;
        RECT  4.045000 70.995000  4.245000 71.195000 ;
        RECT  4.045000 71.405000  4.245000 71.605000 ;
        RECT  4.045000 71.815000  4.245000 72.015000 ;
        RECT  4.045000 72.225000  4.245000 72.425000 ;
        RECT  4.045000 72.635000  4.245000 72.835000 ;
        RECT  4.045000 73.045000  4.245000 73.245000 ;
        RECT  4.045000 73.450000  4.245000 73.650000 ;
        RECT  4.045000 73.855000  4.245000 74.055000 ;
        RECT  4.045000 74.260000  4.245000 74.460000 ;
        RECT  4.045000 74.665000  4.245000 74.865000 ;
        RECT  4.045000 75.070000  4.245000 75.270000 ;
        RECT  4.045000 75.475000  4.245000 75.675000 ;
        RECT  4.045000 75.880000  4.245000 76.080000 ;
        RECT  4.045000 76.285000  4.245000 76.485000 ;
        RECT  4.045000 76.690000  4.245000 76.890000 ;
        RECT  4.045000 77.095000  4.245000 77.295000 ;
        RECT  4.045000 77.500000  4.245000 77.700000 ;
        RECT  4.045000 77.905000  4.245000 78.105000 ;
        RECT  4.045000 78.310000  4.245000 78.510000 ;
        RECT  4.045000 78.715000  4.245000 78.915000 ;
        RECT  4.045000 79.120000  4.245000 79.320000 ;
        RECT  4.045000 79.525000  4.245000 79.725000 ;
        RECT  4.045000 79.930000  4.245000 80.130000 ;
        RECT  4.045000 80.335000  4.245000 80.535000 ;
        RECT  4.045000 80.740000  4.245000 80.940000 ;
        RECT  4.045000 81.145000  4.245000 81.345000 ;
        RECT  4.045000 81.550000  4.245000 81.750000 ;
        RECT  4.045000 81.955000  4.245000 82.155000 ;
        RECT  4.045000 82.360000  4.245000 82.560000 ;
        RECT  4.335000 17.860000  4.535000 18.060000 ;
        RECT  4.335000 18.290000  4.535000 18.490000 ;
        RECT  4.335000 18.720000  4.535000 18.920000 ;
        RECT  4.335000 19.150000  4.535000 19.350000 ;
        RECT  4.335000 19.580000  4.535000 19.780000 ;
        RECT  4.335000 20.010000  4.535000 20.210000 ;
        RECT  4.335000 20.440000  4.535000 20.640000 ;
        RECT  4.335000 20.870000  4.535000 21.070000 ;
        RECT  4.335000 21.300000  4.535000 21.500000 ;
        RECT  4.335000 21.730000  4.535000 21.930000 ;
        RECT  4.335000 22.160000  4.535000 22.360000 ;
        RECT  4.425000 82.855000  4.625000 83.055000 ;
        RECT  4.425000 83.265000  4.625000 83.465000 ;
        RECT  4.425000 83.675000  4.625000 83.875000 ;
        RECT  4.425000 84.085000  4.625000 84.285000 ;
        RECT  4.425000 84.495000  4.625000 84.695000 ;
        RECT  4.425000 84.905000  4.625000 85.105000 ;
        RECT  4.425000 85.315000  4.625000 85.515000 ;
        RECT  4.425000 85.725000  4.625000 85.925000 ;
        RECT  4.425000 86.135000  4.625000 86.335000 ;
        RECT  4.425000 86.545000  4.625000 86.745000 ;
        RECT  4.425000 86.955000  4.625000 87.155000 ;
        RECT  4.425000 87.365000  4.625000 87.565000 ;
        RECT  4.425000 87.775000  4.625000 87.975000 ;
        RECT  4.425000 88.185000  4.625000 88.385000 ;
        RECT  4.425000 88.595000  4.625000 88.795000 ;
        RECT  4.425000 89.005000  4.625000 89.205000 ;
        RECT  4.425000 89.415000  4.625000 89.615000 ;
        RECT  4.425000 89.825000  4.625000 90.025000 ;
        RECT  4.425000 90.235000  4.625000 90.435000 ;
        RECT  4.425000 90.645000  4.625000 90.845000 ;
        RECT  4.425000 91.055000  4.625000 91.255000 ;
        RECT  4.425000 91.465000  4.625000 91.665000 ;
        RECT  4.425000 91.875000  4.625000 92.075000 ;
        RECT  4.425000 92.285000  4.625000 92.485000 ;
        RECT  4.425000 92.695000  4.625000 92.895000 ;
        RECT  4.445000 68.125000  4.645000 68.325000 ;
        RECT  4.445000 68.535000  4.645000 68.735000 ;
        RECT  4.445000 68.945000  4.645000 69.145000 ;
        RECT  4.445000 69.355000  4.645000 69.555000 ;
        RECT  4.445000 69.765000  4.645000 69.965000 ;
        RECT  4.445000 70.175000  4.645000 70.375000 ;
        RECT  4.445000 70.585000  4.645000 70.785000 ;
        RECT  4.445000 70.995000  4.645000 71.195000 ;
        RECT  4.445000 71.405000  4.645000 71.605000 ;
        RECT  4.445000 71.815000  4.645000 72.015000 ;
        RECT  4.445000 72.225000  4.645000 72.425000 ;
        RECT  4.445000 72.635000  4.645000 72.835000 ;
        RECT  4.445000 73.045000  4.645000 73.245000 ;
        RECT  4.445000 73.450000  4.645000 73.650000 ;
        RECT  4.445000 73.855000  4.645000 74.055000 ;
        RECT  4.445000 74.260000  4.645000 74.460000 ;
        RECT  4.445000 74.665000  4.645000 74.865000 ;
        RECT  4.445000 75.070000  4.645000 75.270000 ;
        RECT  4.445000 75.475000  4.645000 75.675000 ;
        RECT  4.445000 75.880000  4.645000 76.080000 ;
        RECT  4.445000 76.285000  4.645000 76.485000 ;
        RECT  4.445000 76.690000  4.645000 76.890000 ;
        RECT  4.445000 77.095000  4.645000 77.295000 ;
        RECT  4.445000 77.500000  4.645000 77.700000 ;
        RECT  4.445000 77.905000  4.645000 78.105000 ;
        RECT  4.445000 78.310000  4.645000 78.510000 ;
        RECT  4.445000 78.715000  4.645000 78.915000 ;
        RECT  4.445000 79.120000  4.645000 79.320000 ;
        RECT  4.445000 79.525000  4.645000 79.725000 ;
        RECT  4.445000 79.930000  4.645000 80.130000 ;
        RECT  4.445000 80.335000  4.645000 80.535000 ;
        RECT  4.445000 80.740000  4.645000 80.940000 ;
        RECT  4.445000 81.145000  4.645000 81.345000 ;
        RECT  4.445000 81.550000  4.645000 81.750000 ;
        RECT  4.445000 81.955000  4.645000 82.155000 ;
        RECT  4.445000 82.360000  4.645000 82.560000 ;
        RECT  4.740000 17.860000  4.940000 18.060000 ;
        RECT  4.740000 18.290000  4.940000 18.490000 ;
        RECT  4.740000 18.720000  4.940000 18.920000 ;
        RECT  4.740000 19.150000  4.940000 19.350000 ;
        RECT  4.740000 19.580000  4.940000 19.780000 ;
        RECT  4.740000 20.010000  4.940000 20.210000 ;
        RECT  4.740000 20.440000  4.940000 20.640000 ;
        RECT  4.740000 20.870000  4.940000 21.070000 ;
        RECT  4.740000 21.300000  4.940000 21.500000 ;
        RECT  4.740000 21.730000  4.940000 21.930000 ;
        RECT  4.740000 22.160000  4.940000 22.360000 ;
        RECT  4.835000 82.855000  5.035000 83.055000 ;
        RECT  4.835000 83.265000  5.035000 83.465000 ;
        RECT  4.835000 83.675000  5.035000 83.875000 ;
        RECT  4.835000 84.085000  5.035000 84.285000 ;
        RECT  4.835000 84.495000  5.035000 84.695000 ;
        RECT  4.835000 84.905000  5.035000 85.105000 ;
        RECT  4.835000 85.315000  5.035000 85.515000 ;
        RECT  4.835000 85.725000  5.035000 85.925000 ;
        RECT  4.835000 86.135000  5.035000 86.335000 ;
        RECT  4.835000 86.545000  5.035000 86.745000 ;
        RECT  4.835000 86.955000  5.035000 87.155000 ;
        RECT  4.835000 87.365000  5.035000 87.565000 ;
        RECT  4.835000 87.775000  5.035000 87.975000 ;
        RECT  4.835000 88.185000  5.035000 88.385000 ;
        RECT  4.835000 88.595000  5.035000 88.795000 ;
        RECT  4.835000 89.005000  5.035000 89.205000 ;
        RECT  4.835000 89.415000  5.035000 89.615000 ;
        RECT  4.835000 89.825000  5.035000 90.025000 ;
        RECT  4.835000 90.235000  5.035000 90.435000 ;
        RECT  4.835000 90.645000  5.035000 90.845000 ;
        RECT  4.835000 91.055000  5.035000 91.255000 ;
        RECT  4.835000 91.465000  5.035000 91.665000 ;
        RECT  4.835000 91.875000  5.035000 92.075000 ;
        RECT  4.835000 92.285000  5.035000 92.485000 ;
        RECT  4.835000 92.695000  5.035000 92.895000 ;
        RECT  4.845000 68.125000  5.045000 68.325000 ;
        RECT  4.845000 68.535000  5.045000 68.735000 ;
        RECT  4.845000 68.945000  5.045000 69.145000 ;
        RECT  4.845000 69.355000  5.045000 69.555000 ;
        RECT  4.845000 69.765000  5.045000 69.965000 ;
        RECT  4.845000 70.175000  5.045000 70.375000 ;
        RECT  4.845000 70.585000  5.045000 70.785000 ;
        RECT  4.845000 70.995000  5.045000 71.195000 ;
        RECT  4.845000 71.405000  5.045000 71.605000 ;
        RECT  4.845000 71.815000  5.045000 72.015000 ;
        RECT  4.845000 72.225000  5.045000 72.425000 ;
        RECT  4.845000 72.635000  5.045000 72.835000 ;
        RECT  4.845000 73.045000  5.045000 73.245000 ;
        RECT  4.845000 73.450000  5.045000 73.650000 ;
        RECT  4.845000 73.855000  5.045000 74.055000 ;
        RECT  4.845000 74.260000  5.045000 74.460000 ;
        RECT  4.845000 74.665000  5.045000 74.865000 ;
        RECT  4.845000 75.070000  5.045000 75.270000 ;
        RECT  4.845000 75.475000  5.045000 75.675000 ;
        RECT  4.845000 75.880000  5.045000 76.080000 ;
        RECT  4.845000 76.285000  5.045000 76.485000 ;
        RECT  4.845000 76.690000  5.045000 76.890000 ;
        RECT  4.845000 77.095000  5.045000 77.295000 ;
        RECT  4.845000 77.500000  5.045000 77.700000 ;
        RECT  4.845000 77.905000  5.045000 78.105000 ;
        RECT  4.845000 78.310000  5.045000 78.510000 ;
        RECT  4.845000 78.715000  5.045000 78.915000 ;
        RECT  4.845000 79.120000  5.045000 79.320000 ;
        RECT  4.845000 79.525000  5.045000 79.725000 ;
        RECT  4.845000 79.930000  5.045000 80.130000 ;
        RECT  4.845000 80.335000  5.045000 80.535000 ;
        RECT  4.845000 80.740000  5.045000 80.940000 ;
        RECT  4.845000 81.145000  5.045000 81.345000 ;
        RECT  4.845000 81.550000  5.045000 81.750000 ;
        RECT  4.845000 81.955000  5.045000 82.155000 ;
        RECT  4.845000 82.360000  5.045000 82.560000 ;
        RECT  5.145000 17.860000  5.345000 18.060000 ;
        RECT  5.145000 18.290000  5.345000 18.490000 ;
        RECT  5.145000 18.720000  5.345000 18.920000 ;
        RECT  5.145000 19.150000  5.345000 19.350000 ;
        RECT  5.145000 19.580000  5.345000 19.780000 ;
        RECT  5.145000 20.010000  5.345000 20.210000 ;
        RECT  5.145000 20.440000  5.345000 20.640000 ;
        RECT  5.145000 20.870000  5.345000 21.070000 ;
        RECT  5.145000 21.300000  5.345000 21.500000 ;
        RECT  5.145000 21.730000  5.345000 21.930000 ;
        RECT  5.145000 22.160000  5.345000 22.360000 ;
        RECT  5.245000 68.125000  5.445000 68.325000 ;
        RECT  5.245000 68.535000  5.445000 68.735000 ;
        RECT  5.245000 68.945000  5.445000 69.145000 ;
        RECT  5.245000 69.355000  5.445000 69.555000 ;
        RECT  5.245000 69.765000  5.445000 69.965000 ;
        RECT  5.245000 70.175000  5.445000 70.375000 ;
        RECT  5.245000 70.585000  5.445000 70.785000 ;
        RECT  5.245000 70.995000  5.445000 71.195000 ;
        RECT  5.245000 71.405000  5.445000 71.605000 ;
        RECT  5.245000 71.815000  5.445000 72.015000 ;
        RECT  5.245000 72.225000  5.445000 72.425000 ;
        RECT  5.245000 72.635000  5.445000 72.835000 ;
        RECT  5.245000 73.045000  5.445000 73.245000 ;
        RECT  5.245000 73.450000  5.445000 73.650000 ;
        RECT  5.245000 73.855000  5.445000 74.055000 ;
        RECT  5.245000 74.260000  5.445000 74.460000 ;
        RECT  5.245000 74.665000  5.445000 74.865000 ;
        RECT  5.245000 75.070000  5.445000 75.270000 ;
        RECT  5.245000 75.475000  5.445000 75.675000 ;
        RECT  5.245000 75.880000  5.445000 76.080000 ;
        RECT  5.245000 76.285000  5.445000 76.485000 ;
        RECT  5.245000 76.690000  5.445000 76.890000 ;
        RECT  5.245000 77.095000  5.445000 77.295000 ;
        RECT  5.245000 77.500000  5.445000 77.700000 ;
        RECT  5.245000 77.905000  5.445000 78.105000 ;
        RECT  5.245000 78.310000  5.445000 78.510000 ;
        RECT  5.245000 78.715000  5.445000 78.915000 ;
        RECT  5.245000 79.120000  5.445000 79.320000 ;
        RECT  5.245000 79.525000  5.445000 79.725000 ;
        RECT  5.245000 79.930000  5.445000 80.130000 ;
        RECT  5.245000 80.335000  5.445000 80.535000 ;
        RECT  5.245000 80.740000  5.445000 80.940000 ;
        RECT  5.245000 81.145000  5.445000 81.345000 ;
        RECT  5.245000 81.550000  5.445000 81.750000 ;
        RECT  5.245000 81.955000  5.445000 82.155000 ;
        RECT  5.245000 82.360000  5.445000 82.560000 ;
        RECT  5.245000 82.855000  5.445000 83.055000 ;
        RECT  5.245000 83.265000  5.445000 83.465000 ;
        RECT  5.245000 83.675000  5.445000 83.875000 ;
        RECT  5.245000 84.085000  5.445000 84.285000 ;
        RECT  5.245000 84.495000  5.445000 84.695000 ;
        RECT  5.245000 84.905000  5.445000 85.105000 ;
        RECT  5.245000 85.315000  5.445000 85.515000 ;
        RECT  5.245000 85.725000  5.445000 85.925000 ;
        RECT  5.245000 86.135000  5.445000 86.335000 ;
        RECT  5.245000 86.545000  5.445000 86.745000 ;
        RECT  5.245000 86.955000  5.445000 87.155000 ;
        RECT  5.245000 87.365000  5.445000 87.565000 ;
        RECT  5.245000 87.775000  5.445000 87.975000 ;
        RECT  5.245000 88.185000  5.445000 88.385000 ;
        RECT  5.245000 88.595000  5.445000 88.795000 ;
        RECT  5.245000 89.005000  5.445000 89.205000 ;
        RECT  5.245000 89.415000  5.445000 89.615000 ;
        RECT  5.245000 89.825000  5.445000 90.025000 ;
        RECT  5.245000 90.235000  5.445000 90.435000 ;
        RECT  5.245000 90.645000  5.445000 90.845000 ;
        RECT  5.245000 91.055000  5.445000 91.255000 ;
        RECT  5.245000 91.465000  5.445000 91.665000 ;
        RECT  5.245000 91.875000  5.445000 92.075000 ;
        RECT  5.245000 92.285000  5.445000 92.485000 ;
        RECT  5.245000 92.695000  5.445000 92.895000 ;
        RECT  5.550000 17.860000  5.750000 18.060000 ;
        RECT  5.550000 18.290000  5.750000 18.490000 ;
        RECT  5.550000 18.720000  5.750000 18.920000 ;
        RECT  5.550000 19.150000  5.750000 19.350000 ;
        RECT  5.550000 19.580000  5.750000 19.780000 ;
        RECT  5.550000 20.010000  5.750000 20.210000 ;
        RECT  5.550000 20.440000  5.750000 20.640000 ;
        RECT  5.550000 20.870000  5.750000 21.070000 ;
        RECT  5.550000 21.300000  5.750000 21.500000 ;
        RECT  5.550000 21.730000  5.750000 21.930000 ;
        RECT  5.550000 22.160000  5.750000 22.360000 ;
        RECT  5.645000 68.125000  5.845000 68.325000 ;
        RECT  5.645000 68.535000  5.845000 68.735000 ;
        RECT  5.645000 68.945000  5.845000 69.145000 ;
        RECT  5.645000 69.355000  5.845000 69.555000 ;
        RECT  5.645000 69.765000  5.845000 69.965000 ;
        RECT  5.645000 70.175000  5.845000 70.375000 ;
        RECT  5.645000 70.585000  5.845000 70.785000 ;
        RECT  5.645000 70.995000  5.845000 71.195000 ;
        RECT  5.645000 71.405000  5.845000 71.605000 ;
        RECT  5.645000 71.815000  5.845000 72.015000 ;
        RECT  5.645000 72.225000  5.845000 72.425000 ;
        RECT  5.645000 72.635000  5.845000 72.835000 ;
        RECT  5.645000 73.045000  5.845000 73.245000 ;
        RECT  5.645000 73.450000  5.845000 73.650000 ;
        RECT  5.645000 73.855000  5.845000 74.055000 ;
        RECT  5.645000 74.260000  5.845000 74.460000 ;
        RECT  5.645000 74.665000  5.845000 74.865000 ;
        RECT  5.645000 75.070000  5.845000 75.270000 ;
        RECT  5.645000 75.475000  5.845000 75.675000 ;
        RECT  5.645000 75.880000  5.845000 76.080000 ;
        RECT  5.645000 76.285000  5.845000 76.485000 ;
        RECT  5.645000 76.690000  5.845000 76.890000 ;
        RECT  5.645000 77.095000  5.845000 77.295000 ;
        RECT  5.645000 77.500000  5.845000 77.700000 ;
        RECT  5.645000 77.905000  5.845000 78.105000 ;
        RECT  5.645000 78.310000  5.845000 78.510000 ;
        RECT  5.645000 78.715000  5.845000 78.915000 ;
        RECT  5.645000 79.120000  5.845000 79.320000 ;
        RECT  5.645000 79.525000  5.845000 79.725000 ;
        RECT  5.645000 79.930000  5.845000 80.130000 ;
        RECT  5.645000 80.335000  5.845000 80.535000 ;
        RECT  5.645000 80.740000  5.845000 80.940000 ;
        RECT  5.645000 81.145000  5.845000 81.345000 ;
        RECT  5.645000 81.550000  5.845000 81.750000 ;
        RECT  5.645000 81.955000  5.845000 82.155000 ;
        RECT  5.645000 82.360000  5.845000 82.560000 ;
        RECT  5.655000 82.855000  5.855000 83.055000 ;
        RECT  5.655000 83.265000  5.855000 83.465000 ;
        RECT  5.655000 83.675000  5.855000 83.875000 ;
        RECT  5.655000 84.085000  5.855000 84.285000 ;
        RECT  5.655000 84.495000  5.855000 84.695000 ;
        RECT  5.655000 84.905000  5.855000 85.105000 ;
        RECT  5.655000 85.315000  5.855000 85.515000 ;
        RECT  5.655000 85.725000  5.855000 85.925000 ;
        RECT  5.655000 86.135000  5.855000 86.335000 ;
        RECT  5.655000 86.545000  5.855000 86.745000 ;
        RECT  5.655000 86.955000  5.855000 87.155000 ;
        RECT  5.655000 87.365000  5.855000 87.565000 ;
        RECT  5.655000 87.775000  5.855000 87.975000 ;
        RECT  5.655000 88.185000  5.855000 88.385000 ;
        RECT  5.655000 88.595000  5.855000 88.795000 ;
        RECT  5.655000 89.005000  5.855000 89.205000 ;
        RECT  5.655000 89.415000  5.855000 89.615000 ;
        RECT  5.655000 89.825000  5.855000 90.025000 ;
        RECT  5.655000 90.235000  5.855000 90.435000 ;
        RECT  5.655000 90.645000  5.855000 90.845000 ;
        RECT  5.655000 91.055000  5.855000 91.255000 ;
        RECT  5.655000 91.465000  5.855000 91.665000 ;
        RECT  5.655000 91.875000  5.855000 92.075000 ;
        RECT  5.655000 92.285000  5.855000 92.485000 ;
        RECT  5.655000 92.695000  5.855000 92.895000 ;
        RECT  5.955000 17.860000  6.155000 18.060000 ;
        RECT  5.955000 18.290000  6.155000 18.490000 ;
        RECT  5.955000 18.720000  6.155000 18.920000 ;
        RECT  5.955000 19.150000  6.155000 19.350000 ;
        RECT  5.955000 19.580000  6.155000 19.780000 ;
        RECT  5.955000 20.010000  6.155000 20.210000 ;
        RECT  5.955000 20.440000  6.155000 20.640000 ;
        RECT  5.955000 20.870000  6.155000 21.070000 ;
        RECT  5.955000 21.300000  6.155000 21.500000 ;
        RECT  5.955000 21.730000  6.155000 21.930000 ;
        RECT  5.955000 22.160000  6.155000 22.360000 ;
        RECT  6.045000 68.125000  6.245000 68.325000 ;
        RECT  6.045000 68.535000  6.245000 68.735000 ;
        RECT  6.045000 68.945000  6.245000 69.145000 ;
        RECT  6.045000 69.355000  6.245000 69.555000 ;
        RECT  6.045000 69.765000  6.245000 69.965000 ;
        RECT  6.045000 70.175000  6.245000 70.375000 ;
        RECT  6.045000 70.585000  6.245000 70.785000 ;
        RECT  6.045000 70.995000  6.245000 71.195000 ;
        RECT  6.045000 71.405000  6.245000 71.605000 ;
        RECT  6.045000 71.815000  6.245000 72.015000 ;
        RECT  6.045000 72.225000  6.245000 72.425000 ;
        RECT  6.045000 72.635000  6.245000 72.835000 ;
        RECT  6.045000 73.045000  6.245000 73.245000 ;
        RECT  6.045000 73.450000  6.245000 73.650000 ;
        RECT  6.045000 73.855000  6.245000 74.055000 ;
        RECT  6.045000 74.260000  6.245000 74.460000 ;
        RECT  6.045000 74.665000  6.245000 74.865000 ;
        RECT  6.045000 75.070000  6.245000 75.270000 ;
        RECT  6.045000 75.475000  6.245000 75.675000 ;
        RECT  6.045000 75.880000  6.245000 76.080000 ;
        RECT  6.045000 76.285000  6.245000 76.485000 ;
        RECT  6.045000 76.690000  6.245000 76.890000 ;
        RECT  6.045000 77.095000  6.245000 77.295000 ;
        RECT  6.045000 77.500000  6.245000 77.700000 ;
        RECT  6.045000 77.905000  6.245000 78.105000 ;
        RECT  6.045000 78.310000  6.245000 78.510000 ;
        RECT  6.045000 78.715000  6.245000 78.915000 ;
        RECT  6.045000 79.120000  6.245000 79.320000 ;
        RECT  6.045000 79.525000  6.245000 79.725000 ;
        RECT  6.045000 79.930000  6.245000 80.130000 ;
        RECT  6.045000 80.335000  6.245000 80.535000 ;
        RECT  6.045000 80.740000  6.245000 80.940000 ;
        RECT  6.045000 81.145000  6.245000 81.345000 ;
        RECT  6.045000 81.550000  6.245000 81.750000 ;
        RECT  6.045000 81.955000  6.245000 82.155000 ;
        RECT  6.045000 82.360000  6.245000 82.560000 ;
        RECT  6.065000 82.855000  6.265000 83.055000 ;
        RECT  6.065000 83.265000  6.265000 83.465000 ;
        RECT  6.065000 83.675000  6.265000 83.875000 ;
        RECT  6.065000 84.085000  6.265000 84.285000 ;
        RECT  6.065000 84.495000  6.265000 84.695000 ;
        RECT  6.065000 84.905000  6.265000 85.105000 ;
        RECT  6.065000 85.315000  6.265000 85.515000 ;
        RECT  6.065000 85.725000  6.265000 85.925000 ;
        RECT  6.065000 86.135000  6.265000 86.335000 ;
        RECT  6.065000 86.545000  6.265000 86.745000 ;
        RECT  6.065000 86.955000  6.265000 87.155000 ;
        RECT  6.065000 87.365000  6.265000 87.565000 ;
        RECT  6.065000 87.775000  6.265000 87.975000 ;
        RECT  6.065000 88.185000  6.265000 88.385000 ;
        RECT  6.065000 88.595000  6.265000 88.795000 ;
        RECT  6.065000 89.005000  6.265000 89.205000 ;
        RECT  6.065000 89.415000  6.265000 89.615000 ;
        RECT  6.065000 89.825000  6.265000 90.025000 ;
        RECT  6.065000 90.235000  6.265000 90.435000 ;
        RECT  6.065000 90.645000  6.265000 90.845000 ;
        RECT  6.065000 91.055000  6.265000 91.255000 ;
        RECT  6.065000 91.465000  6.265000 91.665000 ;
        RECT  6.065000 91.875000  6.265000 92.075000 ;
        RECT  6.065000 92.285000  6.265000 92.485000 ;
        RECT  6.065000 92.695000  6.265000 92.895000 ;
        RECT  6.360000 17.860000  6.560000 18.060000 ;
        RECT  6.360000 18.290000  6.560000 18.490000 ;
        RECT  6.360000 18.720000  6.560000 18.920000 ;
        RECT  6.360000 19.150000  6.560000 19.350000 ;
        RECT  6.360000 19.580000  6.560000 19.780000 ;
        RECT  6.360000 20.010000  6.560000 20.210000 ;
        RECT  6.360000 20.440000  6.560000 20.640000 ;
        RECT  6.360000 20.870000  6.560000 21.070000 ;
        RECT  6.360000 21.300000  6.560000 21.500000 ;
        RECT  6.360000 21.730000  6.560000 21.930000 ;
        RECT  6.360000 22.160000  6.560000 22.360000 ;
        RECT  6.445000 68.125000  6.645000 68.325000 ;
        RECT  6.445000 68.535000  6.645000 68.735000 ;
        RECT  6.445000 68.945000  6.645000 69.145000 ;
        RECT  6.445000 69.355000  6.645000 69.555000 ;
        RECT  6.445000 69.765000  6.645000 69.965000 ;
        RECT  6.445000 70.175000  6.645000 70.375000 ;
        RECT  6.445000 70.585000  6.645000 70.785000 ;
        RECT  6.445000 70.995000  6.645000 71.195000 ;
        RECT  6.445000 71.405000  6.645000 71.605000 ;
        RECT  6.445000 71.815000  6.645000 72.015000 ;
        RECT  6.445000 72.225000  6.645000 72.425000 ;
        RECT  6.445000 72.635000  6.645000 72.835000 ;
        RECT  6.445000 73.045000  6.645000 73.245000 ;
        RECT  6.445000 73.450000  6.645000 73.650000 ;
        RECT  6.445000 73.855000  6.645000 74.055000 ;
        RECT  6.445000 74.260000  6.645000 74.460000 ;
        RECT  6.445000 74.665000  6.645000 74.865000 ;
        RECT  6.445000 75.070000  6.645000 75.270000 ;
        RECT  6.445000 75.475000  6.645000 75.675000 ;
        RECT  6.445000 75.880000  6.645000 76.080000 ;
        RECT  6.445000 76.285000  6.645000 76.485000 ;
        RECT  6.445000 76.690000  6.645000 76.890000 ;
        RECT  6.445000 77.095000  6.645000 77.295000 ;
        RECT  6.445000 77.500000  6.645000 77.700000 ;
        RECT  6.445000 77.905000  6.645000 78.105000 ;
        RECT  6.445000 78.310000  6.645000 78.510000 ;
        RECT  6.445000 78.715000  6.645000 78.915000 ;
        RECT  6.445000 79.120000  6.645000 79.320000 ;
        RECT  6.445000 79.525000  6.645000 79.725000 ;
        RECT  6.445000 79.930000  6.645000 80.130000 ;
        RECT  6.445000 80.335000  6.645000 80.535000 ;
        RECT  6.445000 80.740000  6.645000 80.940000 ;
        RECT  6.445000 81.145000  6.645000 81.345000 ;
        RECT  6.445000 81.550000  6.645000 81.750000 ;
        RECT  6.445000 81.955000  6.645000 82.155000 ;
        RECT  6.445000 82.360000  6.645000 82.560000 ;
        RECT  6.475000 82.855000  6.675000 83.055000 ;
        RECT  6.475000 83.265000  6.675000 83.465000 ;
        RECT  6.475000 83.675000  6.675000 83.875000 ;
        RECT  6.475000 84.085000  6.675000 84.285000 ;
        RECT  6.475000 84.495000  6.675000 84.695000 ;
        RECT  6.475000 84.905000  6.675000 85.105000 ;
        RECT  6.475000 85.315000  6.675000 85.515000 ;
        RECT  6.475000 85.725000  6.675000 85.925000 ;
        RECT  6.475000 86.135000  6.675000 86.335000 ;
        RECT  6.475000 86.545000  6.675000 86.745000 ;
        RECT  6.475000 86.955000  6.675000 87.155000 ;
        RECT  6.475000 87.365000  6.675000 87.565000 ;
        RECT  6.475000 87.775000  6.675000 87.975000 ;
        RECT  6.475000 88.185000  6.675000 88.385000 ;
        RECT  6.475000 88.595000  6.675000 88.795000 ;
        RECT  6.475000 89.005000  6.675000 89.205000 ;
        RECT  6.475000 89.415000  6.675000 89.615000 ;
        RECT  6.475000 89.825000  6.675000 90.025000 ;
        RECT  6.475000 90.235000  6.675000 90.435000 ;
        RECT  6.475000 90.645000  6.675000 90.845000 ;
        RECT  6.475000 91.055000  6.675000 91.255000 ;
        RECT  6.475000 91.465000  6.675000 91.665000 ;
        RECT  6.475000 91.875000  6.675000 92.075000 ;
        RECT  6.475000 92.285000  6.675000 92.485000 ;
        RECT  6.475000 92.695000  6.675000 92.895000 ;
        RECT  6.765000 17.860000  6.965000 18.060000 ;
        RECT  6.765000 18.290000  6.965000 18.490000 ;
        RECT  6.765000 18.720000  6.965000 18.920000 ;
        RECT  6.765000 19.150000  6.965000 19.350000 ;
        RECT  6.765000 19.580000  6.965000 19.780000 ;
        RECT  6.765000 20.010000  6.965000 20.210000 ;
        RECT  6.765000 20.440000  6.965000 20.640000 ;
        RECT  6.765000 20.870000  6.965000 21.070000 ;
        RECT  6.765000 21.300000  6.965000 21.500000 ;
        RECT  6.765000 21.730000  6.965000 21.930000 ;
        RECT  6.765000 22.160000  6.965000 22.360000 ;
        RECT  6.845000 68.125000  7.045000 68.325000 ;
        RECT  6.845000 68.535000  7.045000 68.735000 ;
        RECT  6.845000 68.945000  7.045000 69.145000 ;
        RECT  6.845000 69.355000  7.045000 69.555000 ;
        RECT  6.845000 69.765000  7.045000 69.965000 ;
        RECT  6.845000 70.175000  7.045000 70.375000 ;
        RECT  6.845000 70.585000  7.045000 70.785000 ;
        RECT  6.845000 70.995000  7.045000 71.195000 ;
        RECT  6.845000 71.405000  7.045000 71.605000 ;
        RECT  6.845000 71.815000  7.045000 72.015000 ;
        RECT  6.845000 72.225000  7.045000 72.425000 ;
        RECT  6.845000 72.635000  7.045000 72.835000 ;
        RECT  6.845000 73.045000  7.045000 73.245000 ;
        RECT  6.845000 73.450000  7.045000 73.650000 ;
        RECT  6.845000 73.855000  7.045000 74.055000 ;
        RECT  6.845000 74.260000  7.045000 74.460000 ;
        RECT  6.845000 74.665000  7.045000 74.865000 ;
        RECT  6.845000 75.070000  7.045000 75.270000 ;
        RECT  6.845000 75.475000  7.045000 75.675000 ;
        RECT  6.845000 75.880000  7.045000 76.080000 ;
        RECT  6.845000 76.285000  7.045000 76.485000 ;
        RECT  6.845000 76.690000  7.045000 76.890000 ;
        RECT  6.845000 77.095000  7.045000 77.295000 ;
        RECT  6.845000 77.500000  7.045000 77.700000 ;
        RECT  6.845000 77.905000  7.045000 78.105000 ;
        RECT  6.845000 78.310000  7.045000 78.510000 ;
        RECT  6.845000 78.715000  7.045000 78.915000 ;
        RECT  6.845000 79.120000  7.045000 79.320000 ;
        RECT  6.845000 79.525000  7.045000 79.725000 ;
        RECT  6.845000 79.930000  7.045000 80.130000 ;
        RECT  6.845000 80.335000  7.045000 80.535000 ;
        RECT  6.845000 80.740000  7.045000 80.940000 ;
        RECT  6.845000 81.145000  7.045000 81.345000 ;
        RECT  6.845000 81.550000  7.045000 81.750000 ;
        RECT  6.845000 81.955000  7.045000 82.155000 ;
        RECT  6.845000 82.360000  7.045000 82.560000 ;
        RECT  6.885000 82.855000  7.085000 83.055000 ;
        RECT  6.885000 83.265000  7.085000 83.465000 ;
        RECT  6.885000 83.675000  7.085000 83.875000 ;
        RECT  6.885000 84.085000  7.085000 84.285000 ;
        RECT  6.885000 84.495000  7.085000 84.695000 ;
        RECT  6.885000 84.905000  7.085000 85.105000 ;
        RECT  6.885000 85.315000  7.085000 85.515000 ;
        RECT  6.885000 85.725000  7.085000 85.925000 ;
        RECT  6.885000 86.135000  7.085000 86.335000 ;
        RECT  6.885000 86.545000  7.085000 86.745000 ;
        RECT  6.885000 86.955000  7.085000 87.155000 ;
        RECT  6.885000 87.365000  7.085000 87.565000 ;
        RECT  6.885000 87.775000  7.085000 87.975000 ;
        RECT  6.885000 88.185000  7.085000 88.385000 ;
        RECT  6.885000 88.595000  7.085000 88.795000 ;
        RECT  6.885000 89.005000  7.085000 89.205000 ;
        RECT  6.885000 89.415000  7.085000 89.615000 ;
        RECT  6.885000 89.825000  7.085000 90.025000 ;
        RECT  6.885000 90.235000  7.085000 90.435000 ;
        RECT  6.885000 90.645000  7.085000 90.845000 ;
        RECT  6.885000 91.055000  7.085000 91.255000 ;
        RECT  6.885000 91.465000  7.085000 91.665000 ;
        RECT  6.885000 91.875000  7.085000 92.075000 ;
        RECT  6.885000 92.285000  7.085000 92.485000 ;
        RECT  6.885000 92.695000  7.085000 92.895000 ;
        RECT  7.170000 17.860000  7.370000 18.060000 ;
        RECT  7.170000 18.290000  7.370000 18.490000 ;
        RECT  7.170000 18.720000  7.370000 18.920000 ;
        RECT  7.170000 19.150000  7.370000 19.350000 ;
        RECT  7.170000 19.580000  7.370000 19.780000 ;
        RECT  7.170000 20.010000  7.370000 20.210000 ;
        RECT  7.170000 20.440000  7.370000 20.640000 ;
        RECT  7.170000 20.870000  7.370000 21.070000 ;
        RECT  7.170000 21.300000  7.370000 21.500000 ;
        RECT  7.170000 21.730000  7.370000 21.930000 ;
        RECT  7.170000 22.160000  7.370000 22.360000 ;
        RECT  7.245000 68.125000  7.445000 68.325000 ;
        RECT  7.245000 68.535000  7.445000 68.735000 ;
        RECT  7.245000 68.945000  7.445000 69.145000 ;
        RECT  7.245000 69.355000  7.445000 69.555000 ;
        RECT  7.245000 69.765000  7.445000 69.965000 ;
        RECT  7.245000 70.175000  7.445000 70.375000 ;
        RECT  7.245000 70.585000  7.445000 70.785000 ;
        RECT  7.245000 70.995000  7.445000 71.195000 ;
        RECT  7.245000 71.405000  7.445000 71.605000 ;
        RECT  7.245000 71.815000  7.445000 72.015000 ;
        RECT  7.245000 72.225000  7.445000 72.425000 ;
        RECT  7.245000 72.635000  7.445000 72.835000 ;
        RECT  7.245000 73.045000  7.445000 73.245000 ;
        RECT  7.245000 73.450000  7.445000 73.650000 ;
        RECT  7.245000 73.855000  7.445000 74.055000 ;
        RECT  7.245000 74.260000  7.445000 74.460000 ;
        RECT  7.245000 74.665000  7.445000 74.865000 ;
        RECT  7.245000 75.070000  7.445000 75.270000 ;
        RECT  7.245000 75.475000  7.445000 75.675000 ;
        RECT  7.245000 75.880000  7.445000 76.080000 ;
        RECT  7.245000 76.285000  7.445000 76.485000 ;
        RECT  7.245000 76.690000  7.445000 76.890000 ;
        RECT  7.245000 77.095000  7.445000 77.295000 ;
        RECT  7.245000 77.500000  7.445000 77.700000 ;
        RECT  7.245000 77.905000  7.445000 78.105000 ;
        RECT  7.245000 78.310000  7.445000 78.510000 ;
        RECT  7.245000 78.715000  7.445000 78.915000 ;
        RECT  7.245000 79.120000  7.445000 79.320000 ;
        RECT  7.245000 79.525000  7.445000 79.725000 ;
        RECT  7.245000 79.930000  7.445000 80.130000 ;
        RECT  7.245000 80.335000  7.445000 80.535000 ;
        RECT  7.245000 80.740000  7.445000 80.940000 ;
        RECT  7.245000 81.145000  7.445000 81.345000 ;
        RECT  7.245000 81.550000  7.445000 81.750000 ;
        RECT  7.245000 81.955000  7.445000 82.155000 ;
        RECT  7.245000 82.360000  7.445000 82.560000 ;
        RECT  7.295000 82.855000  7.495000 83.055000 ;
        RECT  7.295000 83.265000  7.495000 83.465000 ;
        RECT  7.295000 83.675000  7.495000 83.875000 ;
        RECT  7.295000 84.085000  7.495000 84.285000 ;
        RECT  7.295000 84.495000  7.495000 84.695000 ;
        RECT  7.295000 84.905000  7.495000 85.105000 ;
        RECT  7.295000 85.315000  7.495000 85.515000 ;
        RECT  7.295000 85.725000  7.495000 85.925000 ;
        RECT  7.295000 86.135000  7.495000 86.335000 ;
        RECT  7.295000 86.545000  7.495000 86.745000 ;
        RECT  7.295000 86.955000  7.495000 87.155000 ;
        RECT  7.295000 87.365000  7.495000 87.565000 ;
        RECT  7.295000 87.775000  7.495000 87.975000 ;
        RECT  7.295000 88.185000  7.495000 88.385000 ;
        RECT  7.295000 88.595000  7.495000 88.795000 ;
        RECT  7.295000 89.005000  7.495000 89.205000 ;
        RECT  7.295000 89.415000  7.495000 89.615000 ;
        RECT  7.295000 89.825000  7.495000 90.025000 ;
        RECT  7.295000 90.235000  7.495000 90.435000 ;
        RECT  7.295000 90.645000  7.495000 90.845000 ;
        RECT  7.295000 91.055000  7.495000 91.255000 ;
        RECT  7.295000 91.465000  7.495000 91.665000 ;
        RECT  7.295000 91.875000  7.495000 92.075000 ;
        RECT  7.295000 92.285000  7.495000 92.485000 ;
        RECT  7.295000 92.695000  7.495000 92.895000 ;
        RECT  7.575000 17.860000  7.775000 18.060000 ;
        RECT  7.575000 18.290000  7.775000 18.490000 ;
        RECT  7.575000 18.720000  7.775000 18.920000 ;
        RECT  7.575000 19.150000  7.775000 19.350000 ;
        RECT  7.575000 19.580000  7.775000 19.780000 ;
        RECT  7.575000 20.010000  7.775000 20.210000 ;
        RECT  7.575000 20.440000  7.775000 20.640000 ;
        RECT  7.575000 20.870000  7.775000 21.070000 ;
        RECT  7.575000 21.300000  7.775000 21.500000 ;
        RECT  7.575000 21.730000  7.775000 21.930000 ;
        RECT  7.575000 22.160000  7.775000 22.360000 ;
        RECT  7.645000 68.125000  7.845000 68.325000 ;
        RECT  7.645000 68.535000  7.845000 68.735000 ;
        RECT  7.645000 68.945000  7.845000 69.145000 ;
        RECT  7.645000 69.355000  7.845000 69.555000 ;
        RECT  7.645000 69.765000  7.845000 69.965000 ;
        RECT  7.645000 70.175000  7.845000 70.375000 ;
        RECT  7.645000 70.585000  7.845000 70.785000 ;
        RECT  7.645000 70.995000  7.845000 71.195000 ;
        RECT  7.645000 71.405000  7.845000 71.605000 ;
        RECT  7.645000 71.815000  7.845000 72.015000 ;
        RECT  7.645000 72.225000  7.845000 72.425000 ;
        RECT  7.645000 72.635000  7.845000 72.835000 ;
        RECT  7.645000 73.045000  7.845000 73.245000 ;
        RECT  7.645000 73.450000  7.845000 73.650000 ;
        RECT  7.645000 73.855000  7.845000 74.055000 ;
        RECT  7.645000 74.260000  7.845000 74.460000 ;
        RECT  7.645000 74.665000  7.845000 74.865000 ;
        RECT  7.645000 75.070000  7.845000 75.270000 ;
        RECT  7.645000 75.475000  7.845000 75.675000 ;
        RECT  7.645000 75.880000  7.845000 76.080000 ;
        RECT  7.645000 76.285000  7.845000 76.485000 ;
        RECT  7.645000 76.690000  7.845000 76.890000 ;
        RECT  7.645000 77.095000  7.845000 77.295000 ;
        RECT  7.645000 77.500000  7.845000 77.700000 ;
        RECT  7.645000 77.905000  7.845000 78.105000 ;
        RECT  7.645000 78.310000  7.845000 78.510000 ;
        RECT  7.645000 78.715000  7.845000 78.915000 ;
        RECT  7.645000 79.120000  7.845000 79.320000 ;
        RECT  7.645000 79.525000  7.845000 79.725000 ;
        RECT  7.645000 79.930000  7.845000 80.130000 ;
        RECT  7.645000 80.335000  7.845000 80.535000 ;
        RECT  7.645000 80.740000  7.845000 80.940000 ;
        RECT  7.645000 81.145000  7.845000 81.345000 ;
        RECT  7.645000 81.550000  7.845000 81.750000 ;
        RECT  7.645000 81.955000  7.845000 82.155000 ;
        RECT  7.645000 82.360000  7.845000 82.560000 ;
        RECT  7.705000 82.855000  7.905000 83.055000 ;
        RECT  7.705000 83.265000  7.905000 83.465000 ;
        RECT  7.705000 83.675000  7.905000 83.875000 ;
        RECT  7.705000 84.085000  7.905000 84.285000 ;
        RECT  7.705000 84.495000  7.905000 84.695000 ;
        RECT  7.705000 84.905000  7.905000 85.105000 ;
        RECT  7.705000 85.315000  7.905000 85.515000 ;
        RECT  7.705000 85.725000  7.905000 85.925000 ;
        RECT  7.705000 86.135000  7.905000 86.335000 ;
        RECT  7.705000 86.545000  7.905000 86.745000 ;
        RECT  7.705000 86.955000  7.905000 87.155000 ;
        RECT  7.705000 87.365000  7.905000 87.565000 ;
        RECT  7.705000 87.775000  7.905000 87.975000 ;
        RECT  7.705000 88.185000  7.905000 88.385000 ;
        RECT  7.705000 88.595000  7.905000 88.795000 ;
        RECT  7.705000 89.005000  7.905000 89.205000 ;
        RECT  7.705000 89.415000  7.905000 89.615000 ;
        RECT  7.705000 89.825000  7.905000 90.025000 ;
        RECT  7.705000 90.235000  7.905000 90.435000 ;
        RECT  7.705000 90.645000  7.905000 90.845000 ;
        RECT  7.705000 91.055000  7.905000 91.255000 ;
        RECT  7.705000 91.465000  7.905000 91.665000 ;
        RECT  7.705000 91.875000  7.905000 92.075000 ;
        RECT  7.705000 92.285000  7.905000 92.485000 ;
        RECT  7.705000 92.695000  7.905000 92.895000 ;
        RECT  7.980000 17.860000  8.180000 18.060000 ;
        RECT  7.980000 18.290000  8.180000 18.490000 ;
        RECT  7.980000 18.720000  8.180000 18.920000 ;
        RECT  7.980000 19.150000  8.180000 19.350000 ;
        RECT  7.980000 19.580000  8.180000 19.780000 ;
        RECT  7.980000 20.010000  8.180000 20.210000 ;
        RECT  7.980000 20.440000  8.180000 20.640000 ;
        RECT  7.980000 20.870000  8.180000 21.070000 ;
        RECT  7.980000 21.300000  8.180000 21.500000 ;
        RECT  7.980000 21.730000  8.180000 21.930000 ;
        RECT  7.980000 22.160000  8.180000 22.360000 ;
        RECT  8.045000 68.125000  8.245000 68.325000 ;
        RECT  8.045000 68.535000  8.245000 68.735000 ;
        RECT  8.045000 68.945000  8.245000 69.145000 ;
        RECT  8.045000 69.355000  8.245000 69.555000 ;
        RECT  8.045000 69.765000  8.245000 69.965000 ;
        RECT  8.045000 70.175000  8.245000 70.375000 ;
        RECT  8.045000 70.585000  8.245000 70.785000 ;
        RECT  8.045000 70.995000  8.245000 71.195000 ;
        RECT  8.045000 71.405000  8.245000 71.605000 ;
        RECT  8.045000 71.815000  8.245000 72.015000 ;
        RECT  8.045000 72.225000  8.245000 72.425000 ;
        RECT  8.045000 72.635000  8.245000 72.835000 ;
        RECT  8.045000 73.045000  8.245000 73.245000 ;
        RECT  8.045000 73.450000  8.245000 73.650000 ;
        RECT  8.045000 73.855000  8.245000 74.055000 ;
        RECT  8.045000 74.260000  8.245000 74.460000 ;
        RECT  8.045000 74.665000  8.245000 74.865000 ;
        RECT  8.045000 75.070000  8.245000 75.270000 ;
        RECT  8.045000 75.475000  8.245000 75.675000 ;
        RECT  8.045000 75.880000  8.245000 76.080000 ;
        RECT  8.045000 76.285000  8.245000 76.485000 ;
        RECT  8.045000 76.690000  8.245000 76.890000 ;
        RECT  8.045000 77.095000  8.245000 77.295000 ;
        RECT  8.045000 77.500000  8.245000 77.700000 ;
        RECT  8.045000 77.905000  8.245000 78.105000 ;
        RECT  8.045000 78.310000  8.245000 78.510000 ;
        RECT  8.045000 78.715000  8.245000 78.915000 ;
        RECT  8.045000 79.120000  8.245000 79.320000 ;
        RECT  8.045000 79.525000  8.245000 79.725000 ;
        RECT  8.045000 79.930000  8.245000 80.130000 ;
        RECT  8.045000 80.335000  8.245000 80.535000 ;
        RECT  8.045000 80.740000  8.245000 80.940000 ;
        RECT  8.045000 81.145000  8.245000 81.345000 ;
        RECT  8.045000 81.550000  8.245000 81.750000 ;
        RECT  8.045000 81.955000  8.245000 82.155000 ;
        RECT  8.045000 82.360000  8.245000 82.560000 ;
        RECT  8.115000 82.855000  8.315000 83.055000 ;
        RECT  8.115000 83.265000  8.315000 83.465000 ;
        RECT  8.115000 83.675000  8.315000 83.875000 ;
        RECT  8.115000 84.085000  8.315000 84.285000 ;
        RECT  8.115000 84.495000  8.315000 84.695000 ;
        RECT  8.115000 84.905000  8.315000 85.105000 ;
        RECT  8.115000 85.315000  8.315000 85.515000 ;
        RECT  8.115000 85.725000  8.315000 85.925000 ;
        RECT  8.115000 86.135000  8.315000 86.335000 ;
        RECT  8.115000 86.545000  8.315000 86.745000 ;
        RECT  8.115000 86.955000  8.315000 87.155000 ;
        RECT  8.115000 87.365000  8.315000 87.565000 ;
        RECT  8.115000 87.775000  8.315000 87.975000 ;
        RECT  8.115000 88.185000  8.315000 88.385000 ;
        RECT  8.115000 88.595000  8.315000 88.795000 ;
        RECT  8.115000 89.005000  8.315000 89.205000 ;
        RECT  8.115000 89.415000  8.315000 89.615000 ;
        RECT  8.115000 89.825000  8.315000 90.025000 ;
        RECT  8.115000 90.235000  8.315000 90.435000 ;
        RECT  8.115000 90.645000  8.315000 90.845000 ;
        RECT  8.115000 91.055000  8.315000 91.255000 ;
        RECT  8.115000 91.465000  8.315000 91.665000 ;
        RECT  8.115000 91.875000  8.315000 92.075000 ;
        RECT  8.115000 92.285000  8.315000 92.485000 ;
        RECT  8.115000 92.695000  8.315000 92.895000 ;
        RECT  8.385000 17.860000  8.585000 18.060000 ;
        RECT  8.385000 18.290000  8.585000 18.490000 ;
        RECT  8.385000 18.720000  8.585000 18.920000 ;
        RECT  8.385000 19.150000  8.585000 19.350000 ;
        RECT  8.385000 19.580000  8.585000 19.780000 ;
        RECT  8.385000 20.010000  8.585000 20.210000 ;
        RECT  8.385000 20.440000  8.585000 20.640000 ;
        RECT  8.385000 20.870000  8.585000 21.070000 ;
        RECT  8.385000 21.300000  8.585000 21.500000 ;
        RECT  8.385000 21.730000  8.585000 21.930000 ;
        RECT  8.385000 22.160000  8.585000 22.360000 ;
        RECT  8.445000 68.125000  8.645000 68.325000 ;
        RECT  8.445000 68.535000  8.645000 68.735000 ;
        RECT  8.445000 68.945000  8.645000 69.145000 ;
        RECT  8.445000 69.355000  8.645000 69.555000 ;
        RECT  8.445000 69.765000  8.645000 69.965000 ;
        RECT  8.445000 70.175000  8.645000 70.375000 ;
        RECT  8.445000 70.585000  8.645000 70.785000 ;
        RECT  8.445000 70.995000  8.645000 71.195000 ;
        RECT  8.445000 71.405000  8.645000 71.605000 ;
        RECT  8.445000 71.815000  8.645000 72.015000 ;
        RECT  8.445000 72.225000  8.645000 72.425000 ;
        RECT  8.445000 72.635000  8.645000 72.835000 ;
        RECT  8.445000 73.045000  8.645000 73.245000 ;
        RECT  8.445000 73.450000  8.645000 73.650000 ;
        RECT  8.445000 73.855000  8.645000 74.055000 ;
        RECT  8.445000 74.260000  8.645000 74.460000 ;
        RECT  8.445000 74.665000  8.645000 74.865000 ;
        RECT  8.445000 75.070000  8.645000 75.270000 ;
        RECT  8.445000 75.475000  8.645000 75.675000 ;
        RECT  8.445000 75.880000  8.645000 76.080000 ;
        RECT  8.445000 76.285000  8.645000 76.485000 ;
        RECT  8.445000 76.690000  8.645000 76.890000 ;
        RECT  8.445000 77.095000  8.645000 77.295000 ;
        RECT  8.445000 77.500000  8.645000 77.700000 ;
        RECT  8.445000 77.905000  8.645000 78.105000 ;
        RECT  8.445000 78.310000  8.645000 78.510000 ;
        RECT  8.445000 78.715000  8.645000 78.915000 ;
        RECT  8.445000 79.120000  8.645000 79.320000 ;
        RECT  8.445000 79.525000  8.645000 79.725000 ;
        RECT  8.445000 79.930000  8.645000 80.130000 ;
        RECT  8.445000 80.335000  8.645000 80.535000 ;
        RECT  8.445000 80.740000  8.645000 80.940000 ;
        RECT  8.445000 81.145000  8.645000 81.345000 ;
        RECT  8.445000 81.550000  8.645000 81.750000 ;
        RECT  8.445000 81.955000  8.645000 82.155000 ;
        RECT  8.445000 82.360000  8.645000 82.560000 ;
        RECT  8.525000 82.855000  8.725000 83.055000 ;
        RECT  8.525000 83.265000  8.725000 83.465000 ;
        RECT  8.525000 83.675000  8.725000 83.875000 ;
        RECT  8.525000 84.085000  8.725000 84.285000 ;
        RECT  8.525000 84.495000  8.725000 84.695000 ;
        RECT  8.525000 84.905000  8.725000 85.105000 ;
        RECT  8.525000 85.315000  8.725000 85.515000 ;
        RECT  8.525000 85.725000  8.725000 85.925000 ;
        RECT  8.525000 86.135000  8.725000 86.335000 ;
        RECT  8.525000 86.545000  8.725000 86.745000 ;
        RECT  8.525000 86.955000  8.725000 87.155000 ;
        RECT  8.525000 87.365000  8.725000 87.565000 ;
        RECT  8.525000 87.775000  8.725000 87.975000 ;
        RECT  8.525000 88.185000  8.725000 88.385000 ;
        RECT  8.525000 88.595000  8.725000 88.795000 ;
        RECT  8.525000 89.005000  8.725000 89.205000 ;
        RECT  8.525000 89.415000  8.725000 89.615000 ;
        RECT  8.525000 89.825000  8.725000 90.025000 ;
        RECT  8.525000 90.235000  8.725000 90.435000 ;
        RECT  8.525000 90.645000  8.725000 90.845000 ;
        RECT  8.525000 91.055000  8.725000 91.255000 ;
        RECT  8.525000 91.465000  8.725000 91.665000 ;
        RECT  8.525000 91.875000  8.725000 92.075000 ;
        RECT  8.525000 92.285000  8.725000 92.485000 ;
        RECT  8.525000 92.695000  8.725000 92.895000 ;
        RECT  8.790000 17.860000  8.990000 18.060000 ;
        RECT  8.790000 18.290000  8.990000 18.490000 ;
        RECT  8.790000 18.720000  8.990000 18.920000 ;
        RECT  8.790000 19.150000  8.990000 19.350000 ;
        RECT  8.790000 19.580000  8.990000 19.780000 ;
        RECT  8.790000 20.010000  8.990000 20.210000 ;
        RECT  8.790000 20.440000  8.990000 20.640000 ;
        RECT  8.790000 20.870000  8.990000 21.070000 ;
        RECT  8.790000 21.300000  8.990000 21.500000 ;
        RECT  8.790000 21.730000  8.990000 21.930000 ;
        RECT  8.790000 22.160000  8.990000 22.360000 ;
        RECT  8.845000 68.125000  9.045000 68.325000 ;
        RECT  8.845000 68.535000  9.045000 68.735000 ;
        RECT  8.845000 68.945000  9.045000 69.145000 ;
        RECT  8.845000 69.355000  9.045000 69.555000 ;
        RECT  8.845000 69.765000  9.045000 69.965000 ;
        RECT  8.845000 70.175000  9.045000 70.375000 ;
        RECT  8.845000 70.585000  9.045000 70.785000 ;
        RECT  8.845000 70.995000  9.045000 71.195000 ;
        RECT  8.845000 71.405000  9.045000 71.605000 ;
        RECT  8.845000 71.815000  9.045000 72.015000 ;
        RECT  8.845000 72.225000  9.045000 72.425000 ;
        RECT  8.845000 72.635000  9.045000 72.835000 ;
        RECT  8.845000 73.045000  9.045000 73.245000 ;
        RECT  8.845000 73.450000  9.045000 73.650000 ;
        RECT  8.845000 73.855000  9.045000 74.055000 ;
        RECT  8.845000 74.260000  9.045000 74.460000 ;
        RECT  8.845000 74.665000  9.045000 74.865000 ;
        RECT  8.845000 75.070000  9.045000 75.270000 ;
        RECT  8.845000 75.475000  9.045000 75.675000 ;
        RECT  8.845000 75.880000  9.045000 76.080000 ;
        RECT  8.845000 76.285000  9.045000 76.485000 ;
        RECT  8.845000 76.690000  9.045000 76.890000 ;
        RECT  8.845000 77.095000  9.045000 77.295000 ;
        RECT  8.845000 77.500000  9.045000 77.700000 ;
        RECT  8.845000 77.905000  9.045000 78.105000 ;
        RECT  8.845000 78.310000  9.045000 78.510000 ;
        RECT  8.845000 78.715000  9.045000 78.915000 ;
        RECT  8.845000 79.120000  9.045000 79.320000 ;
        RECT  8.845000 79.525000  9.045000 79.725000 ;
        RECT  8.845000 79.930000  9.045000 80.130000 ;
        RECT  8.845000 80.335000  9.045000 80.535000 ;
        RECT  8.845000 80.740000  9.045000 80.940000 ;
        RECT  8.845000 81.145000  9.045000 81.345000 ;
        RECT  8.845000 81.550000  9.045000 81.750000 ;
        RECT  8.845000 81.955000  9.045000 82.155000 ;
        RECT  8.845000 82.360000  9.045000 82.560000 ;
        RECT  8.935000 82.855000  9.135000 83.055000 ;
        RECT  8.935000 83.265000  9.135000 83.465000 ;
        RECT  8.935000 83.675000  9.135000 83.875000 ;
        RECT  8.935000 84.085000  9.135000 84.285000 ;
        RECT  8.935000 84.495000  9.135000 84.695000 ;
        RECT  8.935000 84.905000  9.135000 85.105000 ;
        RECT  8.935000 85.315000  9.135000 85.515000 ;
        RECT  8.935000 85.725000  9.135000 85.925000 ;
        RECT  8.935000 86.135000  9.135000 86.335000 ;
        RECT  8.935000 86.545000  9.135000 86.745000 ;
        RECT  8.935000 86.955000  9.135000 87.155000 ;
        RECT  8.935000 87.365000  9.135000 87.565000 ;
        RECT  8.935000 87.775000  9.135000 87.975000 ;
        RECT  8.935000 88.185000  9.135000 88.385000 ;
        RECT  8.935000 88.595000  9.135000 88.795000 ;
        RECT  8.935000 89.005000  9.135000 89.205000 ;
        RECT  8.935000 89.415000  9.135000 89.615000 ;
        RECT  8.935000 89.825000  9.135000 90.025000 ;
        RECT  8.935000 90.235000  9.135000 90.435000 ;
        RECT  8.935000 90.645000  9.135000 90.845000 ;
        RECT  8.935000 91.055000  9.135000 91.255000 ;
        RECT  8.935000 91.465000  9.135000 91.665000 ;
        RECT  8.935000 91.875000  9.135000 92.075000 ;
        RECT  8.935000 92.285000  9.135000 92.485000 ;
        RECT  8.935000 92.695000  9.135000 92.895000 ;
        RECT  9.195000 17.860000  9.395000 18.060000 ;
        RECT  9.195000 18.290000  9.395000 18.490000 ;
        RECT  9.195000 18.720000  9.395000 18.920000 ;
        RECT  9.195000 19.150000  9.395000 19.350000 ;
        RECT  9.195000 19.580000  9.395000 19.780000 ;
        RECT  9.195000 20.010000  9.395000 20.210000 ;
        RECT  9.195000 20.440000  9.395000 20.640000 ;
        RECT  9.195000 20.870000  9.395000 21.070000 ;
        RECT  9.195000 21.300000  9.395000 21.500000 ;
        RECT  9.195000 21.730000  9.395000 21.930000 ;
        RECT  9.195000 22.160000  9.395000 22.360000 ;
        RECT  9.245000 68.125000  9.445000 68.325000 ;
        RECT  9.245000 68.535000  9.445000 68.735000 ;
        RECT  9.245000 68.945000  9.445000 69.145000 ;
        RECT  9.245000 69.355000  9.445000 69.555000 ;
        RECT  9.245000 69.765000  9.445000 69.965000 ;
        RECT  9.245000 70.175000  9.445000 70.375000 ;
        RECT  9.245000 70.585000  9.445000 70.785000 ;
        RECT  9.245000 70.995000  9.445000 71.195000 ;
        RECT  9.245000 71.405000  9.445000 71.605000 ;
        RECT  9.245000 71.815000  9.445000 72.015000 ;
        RECT  9.245000 72.225000  9.445000 72.425000 ;
        RECT  9.245000 72.635000  9.445000 72.835000 ;
        RECT  9.245000 73.045000  9.445000 73.245000 ;
        RECT  9.245000 73.450000  9.445000 73.650000 ;
        RECT  9.245000 73.855000  9.445000 74.055000 ;
        RECT  9.245000 74.260000  9.445000 74.460000 ;
        RECT  9.245000 74.665000  9.445000 74.865000 ;
        RECT  9.245000 75.070000  9.445000 75.270000 ;
        RECT  9.245000 75.475000  9.445000 75.675000 ;
        RECT  9.245000 75.880000  9.445000 76.080000 ;
        RECT  9.245000 76.285000  9.445000 76.485000 ;
        RECT  9.245000 76.690000  9.445000 76.890000 ;
        RECT  9.245000 77.095000  9.445000 77.295000 ;
        RECT  9.245000 77.500000  9.445000 77.700000 ;
        RECT  9.245000 77.905000  9.445000 78.105000 ;
        RECT  9.245000 78.310000  9.445000 78.510000 ;
        RECT  9.245000 78.715000  9.445000 78.915000 ;
        RECT  9.245000 79.120000  9.445000 79.320000 ;
        RECT  9.245000 79.525000  9.445000 79.725000 ;
        RECT  9.245000 79.930000  9.445000 80.130000 ;
        RECT  9.245000 80.335000  9.445000 80.535000 ;
        RECT  9.245000 80.740000  9.445000 80.940000 ;
        RECT  9.245000 81.145000  9.445000 81.345000 ;
        RECT  9.245000 81.550000  9.445000 81.750000 ;
        RECT  9.245000 81.955000  9.445000 82.155000 ;
        RECT  9.245000 82.360000  9.445000 82.560000 ;
        RECT  9.345000 82.855000  9.545000 83.055000 ;
        RECT  9.345000 83.265000  9.545000 83.465000 ;
        RECT  9.345000 83.675000  9.545000 83.875000 ;
        RECT  9.345000 84.085000  9.545000 84.285000 ;
        RECT  9.345000 84.495000  9.545000 84.695000 ;
        RECT  9.345000 84.905000  9.545000 85.105000 ;
        RECT  9.345000 85.315000  9.545000 85.515000 ;
        RECT  9.345000 85.725000  9.545000 85.925000 ;
        RECT  9.345000 86.135000  9.545000 86.335000 ;
        RECT  9.345000 86.545000  9.545000 86.745000 ;
        RECT  9.345000 86.955000  9.545000 87.155000 ;
        RECT  9.345000 87.365000  9.545000 87.565000 ;
        RECT  9.345000 87.775000  9.545000 87.975000 ;
        RECT  9.345000 88.185000  9.545000 88.385000 ;
        RECT  9.345000 88.595000  9.545000 88.795000 ;
        RECT  9.345000 89.005000  9.545000 89.205000 ;
        RECT  9.345000 89.415000  9.545000 89.615000 ;
        RECT  9.345000 89.825000  9.545000 90.025000 ;
        RECT  9.345000 90.235000  9.545000 90.435000 ;
        RECT  9.345000 90.645000  9.545000 90.845000 ;
        RECT  9.345000 91.055000  9.545000 91.255000 ;
        RECT  9.345000 91.465000  9.545000 91.665000 ;
        RECT  9.345000 91.875000  9.545000 92.075000 ;
        RECT  9.345000 92.285000  9.545000 92.485000 ;
        RECT  9.345000 92.695000  9.545000 92.895000 ;
        RECT  9.600000 17.860000  9.800000 18.060000 ;
        RECT  9.600000 18.290000  9.800000 18.490000 ;
        RECT  9.600000 18.720000  9.800000 18.920000 ;
        RECT  9.600000 19.150000  9.800000 19.350000 ;
        RECT  9.600000 19.580000  9.800000 19.780000 ;
        RECT  9.600000 20.010000  9.800000 20.210000 ;
        RECT  9.600000 20.440000  9.800000 20.640000 ;
        RECT  9.600000 20.870000  9.800000 21.070000 ;
        RECT  9.600000 21.300000  9.800000 21.500000 ;
        RECT  9.600000 21.730000  9.800000 21.930000 ;
        RECT  9.600000 22.160000  9.800000 22.360000 ;
        RECT  9.645000 68.125000  9.845000 68.325000 ;
        RECT  9.645000 68.535000  9.845000 68.735000 ;
        RECT  9.645000 68.945000  9.845000 69.145000 ;
        RECT  9.645000 69.355000  9.845000 69.555000 ;
        RECT  9.645000 69.765000  9.845000 69.965000 ;
        RECT  9.645000 70.175000  9.845000 70.375000 ;
        RECT  9.645000 70.585000  9.845000 70.785000 ;
        RECT  9.645000 70.995000  9.845000 71.195000 ;
        RECT  9.645000 71.405000  9.845000 71.605000 ;
        RECT  9.645000 71.815000  9.845000 72.015000 ;
        RECT  9.645000 72.225000  9.845000 72.425000 ;
        RECT  9.645000 72.635000  9.845000 72.835000 ;
        RECT  9.645000 73.045000  9.845000 73.245000 ;
        RECT  9.645000 73.450000  9.845000 73.650000 ;
        RECT  9.645000 73.855000  9.845000 74.055000 ;
        RECT  9.645000 74.260000  9.845000 74.460000 ;
        RECT  9.645000 74.665000  9.845000 74.865000 ;
        RECT  9.645000 75.070000  9.845000 75.270000 ;
        RECT  9.645000 75.475000  9.845000 75.675000 ;
        RECT  9.645000 75.880000  9.845000 76.080000 ;
        RECT  9.645000 76.285000  9.845000 76.485000 ;
        RECT  9.645000 76.690000  9.845000 76.890000 ;
        RECT  9.645000 77.095000  9.845000 77.295000 ;
        RECT  9.645000 77.500000  9.845000 77.700000 ;
        RECT  9.645000 77.905000  9.845000 78.105000 ;
        RECT  9.645000 78.310000  9.845000 78.510000 ;
        RECT  9.645000 78.715000  9.845000 78.915000 ;
        RECT  9.645000 79.120000  9.845000 79.320000 ;
        RECT  9.645000 79.525000  9.845000 79.725000 ;
        RECT  9.645000 79.930000  9.845000 80.130000 ;
        RECT  9.645000 80.335000  9.845000 80.535000 ;
        RECT  9.645000 80.740000  9.845000 80.940000 ;
        RECT  9.645000 81.145000  9.845000 81.345000 ;
        RECT  9.645000 81.550000  9.845000 81.750000 ;
        RECT  9.645000 81.955000  9.845000 82.155000 ;
        RECT  9.645000 82.360000  9.845000 82.560000 ;
        RECT  9.755000 82.855000  9.955000 83.055000 ;
        RECT  9.755000 83.265000  9.955000 83.465000 ;
        RECT  9.755000 83.675000  9.955000 83.875000 ;
        RECT  9.755000 84.085000  9.955000 84.285000 ;
        RECT  9.755000 84.495000  9.955000 84.695000 ;
        RECT  9.755000 84.905000  9.955000 85.105000 ;
        RECT  9.755000 85.315000  9.955000 85.515000 ;
        RECT  9.755000 85.725000  9.955000 85.925000 ;
        RECT  9.755000 86.135000  9.955000 86.335000 ;
        RECT  9.755000 86.545000  9.955000 86.745000 ;
        RECT  9.755000 86.955000  9.955000 87.155000 ;
        RECT  9.755000 87.365000  9.955000 87.565000 ;
        RECT  9.755000 87.775000  9.955000 87.975000 ;
        RECT  9.755000 88.185000  9.955000 88.385000 ;
        RECT  9.755000 88.595000  9.955000 88.795000 ;
        RECT  9.755000 89.005000  9.955000 89.205000 ;
        RECT  9.755000 89.415000  9.955000 89.615000 ;
        RECT  9.755000 89.825000  9.955000 90.025000 ;
        RECT  9.755000 90.235000  9.955000 90.435000 ;
        RECT  9.755000 90.645000  9.955000 90.845000 ;
        RECT  9.755000 91.055000  9.955000 91.255000 ;
        RECT  9.755000 91.465000  9.955000 91.665000 ;
        RECT  9.755000 91.875000  9.955000 92.075000 ;
        RECT  9.755000 92.285000  9.955000 92.485000 ;
        RECT  9.755000 92.695000  9.955000 92.895000 ;
        RECT 10.005000 17.860000 10.205000 18.060000 ;
        RECT 10.005000 18.290000 10.205000 18.490000 ;
        RECT 10.005000 18.720000 10.205000 18.920000 ;
        RECT 10.005000 19.150000 10.205000 19.350000 ;
        RECT 10.005000 19.580000 10.205000 19.780000 ;
        RECT 10.005000 20.010000 10.205000 20.210000 ;
        RECT 10.005000 20.440000 10.205000 20.640000 ;
        RECT 10.005000 20.870000 10.205000 21.070000 ;
        RECT 10.005000 21.300000 10.205000 21.500000 ;
        RECT 10.005000 21.730000 10.205000 21.930000 ;
        RECT 10.005000 22.160000 10.205000 22.360000 ;
        RECT 10.045000 68.125000 10.245000 68.325000 ;
        RECT 10.045000 68.535000 10.245000 68.735000 ;
        RECT 10.045000 68.945000 10.245000 69.145000 ;
        RECT 10.045000 69.355000 10.245000 69.555000 ;
        RECT 10.045000 69.765000 10.245000 69.965000 ;
        RECT 10.045000 70.175000 10.245000 70.375000 ;
        RECT 10.045000 70.585000 10.245000 70.785000 ;
        RECT 10.045000 70.995000 10.245000 71.195000 ;
        RECT 10.045000 71.405000 10.245000 71.605000 ;
        RECT 10.045000 71.815000 10.245000 72.015000 ;
        RECT 10.045000 72.225000 10.245000 72.425000 ;
        RECT 10.045000 72.635000 10.245000 72.835000 ;
        RECT 10.045000 73.045000 10.245000 73.245000 ;
        RECT 10.045000 73.450000 10.245000 73.650000 ;
        RECT 10.045000 73.855000 10.245000 74.055000 ;
        RECT 10.045000 74.260000 10.245000 74.460000 ;
        RECT 10.045000 74.665000 10.245000 74.865000 ;
        RECT 10.045000 75.070000 10.245000 75.270000 ;
        RECT 10.045000 75.475000 10.245000 75.675000 ;
        RECT 10.045000 75.880000 10.245000 76.080000 ;
        RECT 10.045000 76.285000 10.245000 76.485000 ;
        RECT 10.045000 76.690000 10.245000 76.890000 ;
        RECT 10.045000 77.095000 10.245000 77.295000 ;
        RECT 10.045000 77.500000 10.245000 77.700000 ;
        RECT 10.045000 77.905000 10.245000 78.105000 ;
        RECT 10.045000 78.310000 10.245000 78.510000 ;
        RECT 10.045000 78.715000 10.245000 78.915000 ;
        RECT 10.045000 79.120000 10.245000 79.320000 ;
        RECT 10.045000 79.525000 10.245000 79.725000 ;
        RECT 10.045000 79.930000 10.245000 80.130000 ;
        RECT 10.045000 80.335000 10.245000 80.535000 ;
        RECT 10.045000 80.740000 10.245000 80.940000 ;
        RECT 10.045000 81.145000 10.245000 81.345000 ;
        RECT 10.045000 81.550000 10.245000 81.750000 ;
        RECT 10.045000 81.955000 10.245000 82.155000 ;
        RECT 10.045000 82.360000 10.245000 82.560000 ;
        RECT 10.165000 82.855000 10.365000 83.055000 ;
        RECT 10.165000 83.265000 10.365000 83.465000 ;
        RECT 10.165000 83.675000 10.365000 83.875000 ;
        RECT 10.165000 84.085000 10.365000 84.285000 ;
        RECT 10.165000 84.495000 10.365000 84.695000 ;
        RECT 10.165000 84.905000 10.365000 85.105000 ;
        RECT 10.165000 85.315000 10.365000 85.515000 ;
        RECT 10.165000 85.725000 10.365000 85.925000 ;
        RECT 10.165000 86.135000 10.365000 86.335000 ;
        RECT 10.165000 86.545000 10.365000 86.745000 ;
        RECT 10.165000 86.955000 10.365000 87.155000 ;
        RECT 10.165000 87.365000 10.365000 87.565000 ;
        RECT 10.165000 87.775000 10.365000 87.975000 ;
        RECT 10.165000 88.185000 10.365000 88.385000 ;
        RECT 10.165000 88.595000 10.365000 88.795000 ;
        RECT 10.165000 89.005000 10.365000 89.205000 ;
        RECT 10.165000 89.415000 10.365000 89.615000 ;
        RECT 10.165000 89.825000 10.365000 90.025000 ;
        RECT 10.165000 90.235000 10.365000 90.435000 ;
        RECT 10.165000 90.645000 10.365000 90.845000 ;
        RECT 10.165000 91.055000 10.365000 91.255000 ;
        RECT 10.165000 91.465000 10.365000 91.665000 ;
        RECT 10.165000 91.875000 10.365000 92.075000 ;
        RECT 10.165000 92.285000 10.365000 92.485000 ;
        RECT 10.165000 92.695000 10.365000 92.895000 ;
        RECT 10.410000 17.860000 10.610000 18.060000 ;
        RECT 10.410000 18.290000 10.610000 18.490000 ;
        RECT 10.410000 18.720000 10.610000 18.920000 ;
        RECT 10.410000 19.150000 10.610000 19.350000 ;
        RECT 10.410000 19.580000 10.610000 19.780000 ;
        RECT 10.410000 20.010000 10.610000 20.210000 ;
        RECT 10.410000 20.440000 10.610000 20.640000 ;
        RECT 10.410000 20.870000 10.610000 21.070000 ;
        RECT 10.410000 21.300000 10.610000 21.500000 ;
        RECT 10.410000 21.730000 10.610000 21.930000 ;
        RECT 10.410000 22.160000 10.610000 22.360000 ;
        RECT 10.445000 68.125000 10.645000 68.325000 ;
        RECT 10.445000 68.535000 10.645000 68.735000 ;
        RECT 10.445000 68.945000 10.645000 69.145000 ;
        RECT 10.445000 69.355000 10.645000 69.555000 ;
        RECT 10.445000 69.765000 10.645000 69.965000 ;
        RECT 10.445000 70.175000 10.645000 70.375000 ;
        RECT 10.445000 70.585000 10.645000 70.785000 ;
        RECT 10.445000 70.995000 10.645000 71.195000 ;
        RECT 10.445000 71.405000 10.645000 71.605000 ;
        RECT 10.445000 71.815000 10.645000 72.015000 ;
        RECT 10.445000 72.225000 10.645000 72.425000 ;
        RECT 10.445000 72.635000 10.645000 72.835000 ;
        RECT 10.445000 73.045000 10.645000 73.245000 ;
        RECT 10.445000 73.450000 10.645000 73.650000 ;
        RECT 10.445000 73.855000 10.645000 74.055000 ;
        RECT 10.445000 74.260000 10.645000 74.460000 ;
        RECT 10.445000 74.665000 10.645000 74.865000 ;
        RECT 10.445000 75.070000 10.645000 75.270000 ;
        RECT 10.445000 75.475000 10.645000 75.675000 ;
        RECT 10.445000 75.880000 10.645000 76.080000 ;
        RECT 10.445000 76.285000 10.645000 76.485000 ;
        RECT 10.445000 76.690000 10.645000 76.890000 ;
        RECT 10.445000 77.095000 10.645000 77.295000 ;
        RECT 10.445000 77.500000 10.645000 77.700000 ;
        RECT 10.445000 77.905000 10.645000 78.105000 ;
        RECT 10.445000 78.310000 10.645000 78.510000 ;
        RECT 10.445000 78.715000 10.645000 78.915000 ;
        RECT 10.445000 79.120000 10.645000 79.320000 ;
        RECT 10.445000 79.525000 10.645000 79.725000 ;
        RECT 10.445000 79.930000 10.645000 80.130000 ;
        RECT 10.445000 80.335000 10.645000 80.535000 ;
        RECT 10.445000 80.740000 10.645000 80.940000 ;
        RECT 10.445000 81.145000 10.645000 81.345000 ;
        RECT 10.445000 81.550000 10.645000 81.750000 ;
        RECT 10.445000 81.955000 10.645000 82.155000 ;
        RECT 10.445000 82.360000 10.645000 82.560000 ;
        RECT 10.575000 82.855000 10.775000 83.055000 ;
        RECT 10.575000 83.265000 10.775000 83.465000 ;
        RECT 10.575000 83.675000 10.775000 83.875000 ;
        RECT 10.575000 84.085000 10.775000 84.285000 ;
        RECT 10.575000 84.495000 10.775000 84.695000 ;
        RECT 10.575000 84.905000 10.775000 85.105000 ;
        RECT 10.575000 85.315000 10.775000 85.515000 ;
        RECT 10.575000 85.725000 10.775000 85.925000 ;
        RECT 10.575000 86.135000 10.775000 86.335000 ;
        RECT 10.575000 86.545000 10.775000 86.745000 ;
        RECT 10.575000 86.955000 10.775000 87.155000 ;
        RECT 10.575000 87.365000 10.775000 87.565000 ;
        RECT 10.575000 87.775000 10.775000 87.975000 ;
        RECT 10.575000 88.185000 10.775000 88.385000 ;
        RECT 10.575000 88.595000 10.775000 88.795000 ;
        RECT 10.575000 89.005000 10.775000 89.205000 ;
        RECT 10.575000 89.415000 10.775000 89.615000 ;
        RECT 10.575000 89.825000 10.775000 90.025000 ;
        RECT 10.575000 90.235000 10.775000 90.435000 ;
        RECT 10.575000 90.645000 10.775000 90.845000 ;
        RECT 10.575000 91.055000 10.775000 91.255000 ;
        RECT 10.575000 91.465000 10.775000 91.665000 ;
        RECT 10.575000 91.875000 10.775000 92.075000 ;
        RECT 10.575000 92.285000 10.775000 92.485000 ;
        RECT 10.575000 92.695000 10.775000 92.895000 ;
        RECT 10.815000 17.860000 11.015000 18.060000 ;
        RECT 10.815000 18.290000 11.015000 18.490000 ;
        RECT 10.815000 18.720000 11.015000 18.920000 ;
        RECT 10.815000 19.150000 11.015000 19.350000 ;
        RECT 10.815000 19.580000 11.015000 19.780000 ;
        RECT 10.815000 20.010000 11.015000 20.210000 ;
        RECT 10.815000 20.440000 11.015000 20.640000 ;
        RECT 10.815000 20.870000 11.015000 21.070000 ;
        RECT 10.815000 21.300000 11.015000 21.500000 ;
        RECT 10.815000 21.730000 11.015000 21.930000 ;
        RECT 10.815000 22.160000 11.015000 22.360000 ;
        RECT 10.845000 68.125000 11.045000 68.325000 ;
        RECT 10.845000 68.535000 11.045000 68.735000 ;
        RECT 10.845000 68.945000 11.045000 69.145000 ;
        RECT 10.845000 69.355000 11.045000 69.555000 ;
        RECT 10.845000 69.765000 11.045000 69.965000 ;
        RECT 10.845000 70.175000 11.045000 70.375000 ;
        RECT 10.845000 70.585000 11.045000 70.785000 ;
        RECT 10.845000 70.995000 11.045000 71.195000 ;
        RECT 10.845000 71.405000 11.045000 71.605000 ;
        RECT 10.845000 71.815000 11.045000 72.015000 ;
        RECT 10.845000 72.225000 11.045000 72.425000 ;
        RECT 10.845000 72.635000 11.045000 72.835000 ;
        RECT 10.845000 73.045000 11.045000 73.245000 ;
        RECT 10.845000 73.450000 11.045000 73.650000 ;
        RECT 10.845000 73.855000 11.045000 74.055000 ;
        RECT 10.845000 74.260000 11.045000 74.460000 ;
        RECT 10.845000 74.665000 11.045000 74.865000 ;
        RECT 10.845000 75.070000 11.045000 75.270000 ;
        RECT 10.845000 75.475000 11.045000 75.675000 ;
        RECT 10.845000 75.880000 11.045000 76.080000 ;
        RECT 10.845000 76.285000 11.045000 76.485000 ;
        RECT 10.845000 76.690000 11.045000 76.890000 ;
        RECT 10.845000 77.095000 11.045000 77.295000 ;
        RECT 10.845000 77.500000 11.045000 77.700000 ;
        RECT 10.845000 77.905000 11.045000 78.105000 ;
        RECT 10.845000 78.310000 11.045000 78.510000 ;
        RECT 10.845000 78.715000 11.045000 78.915000 ;
        RECT 10.845000 79.120000 11.045000 79.320000 ;
        RECT 10.845000 79.525000 11.045000 79.725000 ;
        RECT 10.845000 79.930000 11.045000 80.130000 ;
        RECT 10.845000 80.335000 11.045000 80.535000 ;
        RECT 10.845000 80.740000 11.045000 80.940000 ;
        RECT 10.845000 81.145000 11.045000 81.345000 ;
        RECT 10.845000 81.550000 11.045000 81.750000 ;
        RECT 10.845000 81.955000 11.045000 82.155000 ;
        RECT 10.845000 82.360000 11.045000 82.560000 ;
        RECT 10.985000 82.855000 11.185000 83.055000 ;
        RECT 10.985000 83.265000 11.185000 83.465000 ;
        RECT 10.985000 83.675000 11.185000 83.875000 ;
        RECT 10.985000 84.085000 11.185000 84.285000 ;
        RECT 10.985000 84.495000 11.185000 84.695000 ;
        RECT 10.985000 84.905000 11.185000 85.105000 ;
        RECT 10.985000 85.315000 11.185000 85.515000 ;
        RECT 10.985000 85.725000 11.185000 85.925000 ;
        RECT 10.985000 86.135000 11.185000 86.335000 ;
        RECT 10.985000 86.545000 11.185000 86.745000 ;
        RECT 10.985000 86.955000 11.185000 87.155000 ;
        RECT 10.985000 87.365000 11.185000 87.565000 ;
        RECT 10.985000 87.775000 11.185000 87.975000 ;
        RECT 10.985000 88.185000 11.185000 88.385000 ;
        RECT 10.985000 88.595000 11.185000 88.795000 ;
        RECT 10.985000 89.005000 11.185000 89.205000 ;
        RECT 10.985000 89.415000 11.185000 89.615000 ;
        RECT 10.985000 89.825000 11.185000 90.025000 ;
        RECT 10.985000 90.235000 11.185000 90.435000 ;
        RECT 10.985000 90.645000 11.185000 90.845000 ;
        RECT 10.985000 91.055000 11.185000 91.255000 ;
        RECT 10.985000 91.465000 11.185000 91.665000 ;
        RECT 10.985000 91.875000 11.185000 92.075000 ;
        RECT 10.985000 92.285000 11.185000 92.485000 ;
        RECT 10.985000 92.695000 11.185000 92.895000 ;
        RECT 11.220000 17.860000 11.420000 18.060000 ;
        RECT 11.220000 18.290000 11.420000 18.490000 ;
        RECT 11.220000 18.720000 11.420000 18.920000 ;
        RECT 11.220000 19.150000 11.420000 19.350000 ;
        RECT 11.220000 19.580000 11.420000 19.780000 ;
        RECT 11.220000 20.010000 11.420000 20.210000 ;
        RECT 11.220000 20.440000 11.420000 20.640000 ;
        RECT 11.220000 20.870000 11.420000 21.070000 ;
        RECT 11.220000 21.300000 11.420000 21.500000 ;
        RECT 11.220000 21.730000 11.420000 21.930000 ;
        RECT 11.220000 22.160000 11.420000 22.360000 ;
        RECT 11.245000 68.125000 11.445000 68.325000 ;
        RECT 11.245000 68.535000 11.445000 68.735000 ;
        RECT 11.245000 68.945000 11.445000 69.145000 ;
        RECT 11.245000 69.355000 11.445000 69.555000 ;
        RECT 11.245000 69.765000 11.445000 69.965000 ;
        RECT 11.245000 70.175000 11.445000 70.375000 ;
        RECT 11.245000 70.585000 11.445000 70.785000 ;
        RECT 11.245000 70.995000 11.445000 71.195000 ;
        RECT 11.245000 71.405000 11.445000 71.605000 ;
        RECT 11.245000 71.815000 11.445000 72.015000 ;
        RECT 11.245000 72.225000 11.445000 72.425000 ;
        RECT 11.245000 72.635000 11.445000 72.835000 ;
        RECT 11.245000 73.045000 11.445000 73.245000 ;
        RECT 11.245000 73.450000 11.445000 73.650000 ;
        RECT 11.245000 73.855000 11.445000 74.055000 ;
        RECT 11.245000 74.260000 11.445000 74.460000 ;
        RECT 11.245000 74.665000 11.445000 74.865000 ;
        RECT 11.245000 75.070000 11.445000 75.270000 ;
        RECT 11.245000 75.475000 11.445000 75.675000 ;
        RECT 11.245000 75.880000 11.445000 76.080000 ;
        RECT 11.245000 76.285000 11.445000 76.485000 ;
        RECT 11.245000 76.690000 11.445000 76.890000 ;
        RECT 11.245000 77.095000 11.445000 77.295000 ;
        RECT 11.245000 77.500000 11.445000 77.700000 ;
        RECT 11.245000 77.905000 11.445000 78.105000 ;
        RECT 11.245000 78.310000 11.445000 78.510000 ;
        RECT 11.245000 78.715000 11.445000 78.915000 ;
        RECT 11.245000 79.120000 11.445000 79.320000 ;
        RECT 11.245000 79.525000 11.445000 79.725000 ;
        RECT 11.245000 79.930000 11.445000 80.130000 ;
        RECT 11.245000 80.335000 11.445000 80.535000 ;
        RECT 11.245000 80.740000 11.445000 80.940000 ;
        RECT 11.245000 81.145000 11.445000 81.345000 ;
        RECT 11.245000 81.550000 11.445000 81.750000 ;
        RECT 11.245000 81.955000 11.445000 82.155000 ;
        RECT 11.245000 82.360000 11.445000 82.560000 ;
        RECT 11.395000 82.855000 11.595000 83.055000 ;
        RECT 11.395000 83.265000 11.595000 83.465000 ;
        RECT 11.395000 83.675000 11.595000 83.875000 ;
        RECT 11.395000 84.085000 11.595000 84.285000 ;
        RECT 11.395000 84.495000 11.595000 84.695000 ;
        RECT 11.395000 84.905000 11.595000 85.105000 ;
        RECT 11.395000 85.315000 11.595000 85.515000 ;
        RECT 11.395000 85.725000 11.595000 85.925000 ;
        RECT 11.395000 86.135000 11.595000 86.335000 ;
        RECT 11.395000 86.545000 11.595000 86.745000 ;
        RECT 11.395000 86.955000 11.595000 87.155000 ;
        RECT 11.395000 87.365000 11.595000 87.565000 ;
        RECT 11.395000 87.775000 11.595000 87.975000 ;
        RECT 11.395000 88.185000 11.595000 88.385000 ;
        RECT 11.395000 88.595000 11.595000 88.795000 ;
        RECT 11.395000 89.005000 11.595000 89.205000 ;
        RECT 11.395000 89.415000 11.595000 89.615000 ;
        RECT 11.395000 89.825000 11.595000 90.025000 ;
        RECT 11.395000 90.235000 11.595000 90.435000 ;
        RECT 11.395000 90.645000 11.595000 90.845000 ;
        RECT 11.395000 91.055000 11.595000 91.255000 ;
        RECT 11.395000 91.465000 11.595000 91.665000 ;
        RECT 11.395000 91.875000 11.595000 92.075000 ;
        RECT 11.395000 92.285000 11.595000 92.485000 ;
        RECT 11.395000 92.695000 11.595000 92.895000 ;
        RECT 11.625000 17.860000 11.825000 18.060000 ;
        RECT 11.625000 18.290000 11.825000 18.490000 ;
        RECT 11.625000 18.720000 11.825000 18.920000 ;
        RECT 11.625000 19.150000 11.825000 19.350000 ;
        RECT 11.625000 19.580000 11.825000 19.780000 ;
        RECT 11.625000 20.010000 11.825000 20.210000 ;
        RECT 11.625000 20.440000 11.825000 20.640000 ;
        RECT 11.625000 20.870000 11.825000 21.070000 ;
        RECT 11.625000 21.300000 11.825000 21.500000 ;
        RECT 11.625000 21.730000 11.825000 21.930000 ;
        RECT 11.625000 22.160000 11.825000 22.360000 ;
        RECT 11.645000 68.125000 11.845000 68.325000 ;
        RECT 11.645000 68.535000 11.845000 68.735000 ;
        RECT 11.645000 68.945000 11.845000 69.145000 ;
        RECT 11.645000 69.355000 11.845000 69.555000 ;
        RECT 11.645000 69.765000 11.845000 69.965000 ;
        RECT 11.645000 70.175000 11.845000 70.375000 ;
        RECT 11.645000 70.585000 11.845000 70.785000 ;
        RECT 11.645000 70.995000 11.845000 71.195000 ;
        RECT 11.645000 71.405000 11.845000 71.605000 ;
        RECT 11.645000 71.815000 11.845000 72.015000 ;
        RECT 11.645000 72.225000 11.845000 72.425000 ;
        RECT 11.645000 72.635000 11.845000 72.835000 ;
        RECT 11.645000 73.045000 11.845000 73.245000 ;
        RECT 11.645000 73.450000 11.845000 73.650000 ;
        RECT 11.645000 73.855000 11.845000 74.055000 ;
        RECT 11.645000 74.260000 11.845000 74.460000 ;
        RECT 11.645000 74.665000 11.845000 74.865000 ;
        RECT 11.645000 75.070000 11.845000 75.270000 ;
        RECT 11.645000 75.475000 11.845000 75.675000 ;
        RECT 11.645000 75.880000 11.845000 76.080000 ;
        RECT 11.645000 76.285000 11.845000 76.485000 ;
        RECT 11.645000 76.690000 11.845000 76.890000 ;
        RECT 11.645000 77.095000 11.845000 77.295000 ;
        RECT 11.645000 77.500000 11.845000 77.700000 ;
        RECT 11.645000 77.905000 11.845000 78.105000 ;
        RECT 11.645000 78.310000 11.845000 78.510000 ;
        RECT 11.645000 78.715000 11.845000 78.915000 ;
        RECT 11.645000 79.120000 11.845000 79.320000 ;
        RECT 11.645000 79.525000 11.845000 79.725000 ;
        RECT 11.645000 79.930000 11.845000 80.130000 ;
        RECT 11.645000 80.335000 11.845000 80.535000 ;
        RECT 11.645000 80.740000 11.845000 80.940000 ;
        RECT 11.645000 81.145000 11.845000 81.345000 ;
        RECT 11.645000 81.550000 11.845000 81.750000 ;
        RECT 11.645000 81.955000 11.845000 82.155000 ;
        RECT 11.645000 82.360000 11.845000 82.560000 ;
        RECT 11.805000 82.855000 12.005000 83.055000 ;
        RECT 11.805000 83.265000 12.005000 83.465000 ;
        RECT 11.805000 83.675000 12.005000 83.875000 ;
        RECT 11.805000 84.085000 12.005000 84.285000 ;
        RECT 11.805000 84.495000 12.005000 84.695000 ;
        RECT 11.805000 84.905000 12.005000 85.105000 ;
        RECT 11.805000 85.315000 12.005000 85.515000 ;
        RECT 11.805000 85.725000 12.005000 85.925000 ;
        RECT 11.805000 86.135000 12.005000 86.335000 ;
        RECT 11.805000 86.545000 12.005000 86.745000 ;
        RECT 11.805000 86.955000 12.005000 87.155000 ;
        RECT 11.805000 87.365000 12.005000 87.565000 ;
        RECT 11.805000 87.775000 12.005000 87.975000 ;
        RECT 11.805000 88.185000 12.005000 88.385000 ;
        RECT 11.805000 88.595000 12.005000 88.795000 ;
        RECT 11.805000 89.005000 12.005000 89.205000 ;
        RECT 11.805000 89.415000 12.005000 89.615000 ;
        RECT 11.805000 89.825000 12.005000 90.025000 ;
        RECT 11.805000 90.235000 12.005000 90.435000 ;
        RECT 11.805000 90.645000 12.005000 90.845000 ;
        RECT 11.805000 91.055000 12.005000 91.255000 ;
        RECT 11.805000 91.465000 12.005000 91.665000 ;
        RECT 11.805000 91.875000 12.005000 92.075000 ;
        RECT 11.805000 92.285000 12.005000 92.485000 ;
        RECT 11.805000 92.695000 12.005000 92.895000 ;
        RECT 12.030000 17.860000 12.230000 18.060000 ;
        RECT 12.030000 18.290000 12.230000 18.490000 ;
        RECT 12.030000 18.720000 12.230000 18.920000 ;
        RECT 12.030000 19.150000 12.230000 19.350000 ;
        RECT 12.030000 19.580000 12.230000 19.780000 ;
        RECT 12.030000 20.010000 12.230000 20.210000 ;
        RECT 12.030000 20.440000 12.230000 20.640000 ;
        RECT 12.030000 20.870000 12.230000 21.070000 ;
        RECT 12.030000 21.300000 12.230000 21.500000 ;
        RECT 12.030000 21.730000 12.230000 21.930000 ;
        RECT 12.030000 22.160000 12.230000 22.360000 ;
        RECT 12.045000 68.125000 12.245000 68.325000 ;
        RECT 12.045000 68.535000 12.245000 68.735000 ;
        RECT 12.045000 68.945000 12.245000 69.145000 ;
        RECT 12.045000 69.355000 12.245000 69.555000 ;
        RECT 12.045000 69.765000 12.245000 69.965000 ;
        RECT 12.045000 70.175000 12.245000 70.375000 ;
        RECT 12.045000 70.585000 12.245000 70.785000 ;
        RECT 12.045000 70.995000 12.245000 71.195000 ;
        RECT 12.045000 71.405000 12.245000 71.605000 ;
        RECT 12.045000 71.815000 12.245000 72.015000 ;
        RECT 12.045000 72.225000 12.245000 72.425000 ;
        RECT 12.045000 72.635000 12.245000 72.835000 ;
        RECT 12.045000 73.045000 12.245000 73.245000 ;
        RECT 12.045000 73.450000 12.245000 73.650000 ;
        RECT 12.045000 73.855000 12.245000 74.055000 ;
        RECT 12.045000 74.260000 12.245000 74.460000 ;
        RECT 12.045000 74.665000 12.245000 74.865000 ;
        RECT 12.045000 75.070000 12.245000 75.270000 ;
        RECT 12.045000 75.475000 12.245000 75.675000 ;
        RECT 12.045000 75.880000 12.245000 76.080000 ;
        RECT 12.045000 76.285000 12.245000 76.485000 ;
        RECT 12.045000 76.690000 12.245000 76.890000 ;
        RECT 12.045000 77.095000 12.245000 77.295000 ;
        RECT 12.045000 77.500000 12.245000 77.700000 ;
        RECT 12.045000 77.905000 12.245000 78.105000 ;
        RECT 12.045000 78.310000 12.245000 78.510000 ;
        RECT 12.045000 78.715000 12.245000 78.915000 ;
        RECT 12.045000 79.120000 12.245000 79.320000 ;
        RECT 12.045000 79.525000 12.245000 79.725000 ;
        RECT 12.045000 79.930000 12.245000 80.130000 ;
        RECT 12.045000 80.335000 12.245000 80.535000 ;
        RECT 12.045000 80.740000 12.245000 80.940000 ;
        RECT 12.045000 81.145000 12.245000 81.345000 ;
        RECT 12.045000 81.550000 12.245000 81.750000 ;
        RECT 12.045000 81.955000 12.245000 82.155000 ;
        RECT 12.045000 82.360000 12.245000 82.560000 ;
        RECT 12.215000 82.855000 12.415000 83.055000 ;
        RECT 12.215000 83.265000 12.415000 83.465000 ;
        RECT 12.215000 83.675000 12.415000 83.875000 ;
        RECT 12.215000 84.085000 12.415000 84.285000 ;
        RECT 12.215000 84.495000 12.415000 84.695000 ;
        RECT 12.215000 84.905000 12.415000 85.105000 ;
        RECT 12.215000 85.315000 12.415000 85.515000 ;
        RECT 12.215000 85.725000 12.415000 85.925000 ;
        RECT 12.215000 86.135000 12.415000 86.335000 ;
        RECT 12.215000 86.545000 12.415000 86.745000 ;
        RECT 12.215000 86.955000 12.415000 87.155000 ;
        RECT 12.215000 87.365000 12.415000 87.565000 ;
        RECT 12.215000 87.775000 12.415000 87.975000 ;
        RECT 12.215000 88.185000 12.415000 88.385000 ;
        RECT 12.215000 88.595000 12.415000 88.795000 ;
        RECT 12.215000 89.005000 12.415000 89.205000 ;
        RECT 12.215000 89.415000 12.415000 89.615000 ;
        RECT 12.215000 89.825000 12.415000 90.025000 ;
        RECT 12.215000 90.235000 12.415000 90.435000 ;
        RECT 12.215000 90.645000 12.415000 90.845000 ;
        RECT 12.215000 91.055000 12.415000 91.255000 ;
        RECT 12.215000 91.465000 12.415000 91.665000 ;
        RECT 12.215000 91.875000 12.415000 92.075000 ;
        RECT 12.215000 92.285000 12.415000 92.485000 ;
        RECT 12.215000 92.695000 12.415000 92.895000 ;
        RECT 12.435000 17.860000 12.635000 18.060000 ;
        RECT 12.435000 18.290000 12.635000 18.490000 ;
        RECT 12.435000 18.720000 12.635000 18.920000 ;
        RECT 12.435000 19.150000 12.635000 19.350000 ;
        RECT 12.435000 19.580000 12.635000 19.780000 ;
        RECT 12.435000 20.010000 12.635000 20.210000 ;
        RECT 12.435000 20.440000 12.635000 20.640000 ;
        RECT 12.435000 20.870000 12.635000 21.070000 ;
        RECT 12.435000 21.300000 12.635000 21.500000 ;
        RECT 12.435000 21.730000 12.635000 21.930000 ;
        RECT 12.435000 22.160000 12.635000 22.360000 ;
        RECT 12.445000 68.125000 12.645000 68.325000 ;
        RECT 12.445000 68.535000 12.645000 68.735000 ;
        RECT 12.445000 68.945000 12.645000 69.145000 ;
        RECT 12.445000 69.355000 12.645000 69.555000 ;
        RECT 12.445000 69.765000 12.645000 69.965000 ;
        RECT 12.445000 70.175000 12.645000 70.375000 ;
        RECT 12.445000 70.585000 12.645000 70.785000 ;
        RECT 12.445000 70.995000 12.645000 71.195000 ;
        RECT 12.445000 71.405000 12.645000 71.605000 ;
        RECT 12.445000 71.815000 12.645000 72.015000 ;
        RECT 12.445000 72.225000 12.645000 72.425000 ;
        RECT 12.445000 72.635000 12.645000 72.835000 ;
        RECT 12.445000 73.045000 12.645000 73.245000 ;
        RECT 12.445000 73.450000 12.645000 73.650000 ;
        RECT 12.445000 73.855000 12.645000 74.055000 ;
        RECT 12.445000 74.260000 12.645000 74.460000 ;
        RECT 12.445000 74.665000 12.645000 74.865000 ;
        RECT 12.445000 75.070000 12.645000 75.270000 ;
        RECT 12.445000 75.475000 12.645000 75.675000 ;
        RECT 12.445000 75.880000 12.645000 76.080000 ;
        RECT 12.445000 76.285000 12.645000 76.485000 ;
        RECT 12.445000 76.690000 12.645000 76.890000 ;
        RECT 12.445000 77.095000 12.645000 77.295000 ;
        RECT 12.445000 77.500000 12.645000 77.700000 ;
        RECT 12.445000 77.905000 12.645000 78.105000 ;
        RECT 12.445000 78.310000 12.645000 78.510000 ;
        RECT 12.445000 78.715000 12.645000 78.915000 ;
        RECT 12.445000 79.120000 12.645000 79.320000 ;
        RECT 12.445000 79.525000 12.645000 79.725000 ;
        RECT 12.445000 79.930000 12.645000 80.130000 ;
        RECT 12.445000 80.335000 12.645000 80.535000 ;
        RECT 12.445000 80.740000 12.645000 80.940000 ;
        RECT 12.445000 81.145000 12.645000 81.345000 ;
        RECT 12.445000 81.550000 12.645000 81.750000 ;
        RECT 12.445000 81.955000 12.645000 82.155000 ;
        RECT 12.445000 82.360000 12.645000 82.560000 ;
        RECT 12.625000 82.855000 12.825000 83.055000 ;
        RECT 12.625000 83.265000 12.825000 83.465000 ;
        RECT 12.625000 83.675000 12.825000 83.875000 ;
        RECT 12.625000 84.085000 12.825000 84.285000 ;
        RECT 12.625000 84.495000 12.825000 84.695000 ;
        RECT 12.625000 84.905000 12.825000 85.105000 ;
        RECT 12.625000 85.315000 12.825000 85.515000 ;
        RECT 12.625000 85.725000 12.825000 85.925000 ;
        RECT 12.625000 86.135000 12.825000 86.335000 ;
        RECT 12.625000 86.545000 12.825000 86.745000 ;
        RECT 12.625000 86.955000 12.825000 87.155000 ;
        RECT 12.625000 87.365000 12.825000 87.565000 ;
        RECT 12.625000 87.775000 12.825000 87.975000 ;
        RECT 12.625000 88.185000 12.825000 88.385000 ;
        RECT 12.625000 88.595000 12.825000 88.795000 ;
        RECT 12.625000 89.005000 12.825000 89.205000 ;
        RECT 12.625000 89.415000 12.825000 89.615000 ;
        RECT 12.625000 89.825000 12.825000 90.025000 ;
        RECT 12.625000 90.235000 12.825000 90.435000 ;
        RECT 12.625000 90.645000 12.825000 90.845000 ;
        RECT 12.625000 91.055000 12.825000 91.255000 ;
        RECT 12.625000 91.465000 12.825000 91.665000 ;
        RECT 12.625000 91.875000 12.825000 92.075000 ;
        RECT 12.625000 92.285000 12.825000 92.485000 ;
        RECT 12.625000 92.695000 12.825000 92.895000 ;
        RECT 12.840000 17.860000 13.040000 18.060000 ;
        RECT 12.840000 18.290000 13.040000 18.490000 ;
        RECT 12.840000 18.720000 13.040000 18.920000 ;
        RECT 12.840000 19.150000 13.040000 19.350000 ;
        RECT 12.840000 19.580000 13.040000 19.780000 ;
        RECT 12.840000 20.010000 13.040000 20.210000 ;
        RECT 12.840000 20.440000 13.040000 20.640000 ;
        RECT 12.840000 20.870000 13.040000 21.070000 ;
        RECT 12.840000 21.300000 13.040000 21.500000 ;
        RECT 12.840000 21.730000 13.040000 21.930000 ;
        RECT 12.840000 22.160000 13.040000 22.360000 ;
        RECT 12.845000 68.125000 13.045000 68.325000 ;
        RECT 12.845000 68.535000 13.045000 68.735000 ;
        RECT 12.845000 68.945000 13.045000 69.145000 ;
        RECT 12.845000 69.355000 13.045000 69.555000 ;
        RECT 12.845000 69.765000 13.045000 69.965000 ;
        RECT 12.845000 70.175000 13.045000 70.375000 ;
        RECT 12.845000 70.585000 13.045000 70.785000 ;
        RECT 12.845000 70.995000 13.045000 71.195000 ;
        RECT 12.845000 71.405000 13.045000 71.605000 ;
        RECT 12.845000 71.815000 13.045000 72.015000 ;
        RECT 12.845000 72.225000 13.045000 72.425000 ;
        RECT 12.845000 72.635000 13.045000 72.835000 ;
        RECT 12.845000 73.045000 13.045000 73.245000 ;
        RECT 12.845000 73.450000 13.045000 73.650000 ;
        RECT 12.845000 73.855000 13.045000 74.055000 ;
        RECT 12.845000 74.260000 13.045000 74.460000 ;
        RECT 12.845000 74.665000 13.045000 74.865000 ;
        RECT 12.845000 75.070000 13.045000 75.270000 ;
        RECT 12.845000 75.475000 13.045000 75.675000 ;
        RECT 12.845000 75.880000 13.045000 76.080000 ;
        RECT 12.845000 76.285000 13.045000 76.485000 ;
        RECT 12.845000 76.690000 13.045000 76.890000 ;
        RECT 12.845000 77.095000 13.045000 77.295000 ;
        RECT 12.845000 77.500000 13.045000 77.700000 ;
        RECT 12.845000 77.905000 13.045000 78.105000 ;
        RECT 12.845000 78.310000 13.045000 78.510000 ;
        RECT 12.845000 78.715000 13.045000 78.915000 ;
        RECT 12.845000 79.120000 13.045000 79.320000 ;
        RECT 12.845000 79.525000 13.045000 79.725000 ;
        RECT 12.845000 79.930000 13.045000 80.130000 ;
        RECT 12.845000 80.335000 13.045000 80.535000 ;
        RECT 12.845000 80.740000 13.045000 80.940000 ;
        RECT 12.845000 81.145000 13.045000 81.345000 ;
        RECT 12.845000 81.550000 13.045000 81.750000 ;
        RECT 12.845000 81.955000 13.045000 82.155000 ;
        RECT 12.845000 82.360000 13.045000 82.560000 ;
        RECT 13.030000 82.855000 13.230000 83.055000 ;
        RECT 13.030000 83.265000 13.230000 83.465000 ;
        RECT 13.030000 83.675000 13.230000 83.875000 ;
        RECT 13.030000 84.085000 13.230000 84.285000 ;
        RECT 13.030000 84.495000 13.230000 84.695000 ;
        RECT 13.030000 84.905000 13.230000 85.105000 ;
        RECT 13.030000 85.315000 13.230000 85.515000 ;
        RECT 13.030000 85.725000 13.230000 85.925000 ;
        RECT 13.030000 86.135000 13.230000 86.335000 ;
        RECT 13.030000 86.545000 13.230000 86.745000 ;
        RECT 13.030000 86.955000 13.230000 87.155000 ;
        RECT 13.030000 87.365000 13.230000 87.565000 ;
        RECT 13.030000 87.775000 13.230000 87.975000 ;
        RECT 13.030000 88.185000 13.230000 88.385000 ;
        RECT 13.030000 88.595000 13.230000 88.795000 ;
        RECT 13.030000 89.005000 13.230000 89.205000 ;
        RECT 13.030000 89.415000 13.230000 89.615000 ;
        RECT 13.030000 89.825000 13.230000 90.025000 ;
        RECT 13.030000 90.235000 13.230000 90.435000 ;
        RECT 13.030000 90.645000 13.230000 90.845000 ;
        RECT 13.030000 91.055000 13.230000 91.255000 ;
        RECT 13.030000 91.465000 13.230000 91.665000 ;
        RECT 13.030000 91.875000 13.230000 92.075000 ;
        RECT 13.030000 92.285000 13.230000 92.485000 ;
        RECT 13.030000 92.695000 13.230000 92.895000 ;
        RECT 13.245000 17.860000 13.445000 18.060000 ;
        RECT 13.245000 18.290000 13.445000 18.490000 ;
        RECT 13.245000 18.720000 13.445000 18.920000 ;
        RECT 13.245000 19.150000 13.445000 19.350000 ;
        RECT 13.245000 19.580000 13.445000 19.780000 ;
        RECT 13.245000 20.010000 13.445000 20.210000 ;
        RECT 13.245000 20.440000 13.445000 20.640000 ;
        RECT 13.245000 20.870000 13.445000 21.070000 ;
        RECT 13.245000 21.300000 13.445000 21.500000 ;
        RECT 13.245000 21.730000 13.445000 21.930000 ;
        RECT 13.245000 22.160000 13.445000 22.360000 ;
        RECT 13.245000 68.125000 13.445000 68.325000 ;
        RECT 13.245000 68.535000 13.445000 68.735000 ;
        RECT 13.245000 68.945000 13.445000 69.145000 ;
        RECT 13.245000 69.355000 13.445000 69.555000 ;
        RECT 13.245000 69.765000 13.445000 69.965000 ;
        RECT 13.245000 70.175000 13.445000 70.375000 ;
        RECT 13.245000 70.585000 13.445000 70.785000 ;
        RECT 13.245000 70.995000 13.445000 71.195000 ;
        RECT 13.245000 71.405000 13.445000 71.605000 ;
        RECT 13.245000 71.815000 13.445000 72.015000 ;
        RECT 13.245000 72.225000 13.445000 72.425000 ;
        RECT 13.245000 72.635000 13.445000 72.835000 ;
        RECT 13.245000 73.045000 13.445000 73.245000 ;
        RECT 13.245000 73.450000 13.445000 73.650000 ;
        RECT 13.245000 73.855000 13.445000 74.055000 ;
        RECT 13.245000 74.260000 13.445000 74.460000 ;
        RECT 13.245000 74.665000 13.445000 74.865000 ;
        RECT 13.245000 75.070000 13.445000 75.270000 ;
        RECT 13.245000 75.475000 13.445000 75.675000 ;
        RECT 13.245000 75.880000 13.445000 76.080000 ;
        RECT 13.245000 76.285000 13.445000 76.485000 ;
        RECT 13.245000 76.690000 13.445000 76.890000 ;
        RECT 13.245000 77.095000 13.445000 77.295000 ;
        RECT 13.245000 77.500000 13.445000 77.700000 ;
        RECT 13.245000 77.905000 13.445000 78.105000 ;
        RECT 13.245000 78.310000 13.445000 78.510000 ;
        RECT 13.245000 78.715000 13.445000 78.915000 ;
        RECT 13.245000 79.120000 13.445000 79.320000 ;
        RECT 13.245000 79.525000 13.445000 79.725000 ;
        RECT 13.245000 79.930000 13.445000 80.130000 ;
        RECT 13.245000 80.335000 13.445000 80.535000 ;
        RECT 13.245000 80.740000 13.445000 80.940000 ;
        RECT 13.245000 81.145000 13.445000 81.345000 ;
        RECT 13.245000 81.550000 13.445000 81.750000 ;
        RECT 13.245000 81.955000 13.445000 82.155000 ;
        RECT 13.245000 82.360000 13.445000 82.560000 ;
        RECT 13.435000 82.855000 13.635000 83.055000 ;
        RECT 13.435000 83.265000 13.635000 83.465000 ;
        RECT 13.435000 83.675000 13.635000 83.875000 ;
        RECT 13.435000 84.085000 13.635000 84.285000 ;
        RECT 13.435000 84.495000 13.635000 84.695000 ;
        RECT 13.435000 84.905000 13.635000 85.105000 ;
        RECT 13.435000 85.315000 13.635000 85.515000 ;
        RECT 13.435000 85.725000 13.635000 85.925000 ;
        RECT 13.435000 86.135000 13.635000 86.335000 ;
        RECT 13.435000 86.545000 13.635000 86.745000 ;
        RECT 13.435000 86.955000 13.635000 87.155000 ;
        RECT 13.435000 87.365000 13.635000 87.565000 ;
        RECT 13.435000 87.775000 13.635000 87.975000 ;
        RECT 13.435000 88.185000 13.635000 88.385000 ;
        RECT 13.435000 88.595000 13.635000 88.795000 ;
        RECT 13.435000 89.005000 13.635000 89.205000 ;
        RECT 13.435000 89.415000 13.635000 89.615000 ;
        RECT 13.435000 89.825000 13.635000 90.025000 ;
        RECT 13.435000 90.235000 13.635000 90.435000 ;
        RECT 13.435000 90.645000 13.635000 90.845000 ;
        RECT 13.435000 91.055000 13.635000 91.255000 ;
        RECT 13.435000 91.465000 13.635000 91.665000 ;
        RECT 13.435000 91.875000 13.635000 92.075000 ;
        RECT 13.435000 92.285000 13.635000 92.485000 ;
        RECT 13.435000 92.695000 13.635000 92.895000 ;
        RECT 13.645000 68.125000 13.845000 68.325000 ;
        RECT 13.645000 68.535000 13.845000 68.735000 ;
        RECT 13.645000 68.945000 13.845000 69.145000 ;
        RECT 13.645000 69.355000 13.845000 69.555000 ;
        RECT 13.645000 69.765000 13.845000 69.965000 ;
        RECT 13.645000 70.175000 13.845000 70.375000 ;
        RECT 13.645000 70.585000 13.845000 70.785000 ;
        RECT 13.645000 70.995000 13.845000 71.195000 ;
        RECT 13.645000 71.405000 13.845000 71.605000 ;
        RECT 13.645000 71.815000 13.845000 72.015000 ;
        RECT 13.645000 72.225000 13.845000 72.425000 ;
        RECT 13.645000 72.635000 13.845000 72.835000 ;
        RECT 13.645000 73.045000 13.845000 73.245000 ;
        RECT 13.645000 73.450000 13.845000 73.650000 ;
        RECT 13.645000 73.855000 13.845000 74.055000 ;
        RECT 13.645000 74.260000 13.845000 74.460000 ;
        RECT 13.645000 74.665000 13.845000 74.865000 ;
        RECT 13.645000 75.070000 13.845000 75.270000 ;
        RECT 13.645000 75.475000 13.845000 75.675000 ;
        RECT 13.645000 75.880000 13.845000 76.080000 ;
        RECT 13.645000 76.285000 13.845000 76.485000 ;
        RECT 13.645000 76.690000 13.845000 76.890000 ;
        RECT 13.645000 77.095000 13.845000 77.295000 ;
        RECT 13.645000 77.500000 13.845000 77.700000 ;
        RECT 13.645000 77.905000 13.845000 78.105000 ;
        RECT 13.645000 78.310000 13.845000 78.510000 ;
        RECT 13.645000 78.715000 13.845000 78.915000 ;
        RECT 13.645000 79.120000 13.845000 79.320000 ;
        RECT 13.645000 79.525000 13.845000 79.725000 ;
        RECT 13.645000 79.930000 13.845000 80.130000 ;
        RECT 13.645000 80.335000 13.845000 80.535000 ;
        RECT 13.645000 80.740000 13.845000 80.940000 ;
        RECT 13.645000 81.145000 13.845000 81.345000 ;
        RECT 13.645000 81.550000 13.845000 81.750000 ;
        RECT 13.645000 81.955000 13.845000 82.155000 ;
        RECT 13.645000 82.360000 13.845000 82.560000 ;
        RECT 13.650000 17.860000 13.850000 18.060000 ;
        RECT 13.650000 18.290000 13.850000 18.490000 ;
        RECT 13.650000 18.720000 13.850000 18.920000 ;
        RECT 13.650000 19.150000 13.850000 19.350000 ;
        RECT 13.650000 19.580000 13.850000 19.780000 ;
        RECT 13.650000 20.010000 13.850000 20.210000 ;
        RECT 13.650000 20.440000 13.850000 20.640000 ;
        RECT 13.650000 20.870000 13.850000 21.070000 ;
        RECT 13.650000 21.300000 13.850000 21.500000 ;
        RECT 13.650000 21.730000 13.850000 21.930000 ;
        RECT 13.650000 22.160000 13.850000 22.360000 ;
        RECT 13.840000 82.855000 14.040000 83.055000 ;
        RECT 13.840000 83.265000 14.040000 83.465000 ;
        RECT 13.840000 83.675000 14.040000 83.875000 ;
        RECT 13.840000 84.085000 14.040000 84.285000 ;
        RECT 13.840000 84.495000 14.040000 84.695000 ;
        RECT 13.840000 84.905000 14.040000 85.105000 ;
        RECT 13.840000 85.315000 14.040000 85.515000 ;
        RECT 13.840000 85.725000 14.040000 85.925000 ;
        RECT 13.840000 86.135000 14.040000 86.335000 ;
        RECT 13.840000 86.545000 14.040000 86.745000 ;
        RECT 13.840000 86.955000 14.040000 87.155000 ;
        RECT 13.840000 87.365000 14.040000 87.565000 ;
        RECT 13.840000 87.775000 14.040000 87.975000 ;
        RECT 13.840000 88.185000 14.040000 88.385000 ;
        RECT 13.840000 88.595000 14.040000 88.795000 ;
        RECT 13.840000 89.005000 14.040000 89.205000 ;
        RECT 13.840000 89.415000 14.040000 89.615000 ;
        RECT 13.840000 89.825000 14.040000 90.025000 ;
        RECT 13.840000 90.235000 14.040000 90.435000 ;
        RECT 13.840000 90.645000 14.040000 90.845000 ;
        RECT 13.840000 91.055000 14.040000 91.255000 ;
        RECT 13.840000 91.465000 14.040000 91.665000 ;
        RECT 13.840000 91.875000 14.040000 92.075000 ;
        RECT 13.840000 92.285000 14.040000 92.485000 ;
        RECT 13.840000 92.695000 14.040000 92.895000 ;
        RECT 14.045000 68.125000 14.245000 68.325000 ;
        RECT 14.045000 68.535000 14.245000 68.735000 ;
        RECT 14.045000 68.945000 14.245000 69.145000 ;
        RECT 14.045000 69.355000 14.245000 69.555000 ;
        RECT 14.045000 69.765000 14.245000 69.965000 ;
        RECT 14.045000 70.175000 14.245000 70.375000 ;
        RECT 14.045000 70.585000 14.245000 70.785000 ;
        RECT 14.045000 70.995000 14.245000 71.195000 ;
        RECT 14.045000 71.405000 14.245000 71.605000 ;
        RECT 14.045000 71.815000 14.245000 72.015000 ;
        RECT 14.045000 72.225000 14.245000 72.425000 ;
        RECT 14.045000 72.635000 14.245000 72.835000 ;
        RECT 14.045000 73.045000 14.245000 73.245000 ;
        RECT 14.045000 73.450000 14.245000 73.650000 ;
        RECT 14.045000 73.855000 14.245000 74.055000 ;
        RECT 14.045000 74.260000 14.245000 74.460000 ;
        RECT 14.045000 74.665000 14.245000 74.865000 ;
        RECT 14.045000 75.070000 14.245000 75.270000 ;
        RECT 14.045000 75.475000 14.245000 75.675000 ;
        RECT 14.045000 75.880000 14.245000 76.080000 ;
        RECT 14.045000 76.285000 14.245000 76.485000 ;
        RECT 14.045000 76.690000 14.245000 76.890000 ;
        RECT 14.045000 77.095000 14.245000 77.295000 ;
        RECT 14.045000 77.500000 14.245000 77.700000 ;
        RECT 14.045000 77.905000 14.245000 78.105000 ;
        RECT 14.045000 78.310000 14.245000 78.510000 ;
        RECT 14.045000 78.715000 14.245000 78.915000 ;
        RECT 14.045000 79.120000 14.245000 79.320000 ;
        RECT 14.045000 79.525000 14.245000 79.725000 ;
        RECT 14.045000 79.930000 14.245000 80.130000 ;
        RECT 14.045000 80.335000 14.245000 80.535000 ;
        RECT 14.045000 80.740000 14.245000 80.940000 ;
        RECT 14.045000 81.145000 14.245000 81.345000 ;
        RECT 14.045000 81.550000 14.245000 81.750000 ;
        RECT 14.045000 81.955000 14.245000 82.155000 ;
        RECT 14.045000 82.360000 14.245000 82.560000 ;
        RECT 14.055000 17.860000 14.255000 18.060000 ;
        RECT 14.055000 18.290000 14.255000 18.490000 ;
        RECT 14.055000 18.720000 14.255000 18.920000 ;
        RECT 14.055000 19.150000 14.255000 19.350000 ;
        RECT 14.055000 19.580000 14.255000 19.780000 ;
        RECT 14.055000 20.010000 14.255000 20.210000 ;
        RECT 14.055000 20.440000 14.255000 20.640000 ;
        RECT 14.055000 20.870000 14.255000 21.070000 ;
        RECT 14.055000 21.300000 14.255000 21.500000 ;
        RECT 14.055000 21.730000 14.255000 21.930000 ;
        RECT 14.055000 22.160000 14.255000 22.360000 ;
        RECT 14.320000 91.015000 14.520000 91.215000 ;
        RECT 14.320000 91.445000 14.520000 91.645000 ;
        RECT 14.340000 88.410000 14.540000 88.610000 ;
        RECT 14.340000 88.835000 14.540000 89.035000 ;
        RECT 14.340000 89.265000 14.540000 89.465000 ;
        RECT 14.340000 89.695000 14.540000 89.895000 ;
        RECT 14.340000 90.125000 14.540000 90.325000 ;
        RECT 14.340000 90.555000 14.540000 90.755000 ;
        RECT 14.445000 68.125000 14.645000 68.325000 ;
        RECT 14.445000 68.535000 14.645000 68.735000 ;
        RECT 14.445000 68.945000 14.645000 69.145000 ;
        RECT 14.445000 69.355000 14.645000 69.555000 ;
        RECT 14.445000 69.765000 14.645000 69.965000 ;
        RECT 14.445000 70.175000 14.645000 70.375000 ;
        RECT 14.445000 70.585000 14.645000 70.785000 ;
        RECT 14.445000 70.995000 14.645000 71.195000 ;
        RECT 14.445000 71.405000 14.645000 71.605000 ;
        RECT 14.445000 71.815000 14.645000 72.015000 ;
        RECT 14.445000 72.225000 14.645000 72.425000 ;
        RECT 14.445000 72.635000 14.645000 72.835000 ;
        RECT 14.445000 73.045000 14.645000 73.245000 ;
        RECT 14.445000 73.450000 14.645000 73.650000 ;
        RECT 14.445000 73.855000 14.645000 74.055000 ;
        RECT 14.445000 74.260000 14.645000 74.460000 ;
        RECT 14.445000 74.665000 14.645000 74.865000 ;
        RECT 14.445000 75.070000 14.645000 75.270000 ;
        RECT 14.445000 75.475000 14.645000 75.675000 ;
        RECT 14.445000 75.880000 14.645000 76.080000 ;
        RECT 14.445000 76.285000 14.645000 76.485000 ;
        RECT 14.445000 76.690000 14.645000 76.890000 ;
        RECT 14.445000 77.095000 14.645000 77.295000 ;
        RECT 14.445000 77.500000 14.645000 77.700000 ;
        RECT 14.445000 77.905000 14.645000 78.105000 ;
        RECT 14.445000 78.310000 14.645000 78.510000 ;
        RECT 14.445000 78.715000 14.645000 78.915000 ;
        RECT 14.445000 79.120000 14.645000 79.320000 ;
        RECT 14.445000 79.525000 14.645000 79.725000 ;
        RECT 14.445000 79.930000 14.645000 80.130000 ;
        RECT 14.445000 80.335000 14.645000 80.535000 ;
        RECT 14.445000 80.740000 14.645000 80.940000 ;
        RECT 14.445000 81.145000 14.645000 81.345000 ;
        RECT 14.445000 81.550000 14.645000 81.750000 ;
        RECT 14.445000 81.955000 14.645000 82.155000 ;
        RECT 14.445000 82.360000 14.645000 82.560000 ;
        RECT 14.460000 17.860000 14.660000 18.060000 ;
        RECT 14.460000 18.290000 14.660000 18.490000 ;
        RECT 14.460000 18.720000 14.660000 18.920000 ;
        RECT 14.460000 19.150000 14.660000 19.350000 ;
        RECT 14.460000 19.580000 14.660000 19.780000 ;
        RECT 14.460000 20.010000 14.660000 20.210000 ;
        RECT 14.460000 20.440000 14.660000 20.640000 ;
        RECT 14.460000 20.870000 14.660000 21.070000 ;
        RECT 14.460000 21.300000 14.660000 21.500000 ;
        RECT 14.460000 21.730000 14.660000 21.930000 ;
        RECT 14.460000 22.160000 14.660000 22.360000 ;
        RECT 14.465000 83.055000 14.665000 83.255000 ;
        RECT 14.465000 83.455000 14.665000 83.655000 ;
        RECT 14.465000 83.855000 14.665000 84.055000 ;
        RECT 14.465000 84.255000 14.665000 84.455000 ;
        RECT 14.465000 84.655000 14.665000 84.855000 ;
        RECT 14.465000 85.055000 14.665000 85.255000 ;
        RECT 14.465000 85.455000 14.665000 85.655000 ;
        RECT 14.465000 85.855000 14.665000 86.055000 ;
        RECT 14.465000 86.255000 14.665000 86.455000 ;
        RECT 14.465000 86.660000 14.665000 86.860000 ;
        RECT 14.465000 87.065000 14.665000 87.265000 ;
        RECT 14.465000 87.470000 14.665000 87.670000 ;
        RECT 14.465000 87.875000 14.665000 88.075000 ;
        RECT 14.750000 88.410000 14.950000 88.610000 ;
        RECT 14.750000 88.835000 14.950000 89.035000 ;
        RECT 14.750000 89.265000 14.950000 89.465000 ;
        RECT 14.750000 89.695000 14.950000 89.895000 ;
        RECT 14.750000 90.125000 14.950000 90.325000 ;
        RECT 14.750000 90.555000 14.950000 90.755000 ;
        RECT 14.845000 68.125000 15.045000 68.325000 ;
        RECT 14.845000 68.535000 15.045000 68.735000 ;
        RECT 14.845000 68.945000 15.045000 69.145000 ;
        RECT 14.845000 69.355000 15.045000 69.555000 ;
        RECT 14.845000 69.765000 15.045000 69.965000 ;
        RECT 14.845000 70.175000 15.045000 70.375000 ;
        RECT 14.845000 70.585000 15.045000 70.785000 ;
        RECT 14.845000 70.995000 15.045000 71.195000 ;
        RECT 14.845000 71.405000 15.045000 71.605000 ;
        RECT 14.845000 71.815000 15.045000 72.015000 ;
        RECT 14.845000 72.225000 15.045000 72.425000 ;
        RECT 14.845000 72.635000 15.045000 72.835000 ;
        RECT 14.845000 73.045000 15.045000 73.245000 ;
        RECT 14.845000 73.450000 15.045000 73.650000 ;
        RECT 14.845000 73.855000 15.045000 74.055000 ;
        RECT 14.845000 74.260000 15.045000 74.460000 ;
        RECT 14.845000 74.665000 15.045000 74.865000 ;
        RECT 14.845000 75.070000 15.045000 75.270000 ;
        RECT 14.845000 75.475000 15.045000 75.675000 ;
        RECT 14.845000 75.880000 15.045000 76.080000 ;
        RECT 14.845000 76.285000 15.045000 76.485000 ;
        RECT 14.845000 76.690000 15.045000 76.890000 ;
        RECT 14.845000 77.095000 15.045000 77.295000 ;
        RECT 14.845000 77.500000 15.045000 77.700000 ;
        RECT 14.845000 77.905000 15.045000 78.105000 ;
        RECT 14.845000 78.310000 15.045000 78.510000 ;
        RECT 14.845000 78.715000 15.045000 78.915000 ;
        RECT 14.845000 79.120000 15.045000 79.320000 ;
        RECT 14.845000 79.525000 15.045000 79.725000 ;
        RECT 14.845000 79.930000 15.045000 80.130000 ;
        RECT 14.845000 80.335000 15.045000 80.535000 ;
        RECT 14.845000 80.740000 15.045000 80.940000 ;
        RECT 14.845000 81.145000 15.045000 81.345000 ;
        RECT 14.845000 81.550000 15.045000 81.750000 ;
        RECT 14.845000 81.955000 15.045000 82.155000 ;
        RECT 14.845000 82.360000 15.045000 82.560000 ;
        RECT 14.865000 17.860000 15.065000 18.060000 ;
        RECT 14.865000 18.290000 15.065000 18.490000 ;
        RECT 14.865000 18.720000 15.065000 18.920000 ;
        RECT 14.865000 19.150000 15.065000 19.350000 ;
        RECT 14.865000 19.580000 15.065000 19.780000 ;
        RECT 14.865000 20.010000 15.065000 20.210000 ;
        RECT 14.865000 20.440000 15.065000 20.640000 ;
        RECT 14.865000 20.870000 15.065000 21.070000 ;
        RECT 14.865000 21.300000 15.065000 21.500000 ;
        RECT 14.865000 21.730000 15.065000 21.930000 ;
        RECT 14.865000 22.160000 15.065000 22.360000 ;
        RECT 14.875000 83.055000 15.075000 83.255000 ;
        RECT 14.875000 83.455000 15.075000 83.655000 ;
        RECT 14.875000 83.855000 15.075000 84.055000 ;
        RECT 14.875000 84.255000 15.075000 84.455000 ;
        RECT 14.875000 84.655000 15.075000 84.855000 ;
        RECT 14.875000 85.055000 15.075000 85.255000 ;
        RECT 14.875000 85.455000 15.075000 85.655000 ;
        RECT 14.875000 85.855000 15.075000 86.055000 ;
        RECT 14.875000 86.255000 15.075000 86.455000 ;
        RECT 14.875000 86.660000 15.075000 86.860000 ;
        RECT 14.875000 87.065000 15.075000 87.265000 ;
        RECT 14.875000 87.470000 15.075000 87.670000 ;
        RECT 14.875000 87.875000 15.075000 88.075000 ;
        RECT 15.100000 91.015000 15.300000 91.215000 ;
        RECT 15.100000 91.445000 15.300000 91.645000 ;
        RECT 15.160000 88.410000 15.360000 88.610000 ;
        RECT 15.160000 88.835000 15.360000 89.035000 ;
        RECT 15.160000 89.265000 15.360000 89.465000 ;
        RECT 15.160000 89.695000 15.360000 89.895000 ;
        RECT 15.160000 90.125000 15.360000 90.325000 ;
        RECT 15.160000 90.555000 15.360000 90.755000 ;
        RECT 15.245000 68.125000 15.445000 68.325000 ;
        RECT 15.245000 68.535000 15.445000 68.735000 ;
        RECT 15.245000 68.945000 15.445000 69.145000 ;
        RECT 15.245000 69.355000 15.445000 69.555000 ;
        RECT 15.245000 69.765000 15.445000 69.965000 ;
        RECT 15.245000 70.175000 15.445000 70.375000 ;
        RECT 15.245000 70.585000 15.445000 70.785000 ;
        RECT 15.245000 70.995000 15.445000 71.195000 ;
        RECT 15.245000 71.405000 15.445000 71.605000 ;
        RECT 15.245000 71.815000 15.445000 72.015000 ;
        RECT 15.245000 72.225000 15.445000 72.425000 ;
        RECT 15.245000 72.635000 15.445000 72.835000 ;
        RECT 15.245000 73.045000 15.445000 73.245000 ;
        RECT 15.245000 73.450000 15.445000 73.650000 ;
        RECT 15.245000 73.855000 15.445000 74.055000 ;
        RECT 15.245000 74.260000 15.445000 74.460000 ;
        RECT 15.245000 74.665000 15.445000 74.865000 ;
        RECT 15.245000 75.070000 15.445000 75.270000 ;
        RECT 15.245000 75.475000 15.445000 75.675000 ;
        RECT 15.245000 75.880000 15.445000 76.080000 ;
        RECT 15.245000 76.285000 15.445000 76.485000 ;
        RECT 15.245000 76.690000 15.445000 76.890000 ;
        RECT 15.245000 77.095000 15.445000 77.295000 ;
        RECT 15.245000 77.500000 15.445000 77.700000 ;
        RECT 15.245000 77.905000 15.445000 78.105000 ;
        RECT 15.245000 78.310000 15.445000 78.510000 ;
        RECT 15.245000 78.715000 15.445000 78.915000 ;
        RECT 15.245000 79.120000 15.445000 79.320000 ;
        RECT 15.245000 79.525000 15.445000 79.725000 ;
        RECT 15.245000 79.930000 15.445000 80.130000 ;
        RECT 15.245000 80.335000 15.445000 80.535000 ;
        RECT 15.245000 80.740000 15.445000 80.940000 ;
        RECT 15.245000 81.145000 15.445000 81.345000 ;
        RECT 15.245000 81.550000 15.445000 81.750000 ;
        RECT 15.245000 81.955000 15.445000 82.155000 ;
        RECT 15.245000 82.360000 15.445000 82.560000 ;
        RECT 15.270000 17.860000 15.470000 18.060000 ;
        RECT 15.270000 18.290000 15.470000 18.490000 ;
        RECT 15.270000 18.720000 15.470000 18.920000 ;
        RECT 15.270000 19.150000 15.470000 19.350000 ;
        RECT 15.270000 19.580000 15.470000 19.780000 ;
        RECT 15.270000 20.010000 15.470000 20.210000 ;
        RECT 15.270000 20.440000 15.470000 20.640000 ;
        RECT 15.270000 20.870000 15.470000 21.070000 ;
        RECT 15.270000 21.300000 15.470000 21.500000 ;
        RECT 15.270000 21.730000 15.470000 21.930000 ;
        RECT 15.270000 22.160000 15.470000 22.360000 ;
        RECT 15.285000 83.055000 15.485000 83.255000 ;
        RECT 15.285000 83.455000 15.485000 83.655000 ;
        RECT 15.285000 83.855000 15.485000 84.055000 ;
        RECT 15.285000 84.255000 15.485000 84.455000 ;
        RECT 15.285000 84.655000 15.485000 84.855000 ;
        RECT 15.285000 85.055000 15.485000 85.255000 ;
        RECT 15.285000 85.455000 15.485000 85.655000 ;
        RECT 15.285000 85.855000 15.485000 86.055000 ;
        RECT 15.285000 86.255000 15.485000 86.455000 ;
        RECT 15.285000 86.660000 15.485000 86.860000 ;
        RECT 15.285000 87.065000 15.485000 87.265000 ;
        RECT 15.285000 87.470000 15.485000 87.670000 ;
        RECT 15.285000 87.875000 15.485000 88.075000 ;
        RECT 15.570000 88.410000 15.770000 88.610000 ;
        RECT 15.570000 88.835000 15.770000 89.035000 ;
        RECT 15.570000 89.265000 15.770000 89.465000 ;
        RECT 15.570000 89.695000 15.770000 89.895000 ;
        RECT 15.570000 90.125000 15.770000 90.325000 ;
        RECT 15.570000 90.555000 15.770000 90.755000 ;
        RECT 15.645000 68.125000 15.845000 68.325000 ;
        RECT 15.645000 68.535000 15.845000 68.735000 ;
        RECT 15.645000 68.945000 15.845000 69.145000 ;
        RECT 15.645000 69.355000 15.845000 69.555000 ;
        RECT 15.645000 69.765000 15.845000 69.965000 ;
        RECT 15.645000 70.175000 15.845000 70.375000 ;
        RECT 15.645000 70.585000 15.845000 70.785000 ;
        RECT 15.645000 70.995000 15.845000 71.195000 ;
        RECT 15.645000 71.405000 15.845000 71.605000 ;
        RECT 15.645000 71.815000 15.845000 72.015000 ;
        RECT 15.645000 72.225000 15.845000 72.425000 ;
        RECT 15.645000 72.635000 15.845000 72.835000 ;
        RECT 15.645000 73.045000 15.845000 73.245000 ;
        RECT 15.645000 73.450000 15.845000 73.650000 ;
        RECT 15.645000 73.855000 15.845000 74.055000 ;
        RECT 15.645000 74.260000 15.845000 74.460000 ;
        RECT 15.645000 74.665000 15.845000 74.865000 ;
        RECT 15.645000 75.070000 15.845000 75.270000 ;
        RECT 15.645000 75.475000 15.845000 75.675000 ;
        RECT 15.645000 75.880000 15.845000 76.080000 ;
        RECT 15.645000 76.285000 15.845000 76.485000 ;
        RECT 15.645000 76.690000 15.845000 76.890000 ;
        RECT 15.645000 77.095000 15.845000 77.295000 ;
        RECT 15.645000 77.500000 15.845000 77.700000 ;
        RECT 15.645000 77.905000 15.845000 78.105000 ;
        RECT 15.645000 78.310000 15.845000 78.510000 ;
        RECT 15.645000 78.715000 15.845000 78.915000 ;
        RECT 15.645000 79.120000 15.845000 79.320000 ;
        RECT 15.645000 79.525000 15.845000 79.725000 ;
        RECT 15.645000 79.930000 15.845000 80.130000 ;
        RECT 15.645000 80.335000 15.845000 80.535000 ;
        RECT 15.645000 80.740000 15.845000 80.940000 ;
        RECT 15.645000 81.145000 15.845000 81.345000 ;
        RECT 15.645000 81.550000 15.845000 81.750000 ;
        RECT 15.645000 81.955000 15.845000 82.155000 ;
        RECT 15.645000 82.360000 15.845000 82.560000 ;
        RECT 15.675000 17.860000 15.875000 18.060000 ;
        RECT 15.675000 18.290000 15.875000 18.490000 ;
        RECT 15.675000 18.720000 15.875000 18.920000 ;
        RECT 15.675000 19.150000 15.875000 19.350000 ;
        RECT 15.675000 19.580000 15.875000 19.780000 ;
        RECT 15.675000 20.010000 15.875000 20.210000 ;
        RECT 15.675000 20.440000 15.875000 20.640000 ;
        RECT 15.675000 20.870000 15.875000 21.070000 ;
        RECT 15.675000 21.300000 15.875000 21.500000 ;
        RECT 15.675000 21.730000 15.875000 21.930000 ;
        RECT 15.675000 22.160000 15.875000 22.360000 ;
        RECT 15.695000 83.055000 15.895000 83.255000 ;
        RECT 15.695000 83.455000 15.895000 83.655000 ;
        RECT 15.695000 83.855000 15.895000 84.055000 ;
        RECT 15.695000 84.255000 15.895000 84.455000 ;
        RECT 15.695000 84.655000 15.895000 84.855000 ;
        RECT 15.695000 85.055000 15.895000 85.255000 ;
        RECT 15.695000 85.455000 15.895000 85.655000 ;
        RECT 15.695000 85.855000 15.895000 86.055000 ;
        RECT 15.695000 86.255000 15.895000 86.455000 ;
        RECT 15.695000 86.660000 15.895000 86.860000 ;
        RECT 15.695000 87.065000 15.895000 87.265000 ;
        RECT 15.695000 87.470000 15.895000 87.670000 ;
        RECT 15.695000 87.875000 15.895000 88.075000 ;
        RECT 15.980000 88.410000 16.180000 88.610000 ;
        RECT 15.980000 88.835000 16.180000 89.035000 ;
        RECT 15.980000 89.265000 16.180000 89.465000 ;
        RECT 15.980000 89.695000 16.180000 89.895000 ;
        RECT 15.980000 90.125000 16.180000 90.325000 ;
        RECT 15.980000 90.555000 16.180000 90.755000 ;
        RECT 16.045000 68.125000 16.245000 68.325000 ;
        RECT 16.045000 68.535000 16.245000 68.735000 ;
        RECT 16.045000 68.945000 16.245000 69.145000 ;
        RECT 16.045000 69.355000 16.245000 69.555000 ;
        RECT 16.045000 69.765000 16.245000 69.965000 ;
        RECT 16.045000 70.175000 16.245000 70.375000 ;
        RECT 16.045000 70.585000 16.245000 70.785000 ;
        RECT 16.045000 70.995000 16.245000 71.195000 ;
        RECT 16.045000 71.405000 16.245000 71.605000 ;
        RECT 16.045000 71.815000 16.245000 72.015000 ;
        RECT 16.045000 72.225000 16.245000 72.425000 ;
        RECT 16.045000 72.635000 16.245000 72.835000 ;
        RECT 16.045000 73.045000 16.245000 73.245000 ;
        RECT 16.045000 73.450000 16.245000 73.650000 ;
        RECT 16.045000 73.855000 16.245000 74.055000 ;
        RECT 16.045000 74.260000 16.245000 74.460000 ;
        RECT 16.045000 74.665000 16.245000 74.865000 ;
        RECT 16.045000 75.070000 16.245000 75.270000 ;
        RECT 16.045000 75.475000 16.245000 75.675000 ;
        RECT 16.045000 75.880000 16.245000 76.080000 ;
        RECT 16.045000 76.285000 16.245000 76.485000 ;
        RECT 16.045000 76.690000 16.245000 76.890000 ;
        RECT 16.045000 77.095000 16.245000 77.295000 ;
        RECT 16.045000 77.500000 16.245000 77.700000 ;
        RECT 16.045000 77.905000 16.245000 78.105000 ;
        RECT 16.045000 78.310000 16.245000 78.510000 ;
        RECT 16.045000 78.715000 16.245000 78.915000 ;
        RECT 16.045000 79.120000 16.245000 79.320000 ;
        RECT 16.045000 79.525000 16.245000 79.725000 ;
        RECT 16.045000 79.930000 16.245000 80.130000 ;
        RECT 16.045000 80.335000 16.245000 80.535000 ;
        RECT 16.045000 80.740000 16.245000 80.940000 ;
        RECT 16.045000 81.145000 16.245000 81.345000 ;
        RECT 16.045000 81.550000 16.245000 81.750000 ;
        RECT 16.045000 81.955000 16.245000 82.155000 ;
        RECT 16.045000 82.360000 16.245000 82.560000 ;
        RECT 16.080000 17.860000 16.280000 18.060000 ;
        RECT 16.080000 18.290000 16.280000 18.490000 ;
        RECT 16.080000 18.720000 16.280000 18.920000 ;
        RECT 16.080000 19.150000 16.280000 19.350000 ;
        RECT 16.080000 19.580000 16.280000 19.780000 ;
        RECT 16.080000 20.010000 16.280000 20.210000 ;
        RECT 16.080000 20.440000 16.280000 20.640000 ;
        RECT 16.080000 20.870000 16.280000 21.070000 ;
        RECT 16.080000 21.300000 16.280000 21.500000 ;
        RECT 16.080000 21.730000 16.280000 21.930000 ;
        RECT 16.080000 22.160000 16.280000 22.360000 ;
        RECT 16.105000 83.055000 16.305000 83.255000 ;
        RECT 16.105000 83.455000 16.305000 83.655000 ;
        RECT 16.105000 83.855000 16.305000 84.055000 ;
        RECT 16.105000 84.255000 16.305000 84.455000 ;
        RECT 16.105000 84.655000 16.305000 84.855000 ;
        RECT 16.105000 85.055000 16.305000 85.255000 ;
        RECT 16.105000 85.455000 16.305000 85.655000 ;
        RECT 16.105000 85.855000 16.305000 86.055000 ;
        RECT 16.105000 86.255000 16.305000 86.455000 ;
        RECT 16.105000 86.660000 16.305000 86.860000 ;
        RECT 16.105000 87.065000 16.305000 87.265000 ;
        RECT 16.105000 87.470000 16.305000 87.670000 ;
        RECT 16.105000 87.875000 16.305000 88.075000 ;
        RECT 16.445000 68.125000 16.645000 68.325000 ;
        RECT 16.445000 68.535000 16.645000 68.735000 ;
        RECT 16.445000 68.945000 16.645000 69.145000 ;
        RECT 16.445000 69.355000 16.645000 69.555000 ;
        RECT 16.445000 69.765000 16.645000 69.965000 ;
        RECT 16.445000 70.175000 16.645000 70.375000 ;
        RECT 16.445000 70.585000 16.645000 70.785000 ;
        RECT 16.445000 70.995000 16.645000 71.195000 ;
        RECT 16.445000 71.405000 16.645000 71.605000 ;
        RECT 16.445000 71.815000 16.645000 72.015000 ;
        RECT 16.445000 72.225000 16.645000 72.425000 ;
        RECT 16.445000 72.635000 16.645000 72.835000 ;
        RECT 16.445000 73.045000 16.645000 73.245000 ;
        RECT 16.445000 73.450000 16.645000 73.650000 ;
        RECT 16.445000 73.855000 16.645000 74.055000 ;
        RECT 16.445000 74.260000 16.645000 74.460000 ;
        RECT 16.445000 74.665000 16.645000 74.865000 ;
        RECT 16.445000 75.070000 16.645000 75.270000 ;
        RECT 16.445000 75.475000 16.645000 75.675000 ;
        RECT 16.445000 75.880000 16.645000 76.080000 ;
        RECT 16.445000 76.285000 16.645000 76.485000 ;
        RECT 16.445000 76.690000 16.645000 76.890000 ;
        RECT 16.445000 77.095000 16.645000 77.295000 ;
        RECT 16.445000 77.500000 16.645000 77.700000 ;
        RECT 16.445000 77.905000 16.645000 78.105000 ;
        RECT 16.445000 78.310000 16.645000 78.510000 ;
        RECT 16.445000 78.715000 16.645000 78.915000 ;
        RECT 16.445000 79.120000 16.645000 79.320000 ;
        RECT 16.445000 79.525000 16.645000 79.725000 ;
        RECT 16.445000 79.930000 16.645000 80.130000 ;
        RECT 16.445000 80.335000 16.645000 80.535000 ;
        RECT 16.445000 80.740000 16.645000 80.940000 ;
        RECT 16.445000 81.145000 16.645000 81.345000 ;
        RECT 16.445000 81.550000 16.645000 81.750000 ;
        RECT 16.445000 81.955000 16.645000 82.155000 ;
        RECT 16.445000 82.360000 16.645000 82.560000 ;
        RECT 16.480000 88.430000 16.680000 88.630000 ;
        RECT 16.480000 88.845000 16.680000 89.045000 ;
        RECT 16.480000 89.265000 16.680000 89.465000 ;
        RECT 16.485000 17.860000 16.685000 18.060000 ;
        RECT 16.485000 18.290000 16.685000 18.490000 ;
        RECT 16.485000 18.720000 16.685000 18.920000 ;
        RECT 16.485000 19.150000 16.685000 19.350000 ;
        RECT 16.485000 19.580000 16.685000 19.780000 ;
        RECT 16.485000 20.010000 16.685000 20.210000 ;
        RECT 16.485000 20.440000 16.685000 20.640000 ;
        RECT 16.485000 20.870000 16.685000 21.070000 ;
        RECT 16.485000 21.300000 16.685000 21.500000 ;
        RECT 16.485000 21.730000 16.685000 21.930000 ;
        RECT 16.485000 22.160000 16.685000 22.360000 ;
        RECT 16.515000 83.055000 16.715000 83.255000 ;
        RECT 16.515000 83.455000 16.715000 83.655000 ;
        RECT 16.515000 83.855000 16.715000 84.055000 ;
        RECT 16.515000 84.255000 16.715000 84.455000 ;
        RECT 16.515000 84.655000 16.715000 84.855000 ;
        RECT 16.515000 85.055000 16.715000 85.255000 ;
        RECT 16.515000 85.455000 16.715000 85.655000 ;
        RECT 16.515000 85.855000 16.715000 86.055000 ;
        RECT 16.515000 86.255000 16.715000 86.455000 ;
        RECT 16.515000 86.660000 16.715000 86.860000 ;
        RECT 16.515000 87.065000 16.715000 87.265000 ;
        RECT 16.515000 87.470000 16.715000 87.670000 ;
        RECT 16.515000 87.875000 16.715000 88.075000 ;
        RECT 16.845000 68.125000 17.045000 68.325000 ;
        RECT 16.845000 68.535000 17.045000 68.735000 ;
        RECT 16.845000 68.945000 17.045000 69.145000 ;
        RECT 16.845000 69.355000 17.045000 69.555000 ;
        RECT 16.845000 69.765000 17.045000 69.965000 ;
        RECT 16.845000 70.175000 17.045000 70.375000 ;
        RECT 16.845000 70.585000 17.045000 70.785000 ;
        RECT 16.845000 70.995000 17.045000 71.195000 ;
        RECT 16.845000 71.405000 17.045000 71.605000 ;
        RECT 16.845000 71.815000 17.045000 72.015000 ;
        RECT 16.845000 72.225000 17.045000 72.425000 ;
        RECT 16.845000 72.635000 17.045000 72.835000 ;
        RECT 16.845000 73.045000 17.045000 73.245000 ;
        RECT 16.845000 73.450000 17.045000 73.650000 ;
        RECT 16.845000 73.855000 17.045000 74.055000 ;
        RECT 16.845000 74.260000 17.045000 74.460000 ;
        RECT 16.845000 74.665000 17.045000 74.865000 ;
        RECT 16.845000 75.070000 17.045000 75.270000 ;
        RECT 16.845000 75.475000 17.045000 75.675000 ;
        RECT 16.845000 75.880000 17.045000 76.080000 ;
        RECT 16.845000 76.285000 17.045000 76.485000 ;
        RECT 16.845000 76.690000 17.045000 76.890000 ;
        RECT 16.845000 77.095000 17.045000 77.295000 ;
        RECT 16.845000 77.500000 17.045000 77.700000 ;
        RECT 16.845000 77.905000 17.045000 78.105000 ;
        RECT 16.845000 78.310000 17.045000 78.510000 ;
        RECT 16.845000 78.715000 17.045000 78.915000 ;
        RECT 16.845000 79.120000 17.045000 79.320000 ;
        RECT 16.845000 79.525000 17.045000 79.725000 ;
        RECT 16.845000 79.930000 17.045000 80.130000 ;
        RECT 16.845000 80.335000 17.045000 80.535000 ;
        RECT 16.845000 80.740000 17.045000 80.940000 ;
        RECT 16.845000 81.145000 17.045000 81.345000 ;
        RECT 16.845000 81.550000 17.045000 81.750000 ;
        RECT 16.845000 81.955000 17.045000 82.155000 ;
        RECT 16.845000 82.360000 17.045000 82.560000 ;
        RECT 16.890000 17.860000 17.090000 18.060000 ;
        RECT 16.890000 18.290000 17.090000 18.490000 ;
        RECT 16.890000 18.720000 17.090000 18.920000 ;
        RECT 16.890000 19.150000 17.090000 19.350000 ;
        RECT 16.890000 19.580000 17.090000 19.780000 ;
        RECT 16.890000 20.010000 17.090000 20.210000 ;
        RECT 16.890000 20.440000 17.090000 20.640000 ;
        RECT 16.890000 20.870000 17.090000 21.070000 ;
        RECT 16.890000 21.300000 17.090000 21.500000 ;
        RECT 16.890000 21.730000 17.090000 21.930000 ;
        RECT 16.890000 22.160000 17.090000 22.360000 ;
        RECT 16.925000 83.055000 17.125000 83.255000 ;
        RECT 16.925000 83.455000 17.125000 83.655000 ;
        RECT 16.925000 83.855000 17.125000 84.055000 ;
        RECT 16.925000 84.255000 17.125000 84.455000 ;
        RECT 16.925000 84.655000 17.125000 84.855000 ;
        RECT 16.925000 85.055000 17.125000 85.255000 ;
        RECT 16.925000 85.455000 17.125000 85.655000 ;
        RECT 16.925000 85.855000 17.125000 86.055000 ;
        RECT 16.925000 86.255000 17.125000 86.455000 ;
        RECT 16.925000 86.660000 17.125000 86.860000 ;
        RECT 16.925000 87.065000 17.125000 87.265000 ;
        RECT 16.925000 87.470000 17.125000 87.670000 ;
        RECT 16.925000 87.875000 17.125000 88.075000 ;
        RECT 17.245000 68.125000 17.445000 68.325000 ;
        RECT 17.245000 68.535000 17.445000 68.735000 ;
        RECT 17.245000 68.945000 17.445000 69.145000 ;
        RECT 17.245000 69.355000 17.445000 69.555000 ;
        RECT 17.245000 69.765000 17.445000 69.965000 ;
        RECT 17.245000 70.175000 17.445000 70.375000 ;
        RECT 17.245000 70.585000 17.445000 70.785000 ;
        RECT 17.245000 70.995000 17.445000 71.195000 ;
        RECT 17.245000 71.405000 17.445000 71.605000 ;
        RECT 17.245000 71.815000 17.445000 72.015000 ;
        RECT 17.245000 72.225000 17.445000 72.425000 ;
        RECT 17.245000 72.635000 17.445000 72.835000 ;
        RECT 17.245000 73.045000 17.445000 73.245000 ;
        RECT 17.245000 73.450000 17.445000 73.650000 ;
        RECT 17.245000 73.855000 17.445000 74.055000 ;
        RECT 17.245000 74.260000 17.445000 74.460000 ;
        RECT 17.245000 74.665000 17.445000 74.865000 ;
        RECT 17.245000 75.070000 17.445000 75.270000 ;
        RECT 17.245000 75.475000 17.445000 75.675000 ;
        RECT 17.245000 75.880000 17.445000 76.080000 ;
        RECT 17.245000 76.285000 17.445000 76.485000 ;
        RECT 17.245000 76.690000 17.445000 76.890000 ;
        RECT 17.245000 77.095000 17.445000 77.295000 ;
        RECT 17.245000 77.500000 17.445000 77.700000 ;
        RECT 17.245000 77.905000 17.445000 78.105000 ;
        RECT 17.245000 78.310000 17.445000 78.510000 ;
        RECT 17.245000 78.715000 17.445000 78.915000 ;
        RECT 17.245000 79.120000 17.445000 79.320000 ;
        RECT 17.245000 79.525000 17.445000 79.725000 ;
        RECT 17.245000 79.930000 17.445000 80.130000 ;
        RECT 17.245000 80.335000 17.445000 80.535000 ;
        RECT 17.245000 80.740000 17.445000 80.940000 ;
        RECT 17.245000 81.145000 17.445000 81.345000 ;
        RECT 17.245000 81.550000 17.445000 81.750000 ;
        RECT 17.245000 81.955000 17.445000 82.155000 ;
        RECT 17.245000 82.360000 17.445000 82.560000 ;
        RECT 17.260000 88.430000 17.460000 88.630000 ;
        RECT 17.260000 88.845000 17.460000 89.045000 ;
        RECT 17.260000 89.265000 17.460000 89.465000 ;
        RECT 17.295000 17.860000 17.495000 18.060000 ;
        RECT 17.295000 18.290000 17.495000 18.490000 ;
        RECT 17.295000 18.720000 17.495000 18.920000 ;
        RECT 17.295000 19.150000 17.495000 19.350000 ;
        RECT 17.295000 19.580000 17.495000 19.780000 ;
        RECT 17.295000 20.010000 17.495000 20.210000 ;
        RECT 17.295000 20.440000 17.495000 20.640000 ;
        RECT 17.295000 20.870000 17.495000 21.070000 ;
        RECT 17.295000 21.300000 17.495000 21.500000 ;
        RECT 17.295000 21.730000 17.495000 21.930000 ;
        RECT 17.295000 22.160000 17.495000 22.360000 ;
        RECT 17.335000 83.055000 17.535000 83.255000 ;
        RECT 17.335000 83.455000 17.535000 83.655000 ;
        RECT 17.335000 83.855000 17.535000 84.055000 ;
        RECT 17.335000 84.255000 17.535000 84.455000 ;
        RECT 17.335000 84.655000 17.535000 84.855000 ;
        RECT 17.335000 85.055000 17.535000 85.255000 ;
        RECT 17.335000 85.455000 17.535000 85.655000 ;
        RECT 17.335000 85.855000 17.535000 86.055000 ;
        RECT 17.335000 86.255000 17.535000 86.455000 ;
        RECT 17.335000 86.660000 17.535000 86.860000 ;
        RECT 17.335000 87.065000 17.535000 87.265000 ;
        RECT 17.335000 87.470000 17.535000 87.670000 ;
        RECT 17.335000 87.875000 17.535000 88.075000 ;
        RECT 17.645000 68.125000 17.845000 68.325000 ;
        RECT 17.645000 68.535000 17.845000 68.735000 ;
        RECT 17.645000 68.945000 17.845000 69.145000 ;
        RECT 17.645000 69.355000 17.845000 69.555000 ;
        RECT 17.645000 69.765000 17.845000 69.965000 ;
        RECT 17.645000 70.175000 17.845000 70.375000 ;
        RECT 17.645000 70.585000 17.845000 70.785000 ;
        RECT 17.645000 70.995000 17.845000 71.195000 ;
        RECT 17.645000 71.405000 17.845000 71.605000 ;
        RECT 17.645000 71.815000 17.845000 72.015000 ;
        RECT 17.645000 72.225000 17.845000 72.425000 ;
        RECT 17.645000 72.635000 17.845000 72.835000 ;
        RECT 17.645000 73.045000 17.845000 73.245000 ;
        RECT 17.645000 73.450000 17.845000 73.650000 ;
        RECT 17.645000 73.855000 17.845000 74.055000 ;
        RECT 17.645000 74.260000 17.845000 74.460000 ;
        RECT 17.645000 74.665000 17.845000 74.865000 ;
        RECT 17.645000 75.070000 17.845000 75.270000 ;
        RECT 17.645000 75.475000 17.845000 75.675000 ;
        RECT 17.645000 75.880000 17.845000 76.080000 ;
        RECT 17.645000 76.285000 17.845000 76.485000 ;
        RECT 17.645000 76.690000 17.845000 76.890000 ;
        RECT 17.645000 77.095000 17.845000 77.295000 ;
        RECT 17.645000 77.500000 17.845000 77.700000 ;
        RECT 17.645000 77.905000 17.845000 78.105000 ;
        RECT 17.645000 78.310000 17.845000 78.510000 ;
        RECT 17.645000 78.715000 17.845000 78.915000 ;
        RECT 17.645000 79.120000 17.845000 79.320000 ;
        RECT 17.645000 79.525000 17.845000 79.725000 ;
        RECT 17.645000 79.930000 17.845000 80.130000 ;
        RECT 17.645000 80.335000 17.845000 80.535000 ;
        RECT 17.645000 80.740000 17.845000 80.940000 ;
        RECT 17.645000 81.145000 17.845000 81.345000 ;
        RECT 17.645000 81.550000 17.845000 81.750000 ;
        RECT 17.645000 81.955000 17.845000 82.155000 ;
        RECT 17.645000 82.360000 17.845000 82.560000 ;
        RECT 17.700000 17.860000 17.900000 18.060000 ;
        RECT 17.700000 18.290000 17.900000 18.490000 ;
        RECT 17.700000 18.720000 17.900000 18.920000 ;
        RECT 17.700000 19.150000 17.900000 19.350000 ;
        RECT 17.700000 19.580000 17.900000 19.780000 ;
        RECT 17.700000 20.010000 17.900000 20.210000 ;
        RECT 17.700000 20.440000 17.900000 20.640000 ;
        RECT 17.700000 20.870000 17.900000 21.070000 ;
        RECT 17.700000 21.300000 17.900000 21.500000 ;
        RECT 17.700000 21.730000 17.900000 21.930000 ;
        RECT 17.700000 22.160000 17.900000 22.360000 ;
        RECT 17.745000 83.055000 17.945000 83.255000 ;
        RECT 17.745000 83.455000 17.945000 83.655000 ;
        RECT 17.745000 83.855000 17.945000 84.055000 ;
        RECT 17.745000 84.255000 17.945000 84.455000 ;
        RECT 17.745000 84.655000 17.945000 84.855000 ;
        RECT 17.745000 85.055000 17.945000 85.255000 ;
        RECT 17.745000 85.455000 17.945000 85.655000 ;
        RECT 17.745000 85.855000 17.945000 86.055000 ;
        RECT 17.745000 86.255000 17.945000 86.455000 ;
        RECT 17.745000 86.660000 17.945000 86.860000 ;
        RECT 17.745000 87.065000 17.945000 87.265000 ;
        RECT 17.745000 87.470000 17.945000 87.670000 ;
        RECT 17.745000 87.875000 17.945000 88.075000 ;
        RECT 18.045000 68.125000 18.245000 68.325000 ;
        RECT 18.045000 68.535000 18.245000 68.735000 ;
        RECT 18.045000 68.945000 18.245000 69.145000 ;
        RECT 18.045000 69.355000 18.245000 69.555000 ;
        RECT 18.045000 69.765000 18.245000 69.965000 ;
        RECT 18.045000 70.175000 18.245000 70.375000 ;
        RECT 18.045000 70.585000 18.245000 70.785000 ;
        RECT 18.045000 70.995000 18.245000 71.195000 ;
        RECT 18.045000 71.405000 18.245000 71.605000 ;
        RECT 18.045000 71.815000 18.245000 72.015000 ;
        RECT 18.045000 72.225000 18.245000 72.425000 ;
        RECT 18.045000 72.635000 18.245000 72.835000 ;
        RECT 18.045000 73.045000 18.245000 73.245000 ;
        RECT 18.045000 73.450000 18.245000 73.650000 ;
        RECT 18.045000 73.855000 18.245000 74.055000 ;
        RECT 18.045000 74.260000 18.245000 74.460000 ;
        RECT 18.045000 74.665000 18.245000 74.865000 ;
        RECT 18.045000 75.070000 18.245000 75.270000 ;
        RECT 18.045000 75.475000 18.245000 75.675000 ;
        RECT 18.045000 75.880000 18.245000 76.080000 ;
        RECT 18.045000 76.285000 18.245000 76.485000 ;
        RECT 18.045000 76.690000 18.245000 76.890000 ;
        RECT 18.045000 77.095000 18.245000 77.295000 ;
        RECT 18.045000 77.500000 18.245000 77.700000 ;
        RECT 18.045000 77.905000 18.245000 78.105000 ;
        RECT 18.045000 78.310000 18.245000 78.510000 ;
        RECT 18.045000 78.715000 18.245000 78.915000 ;
        RECT 18.045000 79.120000 18.245000 79.320000 ;
        RECT 18.045000 79.525000 18.245000 79.725000 ;
        RECT 18.045000 79.930000 18.245000 80.130000 ;
        RECT 18.045000 80.335000 18.245000 80.535000 ;
        RECT 18.045000 80.740000 18.245000 80.940000 ;
        RECT 18.045000 81.145000 18.245000 81.345000 ;
        RECT 18.045000 81.550000 18.245000 81.750000 ;
        RECT 18.045000 81.955000 18.245000 82.155000 ;
        RECT 18.045000 82.360000 18.245000 82.560000 ;
        RECT 18.105000 17.860000 18.305000 18.060000 ;
        RECT 18.105000 18.290000 18.305000 18.490000 ;
        RECT 18.105000 18.720000 18.305000 18.920000 ;
        RECT 18.105000 19.150000 18.305000 19.350000 ;
        RECT 18.105000 19.580000 18.305000 19.780000 ;
        RECT 18.105000 20.010000 18.305000 20.210000 ;
        RECT 18.105000 20.440000 18.305000 20.640000 ;
        RECT 18.105000 20.870000 18.305000 21.070000 ;
        RECT 18.105000 21.300000 18.305000 21.500000 ;
        RECT 18.105000 21.730000 18.305000 21.930000 ;
        RECT 18.105000 22.160000 18.305000 22.360000 ;
        RECT 18.155000 83.055000 18.355000 83.255000 ;
        RECT 18.155000 83.455000 18.355000 83.655000 ;
        RECT 18.155000 83.855000 18.355000 84.055000 ;
        RECT 18.155000 84.255000 18.355000 84.455000 ;
        RECT 18.155000 84.655000 18.355000 84.855000 ;
        RECT 18.155000 85.055000 18.355000 85.255000 ;
        RECT 18.155000 85.455000 18.355000 85.655000 ;
        RECT 18.155000 85.855000 18.355000 86.055000 ;
        RECT 18.155000 86.255000 18.355000 86.455000 ;
        RECT 18.155000 86.660000 18.355000 86.860000 ;
        RECT 18.155000 87.065000 18.355000 87.265000 ;
        RECT 18.155000 87.470000 18.355000 87.670000 ;
        RECT 18.155000 87.875000 18.355000 88.075000 ;
        RECT 18.445000 68.125000 18.645000 68.325000 ;
        RECT 18.445000 68.535000 18.645000 68.735000 ;
        RECT 18.445000 68.945000 18.645000 69.145000 ;
        RECT 18.445000 69.355000 18.645000 69.555000 ;
        RECT 18.445000 69.765000 18.645000 69.965000 ;
        RECT 18.445000 70.175000 18.645000 70.375000 ;
        RECT 18.445000 70.585000 18.645000 70.785000 ;
        RECT 18.445000 70.995000 18.645000 71.195000 ;
        RECT 18.445000 71.405000 18.645000 71.605000 ;
        RECT 18.445000 71.815000 18.645000 72.015000 ;
        RECT 18.445000 72.225000 18.645000 72.425000 ;
        RECT 18.445000 72.635000 18.645000 72.835000 ;
        RECT 18.445000 73.045000 18.645000 73.245000 ;
        RECT 18.445000 73.450000 18.645000 73.650000 ;
        RECT 18.445000 73.855000 18.645000 74.055000 ;
        RECT 18.445000 74.260000 18.645000 74.460000 ;
        RECT 18.445000 74.665000 18.645000 74.865000 ;
        RECT 18.445000 75.070000 18.645000 75.270000 ;
        RECT 18.445000 75.475000 18.645000 75.675000 ;
        RECT 18.445000 75.880000 18.645000 76.080000 ;
        RECT 18.445000 76.285000 18.645000 76.485000 ;
        RECT 18.445000 76.690000 18.645000 76.890000 ;
        RECT 18.445000 77.095000 18.645000 77.295000 ;
        RECT 18.445000 77.500000 18.645000 77.700000 ;
        RECT 18.445000 77.905000 18.645000 78.105000 ;
        RECT 18.445000 78.310000 18.645000 78.510000 ;
        RECT 18.445000 78.715000 18.645000 78.915000 ;
        RECT 18.445000 79.120000 18.645000 79.320000 ;
        RECT 18.445000 79.525000 18.645000 79.725000 ;
        RECT 18.445000 79.930000 18.645000 80.130000 ;
        RECT 18.445000 80.335000 18.645000 80.535000 ;
        RECT 18.445000 80.740000 18.645000 80.940000 ;
        RECT 18.445000 81.145000 18.645000 81.345000 ;
        RECT 18.445000 81.550000 18.645000 81.750000 ;
        RECT 18.445000 81.955000 18.645000 82.155000 ;
        RECT 18.445000 82.360000 18.645000 82.560000 ;
        RECT 18.510000 17.860000 18.710000 18.060000 ;
        RECT 18.510000 18.290000 18.710000 18.490000 ;
        RECT 18.510000 18.720000 18.710000 18.920000 ;
        RECT 18.510000 19.150000 18.710000 19.350000 ;
        RECT 18.510000 19.580000 18.710000 19.780000 ;
        RECT 18.510000 20.010000 18.710000 20.210000 ;
        RECT 18.510000 20.440000 18.710000 20.640000 ;
        RECT 18.510000 20.870000 18.710000 21.070000 ;
        RECT 18.510000 21.300000 18.710000 21.500000 ;
        RECT 18.510000 21.730000 18.710000 21.930000 ;
        RECT 18.510000 22.160000 18.710000 22.360000 ;
        RECT 18.565000 83.055000 18.765000 83.255000 ;
        RECT 18.565000 83.455000 18.765000 83.655000 ;
        RECT 18.565000 83.855000 18.765000 84.055000 ;
        RECT 18.565000 84.255000 18.765000 84.455000 ;
        RECT 18.565000 84.655000 18.765000 84.855000 ;
        RECT 18.565000 85.055000 18.765000 85.255000 ;
        RECT 18.565000 85.455000 18.765000 85.655000 ;
        RECT 18.565000 85.855000 18.765000 86.055000 ;
        RECT 18.565000 86.255000 18.765000 86.455000 ;
        RECT 18.565000 86.660000 18.765000 86.860000 ;
        RECT 18.565000 87.065000 18.765000 87.265000 ;
        RECT 18.565000 87.470000 18.765000 87.670000 ;
        RECT 18.565000 87.875000 18.765000 88.075000 ;
        RECT 18.845000 68.125000 19.045000 68.325000 ;
        RECT 18.845000 68.535000 19.045000 68.735000 ;
        RECT 18.845000 68.945000 19.045000 69.145000 ;
        RECT 18.845000 69.355000 19.045000 69.555000 ;
        RECT 18.845000 69.765000 19.045000 69.965000 ;
        RECT 18.845000 70.175000 19.045000 70.375000 ;
        RECT 18.845000 70.585000 19.045000 70.785000 ;
        RECT 18.845000 70.995000 19.045000 71.195000 ;
        RECT 18.845000 71.405000 19.045000 71.605000 ;
        RECT 18.845000 71.815000 19.045000 72.015000 ;
        RECT 18.845000 72.225000 19.045000 72.425000 ;
        RECT 18.845000 72.635000 19.045000 72.835000 ;
        RECT 18.845000 73.045000 19.045000 73.245000 ;
        RECT 18.845000 73.450000 19.045000 73.650000 ;
        RECT 18.845000 73.855000 19.045000 74.055000 ;
        RECT 18.845000 74.260000 19.045000 74.460000 ;
        RECT 18.845000 74.665000 19.045000 74.865000 ;
        RECT 18.845000 75.070000 19.045000 75.270000 ;
        RECT 18.845000 75.475000 19.045000 75.675000 ;
        RECT 18.845000 75.880000 19.045000 76.080000 ;
        RECT 18.845000 76.285000 19.045000 76.485000 ;
        RECT 18.845000 76.690000 19.045000 76.890000 ;
        RECT 18.845000 77.095000 19.045000 77.295000 ;
        RECT 18.845000 77.500000 19.045000 77.700000 ;
        RECT 18.845000 77.905000 19.045000 78.105000 ;
        RECT 18.845000 78.310000 19.045000 78.510000 ;
        RECT 18.845000 78.715000 19.045000 78.915000 ;
        RECT 18.845000 79.120000 19.045000 79.320000 ;
        RECT 18.845000 79.525000 19.045000 79.725000 ;
        RECT 18.845000 79.930000 19.045000 80.130000 ;
        RECT 18.845000 80.335000 19.045000 80.535000 ;
        RECT 18.845000 80.740000 19.045000 80.940000 ;
        RECT 18.845000 81.145000 19.045000 81.345000 ;
        RECT 18.845000 81.550000 19.045000 81.750000 ;
        RECT 18.845000 81.955000 19.045000 82.155000 ;
        RECT 18.845000 82.360000 19.045000 82.560000 ;
        RECT 18.915000 17.860000 19.115000 18.060000 ;
        RECT 18.915000 18.290000 19.115000 18.490000 ;
        RECT 18.915000 18.720000 19.115000 18.920000 ;
        RECT 18.915000 19.150000 19.115000 19.350000 ;
        RECT 18.915000 19.580000 19.115000 19.780000 ;
        RECT 18.915000 20.010000 19.115000 20.210000 ;
        RECT 18.915000 20.440000 19.115000 20.640000 ;
        RECT 18.915000 20.870000 19.115000 21.070000 ;
        RECT 18.915000 21.300000 19.115000 21.500000 ;
        RECT 18.915000 21.730000 19.115000 21.930000 ;
        RECT 18.915000 22.160000 19.115000 22.360000 ;
        RECT 19.060000 85.875000 19.260000 86.075000 ;
        RECT 19.060000 86.310000 19.260000 86.510000 ;
        RECT 19.060000 86.750000 19.260000 86.950000 ;
        RECT 19.245000 68.125000 19.445000 68.325000 ;
        RECT 19.245000 68.535000 19.445000 68.735000 ;
        RECT 19.245000 68.945000 19.445000 69.145000 ;
        RECT 19.245000 69.355000 19.445000 69.555000 ;
        RECT 19.245000 69.765000 19.445000 69.965000 ;
        RECT 19.245000 70.175000 19.445000 70.375000 ;
        RECT 19.245000 70.585000 19.445000 70.785000 ;
        RECT 19.245000 70.995000 19.445000 71.195000 ;
        RECT 19.245000 71.405000 19.445000 71.605000 ;
        RECT 19.245000 71.815000 19.445000 72.015000 ;
        RECT 19.245000 72.225000 19.445000 72.425000 ;
        RECT 19.245000 72.635000 19.445000 72.835000 ;
        RECT 19.245000 73.045000 19.445000 73.245000 ;
        RECT 19.245000 73.450000 19.445000 73.650000 ;
        RECT 19.245000 73.855000 19.445000 74.055000 ;
        RECT 19.245000 74.260000 19.445000 74.460000 ;
        RECT 19.245000 74.665000 19.445000 74.865000 ;
        RECT 19.245000 75.070000 19.445000 75.270000 ;
        RECT 19.245000 75.475000 19.445000 75.675000 ;
        RECT 19.245000 75.880000 19.445000 76.080000 ;
        RECT 19.245000 76.285000 19.445000 76.485000 ;
        RECT 19.245000 76.690000 19.445000 76.890000 ;
        RECT 19.245000 77.095000 19.445000 77.295000 ;
        RECT 19.245000 77.500000 19.445000 77.700000 ;
        RECT 19.245000 77.905000 19.445000 78.105000 ;
        RECT 19.245000 78.310000 19.445000 78.510000 ;
        RECT 19.245000 78.715000 19.445000 78.915000 ;
        RECT 19.245000 79.120000 19.445000 79.320000 ;
        RECT 19.245000 79.525000 19.445000 79.725000 ;
        RECT 19.245000 79.930000 19.445000 80.130000 ;
        RECT 19.245000 80.335000 19.445000 80.535000 ;
        RECT 19.245000 80.740000 19.445000 80.940000 ;
        RECT 19.245000 81.145000 19.445000 81.345000 ;
        RECT 19.245000 81.550000 19.445000 81.750000 ;
        RECT 19.245000 81.955000 19.445000 82.155000 ;
        RECT 19.245000 82.360000 19.445000 82.560000 ;
        RECT 19.250000 83.010000 19.450000 83.210000 ;
        RECT 19.250000 83.470000 19.450000 83.670000 ;
        RECT 19.250000 83.930000 19.450000 84.130000 ;
        RECT 19.250000 84.395000 19.450000 84.595000 ;
        RECT 19.250000 84.860000 19.450000 85.060000 ;
        RECT 19.250000 85.325000 19.450000 85.525000 ;
        RECT 19.320000 17.860000 19.520000 18.060000 ;
        RECT 19.320000 18.290000 19.520000 18.490000 ;
        RECT 19.320000 18.720000 19.520000 18.920000 ;
        RECT 19.320000 19.150000 19.520000 19.350000 ;
        RECT 19.320000 19.580000 19.520000 19.780000 ;
        RECT 19.320000 20.010000 19.520000 20.210000 ;
        RECT 19.320000 20.440000 19.520000 20.640000 ;
        RECT 19.320000 20.870000 19.520000 21.070000 ;
        RECT 19.320000 21.300000 19.520000 21.500000 ;
        RECT 19.320000 21.730000 19.520000 21.930000 ;
        RECT 19.320000 22.160000 19.520000 22.360000 ;
        RECT 19.645000 68.125000 19.845000 68.325000 ;
        RECT 19.645000 68.535000 19.845000 68.735000 ;
        RECT 19.645000 68.945000 19.845000 69.145000 ;
        RECT 19.645000 69.355000 19.845000 69.555000 ;
        RECT 19.645000 69.765000 19.845000 69.965000 ;
        RECT 19.645000 70.175000 19.845000 70.375000 ;
        RECT 19.645000 70.585000 19.845000 70.785000 ;
        RECT 19.645000 70.995000 19.845000 71.195000 ;
        RECT 19.645000 71.405000 19.845000 71.605000 ;
        RECT 19.645000 71.815000 19.845000 72.015000 ;
        RECT 19.645000 72.225000 19.845000 72.425000 ;
        RECT 19.645000 72.635000 19.845000 72.835000 ;
        RECT 19.645000 73.045000 19.845000 73.245000 ;
        RECT 19.645000 73.450000 19.845000 73.650000 ;
        RECT 19.645000 73.855000 19.845000 74.055000 ;
        RECT 19.645000 74.260000 19.845000 74.460000 ;
        RECT 19.645000 74.665000 19.845000 74.865000 ;
        RECT 19.645000 75.070000 19.845000 75.270000 ;
        RECT 19.645000 75.475000 19.845000 75.675000 ;
        RECT 19.645000 75.880000 19.845000 76.080000 ;
        RECT 19.645000 76.285000 19.845000 76.485000 ;
        RECT 19.645000 76.690000 19.845000 76.890000 ;
        RECT 19.645000 77.095000 19.845000 77.295000 ;
        RECT 19.645000 77.500000 19.845000 77.700000 ;
        RECT 19.645000 77.905000 19.845000 78.105000 ;
        RECT 19.645000 78.310000 19.845000 78.510000 ;
        RECT 19.645000 78.715000 19.845000 78.915000 ;
        RECT 19.645000 79.120000 19.845000 79.320000 ;
        RECT 19.645000 79.525000 19.845000 79.725000 ;
        RECT 19.645000 79.930000 19.845000 80.130000 ;
        RECT 19.645000 80.335000 19.845000 80.535000 ;
        RECT 19.645000 80.740000 19.845000 80.940000 ;
        RECT 19.645000 81.145000 19.845000 81.345000 ;
        RECT 19.645000 81.550000 19.845000 81.750000 ;
        RECT 19.645000 81.955000 19.845000 82.155000 ;
        RECT 19.645000 82.360000 19.845000 82.560000 ;
        RECT 19.725000 17.860000 19.925000 18.060000 ;
        RECT 19.725000 18.290000 19.925000 18.490000 ;
        RECT 19.725000 18.720000 19.925000 18.920000 ;
        RECT 19.725000 19.150000 19.925000 19.350000 ;
        RECT 19.725000 19.580000 19.925000 19.780000 ;
        RECT 19.725000 20.010000 19.925000 20.210000 ;
        RECT 19.725000 20.440000 19.925000 20.640000 ;
        RECT 19.725000 20.870000 19.925000 21.070000 ;
        RECT 19.725000 21.300000 19.925000 21.500000 ;
        RECT 19.725000 21.730000 19.925000 21.930000 ;
        RECT 19.725000 22.160000 19.925000 22.360000 ;
        RECT 19.730000 83.010000 19.930000 83.210000 ;
        RECT 19.730000 83.470000 19.930000 83.670000 ;
        RECT 19.730000 83.930000 19.930000 84.130000 ;
        RECT 19.730000 84.395000 19.930000 84.595000 ;
        RECT 19.730000 84.860000 19.930000 85.060000 ;
        RECT 19.730000 85.325000 19.930000 85.525000 ;
        RECT 19.800000 85.875000 20.000000 86.075000 ;
        RECT 19.800000 86.310000 20.000000 86.510000 ;
        RECT 19.800000 86.750000 20.000000 86.950000 ;
        RECT 20.045000 68.125000 20.245000 68.325000 ;
        RECT 20.045000 68.535000 20.245000 68.735000 ;
        RECT 20.045000 68.945000 20.245000 69.145000 ;
        RECT 20.045000 69.355000 20.245000 69.555000 ;
        RECT 20.045000 69.765000 20.245000 69.965000 ;
        RECT 20.045000 70.175000 20.245000 70.375000 ;
        RECT 20.045000 70.585000 20.245000 70.785000 ;
        RECT 20.045000 70.995000 20.245000 71.195000 ;
        RECT 20.045000 71.405000 20.245000 71.605000 ;
        RECT 20.045000 71.815000 20.245000 72.015000 ;
        RECT 20.045000 72.225000 20.245000 72.425000 ;
        RECT 20.045000 72.635000 20.245000 72.835000 ;
        RECT 20.045000 73.045000 20.245000 73.245000 ;
        RECT 20.045000 73.450000 20.245000 73.650000 ;
        RECT 20.045000 73.855000 20.245000 74.055000 ;
        RECT 20.045000 74.260000 20.245000 74.460000 ;
        RECT 20.045000 74.665000 20.245000 74.865000 ;
        RECT 20.045000 75.070000 20.245000 75.270000 ;
        RECT 20.045000 75.475000 20.245000 75.675000 ;
        RECT 20.045000 75.880000 20.245000 76.080000 ;
        RECT 20.045000 76.285000 20.245000 76.485000 ;
        RECT 20.045000 76.690000 20.245000 76.890000 ;
        RECT 20.045000 77.095000 20.245000 77.295000 ;
        RECT 20.045000 77.500000 20.245000 77.700000 ;
        RECT 20.045000 77.905000 20.245000 78.105000 ;
        RECT 20.045000 78.310000 20.245000 78.510000 ;
        RECT 20.045000 78.715000 20.245000 78.915000 ;
        RECT 20.045000 79.120000 20.245000 79.320000 ;
        RECT 20.045000 79.525000 20.245000 79.725000 ;
        RECT 20.045000 79.930000 20.245000 80.130000 ;
        RECT 20.045000 80.335000 20.245000 80.535000 ;
        RECT 20.045000 80.740000 20.245000 80.940000 ;
        RECT 20.045000 81.145000 20.245000 81.345000 ;
        RECT 20.045000 81.550000 20.245000 81.750000 ;
        RECT 20.045000 81.955000 20.245000 82.155000 ;
        RECT 20.045000 82.360000 20.245000 82.560000 ;
        RECT 20.130000 17.860000 20.330000 18.060000 ;
        RECT 20.130000 18.290000 20.330000 18.490000 ;
        RECT 20.130000 18.720000 20.330000 18.920000 ;
        RECT 20.130000 19.150000 20.330000 19.350000 ;
        RECT 20.130000 19.580000 20.330000 19.780000 ;
        RECT 20.130000 20.010000 20.330000 20.210000 ;
        RECT 20.130000 20.440000 20.330000 20.640000 ;
        RECT 20.130000 20.870000 20.330000 21.070000 ;
        RECT 20.130000 21.300000 20.330000 21.500000 ;
        RECT 20.130000 21.730000 20.330000 21.930000 ;
        RECT 20.130000 22.160000 20.330000 22.360000 ;
        RECT 20.210000 83.010000 20.410000 83.210000 ;
        RECT 20.210000 83.470000 20.410000 83.670000 ;
        RECT 20.210000 83.930000 20.410000 84.130000 ;
        RECT 20.210000 84.395000 20.410000 84.595000 ;
        RECT 20.210000 84.860000 20.410000 85.060000 ;
        RECT 20.210000 85.325000 20.410000 85.525000 ;
        RECT 20.445000 68.125000 20.645000 68.325000 ;
        RECT 20.445000 68.535000 20.645000 68.735000 ;
        RECT 20.445000 68.945000 20.645000 69.145000 ;
        RECT 20.445000 69.355000 20.645000 69.555000 ;
        RECT 20.445000 69.765000 20.645000 69.965000 ;
        RECT 20.445000 70.175000 20.645000 70.375000 ;
        RECT 20.445000 70.585000 20.645000 70.785000 ;
        RECT 20.445000 70.995000 20.645000 71.195000 ;
        RECT 20.445000 71.405000 20.645000 71.605000 ;
        RECT 20.445000 71.815000 20.645000 72.015000 ;
        RECT 20.445000 72.225000 20.645000 72.425000 ;
        RECT 20.445000 72.635000 20.645000 72.835000 ;
        RECT 20.445000 73.045000 20.645000 73.245000 ;
        RECT 20.445000 73.450000 20.645000 73.650000 ;
        RECT 20.445000 73.855000 20.645000 74.055000 ;
        RECT 20.445000 74.260000 20.645000 74.460000 ;
        RECT 20.445000 74.665000 20.645000 74.865000 ;
        RECT 20.445000 75.070000 20.645000 75.270000 ;
        RECT 20.445000 75.475000 20.645000 75.675000 ;
        RECT 20.445000 75.880000 20.645000 76.080000 ;
        RECT 20.445000 76.285000 20.645000 76.485000 ;
        RECT 20.445000 76.690000 20.645000 76.890000 ;
        RECT 20.445000 77.095000 20.645000 77.295000 ;
        RECT 20.445000 77.500000 20.645000 77.700000 ;
        RECT 20.445000 77.905000 20.645000 78.105000 ;
        RECT 20.445000 78.310000 20.645000 78.510000 ;
        RECT 20.445000 78.715000 20.645000 78.915000 ;
        RECT 20.445000 79.120000 20.645000 79.320000 ;
        RECT 20.445000 79.525000 20.645000 79.725000 ;
        RECT 20.445000 79.930000 20.645000 80.130000 ;
        RECT 20.445000 80.335000 20.645000 80.535000 ;
        RECT 20.445000 80.740000 20.645000 80.940000 ;
        RECT 20.445000 81.145000 20.645000 81.345000 ;
        RECT 20.445000 81.550000 20.645000 81.750000 ;
        RECT 20.445000 81.955000 20.645000 82.155000 ;
        RECT 20.445000 82.360000 20.645000 82.560000 ;
        RECT 20.535000 17.860000 20.735000 18.060000 ;
        RECT 20.535000 18.290000 20.735000 18.490000 ;
        RECT 20.535000 18.720000 20.735000 18.920000 ;
        RECT 20.535000 19.150000 20.735000 19.350000 ;
        RECT 20.535000 19.580000 20.735000 19.780000 ;
        RECT 20.535000 20.010000 20.735000 20.210000 ;
        RECT 20.535000 20.440000 20.735000 20.640000 ;
        RECT 20.535000 20.870000 20.735000 21.070000 ;
        RECT 20.535000 21.300000 20.735000 21.500000 ;
        RECT 20.535000 21.730000 20.735000 21.930000 ;
        RECT 20.535000 22.160000 20.735000 22.360000 ;
        RECT 20.690000 83.010000 20.890000 83.210000 ;
        RECT 20.690000 83.470000 20.890000 83.670000 ;
        RECT 20.690000 83.930000 20.890000 84.130000 ;
        RECT 20.690000 84.395000 20.890000 84.595000 ;
        RECT 20.690000 84.860000 20.890000 85.060000 ;
        RECT 20.690000 85.325000 20.890000 85.525000 ;
        RECT 20.845000 68.125000 21.045000 68.325000 ;
        RECT 20.845000 68.535000 21.045000 68.735000 ;
        RECT 20.845000 68.945000 21.045000 69.145000 ;
        RECT 20.845000 69.355000 21.045000 69.555000 ;
        RECT 20.845000 69.765000 21.045000 69.965000 ;
        RECT 20.845000 70.175000 21.045000 70.375000 ;
        RECT 20.845000 70.585000 21.045000 70.785000 ;
        RECT 20.845000 70.995000 21.045000 71.195000 ;
        RECT 20.845000 71.405000 21.045000 71.605000 ;
        RECT 20.845000 71.815000 21.045000 72.015000 ;
        RECT 20.845000 72.225000 21.045000 72.425000 ;
        RECT 20.845000 72.635000 21.045000 72.835000 ;
        RECT 20.845000 73.045000 21.045000 73.245000 ;
        RECT 20.845000 73.450000 21.045000 73.650000 ;
        RECT 20.845000 73.855000 21.045000 74.055000 ;
        RECT 20.845000 74.260000 21.045000 74.460000 ;
        RECT 20.845000 74.665000 21.045000 74.865000 ;
        RECT 20.845000 75.070000 21.045000 75.270000 ;
        RECT 20.845000 75.475000 21.045000 75.675000 ;
        RECT 20.845000 75.880000 21.045000 76.080000 ;
        RECT 20.845000 76.285000 21.045000 76.485000 ;
        RECT 20.845000 76.690000 21.045000 76.890000 ;
        RECT 20.845000 77.095000 21.045000 77.295000 ;
        RECT 20.845000 77.500000 21.045000 77.700000 ;
        RECT 20.845000 77.905000 21.045000 78.105000 ;
        RECT 20.845000 78.310000 21.045000 78.510000 ;
        RECT 20.845000 78.715000 21.045000 78.915000 ;
        RECT 20.845000 79.120000 21.045000 79.320000 ;
        RECT 20.845000 79.525000 21.045000 79.725000 ;
        RECT 20.845000 79.930000 21.045000 80.130000 ;
        RECT 20.845000 80.335000 21.045000 80.535000 ;
        RECT 20.845000 80.740000 21.045000 80.940000 ;
        RECT 20.845000 81.145000 21.045000 81.345000 ;
        RECT 20.845000 81.550000 21.045000 81.750000 ;
        RECT 20.845000 81.955000 21.045000 82.155000 ;
        RECT 20.845000 82.360000 21.045000 82.560000 ;
        RECT 20.940000 17.860000 21.140000 18.060000 ;
        RECT 20.940000 18.290000 21.140000 18.490000 ;
        RECT 20.940000 18.720000 21.140000 18.920000 ;
        RECT 20.940000 19.150000 21.140000 19.350000 ;
        RECT 20.940000 19.580000 21.140000 19.780000 ;
        RECT 20.940000 20.010000 21.140000 20.210000 ;
        RECT 20.940000 20.440000 21.140000 20.640000 ;
        RECT 20.940000 20.870000 21.140000 21.070000 ;
        RECT 20.940000 21.300000 21.140000 21.500000 ;
        RECT 20.940000 21.730000 21.140000 21.930000 ;
        RECT 20.940000 22.160000 21.140000 22.360000 ;
        RECT 21.170000 83.010000 21.370000 83.210000 ;
        RECT 21.170000 83.470000 21.370000 83.670000 ;
        RECT 21.170000 83.930000 21.370000 84.130000 ;
        RECT 21.170000 84.395000 21.370000 84.595000 ;
        RECT 21.170000 84.860000 21.370000 85.060000 ;
        RECT 21.170000 85.325000 21.370000 85.525000 ;
        RECT 21.245000 68.125000 21.445000 68.325000 ;
        RECT 21.245000 68.535000 21.445000 68.735000 ;
        RECT 21.245000 68.945000 21.445000 69.145000 ;
        RECT 21.245000 69.355000 21.445000 69.555000 ;
        RECT 21.245000 69.765000 21.445000 69.965000 ;
        RECT 21.245000 70.175000 21.445000 70.375000 ;
        RECT 21.245000 70.585000 21.445000 70.785000 ;
        RECT 21.245000 70.995000 21.445000 71.195000 ;
        RECT 21.245000 71.405000 21.445000 71.605000 ;
        RECT 21.245000 71.815000 21.445000 72.015000 ;
        RECT 21.245000 72.225000 21.445000 72.425000 ;
        RECT 21.245000 72.635000 21.445000 72.835000 ;
        RECT 21.245000 73.045000 21.445000 73.245000 ;
        RECT 21.245000 73.450000 21.445000 73.650000 ;
        RECT 21.245000 73.855000 21.445000 74.055000 ;
        RECT 21.245000 74.260000 21.445000 74.460000 ;
        RECT 21.245000 74.665000 21.445000 74.865000 ;
        RECT 21.245000 75.070000 21.445000 75.270000 ;
        RECT 21.245000 75.475000 21.445000 75.675000 ;
        RECT 21.245000 75.880000 21.445000 76.080000 ;
        RECT 21.245000 76.285000 21.445000 76.485000 ;
        RECT 21.245000 76.690000 21.445000 76.890000 ;
        RECT 21.245000 77.095000 21.445000 77.295000 ;
        RECT 21.245000 77.500000 21.445000 77.700000 ;
        RECT 21.245000 77.905000 21.445000 78.105000 ;
        RECT 21.245000 78.310000 21.445000 78.510000 ;
        RECT 21.245000 78.715000 21.445000 78.915000 ;
        RECT 21.245000 79.120000 21.445000 79.320000 ;
        RECT 21.245000 79.525000 21.445000 79.725000 ;
        RECT 21.245000 79.930000 21.445000 80.130000 ;
        RECT 21.245000 80.335000 21.445000 80.535000 ;
        RECT 21.245000 80.740000 21.445000 80.940000 ;
        RECT 21.245000 81.145000 21.445000 81.345000 ;
        RECT 21.245000 81.550000 21.445000 81.750000 ;
        RECT 21.245000 81.955000 21.445000 82.155000 ;
        RECT 21.245000 82.360000 21.445000 82.560000 ;
        RECT 21.345000 17.860000 21.545000 18.060000 ;
        RECT 21.345000 18.290000 21.545000 18.490000 ;
        RECT 21.345000 18.720000 21.545000 18.920000 ;
        RECT 21.345000 19.150000 21.545000 19.350000 ;
        RECT 21.345000 19.580000 21.545000 19.780000 ;
        RECT 21.345000 20.010000 21.545000 20.210000 ;
        RECT 21.345000 20.440000 21.545000 20.640000 ;
        RECT 21.345000 20.870000 21.545000 21.070000 ;
        RECT 21.345000 21.300000 21.545000 21.500000 ;
        RECT 21.345000 21.730000 21.545000 21.930000 ;
        RECT 21.345000 22.160000 21.545000 22.360000 ;
        RECT 21.645000 68.125000 21.845000 68.325000 ;
        RECT 21.645000 68.535000 21.845000 68.735000 ;
        RECT 21.645000 68.945000 21.845000 69.145000 ;
        RECT 21.645000 69.355000 21.845000 69.555000 ;
        RECT 21.645000 69.765000 21.845000 69.965000 ;
        RECT 21.645000 70.175000 21.845000 70.375000 ;
        RECT 21.645000 70.585000 21.845000 70.785000 ;
        RECT 21.645000 70.995000 21.845000 71.195000 ;
        RECT 21.645000 71.405000 21.845000 71.605000 ;
        RECT 21.645000 71.815000 21.845000 72.015000 ;
        RECT 21.645000 72.225000 21.845000 72.425000 ;
        RECT 21.645000 72.635000 21.845000 72.835000 ;
        RECT 21.645000 73.045000 21.845000 73.245000 ;
        RECT 21.645000 73.450000 21.845000 73.650000 ;
        RECT 21.645000 73.855000 21.845000 74.055000 ;
        RECT 21.645000 74.260000 21.845000 74.460000 ;
        RECT 21.645000 74.665000 21.845000 74.865000 ;
        RECT 21.645000 75.070000 21.845000 75.270000 ;
        RECT 21.645000 75.475000 21.845000 75.675000 ;
        RECT 21.645000 75.880000 21.845000 76.080000 ;
        RECT 21.645000 76.285000 21.845000 76.485000 ;
        RECT 21.645000 76.690000 21.845000 76.890000 ;
        RECT 21.645000 77.095000 21.845000 77.295000 ;
        RECT 21.645000 77.500000 21.845000 77.700000 ;
        RECT 21.645000 77.905000 21.845000 78.105000 ;
        RECT 21.645000 78.310000 21.845000 78.510000 ;
        RECT 21.645000 78.715000 21.845000 78.915000 ;
        RECT 21.645000 79.120000 21.845000 79.320000 ;
        RECT 21.645000 79.525000 21.845000 79.725000 ;
        RECT 21.645000 79.930000 21.845000 80.130000 ;
        RECT 21.645000 80.335000 21.845000 80.535000 ;
        RECT 21.645000 80.740000 21.845000 80.940000 ;
        RECT 21.645000 81.145000 21.845000 81.345000 ;
        RECT 21.645000 81.550000 21.845000 81.750000 ;
        RECT 21.645000 81.955000 21.845000 82.155000 ;
        RECT 21.645000 82.360000 21.845000 82.560000 ;
        RECT 21.715000 82.920000 21.915000 83.120000 ;
        RECT 21.715000 83.470000 21.915000 83.670000 ;
        RECT 21.715000 84.020000 21.915000 84.220000 ;
        RECT 21.750000 17.860000 21.950000 18.060000 ;
        RECT 21.750000 18.290000 21.950000 18.490000 ;
        RECT 21.750000 18.720000 21.950000 18.920000 ;
        RECT 21.750000 19.150000 21.950000 19.350000 ;
        RECT 21.750000 19.580000 21.950000 19.780000 ;
        RECT 21.750000 20.010000 21.950000 20.210000 ;
        RECT 21.750000 20.440000 21.950000 20.640000 ;
        RECT 21.750000 20.870000 21.950000 21.070000 ;
        RECT 21.750000 21.300000 21.950000 21.500000 ;
        RECT 21.750000 21.730000 21.950000 21.930000 ;
        RECT 21.750000 22.160000 21.950000 22.360000 ;
        RECT 22.045000 68.125000 22.245000 68.325000 ;
        RECT 22.045000 68.535000 22.245000 68.735000 ;
        RECT 22.045000 68.945000 22.245000 69.145000 ;
        RECT 22.045000 69.355000 22.245000 69.555000 ;
        RECT 22.045000 69.765000 22.245000 69.965000 ;
        RECT 22.045000 70.175000 22.245000 70.375000 ;
        RECT 22.045000 70.585000 22.245000 70.785000 ;
        RECT 22.045000 70.995000 22.245000 71.195000 ;
        RECT 22.045000 71.405000 22.245000 71.605000 ;
        RECT 22.045000 71.815000 22.245000 72.015000 ;
        RECT 22.045000 72.225000 22.245000 72.425000 ;
        RECT 22.045000 72.635000 22.245000 72.835000 ;
        RECT 22.045000 73.045000 22.245000 73.245000 ;
        RECT 22.045000 73.450000 22.245000 73.650000 ;
        RECT 22.045000 73.855000 22.245000 74.055000 ;
        RECT 22.045000 74.260000 22.245000 74.460000 ;
        RECT 22.045000 74.665000 22.245000 74.865000 ;
        RECT 22.045000 75.070000 22.245000 75.270000 ;
        RECT 22.045000 75.475000 22.245000 75.675000 ;
        RECT 22.045000 75.880000 22.245000 76.080000 ;
        RECT 22.045000 76.285000 22.245000 76.485000 ;
        RECT 22.045000 76.690000 22.245000 76.890000 ;
        RECT 22.045000 77.095000 22.245000 77.295000 ;
        RECT 22.045000 77.500000 22.245000 77.700000 ;
        RECT 22.045000 77.905000 22.245000 78.105000 ;
        RECT 22.045000 78.310000 22.245000 78.510000 ;
        RECT 22.045000 78.715000 22.245000 78.915000 ;
        RECT 22.045000 79.120000 22.245000 79.320000 ;
        RECT 22.045000 79.525000 22.245000 79.725000 ;
        RECT 22.045000 79.930000 22.245000 80.130000 ;
        RECT 22.045000 80.335000 22.245000 80.535000 ;
        RECT 22.045000 80.740000 22.245000 80.940000 ;
        RECT 22.045000 81.145000 22.245000 81.345000 ;
        RECT 22.045000 81.550000 22.245000 81.750000 ;
        RECT 22.045000 81.955000 22.245000 82.155000 ;
        RECT 22.045000 82.360000 22.245000 82.560000 ;
        RECT 22.160000 17.860000 22.360000 18.060000 ;
        RECT 22.160000 18.290000 22.360000 18.490000 ;
        RECT 22.160000 18.720000 22.360000 18.920000 ;
        RECT 22.160000 19.150000 22.360000 19.350000 ;
        RECT 22.160000 19.580000 22.360000 19.780000 ;
        RECT 22.160000 20.010000 22.360000 20.210000 ;
        RECT 22.160000 20.440000 22.360000 20.640000 ;
        RECT 22.160000 20.870000 22.360000 21.070000 ;
        RECT 22.160000 21.300000 22.360000 21.500000 ;
        RECT 22.160000 21.730000 22.360000 21.930000 ;
        RECT 22.160000 22.160000 22.360000 22.360000 ;
        RECT 22.445000 68.125000 22.645000 68.325000 ;
        RECT 22.445000 68.535000 22.645000 68.735000 ;
        RECT 22.445000 68.945000 22.645000 69.145000 ;
        RECT 22.445000 69.355000 22.645000 69.555000 ;
        RECT 22.445000 69.765000 22.645000 69.965000 ;
        RECT 22.445000 70.175000 22.645000 70.375000 ;
        RECT 22.445000 70.585000 22.645000 70.785000 ;
        RECT 22.445000 70.995000 22.645000 71.195000 ;
        RECT 22.445000 71.405000 22.645000 71.605000 ;
        RECT 22.445000 71.815000 22.645000 72.015000 ;
        RECT 22.445000 72.225000 22.645000 72.425000 ;
        RECT 22.445000 72.635000 22.645000 72.835000 ;
        RECT 22.445000 73.045000 22.645000 73.245000 ;
        RECT 22.445000 73.450000 22.645000 73.650000 ;
        RECT 22.445000 73.855000 22.645000 74.055000 ;
        RECT 22.445000 74.260000 22.645000 74.460000 ;
        RECT 22.445000 74.665000 22.645000 74.865000 ;
        RECT 22.445000 75.070000 22.645000 75.270000 ;
        RECT 22.445000 75.475000 22.645000 75.675000 ;
        RECT 22.445000 75.880000 22.645000 76.080000 ;
        RECT 22.445000 76.285000 22.645000 76.485000 ;
        RECT 22.445000 76.690000 22.645000 76.890000 ;
        RECT 22.445000 77.095000 22.645000 77.295000 ;
        RECT 22.445000 77.500000 22.645000 77.700000 ;
        RECT 22.445000 77.905000 22.645000 78.105000 ;
        RECT 22.445000 78.310000 22.645000 78.510000 ;
        RECT 22.445000 78.715000 22.645000 78.915000 ;
        RECT 22.445000 79.120000 22.645000 79.320000 ;
        RECT 22.445000 79.525000 22.645000 79.725000 ;
        RECT 22.445000 79.930000 22.645000 80.130000 ;
        RECT 22.445000 80.335000 22.645000 80.535000 ;
        RECT 22.445000 80.740000 22.645000 80.940000 ;
        RECT 22.445000 81.145000 22.645000 81.345000 ;
        RECT 22.445000 81.550000 22.645000 81.750000 ;
        RECT 22.445000 81.955000 22.645000 82.155000 ;
        RECT 22.445000 82.360000 22.645000 82.560000 ;
        RECT 22.505000 82.920000 22.705000 83.120000 ;
        RECT 22.505000 83.470000 22.705000 83.670000 ;
        RECT 22.505000 84.020000 22.705000 84.220000 ;
        RECT 22.570000 17.860000 22.770000 18.060000 ;
        RECT 22.570000 18.290000 22.770000 18.490000 ;
        RECT 22.570000 18.720000 22.770000 18.920000 ;
        RECT 22.570000 19.150000 22.770000 19.350000 ;
        RECT 22.570000 19.580000 22.770000 19.780000 ;
        RECT 22.570000 20.010000 22.770000 20.210000 ;
        RECT 22.570000 20.440000 22.770000 20.640000 ;
        RECT 22.570000 20.870000 22.770000 21.070000 ;
        RECT 22.570000 21.300000 22.770000 21.500000 ;
        RECT 22.570000 21.730000 22.770000 21.930000 ;
        RECT 22.570000 22.160000 22.770000 22.360000 ;
        RECT 22.845000 68.125000 23.045000 68.325000 ;
        RECT 22.845000 68.535000 23.045000 68.735000 ;
        RECT 22.845000 68.945000 23.045000 69.145000 ;
        RECT 22.845000 69.355000 23.045000 69.555000 ;
        RECT 22.845000 69.765000 23.045000 69.965000 ;
        RECT 22.845000 70.175000 23.045000 70.375000 ;
        RECT 22.845000 70.585000 23.045000 70.785000 ;
        RECT 22.845000 70.995000 23.045000 71.195000 ;
        RECT 22.845000 71.405000 23.045000 71.605000 ;
        RECT 22.845000 71.815000 23.045000 72.015000 ;
        RECT 22.845000 72.225000 23.045000 72.425000 ;
        RECT 22.845000 72.635000 23.045000 72.835000 ;
        RECT 22.845000 73.045000 23.045000 73.245000 ;
        RECT 22.845000 73.450000 23.045000 73.650000 ;
        RECT 22.845000 73.855000 23.045000 74.055000 ;
        RECT 22.845000 74.260000 23.045000 74.460000 ;
        RECT 22.845000 74.665000 23.045000 74.865000 ;
        RECT 22.845000 75.070000 23.045000 75.270000 ;
        RECT 22.845000 75.475000 23.045000 75.675000 ;
        RECT 22.845000 75.880000 23.045000 76.080000 ;
        RECT 22.845000 76.285000 23.045000 76.485000 ;
        RECT 22.845000 76.690000 23.045000 76.890000 ;
        RECT 22.845000 77.095000 23.045000 77.295000 ;
        RECT 22.845000 77.500000 23.045000 77.700000 ;
        RECT 22.845000 77.905000 23.045000 78.105000 ;
        RECT 22.845000 78.310000 23.045000 78.510000 ;
        RECT 22.845000 78.715000 23.045000 78.915000 ;
        RECT 22.845000 79.120000 23.045000 79.320000 ;
        RECT 22.845000 79.525000 23.045000 79.725000 ;
        RECT 22.845000 79.930000 23.045000 80.130000 ;
        RECT 22.845000 80.335000 23.045000 80.535000 ;
        RECT 22.845000 80.740000 23.045000 80.940000 ;
        RECT 22.845000 81.145000 23.045000 81.345000 ;
        RECT 22.845000 81.550000 23.045000 81.750000 ;
        RECT 22.845000 81.955000 23.045000 82.155000 ;
        RECT 22.845000 82.360000 23.045000 82.560000 ;
        RECT 22.980000 17.860000 23.180000 18.060000 ;
        RECT 22.980000 18.290000 23.180000 18.490000 ;
        RECT 22.980000 18.720000 23.180000 18.920000 ;
        RECT 22.980000 19.150000 23.180000 19.350000 ;
        RECT 22.980000 19.580000 23.180000 19.780000 ;
        RECT 22.980000 20.010000 23.180000 20.210000 ;
        RECT 22.980000 20.440000 23.180000 20.640000 ;
        RECT 22.980000 20.870000 23.180000 21.070000 ;
        RECT 22.980000 21.300000 23.180000 21.500000 ;
        RECT 22.980000 21.730000 23.180000 21.930000 ;
        RECT 22.980000 22.160000 23.180000 22.360000 ;
        RECT 23.245000 68.125000 23.445000 68.325000 ;
        RECT 23.245000 68.535000 23.445000 68.735000 ;
        RECT 23.245000 68.945000 23.445000 69.145000 ;
        RECT 23.245000 69.355000 23.445000 69.555000 ;
        RECT 23.245000 69.765000 23.445000 69.965000 ;
        RECT 23.245000 70.175000 23.445000 70.375000 ;
        RECT 23.245000 70.585000 23.445000 70.785000 ;
        RECT 23.245000 70.995000 23.445000 71.195000 ;
        RECT 23.245000 71.405000 23.445000 71.605000 ;
        RECT 23.245000 71.815000 23.445000 72.015000 ;
        RECT 23.245000 72.225000 23.445000 72.425000 ;
        RECT 23.245000 72.635000 23.445000 72.835000 ;
        RECT 23.245000 73.045000 23.445000 73.245000 ;
        RECT 23.245000 73.450000 23.445000 73.650000 ;
        RECT 23.245000 73.855000 23.445000 74.055000 ;
        RECT 23.245000 74.260000 23.445000 74.460000 ;
        RECT 23.245000 74.665000 23.445000 74.865000 ;
        RECT 23.245000 75.070000 23.445000 75.270000 ;
        RECT 23.245000 75.475000 23.445000 75.675000 ;
        RECT 23.245000 75.880000 23.445000 76.080000 ;
        RECT 23.245000 76.285000 23.445000 76.485000 ;
        RECT 23.245000 76.690000 23.445000 76.890000 ;
        RECT 23.245000 77.095000 23.445000 77.295000 ;
        RECT 23.245000 77.500000 23.445000 77.700000 ;
        RECT 23.245000 77.905000 23.445000 78.105000 ;
        RECT 23.245000 78.310000 23.445000 78.510000 ;
        RECT 23.245000 78.715000 23.445000 78.915000 ;
        RECT 23.245000 79.120000 23.445000 79.320000 ;
        RECT 23.245000 79.525000 23.445000 79.725000 ;
        RECT 23.245000 79.930000 23.445000 80.130000 ;
        RECT 23.245000 80.335000 23.445000 80.535000 ;
        RECT 23.245000 80.740000 23.445000 80.940000 ;
        RECT 23.245000 81.145000 23.445000 81.345000 ;
        RECT 23.245000 81.550000 23.445000 81.750000 ;
        RECT 23.245000 81.955000 23.445000 82.155000 ;
        RECT 23.245000 82.360000 23.445000 82.560000 ;
        RECT 23.390000 17.860000 23.590000 18.060000 ;
        RECT 23.390000 18.290000 23.590000 18.490000 ;
        RECT 23.390000 18.720000 23.590000 18.920000 ;
        RECT 23.390000 19.150000 23.590000 19.350000 ;
        RECT 23.390000 19.580000 23.590000 19.780000 ;
        RECT 23.390000 20.010000 23.590000 20.210000 ;
        RECT 23.390000 20.440000 23.590000 20.640000 ;
        RECT 23.390000 20.870000 23.590000 21.070000 ;
        RECT 23.390000 21.300000 23.590000 21.500000 ;
        RECT 23.390000 21.730000 23.590000 21.930000 ;
        RECT 23.390000 22.160000 23.590000 22.360000 ;
        RECT 23.645000 68.125000 23.845000 68.325000 ;
        RECT 23.645000 68.535000 23.845000 68.735000 ;
        RECT 23.645000 68.945000 23.845000 69.145000 ;
        RECT 23.645000 69.355000 23.845000 69.555000 ;
        RECT 23.645000 69.765000 23.845000 69.965000 ;
        RECT 23.645000 70.175000 23.845000 70.375000 ;
        RECT 23.645000 70.585000 23.845000 70.785000 ;
        RECT 23.645000 70.995000 23.845000 71.195000 ;
        RECT 23.645000 71.405000 23.845000 71.605000 ;
        RECT 23.645000 71.815000 23.845000 72.015000 ;
        RECT 23.645000 72.225000 23.845000 72.425000 ;
        RECT 23.645000 72.635000 23.845000 72.835000 ;
        RECT 23.645000 73.045000 23.845000 73.245000 ;
        RECT 23.645000 73.450000 23.845000 73.650000 ;
        RECT 23.645000 73.855000 23.845000 74.055000 ;
        RECT 23.645000 74.260000 23.845000 74.460000 ;
        RECT 23.645000 74.665000 23.845000 74.865000 ;
        RECT 23.645000 75.070000 23.845000 75.270000 ;
        RECT 23.645000 75.475000 23.845000 75.675000 ;
        RECT 23.645000 75.880000 23.845000 76.080000 ;
        RECT 23.645000 76.285000 23.845000 76.485000 ;
        RECT 23.645000 76.690000 23.845000 76.890000 ;
        RECT 23.645000 77.095000 23.845000 77.295000 ;
        RECT 23.645000 77.500000 23.845000 77.700000 ;
        RECT 23.645000 77.905000 23.845000 78.105000 ;
        RECT 23.645000 78.310000 23.845000 78.510000 ;
        RECT 23.645000 78.715000 23.845000 78.915000 ;
        RECT 23.645000 79.120000 23.845000 79.320000 ;
        RECT 23.645000 79.525000 23.845000 79.725000 ;
        RECT 23.645000 79.930000 23.845000 80.130000 ;
        RECT 23.645000 80.335000 23.845000 80.535000 ;
        RECT 23.645000 80.740000 23.845000 80.940000 ;
        RECT 23.645000 81.145000 23.845000 81.345000 ;
        RECT 23.645000 81.550000 23.845000 81.750000 ;
        RECT 23.645000 81.955000 23.845000 82.155000 ;
        RECT 23.645000 82.360000 23.845000 82.560000 ;
        RECT 23.800000 17.860000 24.000000 18.060000 ;
        RECT 23.800000 18.290000 24.000000 18.490000 ;
        RECT 23.800000 18.720000 24.000000 18.920000 ;
        RECT 23.800000 19.150000 24.000000 19.350000 ;
        RECT 23.800000 19.580000 24.000000 19.780000 ;
        RECT 23.800000 20.010000 24.000000 20.210000 ;
        RECT 23.800000 20.440000 24.000000 20.640000 ;
        RECT 23.800000 20.870000 24.000000 21.070000 ;
        RECT 23.800000 21.300000 24.000000 21.500000 ;
        RECT 23.800000 21.730000 24.000000 21.930000 ;
        RECT 23.800000 22.160000 24.000000 22.360000 ;
        RECT 24.045000 68.125000 24.245000 68.325000 ;
        RECT 24.045000 68.535000 24.245000 68.735000 ;
        RECT 24.045000 68.945000 24.245000 69.145000 ;
        RECT 24.045000 69.355000 24.245000 69.555000 ;
        RECT 24.045000 69.765000 24.245000 69.965000 ;
        RECT 24.045000 70.175000 24.245000 70.375000 ;
        RECT 24.045000 70.585000 24.245000 70.785000 ;
        RECT 24.045000 70.995000 24.245000 71.195000 ;
        RECT 24.045000 71.405000 24.245000 71.605000 ;
        RECT 24.045000 71.815000 24.245000 72.015000 ;
        RECT 24.045000 72.225000 24.245000 72.425000 ;
        RECT 24.045000 72.635000 24.245000 72.835000 ;
        RECT 24.045000 73.045000 24.245000 73.245000 ;
        RECT 24.045000 73.450000 24.245000 73.650000 ;
        RECT 24.045000 73.855000 24.245000 74.055000 ;
        RECT 24.045000 74.260000 24.245000 74.460000 ;
        RECT 24.045000 74.665000 24.245000 74.865000 ;
        RECT 24.045000 75.070000 24.245000 75.270000 ;
        RECT 24.045000 75.475000 24.245000 75.675000 ;
        RECT 24.045000 75.880000 24.245000 76.080000 ;
        RECT 24.045000 76.285000 24.245000 76.485000 ;
        RECT 24.045000 76.690000 24.245000 76.890000 ;
        RECT 24.045000 77.095000 24.245000 77.295000 ;
        RECT 24.045000 77.500000 24.245000 77.700000 ;
        RECT 24.045000 77.905000 24.245000 78.105000 ;
        RECT 24.045000 78.310000 24.245000 78.510000 ;
        RECT 24.045000 78.715000 24.245000 78.915000 ;
        RECT 24.045000 79.120000 24.245000 79.320000 ;
        RECT 24.045000 79.525000 24.245000 79.725000 ;
        RECT 24.045000 79.930000 24.245000 80.130000 ;
        RECT 24.045000 80.335000 24.245000 80.535000 ;
        RECT 24.045000 80.740000 24.245000 80.940000 ;
        RECT 24.045000 81.145000 24.245000 81.345000 ;
        RECT 24.045000 81.550000 24.245000 81.750000 ;
        RECT 24.045000 81.955000 24.245000 82.155000 ;
        RECT 24.045000 82.360000 24.245000 82.560000 ;
        RECT 24.210000 17.860000 24.410000 18.060000 ;
        RECT 24.210000 18.290000 24.410000 18.490000 ;
        RECT 24.210000 18.720000 24.410000 18.920000 ;
        RECT 24.210000 19.150000 24.410000 19.350000 ;
        RECT 24.210000 19.580000 24.410000 19.780000 ;
        RECT 24.210000 20.010000 24.410000 20.210000 ;
        RECT 24.210000 20.440000 24.410000 20.640000 ;
        RECT 24.210000 20.870000 24.410000 21.070000 ;
        RECT 24.210000 21.300000 24.410000 21.500000 ;
        RECT 24.210000 21.730000 24.410000 21.930000 ;
        RECT 24.210000 22.160000 24.410000 22.360000 ;
        RECT 50.845000 17.860000 51.045000 18.060000 ;
        RECT 50.845000 18.290000 51.045000 18.490000 ;
        RECT 50.845000 18.720000 51.045000 18.920000 ;
        RECT 50.845000 19.150000 51.045000 19.350000 ;
        RECT 50.845000 19.580000 51.045000 19.780000 ;
        RECT 50.845000 20.010000 51.045000 20.210000 ;
        RECT 50.845000 20.440000 51.045000 20.640000 ;
        RECT 50.845000 20.870000 51.045000 21.070000 ;
        RECT 50.845000 21.300000 51.045000 21.500000 ;
        RECT 50.845000 21.730000 51.045000 21.930000 ;
        RECT 50.845000 22.160000 51.045000 22.360000 ;
        RECT 51.010000 68.125000 51.210000 68.325000 ;
        RECT 51.010000 68.535000 51.210000 68.735000 ;
        RECT 51.010000 68.945000 51.210000 69.145000 ;
        RECT 51.010000 69.355000 51.210000 69.555000 ;
        RECT 51.010000 69.765000 51.210000 69.965000 ;
        RECT 51.010000 70.175000 51.210000 70.375000 ;
        RECT 51.010000 70.585000 51.210000 70.785000 ;
        RECT 51.010000 70.995000 51.210000 71.195000 ;
        RECT 51.010000 71.405000 51.210000 71.605000 ;
        RECT 51.010000 71.815000 51.210000 72.015000 ;
        RECT 51.010000 72.225000 51.210000 72.425000 ;
        RECT 51.010000 72.635000 51.210000 72.835000 ;
        RECT 51.010000 73.045000 51.210000 73.245000 ;
        RECT 51.010000 73.450000 51.210000 73.650000 ;
        RECT 51.010000 73.855000 51.210000 74.055000 ;
        RECT 51.010000 74.260000 51.210000 74.460000 ;
        RECT 51.010000 74.665000 51.210000 74.865000 ;
        RECT 51.010000 75.070000 51.210000 75.270000 ;
        RECT 51.010000 75.475000 51.210000 75.675000 ;
        RECT 51.010000 75.880000 51.210000 76.080000 ;
        RECT 51.010000 76.285000 51.210000 76.485000 ;
        RECT 51.010000 76.690000 51.210000 76.890000 ;
        RECT 51.010000 77.095000 51.210000 77.295000 ;
        RECT 51.010000 77.500000 51.210000 77.700000 ;
        RECT 51.010000 77.905000 51.210000 78.105000 ;
        RECT 51.010000 78.310000 51.210000 78.510000 ;
        RECT 51.010000 78.715000 51.210000 78.915000 ;
        RECT 51.010000 79.120000 51.210000 79.320000 ;
        RECT 51.010000 79.525000 51.210000 79.725000 ;
        RECT 51.010000 79.930000 51.210000 80.130000 ;
        RECT 51.010000 80.335000 51.210000 80.535000 ;
        RECT 51.010000 80.740000 51.210000 80.940000 ;
        RECT 51.010000 81.145000 51.210000 81.345000 ;
        RECT 51.010000 81.550000 51.210000 81.750000 ;
        RECT 51.010000 81.955000 51.210000 82.155000 ;
        RECT 51.010000 82.360000 51.210000 82.560000 ;
        RECT 51.250000 17.860000 51.450000 18.060000 ;
        RECT 51.250000 18.290000 51.450000 18.490000 ;
        RECT 51.250000 18.720000 51.450000 18.920000 ;
        RECT 51.250000 19.150000 51.450000 19.350000 ;
        RECT 51.250000 19.580000 51.450000 19.780000 ;
        RECT 51.250000 20.010000 51.450000 20.210000 ;
        RECT 51.250000 20.440000 51.450000 20.640000 ;
        RECT 51.250000 20.870000 51.450000 21.070000 ;
        RECT 51.250000 21.300000 51.450000 21.500000 ;
        RECT 51.250000 21.730000 51.450000 21.930000 ;
        RECT 51.250000 22.160000 51.450000 22.360000 ;
        RECT 51.410000 68.125000 51.610000 68.325000 ;
        RECT 51.410000 68.535000 51.610000 68.735000 ;
        RECT 51.410000 68.945000 51.610000 69.145000 ;
        RECT 51.410000 69.355000 51.610000 69.555000 ;
        RECT 51.410000 69.765000 51.610000 69.965000 ;
        RECT 51.410000 70.175000 51.610000 70.375000 ;
        RECT 51.410000 70.585000 51.610000 70.785000 ;
        RECT 51.410000 70.995000 51.610000 71.195000 ;
        RECT 51.410000 71.405000 51.610000 71.605000 ;
        RECT 51.410000 71.815000 51.610000 72.015000 ;
        RECT 51.410000 72.225000 51.610000 72.425000 ;
        RECT 51.410000 72.635000 51.610000 72.835000 ;
        RECT 51.410000 73.045000 51.610000 73.245000 ;
        RECT 51.410000 73.450000 51.610000 73.650000 ;
        RECT 51.410000 73.855000 51.610000 74.055000 ;
        RECT 51.410000 74.260000 51.610000 74.460000 ;
        RECT 51.410000 74.665000 51.610000 74.865000 ;
        RECT 51.410000 75.070000 51.610000 75.270000 ;
        RECT 51.410000 75.475000 51.610000 75.675000 ;
        RECT 51.410000 75.880000 51.610000 76.080000 ;
        RECT 51.410000 76.285000 51.610000 76.485000 ;
        RECT 51.410000 76.690000 51.610000 76.890000 ;
        RECT 51.410000 77.095000 51.610000 77.295000 ;
        RECT 51.410000 77.500000 51.610000 77.700000 ;
        RECT 51.410000 77.905000 51.610000 78.105000 ;
        RECT 51.410000 78.310000 51.610000 78.510000 ;
        RECT 51.410000 78.715000 51.610000 78.915000 ;
        RECT 51.410000 79.120000 51.610000 79.320000 ;
        RECT 51.410000 79.525000 51.610000 79.725000 ;
        RECT 51.410000 79.930000 51.610000 80.130000 ;
        RECT 51.410000 80.335000 51.610000 80.535000 ;
        RECT 51.410000 80.740000 51.610000 80.940000 ;
        RECT 51.410000 81.145000 51.610000 81.345000 ;
        RECT 51.410000 81.550000 51.610000 81.750000 ;
        RECT 51.410000 81.955000 51.610000 82.155000 ;
        RECT 51.410000 82.360000 51.610000 82.560000 ;
        RECT 51.655000 17.860000 51.855000 18.060000 ;
        RECT 51.655000 18.290000 51.855000 18.490000 ;
        RECT 51.655000 18.720000 51.855000 18.920000 ;
        RECT 51.655000 19.150000 51.855000 19.350000 ;
        RECT 51.655000 19.580000 51.855000 19.780000 ;
        RECT 51.655000 20.010000 51.855000 20.210000 ;
        RECT 51.655000 20.440000 51.855000 20.640000 ;
        RECT 51.655000 20.870000 51.855000 21.070000 ;
        RECT 51.655000 21.300000 51.855000 21.500000 ;
        RECT 51.655000 21.730000 51.855000 21.930000 ;
        RECT 51.655000 22.160000 51.855000 22.360000 ;
        RECT 51.810000 68.125000 52.010000 68.325000 ;
        RECT 51.810000 68.535000 52.010000 68.735000 ;
        RECT 51.810000 68.945000 52.010000 69.145000 ;
        RECT 51.810000 69.355000 52.010000 69.555000 ;
        RECT 51.810000 69.765000 52.010000 69.965000 ;
        RECT 51.810000 70.175000 52.010000 70.375000 ;
        RECT 51.810000 70.585000 52.010000 70.785000 ;
        RECT 51.810000 70.995000 52.010000 71.195000 ;
        RECT 51.810000 71.405000 52.010000 71.605000 ;
        RECT 51.810000 71.815000 52.010000 72.015000 ;
        RECT 51.810000 72.225000 52.010000 72.425000 ;
        RECT 51.810000 72.635000 52.010000 72.835000 ;
        RECT 51.810000 73.045000 52.010000 73.245000 ;
        RECT 51.810000 73.450000 52.010000 73.650000 ;
        RECT 51.810000 73.855000 52.010000 74.055000 ;
        RECT 51.810000 74.260000 52.010000 74.460000 ;
        RECT 51.810000 74.665000 52.010000 74.865000 ;
        RECT 51.810000 75.070000 52.010000 75.270000 ;
        RECT 51.810000 75.475000 52.010000 75.675000 ;
        RECT 51.810000 75.880000 52.010000 76.080000 ;
        RECT 51.810000 76.285000 52.010000 76.485000 ;
        RECT 51.810000 76.690000 52.010000 76.890000 ;
        RECT 51.810000 77.095000 52.010000 77.295000 ;
        RECT 51.810000 77.500000 52.010000 77.700000 ;
        RECT 51.810000 77.905000 52.010000 78.105000 ;
        RECT 51.810000 78.310000 52.010000 78.510000 ;
        RECT 51.810000 78.715000 52.010000 78.915000 ;
        RECT 51.810000 79.120000 52.010000 79.320000 ;
        RECT 51.810000 79.525000 52.010000 79.725000 ;
        RECT 51.810000 79.930000 52.010000 80.130000 ;
        RECT 51.810000 80.335000 52.010000 80.535000 ;
        RECT 51.810000 80.740000 52.010000 80.940000 ;
        RECT 51.810000 81.145000 52.010000 81.345000 ;
        RECT 51.810000 81.550000 52.010000 81.750000 ;
        RECT 51.810000 81.955000 52.010000 82.155000 ;
        RECT 51.810000 82.360000 52.010000 82.560000 ;
        RECT 52.060000 17.860000 52.260000 18.060000 ;
        RECT 52.060000 18.290000 52.260000 18.490000 ;
        RECT 52.060000 18.720000 52.260000 18.920000 ;
        RECT 52.060000 19.150000 52.260000 19.350000 ;
        RECT 52.060000 19.580000 52.260000 19.780000 ;
        RECT 52.060000 20.010000 52.260000 20.210000 ;
        RECT 52.060000 20.440000 52.260000 20.640000 ;
        RECT 52.060000 20.870000 52.260000 21.070000 ;
        RECT 52.060000 21.300000 52.260000 21.500000 ;
        RECT 52.060000 21.730000 52.260000 21.930000 ;
        RECT 52.060000 22.160000 52.260000 22.360000 ;
        RECT 52.210000 68.125000 52.410000 68.325000 ;
        RECT 52.210000 68.535000 52.410000 68.735000 ;
        RECT 52.210000 68.945000 52.410000 69.145000 ;
        RECT 52.210000 69.355000 52.410000 69.555000 ;
        RECT 52.210000 69.765000 52.410000 69.965000 ;
        RECT 52.210000 70.175000 52.410000 70.375000 ;
        RECT 52.210000 70.585000 52.410000 70.785000 ;
        RECT 52.210000 70.995000 52.410000 71.195000 ;
        RECT 52.210000 71.405000 52.410000 71.605000 ;
        RECT 52.210000 71.815000 52.410000 72.015000 ;
        RECT 52.210000 72.225000 52.410000 72.425000 ;
        RECT 52.210000 72.635000 52.410000 72.835000 ;
        RECT 52.210000 73.045000 52.410000 73.245000 ;
        RECT 52.210000 73.450000 52.410000 73.650000 ;
        RECT 52.210000 73.855000 52.410000 74.055000 ;
        RECT 52.210000 74.260000 52.410000 74.460000 ;
        RECT 52.210000 74.665000 52.410000 74.865000 ;
        RECT 52.210000 75.070000 52.410000 75.270000 ;
        RECT 52.210000 75.475000 52.410000 75.675000 ;
        RECT 52.210000 75.880000 52.410000 76.080000 ;
        RECT 52.210000 76.285000 52.410000 76.485000 ;
        RECT 52.210000 76.690000 52.410000 76.890000 ;
        RECT 52.210000 77.095000 52.410000 77.295000 ;
        RECT 52.210000 77.500000 52.410000 77.700000 ;
        RECT 52.210000 77.905000 52.410000 78.105000 ;
        RECT 52.210000 78.310000 52.410000 78.510000 ;
        RECT 52.210000 78.715000 52.410000 78.915000 ;
        RECT 52.210000 79.120000 52.410000 79.320000 ;
        RECT 52.210000 79.525000 52.410000 79.725000 ;
        RECT 52.210000 79.930000 52.410000 80.130000 ;
        RECT 52.210000 80.335000 52.410000 80.535000 ;
        RECT 52.210000 80.740000 52.410000 80.940000 ;
        RECT 52.210000 81.145000 52.410000 81.345000 ;
        RECT 52.210000 81.550000 52.410000 81.750000 ;
        RECT 52.210000 81.955000 52.410000 82.155000 ;
        RECT 52.210000 82.360000 52.410000 82.560000 ;
        RECT 52.465000 17.860000 52.665000 18.060000 ;
        RECT 52.465000 18.290000 52.665000 18.490000 ;
        RECT 52.465000 18.720000 52.665000 18.920000 ;
        RECT 52.465000 19.150000 52.665000 19.350000 ;
        RECT 52.465000 19.580000 52.665000 19.780000 ;
        RECT 52.465000 20.010000 52.665000 20.210000 ;
        RECT 52.465000 20.440000 52.665000 20.640000 ;
        RECT 52.465000 20.870000 52.665000 21.070000 ;
        RECT 52.465000 21.300000 52.665000 21.500000 ;
        RECT 52.465000 21.730000 52.665000 21.930000 ;
        RECT 52.465000 22.160000 52.665000 22.360000 ;
        RECT 52.550000 82.920000 52.750000 83.120000 ;
        RECT 52.550000 83.470000 52.750000 83.670000 ;
        RECT 52.550000 84.020000 52.750000 84.220000 ;
        RECT 52.610000 68.125000 52.810000 68.325000 ;
        RECT 52.610000 68.535000 52.810000 68.735000 ;
        RECT 52.610000 68.945000 52.810000 69.145000 ;
        RECT 52.610000 69.355000 52.810000 69.555000 ;
        RECT 52.610000 69.765000 52.810000 69.965000 ;
        RECT 52.610000 70.175000 52.810000 70.375000 ;
        RECT 52.610000 70.585000 52.810000 70.785000 ;
        RECT 52.610000 70.995000 52.810000 71.195000 ;
        RECT 52.610000 71.405000 52.810000 71.605000 ;
        RECT 52.610000 71.815000 52.810000 72.015000 ;
        RECT 52.610000 72.225000 52.810000 72.425000 ;
        RECT 52.610000 72.635000 52.810000 72.835000 ;
        RECT 52.610000 73.045000 52.810000 73.245000 ;
        RECT 52.610000 73.450000 52.810000 73.650000 ;
        RECT 52.610000 73.855000 52.810000 74.055000 ;
        RECT 52.610000 74.260000 52.810000 74.460000 ;
        RECT 52.610000 74.665000 52.810000 74.865000 ;
        RECT 52.610000 75.070000 52.810000 75.270000 ;
        RECT 52.610000 75.475000 52.810000 75.675000 ;
        RECT 52.610000 75.880000 52.810000 76.080000 ;
        RECT 52.610000 76.285000 52.810000 76.485000 ;
        RECT 52.610000 76.690000 52.810000 76.890000 ;
        RECT 52.610000 77.095000 52.810000 77.295000 ;
        RECT 52.610000 77.500000 52.810000 77.700000 ;
        RECT 52.610000 77.905000 52.810000 78.105000 ;
        RECT 52.610000 78.310000 52.810000 78.510000 ;
        RECT 52.610000 78.715000 52.810000 78.915000 ;
        RECT 52.610000 79.120000 52.810000 79.320000 ;
        RECT 52.610000 79.525000 52.810000 79.725000 ;
        RECT 52.610000 79.930000 52.810000 80.130000 ;
        RECT 52.610000 80.335000 52.810000 80.535000 ;
        RECT 52.610000 80.740000 52.810000 80.940000 ;
        RECT 52.610000 81.145000 52.810000 81.345000 ;
        RECT 52.610000 81.550000 52.810000 81.750000 ;
        RECT 52.610000 81.955000 52.810000 82.155000 ;
        RECT 52.610000 82.360000 52.810000 82.560000 ;
        RECT 52.870000 17.860000 53.070000 18.060000 ;
        RECT 52.870000 18.290000 53.070000 18.490000 ;
        RECT 52.870000 18.720000 53.070000 18.920000 ;
        RECT 52.870000 19.150000 53.070000 19.350000 ;
        RECT 52.870000 19.580000 53.070000 19.780000 ;
        RECT 52.870000 20.010000 53.070000 20.210000 ;
        RECT 52.870000 20.440000 53.070000 20.640000 ;
        RECT 52.870000 20.870000 53.070000 21.070000 ;
        RECT 52.870000 21.300000 53.070000 21.500000 ;
        RECT 52.870000 21.730000 53.070000 21.930000 ;
        RECT 52.870000 22.160000 53.070000 22.360000 ;
        RECT 53.010000 68.125000 53.210000 68.325000 ;
        RECT 53.010000 68.535000 53.210000 68.735000 ;
        RECT 53.010000 68.945000 53.210000 69.145000 ;
        RECT 53.010000 69.355000 53.210000 69.555000 ;
        RECT 53.010000 69.765000 53.210000 69.965000 ;
        RECT 53.010000 70.175000 53.210000 70.375000 ;
        RECT 53.010000 70.585000 53.210000 70.785000 ;
        RECT 53.010000 70.995000 53.210000 71.195000 ;
        RECT 53.010000 71.405000 53.210000 71.605000 ;
        RECT 53.010000 71.815000 53.210000 72.015000 ;
        RECT 53.010000 72.225000 53.210000 72.425000 ;
        RECT 53.010000 72.635000 53.210000 72.835000 ;
        RECT 53.010000 73.045000 53.210000 73.245000 ;
        RECT 53.010000 73.450000 53.210000 73.650000 ;
        RECT 53.010000 73.855000 53.210000 74.055000 ;
        RECT 53.010000 74.260000 53.210000 74.460000 ;
        RECT 53.010000 74.665000 53.210000 74.865000 ;
        RECT 53.010000 75.070000 53.210000 75.270000 ;
        RECT 53.010000 75.475000 53.210000 75.675000 ;
        RECT 53.010000 75.880000 53.210000 76.080000 ;
        RECT 53.010000 76.285000 53.210000 76.485000 ;
        RECT 53.010000 76.690000 53.210000 76.890000 ;
        RECT 53.010000 77.095000 53.210000 77.295000 ;
        RECT 53.010000 77.500000 53.210000 77.700000 ;
        RECT 53.010000 77.905000 53.210000 78.105000 ;
        RECT 53.010000 78.310000 53.210000 78.510000 ;
        RECT 53.010000 78.715000 53.210000 78.915000 ;
        RECT 53.010000 79.120000 53.210000 79.320000 ;
        RECT 53.010000 79.525000 53.210000 79.725000 ;
        RECT 53.010000 79.930000 53.210000 80.130000 ;
        RECT 53.010000 80.335000 53.210000 80.535000 ;
        RECT 53.010000 80.740000 53.210000 80.940000 ;
        RECT 53.010000 81.145000 53.210000 81.345000 ;
        RECT 53.010000 81.550000 53.210000 81.750000 ;
        RECT 53.010000 81.955000 53.210000 82.155000 ;
        RECT 53.010000 82.360000 53.210000 82.560000 ;
        RECT 53.275000 17.860000 53.475000 18.060000 ;
        RECT 53.275000 18.290000 53.475000 18.490000 ;
        RECT 53.275000 18.720000 53.475000 18.920000 ;
        RECT 53.275000 19.150000 53.475000 19.350000 ;
        RECT 53.275000 19.580000 53.475000 19.780000 ;
        RECT 53.275000 20.010000 53.475000 20.210000 ;
        RECT 53.275000 20.440000 53.475000 20.640000 ;
        RECT 53.275000 20.870000 53.475000 21.070000 ;
        RECT 53.275000 21.300000 53.475000 21.500000 ;
        RECT 53.275000 21.730000 53.475000 21.930000 ;
        RECT 53.275000 22.160000 53.475000 22.360000 ;
        RECT 53.340000 82.920000 53.540000 83.120000 ;
        RECT 53.340000 83.470000 53.540000 83.670000 ;
        RECT 53.340000 84.020000 53.540000 84.220000 ;
        RECT 53.410000 68.125000 53.610000 68.325000 ;
        RECT 53.410000 68.535000 53.610000 68.735000 ;
        RECT 53.410000 68.945000 53.610000 69.145000 ;
        RECT 53.410000 69.355000 53.610000 69.555000 ;
        RECT 53.410000 69.765000 53.610000 69.965000 ;
        RECT 53.410000 70.175000 53.610000 70.375000 ;
        RECT 53.410000 70.585000 53.610000 70.785000 ;
        RECT 53.410000 70.995000 53.610000 71.195000 ;
        RECT 53.410000 71.405000 53.610000 71.605000 ;
        RECT 53.410000 71.815000 53.610000 72.015000 ;
        RECT 53.410000 72.225000 53.610000 72.425000 ;
        RECT 53.410000 72.635000 53.610000 72.835000 ;
        RECT 53.410000 73.045000 53.610000 73.245000 ;
        RECT 53.410000 73.450000 53.610000 73.650000 ;
        RECT 53.410000 73.855000 53.610000 74.055000 ;
        RECT 53.410000 74.260000 53.610000 74.460000 ;
        RECT 53.410000 74.665000 53.610000 74.865000 ;
        RECT 53.410000 75.070000 53.610000 75.270000 ;
        RECT 53.410000 75.475000 53.610000 75.675000 ;
        RECT 53.410000 75.880000 53.610000 76.080000 ;
        RECT 53.410000 76.285000 53.610000 76.485000 ;
        RECT 53.410000 76.690000 53.610000 76.890000 ;
        RECT 53.410000 77.095000 53.610000 77.295000 ;
        RECT 53.410000 77.500000 53.610000 77.700000 ;
        RECT 53.410000 77.905000 53.610000 78.105000 ;
        RECT 53.410000 78.310000 53.610000 78.510000 ;
        RECT 53.410000 78.715000 53.610000 78.915000 ;
        RECT 53.410000 79.120000 53.610000 79.320000 ;
        RECT 53.410000 79.525000 53.610000 79.725000 ;
        RECT 53.410000 79.930000 53.610000 80.130000 ;
        RECT 53.410000 80.335000 53.610000 80.535000 ;
        RECT 53.410000 80.740000 53.610000 80.940000 ;
        RECT 53.410000 81.145000 53.610000 81.345000 ;
        RECT 53.410000 81.550000 53.610000 81.750000 ;
        RECT 53.410000 81.955000 53.610000 82.155000 ;
        RECT 53.410000 82.360000 53.610000 82.560000 ;
        RECT 53.680000 17.860000 53.880000 18.060000 ;
        RECT 53.680000 18.290000 53.880000 18.490000 ;
        RECT 53.680000 18.720000 53.880000 18.920000 ;
        RECT 53.680000 19.150000 53.880000 19.350000 ;
        RECT 53.680000 19.580000 53.880000 19.780000 ;
        RECT 53.680000 20.010000 53.880000 20.210000 ;
        RECT 53.680000 20.440000 53.880000 20.640000 ;
        RECT 53.680000 20.870000 53.880000 21.070000 ;
        RECT 53.680000 21.300000 53.880000 21.500000 ;
        RECT 53.680000 21.730000 53.880000 21.930000 ;
        RECT 53.680000 22.160000 53.880000 22.360000 ;
        RECT 53.810000 68.125000 54.010000 68.325000 ;
        RECT 53.810000 68.535000 54.010000 68.735000 ;
        RECT 53.810000 68.945000 54.010000 69.145000 ;
        RECT 53.810000 69.355000 54.010000 69.555000 ;
        RECT 53.810000 69.765000 54.010000 69.965000 ;
        RECT 53.810000 70.175000 54.010000 70.375000 ;
        RECT 53.810000 70.585000 54.010000 70.785000 ;
        RECT 53.810000 70.995000 54.010000 71.195000 ;
        RECT 53.810000 71.405000 54.010000 71.605000 ;
        RECT 53.810000 71.815000 54.010000 72.015000 ;
        RECT 53.810000 72.225000 54.010000 72.425000 ;
        RECT 53.810000 72.635000 54.010000 72.835000 ;
        RECT 53.810000 73.045000 54.010000 73.245000 ;
        RECT 53.810000 73.450000 54.010000 73.650000 ;
        RECT 53.810000 73.855000 54.010000 74.055000 ;
        RECT 53.810000 74.260000 54.010000 74.460000 ;
        RECT 53.810000 74.665000 54.010000 74.865000 ;
        RECT 53.810000 75.070000 54.010000 75.270000 ;
        RECT 53.810000 75.475000 54.010000 75.675000 ;
        RECT 53.810000 75.880000 54.010000 76.080000 ;
        RECT 53.810000 76.285000 54.010000 76.485000 ;
        RECT 53.810000 76.690000 54.010000 76.890000 ;
        RECT 53.810000 77.095000 54.010000 77.295000 ;
        RECT 53.810000 77.500000 54.010000 77.700000 ;
        RECT 53.810000 77.905000 54.010000 78.105000 ;
        RECT 53.810000 78.310000 54.010000 78.510000 ;
        RECT 53.810000 78.715000 54.010000 78.915000 ;
        RECT 53.810000 79.120000 54.010000 79.320000 ;
        RECT 53.810000 79.525000 54.010000 79.725000 ;
        RECT 53.810000 79.930000 54.010000 80.130000 ;
        RECT 53.810000 80.335000 54.010000 80.535000 ;
        RECT 53.810000 80.740000 54.010000 80.940000 ;
        RECT 53.810000 81.145000 54.010000 81.345000 ;
        RECT 53.810000 81.550000 54.010000 81.750000 ;
        RECT 53.810000 81.955000 54.010000 82.155000 ;
        RECT 53.810000 82.360000 54.010000 82.560000 ;
        RECT 53.885000 83.010000 54.085000 83.210000 ;
        RECT 53.885000 83.470000 54.085000 83.670000 ;
        RECT 53.885000 83.930000 54.085000 84.130000 ;
        RECT 53.885000 84.395000 54.085000 84.595000 ;
        RECT 53.885000 84.860000 54.085000 85.060000 ;
        RECT 53.885000 85.325000 54.085000 85.525000 ;
        RECT 54.085000 17.860000 54.285000 18.060000 ;
        RECT 54.085000 18.290000 54.285000 18.490000 ;
        RECT 54.085000 18.720000 54.285000 18.920000 ;
        RECT 54.085000 19.150000 54.285000 19.350000 ;
        RECT 54.085000 19.580000 54.285000 19.780000 ;
        RECT 54.085000 20.010000 54.285000 20.210000 ;
        RECT 54.085000 20.440000 54.285000 20.640000 ;
        RECT 54.085000 20.870000 54.285000 21.070000 ;
        RECT 54.085000 21.300000 54.285000 21.500000 ;
        RECT 54.085000 21.730000 54.285000 21.930000 ;
        RECT 54.085000 22.160000 54.285000 22.360000 ;
        RECT 54.210000 68.125000 54.410000 68.325000 ;
        RECT 54.210000 68.535000 54.410000 68.735000 ;
        RECT 54.210000 68.945000 54.410000 69.145000 ;
        RECT 54.210000 69.355000 54.410000 69.555000 ;
        RECT 54.210000 69.765000 54.410000 69.965000 ;
        RECT 54.210000 70.175000 54.410000 70.375000 ;
        RECT 54.210000 70.585000 54.410000 70.785000 ;
        RECT 54.210000 70.995000 54.410000 71.195000 ;
        RECT 54.210000 71.405000 54.410000 71.605000 ;
        RECT 54.210000 71.815000 54.410000 72.015000 ;
        RECT 54.210000 72.225000 54.410000 72.425000 ;
        RECT 54.210000 72.635000 54.410000 72.835000 ;
        RECT 54.210000 73.045000 54.410000 73.245000 ;
        RECT 54.210000 73.450000 54.410000 73.650000 ;
        RECT 54.210000 73.855000 54.410000 74.055000 ;
        RECT 54.210000 74.260000 54.410000 74.460000 ;
        RECT 54.210000 74.665000 54.410000 74.865000 ;
        RECT 54.210000 75.070000 54.410000 75.270000 ;
        RECT 54.210000 75.475000 54.410000 75.675000 ;
        RECT 54.210000 75.880000 54.410000 76.080000 ;
        RECT 54.210000 76.285000 54.410000 76.485000 ;
        RECT 54.210000 76.690000 54.410000 76.890000 ;
        RECT 54.210000 77.095000 54.410000 77.295000 ;
        RECT 54.210000 77.500000 54.410000 77.700000 ;
        RECT 54.210000 77.905000 54.410000 78.105000 ;
        RECT 54.210000 78.310000 54.410000 78.510000 ;
        RECT 54.210000 78.715000 54.410000 78.915000 ;
        RECT 54.210000 79.120000 54.410000 79.320000 ;
        RECT 54.210000 79.525000 54.410000 79.725000 ;
        RECT 54.210000 79.930000 54.410000 80.130000 ;
        RECT 54.210000 80.335000 54.410000 80.535000 ;
        RECT 54.210000 80.740000 54.410000 80.940000 ;
        RECT 54.210000 81.145000 54.410000 81.345000 ;
        RECT 54.210000 81.550000 54.410000 81.750000 ;
        RECT 54.210000 81.955000 54.410000 82.155000 ;
        RECT 54.210000 82.360000 54.410000 82.560000 ;
        RECT 54.365000 83.010000 54.565000 83.210000 ;
        RECT 54.365000 83.470000 54.565000 83.670000 ;
        RECT 54.365000 83.930000 54.565000 84.130000 ;
        RECT 54.365000 84.395000 54.565000 84.595000 ;
        RECT 54.365000 84.860000 54.565000 85.060000 ;
        RECT 54.365000 85.325000 54.565000 85.525000 ;
        RECT 54.490000 17.860000 54.690000 18.060000 ;
        RECT 54.490000 18.290000 54.690000 18.490000 ;
        RECT 54.490000 18.720000 54.690000 18.920000 ;
        RECT 54.490000 19.150000 54.690000 19.350000 ;
        RECT 54.490000 19.580000 54.690000 19.780000 ;
        RECT 54.490000 20.010000 54.690000 20.210000 ;
        RECT 54.490000 20.440000 54.690000 20.640000 ;
        RECT 54.490000 20.870000 54.690000 21.070000 ;
        RECT 54.490000 21.300000 54.690000 21.500000 ;
        RECT 54.490000 21.730000 54.690000 21.930000 ;
        RECT 54.490000 22.160000 54.690000 22.360000 ;
        RECT 54.610000 68.125000 54.810000 68.325000 ;
        RECT 54.610000 68.535000 54.810000 68.735000 ;
        RECT 54.610000 68.945000 54.810000 69.145000 ;
        RECT 54.610000 69.355000 54.810000 69.555000 ;
        RECT 54.610000 69.765000 54.810000 69.965000 ;
        RECT 54.610000 70.175000 54.810000 70.375000 ;
        RECT 54.610000 70.585000 54.810000 70.785000 ;
        RECT 54.610000 70.995000 54.810000 71.195000 ;
        RECT 54.610000 71.405000 54.810000 71.605000 ;
        RECT 54.610000 71.815000 54.810000 72.015000 ;
        RECT 54.610000 72.225000 54.810000 72.425000 ;
        RECT 54.610000 72.635000 54.810000 72.835000 ;
        RECT 54.610000 73.045000 54.810000 73.245000 ;
        RECT 54.610000 73.450000 54.810000 73.650000 ;
        RECT 54.610000 73.855000 54.810000 74.055000 ;
        RECT 54.610000 74.260000 54.810000 74.460000 ;
        RECT 54.610000 74.665000 54.810000 74.865000 ;
        RECT 54.610000 75.070000 54.810000 75.270000 ;
        RECT 54.610000 75.475000 54.810000 75.675000 ;
        RECT 54.610000 75.880000 54.810000 76.080000 ;
        RECT 54.610000 76.285000 54.810000 76.485000 ;
        RECT 54.610000 76.690000 54.810000 76.890000 ;
        RECT 54.610000 77.095000 54.810000 77.295000 ;
        RECT 54.610000 77.500000 54.810000 77.700000 ;
        RECT 54.610000 77.905000 54.810000 78.105000 ;
        RECT 54.610000 78.310000 54.810000 78.510000 ;
        RECT 54.610000 78.715000 54.810000 78.915000 ;
        RECT 54.610000 79.120000 54.810000 79.320000 ;
        RECT 54.610000 79.525000 54.810000 79.725000 ;
        RECT 54.610000 79.930000 54.810000 80.130000 ;
        RECT 54.610000 80.335000 54.810000 80.535000 ;
        RECT 54.610000 80.740000 54.810000 80.940000 ;
        RECT 54.610000 81.145000 54.810000 81.345000 ;
        RECT 54.610000 81.550000 54.810000 81.750000 ;
        RECT 54.610000 81.955000 54.810000 82.155000 ;
        RECT 54.610000 82.360000 54.810000 82.560000 ;
        RECT 54.845000 83.010000 55.045000 83.210000 ;
        RECT 54.845000 83.470000 55.045000 83.670000 ;
        RECT 54.845000 83.930000 55.045000 84.130000 ;
        RECT 54.845000 84.395000 55.045000 84.595000 ;
        RECT 54.845000 84.860000 55.045000 85.060000 ;
        RECT 54.845000 85.325000 55.045000 85.525000 ;
        RECT 54.895000 17.860000 55.095000 18.060000 ;
        RECT 54.895000 18.290000 55.095000 18.490000 ;
        RECT 54.895000 18.720000 55.095000 18.920000 ;
        RECT 54.895000 19.150000 55.095000 19.350000 ;
        RECT 54.895000 19.580000 55.095000 19.780000 ;
        RECT 54.895000 20.010000 55.095000 20.210000 ;
        RECT 54.895000 20.440000 55.095000 20.640000 ;
        RECT 54.895000 20.870000 55.095000 21.070000 ;
        RECT 54.895000 21.300000 55.095000 21.500000 ;
        RECT 54.895000 21.730000 55.095000 21.930000 ;
        RECT 54.895000 22.160000 55.095000 22.360000 ;
        RECT 55.010000 68.125000 55.210000 68.325000 ;
        RECT 55.010000 68.535000 55.210000 68.735000 ;
        RECT 55.010000 68.945000 55.210000 69.145000 ;
        RECT 55.010000 69.355000 55.210000 69.555000 ;
        RECT 55.010000 69.765000 55.210000 69.965000 ;
        RECT 55.010000 70.175000 55.210000 70.375000 ;
        RECT 55.010000 70.585000 55.210000 70.785000 ;
        RECT 55.010000 70.995000 55.210000 71.195000 ;
        RECT 55.010000 71.405000 55.210000 71.605000 ;
        RECT 55.010000 71.815000 55.210000 72.015000 ;
        RECT 55.010000 72.225000 55.210000 72.425000 ;
        RECT 55.010000 72.635000 55.210000 72.835000 ;
        RECT 55.010000 73.045000 55.210000 73.245000 ;
        RECT 55.010000 73.450000 55.210000 73.650000 ;
        RECT 55.010000 73.855000 55.210000 74.055000 ;
        RECT 55.010000 74.260000 55.210000 74.460000 ;
        RECT 55.010000 74.665000 55.210000 74.865000 ;
        RECT 55.010000 75.070000 55.210000 75.270000 ;
        RECT 55.010000 75.475000 55.210000 75.675000 ;
        RECT 55.010000 75.880000 55.210000 76.080000 ;
        RECT 55.010000 76.285000 55.210000 76.485000 ;
        RECT 55.010000 76.690000 55.210000 76.890000 ;
        RECT 55.010000 77.095000 55.210000 77.295000 ;
        RECT 55.010000 77.500000 55.210000 77.700000 ;
        RECT 55.010000 77.905000 55.210000 78.105000 ;
        RECT 55.010000 78.310000 55.210000 78.510000 ;
        RECT 55.010000 78.715000 55.210000 78.915000 ;
        RECT 55.010000 79.120000 55.210000 79.320000 ;
        RECT 55.010000 79.525000 55.210000 79.725000 ;
        RECT 55.010000 79.930000 55.210000 80.130000 ;
        RECT 55.010000 80.335000 55.210000 80.535000 ;
        RECT 55.010000 80.740000 55.210000 80.940000 ;
        RECT 55.010000 81.145000 55.210000 81.345000 ;
        RECT 55.010000 81.550000 55.210000 81.750000 ;
        RECT 55.010000 81.955000 55.210000 82.155000 ;
        RECT 55.010000 82.360000 55.210000 82.560000 ;
        RECT 55.255000 85.875000 55.455000 86.075000 ;
        RECT 55.255000 86.310000 55.455000 86.510000 ;
        RECT 55.255000 86.750000 55.455000 86.950000 ;
        RECT 55.300000 17.860000 55.500000 18.060000 ;
        RECT 55.300000 18.290000 55.500000 18.490000 ;
        RECT 55.300000 18.720000 55.500000 18.920000 ;
        RECT 55.300000 19.150000 55.500000 19.350000 ;
        RECT 55.300000 19.580000 55.500000 19.780000 ;
        RECT 55.300000 20.010000 55.500000 20.210000 ;
        RECT 55.300000 20.440000 55.500000 20.640000 ;
        RECT 55.300000 20.870000 55.500000 21.070000 ;
        RECT 55.300000 21.300000 55.500000 21.500000 ;
        RECT 55.300000 21.730000 55.500000 21.930000 ;
        RECT 55.300000 22.160000 55.500000 22.360000 ;
        RECT 55.325000 83.010000 55.525000 83.210000 ;
        RECT 55.325000 83.470000 55.525000 83.670000 ;
        RECT 55.325000 83.930000 55.525000 84.130000 ;
        RECT 55.325000 84.395000 55.525000 84.595000 ;
        RECT 55.325000 84.860000 55.525000 85.060000 ;
        RECT 55.325000 85.325000 55.525000 85.525000 ;
        RECT 55.410000 68.125000 55.610000 68.325000 ;
        RECT 55.410000 68.535000 55.610000 68.735000 ;
        RECT 55.410000 68.945000 55.610000 69.145000 ;
        RECT 55.410000 69.355000 55.610000 69.555000 ;
        RECT 55.410000 69.765000 55.610000 69.965000 ;
        RECT 55.410000 70.175000 55.610000 70.375000 ;
        RECT 55.410000 70.585000 55.610000 70.785000 ;
        RECT 55.410000 70.995000 55.610000 71.195000 ;
        RECT 55.410000 71.405000 55.610000 71.605000 ;
        RECT 55.410000 71.815000 55.610000 72.015000 ;
        RECT 55.410000 72.225000 55.610000 72.425000 ;
        RECT 55.410000 72.635000 55.610000 72.835000 ;
        RECT 55.410000 73.045000 55.610000 73.245000 ;
        RECT 55.410000 73.450000 55.610000 73.650000 ;
        RECT 55.410000 73.855000 55.610000 74.055000 ;
        RECT 55.410000 74.260000 55.610000 74.460000 ;
        RECT 55.410000 74.665000 55.610000 74.865000 ;
        RECT 55.410000 75.070000 55.610000 75.270000 ;
        RECT 55.410000 75.475000 55.610000 75.675000 ;
        RECT 55.410000 75.880000 55.610000 76.080000 ;
        RECT 55.410000 76.285000 55.610000 76.485000 ;
        RECT 55.410000 76.690000 55.610000 76.890000 ;
        RECT 55.410000 77.095000 55.610000 77.295000 ;
        RECT 55.410000 77.500000 55.610000 77.700000 ;
        RECT 55.410000 77.905000 55.610000 78.105000 ;
        RECT 55.410000 78.310000 55.610000 78.510000 ;
        RECT 55.410000 78.715000 55.610000 78.915000 ;
        RECT 55.410000 79.120000 55.610000 79.320000 ;
        RECT 55.410000 79.525000 55.610000 79.725000 ;
        RECT 55.410000 79.930000 55.610000 80.130000 ;
        RECT 55.410000 80.335000 55.610000 80.535000 ;
        RECT 55.410000 80.740000 55.610000 80.940000 ;
        RECT 55.410000 81.145000 55.610000 81.345000 ;
        RECT 55.410000 81.550000 55.610000 81.750000 ;
        RECT 55.410000 81.955000 55.610000 82.155000 ;
        RECT 55.410000 82.360000 55.610000 82.560000 ;
        RECT 55.705000 17.860000 55.905000 18.060000 ;
        RECT 55.705000 18.290000 55.905000 18.490000 ;
        RECT 55.705000 18.720000 55.905000 18.920000 ;
        RECT 55.705000 19.150000 55.905000 19.350000 ;
        RECT 55.705000 19.580000 55.905000 19.780000 ;
        RECT 55.705000 20.010000 55.905000 20.210000 ;
        RECT 55.705000 20.440000 55.905000 20.640000 ;
        RECT 55.705000 20.870000 55.905000 21.070000 ;
        RECT 55.705000 21.300000 55.905000 21.500000 ;
        RECT 55.705000 21.730000 55.905000 21.930000 ;
        RECT 55.705000 22.160000 55.905000 22.360000 ;
        RECT 55.805000 83.010000 56.005000 83.210000 ;
        RECT 55.805000 83.470000 56.005000 83.670000 ;
        RECT 55.805000 83.930000 56.005000 84.130000 ;
        RECT 55.805000 84.395000 56.005000 84.595000 ;
        RECT 55.805000 84.860000 56.005000 85.060000 ;
        RECT 55.805000 85.325000 56.005000 85.525000 ;
        RECT 55.810000 68.125000 56.010000 68.325000 ;
        RECT 55.810000 68.535000 56.010000 68.735000 ;
        RECT 55.810000 68.945000 56.010000 69.145000 ;
        RECT 55.810000 69.355000 56.010000 69.555000 ;
        RECT 55.810000 69.765000 56.010000 69.965000 ;
        RECT 55.810000 70.175000 56.010000 70.375000 ;
        RECT 55.810000 70.585000 56.010000 70.785000 ;
        RECT 55.810000 70.995000 56.010000 71.195000 ;
        RECT 55.810000 71.405000 56.010000 71.605000 ;
        RECT 55.810000 71.815000 56.010000 72.015000 ;
        RECT 55.810000 72.225000 56.010000 72.425000 ;
        RECT 55.810000 72.635000 56.010000 72.835000 ;
        RECT 55.810000 73.045000 56.010000 73.245000 ;
        RECT 55.810000 73.450000 56.010000 73.650000 ;
        RECT 55.810000 73.855000 56.010000 74.055000 ;
        RECT 55.810000 74.260000 56.010000 74.460000 ;
        RECT 55.810000 74.665000 56.010000 74.865000 ;
        RECT 55.810000 75.070000 56.010000 75.270000 ;
        RECT 55.810000 75.475000 56.010000 75.675000 ;
        RECT 55.810000 75.880000 56.010000 76.080000 ;
        RECT 55.810000 76.285000 56.010000 76.485000 ;
        RECT 55.810000 76.690000 56.010000 76.890000 ;
        RECT 55.810000 77.095000 56.010000 77.295000 ;
        RECT 55.810000 77.500000 56.010000 77.700000 ;
        RECT 55.810000 77.905000 56.010000 78.105000 ;
        RECT 55.810000 78.310000 56.010000 78.510000 ;
        RECT 55.810000 78.715000 56.010000 78.915000 ;
        RECT 55.810000 79.120000 56.010000 79.320000 ;
        RECT 55.810000 79.525000 56.010000 79.725000 ;
        RECT 55.810000 79.930000 56.010000 80.130000 ;
        RECT 55.810000 80.335000 56.010000 80.535000 ;
        RECT 55.810000 80.740000 56.010000 80.940000 ;
        RECT 55.810000 81.145000 56.010000 81.345000 ;
        RECT 55.810000 81.550000 56.010000 81.750000 ;
        RECT 55.810000 81.955000 56.010000 82.155000 ;
        RECT 55.810000 82.360000 56.010000 82.560000 ;
        RECT 55.995000 85.875000 56.195000 86.075000 ;
        RECT 55.995000 86.310000 56.195000 86.510000 ;
        RECT 55.995000 86.750000 56.195000 86.950000 ;
        RECT 56.110000 17.860000 56.310000 18.060000 ;
        RECT 56.110000 18.290000 56.310000 18.490000 ;
        RECT 56.110000 18.720000 56.310000 18.920000 ;
        RECT 56.110000 19.150000 56.310000 19.350000 ;
        RECT 56.110000 19.580000 56.310000 19.780000 ;
        RECT 56.110000 20.010000 56.310000 20.210000 ;
        RECT 56.110000 20.440000 56.310000 20.640000 ;
        RECT 56.110000 20.870000 56.310000 21.070000 ;
        RECT 56.110000 21.300000 56.310000 21.500000 ;
        RECT 56.110000 21.730000 56.310000 21.930000 ;
        RECT 56.110000 22.160000 56.310000 22.360000 ;
        RECT 56.210000 68.125000 56.410000 68.325000 ;
        RECT 56.210000 68.535000 56.410000 68.735000 ;
        RECT 56.210000 68.945000 56.410000 69.145000 ;
        RECT 56.210000 69.355000 56.410000 69.555000 ;
        RECT 56.210000 69.765000 56.410000 69.965000 ;
        RECT 56.210000 70.175000 56.410000 70.375000 ;
        RECT 56.210000 70.585000 56.410000 70.785000 ;
        RECT 56.210000 70.995000 56.410000 71.195000 ;
        RECT 56.210000 71.405000 56.410000 71.605000 ;
        RECT 56.210000 71.815000 56.410000 72.015000 ;
        RECT 56.210000 72.225000 56.410000 72.425000 ;
        RECT 56.210000 72.635000 56.410000 72.835000 ;
        RECT 56.210000 73.045000 56.410000 73.245000 ;
        RECT 56.210000 73.450000 56.410000 73.650000 ;
        RECT 56.210000 73.855000 56.410000 74.055000 ;
        RECT 56.210000 74.260000 56.410000 74.460000 ;
        RECT 56.210000 74.665000 56.410000 74.865000 ;
        RECT 56.210000 75.070000 56.410000 75.270000 ;
        RECT 56.210000 75.475000 56.410000 75.675000 ;
        RECT 56.210000 75.880000 56.410000 76.080000 ;
        RECT 56.210000 76.285000 56.410000 76.485000 ;
        RECT 56.210000 76.690000 56.410000 76.890000 ;
        RECT 56.210000 77.095000 56.410000 77.295000 ;
        RECT 56.210000 77.500000 56.410000 77.700000 ;
        RECT 56.210000 77.905000 56.410000 78.105000 ;
        RECT 56.210000 78.310000 56.410000 78.510000 ;
        RECT 56.210000 78.715000 56.410000 78.915000 ;
        RECT 56.210000 79.120000 56.410000 79.320000 ;
        RECT 56.210000 79.525000 56.410000 79.725000 ;
        RECT 56.210000 79.930000 56.410000 80.130000 ;
        RECT 56.210000 80.335000 56.410000 80.535000 ;
        RECT 56.210000 80.740000 56.410000 80.940000 ;
        RECT 56.210000 81.145000 56.410000 81.345000 ;
        RECT 56.210000 81.550000 56.410000 81.750000 ;
        RECT 56.210000 81.955000 56.410000 82.155000 ;
        RECT 56.210000 82.360000 56.410000 82.560000 ;
        RECT 56.490000 83.055000 56.690000 83.255000 ;
        RECT 56.490000 83.455000 56.690000 83.655000 ;
        RECT 56.490000 83.855000 56.690000 84.055000 ;
        RECT 56.490000 84.255000 56.690000 84.455000 ;
        RECT 56.490000 84.655000 56.690000 84.855000 ;
        RECT 56.490000 85.055000 56.690000 85.255000 ;
        RECT 56.490000 85.455000 56.690000 85.655000 ;
        RECT 56.490000 85.855000 56.690000 86.055000 ;
        RECT 56.490000 86.255000 56.690000 86.455000 ;
        RECT 56.490000 86.660000 56.690000 86.860000 ;
        RECT 56.490000 87.065000 56.690000 87.265000 ;
        RECT 56.490000 87.470000 56.690000 87.670000 ;
        RECT 56.490000 87.875000 56.690000 88.075000 ;
        RECT 56.515000 17.860000 56.715000 18.060000 ;
        RECT 56.515000 18.290000 56.715000 18.490000 ;
        RECT 56.515000 18.720000 56.715000 18.920000 ;
        RECT 56.515000 19.150000 56.715000 19.350000 ;
        RECT 56.515000 19.580000 56.715000 19.780000 ;
        RECT 56.515000 20.010000 56.715000 20.210000 ;
        RECT 56.515000 20.440000 56.715000 20.640000 ;
        RECT 56.515000 20.870000 56.715000 21.070000 ;
        RECT 56.515000 21.300000 56.715000 21.500000 ;
        RECT 56.515000 21.730000 56.715000 21.930000 ;
        RECT 56.515000 22.160000 56.715000 22.360000 ;
        RECT 56.610000 68.125000 56.810000 68.325000 ;
        RECT 56.610000 68.535000 56.810000 68.735000 ;
        RECT 56.610000 68.945000 56.810000 69.145000 ;
        RECT 56.610000 69.355000 56.810000 69.555000 ;
        RECT 56.610000 69.765000 56.810000 69.965000 ;
        RECT 56.610000 70.175000 56.810000 70.375000 ;
        RECT 56.610000 70.585000 56.810000 70.785000 ;
        RECT 56.610000 70.995000 56.810000 71.195000 ;
        RECT 56.610000 71.405000 56.810000 71.605000 ;
        RECT 56.610000 71.815000 56.810000 72.015000 ;
        RECT 56.610000 72.225000 56.810000 72.425000 ;
        RECT 56.610000 72.635000 56.810000 72.835000 ;
        RECT 56.610000 73.045000 56.810000 73.245000 ;
        RECT 56.610000 73.450000 56.810000 73.650000 ;
        RECT 56.610000 73.855000 56.810000 74.055000 ;
        RECT 56.610000 74.260000 56.810000 74.460000 ;
        RECT 56.610000 74.665000 56.810000 74.865000 ;
        RECT 56.610000 75.070000 56.810000 75.270000 ;
        RECT 56.610000 75.475000 56.810000 75.675000 ;
        RECT 56.610000 75.880000 56.810000 76.080000 ;
        RECT 56.610000 76.285000 56.810000 76.485000 ;
        RECT 56.610000 76.690000 56.810000 76.890000 ;
        RECT 56.610000 77.095000 56.810000 77.295000 ;
        RECT 56.610000 77.500000 56.810000 77.700000 ;
        RECT 56.610000 77.905000 56.810000 78.105000 ;
        RECT 56.610000 78.310000 56.810000 78.510000 ;
        RECT 56.610000 78.715000 56.810000 78.915000 ;
        RECT 56.610000 79.120000 56.810000 79.320000 ;
        RECT 56.610000 79.525000 56.810000 79.725000 ;
        RECT 56.610000 79.930000 56.810000 80.130000 ;
        RECT 56.610000 80.335000 56.810000 80.535000 ;
        RECT 56.610000 80.740000 56.810000 80.940000 ;
        RECT 56.610000 81.145000 56.810000 81.345000 ;
        RECT 56.610000 81.550000 56.810000 81.750000 ;
        RECT 56.610000 81.955000 56.810000 82.155000 ;
        RECT 56.610000 82.360000 56.810000 82.560000 ;
        RECT 56.900000 83.055000 57.100000 83.255000 ;
        RECT 56.900000 83.455000 57.100000 83.655000 ;
        RECT 56.900000 83.855000 57.100000 84.055000 ;
        RECT 56.900000 84.255000 57.100000 84.455000 ;
        RECT 56.900000 84.655000 57.100000 84.855000 ;
        RECT 56.900000 85.055000 57.100000 85.255000 ;
        RECT 56.900000 85.455000 57.100000 85.655000 ;
        RECT 56.900000 85.855000 57.100000 86.055000 ;
        RECT 56.900000 86.255000 57.100000 86.455000 ;
        RECT 56.900000 86.660000 57.100000 86.860000 ;
        RECT 56.900000 87.065000 57.100000 87.265000 ;
        RECT 56.900000 87.470000 57.100000 87.670000 ;
        RECT 56.900000 87.875000 57.100000 88.075000 ;
        RECT 56.920000 17.860000 57.120000 18.060000 ;
        RECT 56.920000 18.290000 57.120000 18.490000 ;
        RECT 56.920000 18.720000 57.120000 18.920000 ;
        RECT 56.920000 19.150000 57.120000 19.350000 ;
        RECT 56.920000 19.580000 57.120000 19.780000 ;
        RECT 56.920000 20.010000 57.120000 20.210000 ;
        RECT 56.920000 20.440000 57.120000 20.640000 ;
        RECT 56.920000 20.870000 57.120000 21.070000 ;
        RECT 56.920000 21.300000 57.120000 21.500000 ;
        RECT 56.920000 21.730000 57.120000 21.930000 ;
        RECT 56.920000 22.160000 57.120000 22.360000 ;
        RECT 57.010000 68.125000 57.210000 68.325000 ;
        RECT 57.010000 68.535000 57.210000 68.735000 ;
        RECT 57.010000 68.945000 57.210000 69.145000 ;
        RECT 57.010000 69.355000 57.210000 69.555000 ;
        RECT 57.010000 69.765000 57.210000 69.965000 ;
        RECT 57.010000 70.175000 57.210000 70.375000 ;
        RECT 57.010000 70.585000 57.210000 70.785000 ;
        RECT 57.010000 70.995000 57.210000 71.195000 ;
        RECT 57.010000 71.405000 57.210000 71.605000 ;
        RECT 57.010000 71.815000 57.210000 72.015000 ;
        RECT 57.010000 72.225000 57.210000 72.425000 ;
        RECT 57.010000 72.635000 57.210000 72.835000 ;
        RECT 57.010000 73.045000 57.210000 73.245000 ;
        RECT 57.010000 73.450000 57.210000 73.650000 ;
        RECT 57.010000 73.855000 57.210000 74.055000 ;
        RECT 57.010000 74.260000 57.210000 74.460000 ;
        RECT 57.010000 74.665000 57.210000 74.865000 ;
        RECT 57.010000 75.070000 57.210000 75.270000 ;
        RECT 57.010000 75.475000 57.210000 75.675000 ;
        RECT 57.010000 75.880000 57.210000 76.080000 ;
        RECT 57.010000 76.285000 57.210000 76.485000 ;
        RECT 57.010000 76.690000 57.210000 76.890000 ;
        RECT 57.010000 77.095000 57.210000 77.295000 ;
        RECT 57.010000 77.500000 57.210000 77.700000 ;
        RECT 57.010000 77.905000 57.210000 78.105000 ;
        RECT 57.010000 78.310000 57.210000 78.510000 ;
        RECT 57.010000 78.715000 57.210000 78.915000 ;
        RECT 57.010000 79.120000 57.210000 79.320000 ;
        RECT 57.010000 79.525000 57.210000 79.725000 ;
        RECT 57.010000 79.930000 57.210000 80.130000 ;
        RECT 57.010000 80.335000 57.210000 80.535000 ;
        RECT 57.010000 80.740000 57.210000 80.940000 ;
        RECT 57.010000 81.145000 57.210000 81.345000 ;
        RECT 57.010000 81.550000 57.210000 81.750000 ;
        RECT 57.010000 81.955000 57.210000 82.155000 ;
        RECT 57.010000 82.360000 57.210000 82.560000 ;
        RECT 57.310000 83.055000 57.510000 83.255000 ;
        RECT 57.310000 83.455000 57.510000 83.655000 ;
        RECT 57.310000 83.855000 57.510000 84.055000 ;
        RECT 57.310000 84.255000 57.510000 84.455000 ;
        RECT 57.310000 84.655000 57.510000 84.855000 ;
        RECT 57.310000 85.055000 57.510000 85.255000 ;
        RECT 57.310000 85.455000 57.510000 85.655000 ;
        RECT 57.310000 85.855000 57.510000 86.055000 ;
        RECT 57.310000 86.255000 57.510000 86.455000 ;
        RECT 57.310000 86.660000 57.510000 86.860000 ;
        RECT 57.310000 87.065000 57.510000 87.265000 ;
        RECT 57.310000 87.470000 57.510000 87.670000 ;
        RECT 57.310000 87.875000 57.510000 88.075000 ;
        RECT 57.325000 17.860000 57.525000 18.060000 ;
        RECT 57.325000 18.290000 57.525000 18.490000 ;
        RECT 57.325000 18.720000 57.525000 18.920000 ;
        RECT 57.325000 19.150000 57.525000 19.350000 ;
        RECT 57.325000 19.580000 57.525000 19.780000 ;
        RECT 57.325000 20.010000 57.525000 20.210000 ;
        RECT 57.325000 20.440000 57.525000 20.640000 ;
        RECT 57.325000 20.870000 57.525000 21.070000 ;
        RECT 57.325000 21.300000 57.525000 21.500000 ;
        RECT 57.325000 21.730000 57.525000 21.930000 ;
        RECT 57.325000 22.160000 57.525000 22.360000 ;
        RECT 57.410000 68.125000 57.610000 68.325000 ;
        RECT 57.410000 68.535000 57.610000 68.735000 ;
        RECT 57.410000 68.945000 57.610000 69.145000 ;
        RECT 57.410000 69.355000 57.610000 69.555000 ;
        RECT 57.410000 69.765000 57.610000 69.965000 ;
        RECT 57.410000 70.175000 57.610000 70.375000 ;
        RECT 57.410000 70.585000 57.610000 70.785000 ;
        RECT 57.410000 70.995000 57.610000 71.195000 ;
        RECT 57.410000 71.405000 57.610000 71.605000 ;
        RECT 57.410000 71.815000 57.610000 72.015000 ;
        RECT 57.410000 72.225000 57.610000 72.425000 ;
        RECT 57.410000 72.635000 57.610000 72.835000 ;
        RECT 57.410000 73.045000 57.610000 73.245000 ;
        RECT 57.410000 73.450000 57.610000 73.650000 ;
        RECT 57.410000 73.855000 57.610000 74.055000 ;
        RECT 57.410000 74.260000 57.610000 74.460000 ;
        RECT 57.410000 74.665000 57.610000 74.865000 ;
        RECT 57.410000 75.070000 57.610000 75.270000 ;
        RECT 57.410000 75.475000 57.610000 75.675000 ;
        RECT 57.410000 75.880000 57.610000 76.080000 ;
        RECT 57.410000 76.285000 57.610000 76.485000 ;
        RECT 57.410000 76.690000 57.610000 76.890000 ;
        RECT 57.410000 77.095000 57.610000 77.295000 ;
        RECT 57.410000 77.500000 57.610000 77.700000 ;
        RECT 57.410000 77.905000 57.610000 78.105000 ;
        RECT 57.410000 78.310000 57.610000 78.510000 ;
        RECT 57.410000 78.715000 57.610000 78.915000 ;
        RECT 57.410000 79.120000 57.610000 79.320000 ;
        RECT 57.410000 79.525000 57.610000 79.725000 ;
        RECT 57.410000 79.930000 57.610000 80.130000 ;
        RECT 57.410000 80.335000 57.610000 80.535000 ;
        RECT 57.410000 80.740000 57.610000 80.940000 ;
        RECT 57.410000 81.145000 57.610000 81.345000 ;
        RECT 57.410000 81.550000 57.610000 81.750000 ;
        RECT 57.410000 81.955000 57.610000 82.155000 ;
        RECT 57.410000 82.360000 57.610000 82.560000 ;
        RECT 57.720000 83.055000 57.920000 83.255000 ;
        RECT 57.720000 83.455000 57.920000 83.655000 ;
        RECT 57.720000 83.855000 57.920000 84.055000 ;
        RECT 57.720000 84.255000 57.920000 84.455000 ;
        RECT 57.720000 84.655000 57.920000 84.855000 ;
        RECT 57.720000 85.055000 57.920000 85.255000 ;
        RECT 57.720000 85.455000 57.920000 85.655000 ;
        RECT 57.720000 85.855000 57.920000 86.055000 ;
        RECT 57.720000 86.255000 57.920000 86.455000 ;
        RECT 57.720000 86.660000 57.920000 86.860000 ;
        RECT 57.720000 87.065000 57.920000 87.265000 ;
        RECT 57.720000 87.470000 57.920000 87.670000 ;
        RECT 57.720000 87.875000 57.920000 88.075000 ;
        RECT 57.730000 17.860000 57.930000 18.060000 ;
        RECT 57.730000 18.290000 57.930000 18.490000 ;
        RECT 57.730000 18.720000 57.930000 18.920000 ;
        RECT 57.730000 19.150000 57.930000 19.350000 ;
        RECT 57.730000 19.580000 57.930000 19.780000 ;
        RECT 57.730000 20.010000 57.930000 20.210000 ;
        RECT 57.730000 20.440000 57.930000 20.640000 ;
        RECT 57.730000 20.870000 57.930000 21.070000 ;
        RECT 57.730000 21.300000 57.930000 21.500000 ;
        RECT 57.730000 21.730000 57.930000 21.930000 ;
        RECT 57.730000 22.160000 57.930000 22.360000 ;
        RECT 57.795000 88.430000 57.995000 88.630000 ;
        RECT 57.795000 88.845000 57.995000 89.045000 ;
        RECT 57.795000 89.265000 57.995000 89.465000 ;
        RECT 57.810000 68.125000 58.010000 68.325000 ;
        RECT 57.810000 68.535000 58.010000 68.735000 ;
        RECT 57.810000 68.945000 58.010000 69.145000 ;
        RECT 57.810000 69.355000 58.010000 69.555000 ;
        RECT 57.810000 69.765000 58.010000 69.965000 ;
        RECT 57.810000 70.175000 58.010000 70.375000 ;
        RECT 57.810000 70.585000 58.010000 70.785000 ;
        RECT 57.810000 70.995000 58.010000 71.195000 ;
        RECT 57.810000 71.405000 58.010000 71.605000 ;
        RECT 57.810000 71.815000 58.010000 72.015000 ;
        RECT 57.810000 72.225000 58.010000 72.425000 ;
        RECT 57.810000 72.635000 58.010000 72.835000 ;
        RECT 57.810000 73.045000 58.010000 73.245000 ;
        RECT 57.810000 73.450000 58.010000 73.650000 ;
        RECT 57.810000 73.855000 58.010000 74.055000 ;
        RECT 57.810000 74.260000 58.010000 74.460000 ;
        RECT 57.810000 74.665000 58.010000 74.865000 ;
        RECT 57.810000 75.070000 58.010000 75.270000 ;
        RECT 57.810000 75.475000 58.010000 75.675000 ;
        RECT 57.810000 75.880000 58.010000 76.080000 ;
        RECT 57.810000 76.285000 58.010000 76.485000 ;
        RECT 57.810000 76.690000 58.010000 76.890000 ;
        RECT 57.810000 77.095000 58.010000 77.295000 ;
        RECT 57.810000 77.500000 58.010000 77.700000 ;
        RECT 57.810000 77.905000 58.010000 78.105000 ;
        RECT 57.810000 78.310000 58.010000 78.510000 ;
        RECT 57.810000 78.715000 58.010000 78.915000 ;
        RECT 57.810000 79.120000 58.010000 79.320000 ;
        RECT 57.810000 79.525000 58.010000 79.725000 ;
        RECT 57.810000 79.930000 58.010000 80.130000 ;
        RECT 57.810000 80.335000 58.010000 80.535000 ;
        RECT 57.810000 80.740000 58.010000 80.940000 ;
        RECT 57.810000 81.145000 58.010000 81.345000 ;
        RECT 57.810000 81.550000 58.010000 81.750000 ;
        RECT 57.810000 81.955000 58.010000 82.155000 ;
        RECT 57.810000 82.360000 58.010000 82.560000 ;
        RECT 58.130000 83.055000 58.330000 83.255000 ;
        RECT 58.130000 83.455000 58.330000 83.655000 ;
        RECT 58.130000 83.855000 58.330000 84.055000 ;
        RECT 58.130000 84.255000 58.330000 84.455000 ;
        RECT 58.130000 84.655000 58.330000 84.855000 ;
        RECT 58.130000 85.055000 58.330000 85.255000 ;
        RECT 58.130000 85.455000 58.330000 85.655000 ;
        RECT 58.130000 85.855000 58.330000 86.055000 ;
        RECT 58.130000 86.255000 58.330000 86.455000 ;
        RECT 58.130000 86.660000 58.330000 86.860000 ;
        RECT 58.130000 87.065000 58.330000 87.265000 ;
        RECT 58.130000 87.470000 58.330000 87.670000 ;
        RECT 58.130000 87.875000 58.330000 88.075000 ;
        RECT 58.135000 17.860000 58.335000 18.060000 ;
        RECT 58.135000 18.290000 58.335000 18.490000 ;
        RECT 58.135000 18.720000 58.335000 18.920000 ;
        RECT 58.135000 19.150000 58.335000 19.350000 ;
        RECT 58.135000 19.580000 58.335000 19.780000 ;
        RECT 58.135000 20.010000 58.335000 20.210000 ;
        RECT 58.135000 20.440000 58.335000 20.640000 ;
        RECT 58.135000 20.870000 58.335000 21.070000 ;
        RECT 58.135000 21.300000 58.335000 21.500000 ;
        RECT 58.135000 21.730000 58.335000 21.930000 ;
        RECT 58.135000 22.160000 58.335000 22.360000 ;
        RECT 58.210000 68.125000 58.410000 68.325000 ;
        RECT 58.210000 68.535000 58.410000 68.735000 ;
        RECT 58.210000 68.945000 58.410000 69.145000 ;
        RECT 58.210000 69.355000 58.410000 69.555000 ;
        RECT 58.210000 69.765000 58.410000 69.965000 ;
        RECT 58.210000 70.175000 58.410000 70.375000 ;
        RECT 58.210000 70.585000 58.410000 70.785000 ;
        RECT 58.210000 70.995000 58.410000 71.195000 ;
        RECT 58.210000 71.405000 58.410000 71.605000 ;
        RECT 58.210000 71.815000 58.410000 72.015000 ;
        RECT 58.210000 72.225000 58.410000 72.425000 ;
        RECT 58.210000 72.635000 58.410000 72.835000 ;
        RECT 58.210000 73.045000 58.410000 73.245000 ;
        RECT 58.210000 73.450000 58.410000 73.650000 ;
        RECT 58.210000 73.855000 58.410000 74.055000 ;
        RECT 58.210000 74.260000 58.410000 74.460000 ;
        RECT 58.210000 74.665000 58.410000 74.865000 ;
        RECT 58.210000 75.070000 58.410000 75.270000 ;
        RECT 58.210000 75.475000 58.410000 75.675000 ;
        RECT 58.210000 75.880000 58.410000 76.080000 ;
        RECT 58.210000 76.285000 58.410000 76.485000 ;
        RECT 58.210000 76.690000 58.410000 76.890000 ;
        RECT 58.210000 77.095000 58.410000 77.295000 ;
        RECT 58.210000 77.500000 58.410000 77.700000 ;
        RECT 58.210000 77.905000 58.410000 78.105000 ;
        RECT 58.210000 78.310000 58.410000 78.510000 ;
        RECT 58.210000 78.715000 58.410000 78.915000 ;
        RECT 58.210000 79.120000 58.410000 79.320000 ;
        RECT 58.210000 79.525000 58.410000 79.725000 ;
        RECT 58.210000 79.930000 58.410000 80.130000 ;
        RECT 58.210000 80.335000 58.410000 80.535000 ;
        RECT 58.210000 80.740000 58.410000 80.940000 ;
        RECT 58.210000 81.145000 58.410000 81.345000 ;
        RECT 58.210000 81.550000 58.410000 81.750000 ;
        RECT 58.210000 81.955000 58.410000 82.155000 ;
        RECT 58.210000 82.360000 58.410000 82.560000 ;
        RECT 58.540000 17.860000 58.740000 18.060000 ;
        RECT 58.540000 18.290000 58.740000 18.490000 ;
        RECT 58.540000 18.720000 58.740000 18.920000 ;
        RECT 58.540000 19.150000 58.740000 19.350000 ;
        RECT 58.540000 19.580000 58.740000 19.780000 ;
        RECT 58.540000 20.010000 58.740000 20.210000 ;
        RECT 58.540000 20.440000 58.740000 20.640000 ;
        RECT 58.540000 20.870000 58.740000 21.070000 ;
        RECT 58.540000 21.300000 58.740000 21.500000 ;
        RECT 58.540000 21.730000 58.740000 21.930000 ;
        RECT 58.540000 22.160000 58.740000 22.360000 ;
        RECT 58.540000 83.055000 58.740000 83.255000 ;
        RECT 58.540000 83.455000 58.740000 83.655000 ;
        RECT 58.540000 83.855000 58.740000 84.055000 ;
        RECT 58.540000 84.255000 58.740000 84.455000 ;
        RECT 58.540000 84.655000 58.740000 84.855000 ;
        RECT 58.540000 85.055000 58.740000 85.255000 ;
        RECT 58.540000 85.455000 58.740000 85.655000 ;
        RECT 58.540000 85.855000 58.740000 86.055000 ;
        RECT 58.540000 86.255000 58.740000 86.455000 ;
        RECT 58.540000 86.660000 58.740000 86.860000 ;
        RECT 58.540000 87.065000 58.740000 87.265000 ;
        RECT 58.540000 87.470000 58.740000 87.670000 ;
        RECT 58.540000 87.875000 58.740000 88.075000 ;
        RECT 58.575000 88.430000 58.775000 88.630000 ;
        RECT 58.575000 88.845000 58.775000 89.045000 ;
        RECT 58.575000 89.265000 58.775000 89.465000 ;
        RECT 58.610000 68.125000 58.810000 68.325000 ;
        RECT 58.610000 68.535000 58.810000 68.735000 ;
        RECT 58.610000 68.945000 58.810000 69.145000 ;
        RECT 58.610000 69.355000 58.810000 69.555000 ;
        RECT 58.610000 69.765000 58.810000 69.965000 ;
        RECT 58.610000 70.175000 58.810000 70.375000 ;
        RECT 58.610000 70.585000 58.810000 70.785000 ;
        RECT 58.610000 70.995000 58.810000 71.195000 ;
        RECT 58.610000 71.405000 58.810000 71.605000 ;
        RECT 58.610000 71.815000 58.810000 72.015000 ;
        RECT 58.610000 72.225000 58.810000 72.425000 ;
        RECT 58.610000 72.635000 58.810000 72.835000 ;
        RECT 58.610000 73.045000 58.810000 73.245000 ;
        RECT 58.610000 73.450000 58.810000 73.650000 ;
        RECT 58.610000 73.855000 58.810000 74.055000 ;
        RECT 58.610000 74.260000 58.810000 74.460000 ;
        RECT 58.610000 74.665000 58.810000 74.865000 ;
        RECT 58.610000 75.070000 58.810000 75.270000 ;
        RECT 58.610000 75.475000 58.810000 75.675000 ;
        RECT 58.610000 75.880000 58.810000 76.080000 ;
        RECT 58.610000 76.285000 58.810000 76.485000 ;
        RECT 58.610000 76.690000 58.810000 76.890000 ;
        RECT 58.610000 77.095000 58.810000 77.295000 ;
        RECT 58.610000 77.500000 58.810000 77.700000 ;
        RECT 58.610000 77.905000 58.810000 78.105000 ;
        RECT 58.610000 78.310000 58.810000 78.510000 ;
        RECT 58.610000 78.715000 58.810000 78.915000 ;
        RECT 58.610000 79.120000 58.810000 79.320000 ;
        RECT 58.610000 79.525000 58.810000 79.725000 ;
        RECT 58.610000 79.930000 58.810000 80.130000 ;
        RECT 58.610000 80.335000 58.810000 80.535000 ;
        RECT 58.610000 80.740000 58.810000 80.940000 ;
        RECT 58.610000 81.145000 58.810000 81.345000 ;
        RECT 58.610000 81.550000 58.810000 81.750000 ;
        RECT 58.610000 81.955000 58.810000 82.155000 ;
        RECT 58.610000 82.360000 58.810000 82.560000 ;
        RECT 58.945000 17.860000 59.145000 18.060000 ;
        RECT 58.945000 18.290000 59.145000 18.490000 ;
        RECT 58.945000 18.720000 59.145000 18.920000 ;
        RECT 58.945000 19.150000 59.145000 19.350000 ;
        RECT 58.945000 19.580000 59.145000 19.780000 ;
        RECT 58.945000 20.010000 59.145000 20.210000 ;
        RECT 58.945000 20.440000 59.145000 20.640000 ;
        RECT 58.945000 20.870000 59.145000 21.070000 ;
        RECT 58.945000 21.300000 59.145000 21.500000 ;
        RECT 58.945000 21.730000 59.145000 21.930000 ;
        RECT 58.945000 22.160000 59.145000 22.360000 ;
        RECT 58.950000 83.055000 59.150000 83.255000 ;
        RECT 58.950000 83.455000 59.150000 83.655000 ;
        RECT 58.950000 83.855000 59.150000 84.055000 ;
        RECT 58.950000 84.255000 59.150000 84.455000 ;
        RECT 58.950000 84.655000 59.150000 84.855000 ;
        RECT 58.950000 85.055000 59.150000 85.255000 ;
        RECT 58.950000 85.455000 59.150000 85.655000 ;
        RECT 58.950000 85.855000 59.150000 86.055000 ;
        RECT 58.950000 86.255000 59.150000 86.455000 ;
        RECT 58.950000 86.660000 59.150000 86.860000 ;
        RECT 58.950000 87.065000 59.150000 87.265000 ;
        RECT 58.950000 87.470000 59.150000 87.670000 ;
        RECT 58.950000 87.875000 59.150000 88.075000 ;
        RECT 59.010000 68.125000 59.210000 68.325000 ;
        RECT 59.010000 68.535000 59.210000 68.735000 ;
        RECT 59.010000 68.945000 59.210000 69.145000 ;
        RECT 59.010000 69.355000 59.210000 69.555000 ;
        RECT 59.010000 69.765000 59.210000 69.965000 ;
        RECT 59.010000 70.175000 59.210000 70.375000 ;
        RECT 59.010000 70.585000 59.210000 70.785000 ;
        RECT 59.010000 70.995000 59.210000 71.195000 ;
        RECT 59.010000 71.405000 59.210000 71.605000 ;
        RECT 59.010000 71.815000 59.210000 72.015000 ;
        RECT 59.010000 72.225000 59.210000 72.425000 ;
        RECT 59.010000 72.635000 59.210000 72.835000 ;
        RECT 59.010000 73.045000 59.210000 73.245000 ;
        RECT 59.010000 73.450000 59.210000 73.650000 ;
        RECT 59.010000 73.855000 59.210000 74.055000 ;
        RECT 59.010000 74.260000 59.210000 74.460000 ;
        RECT 59.010000 74.665000 59.210000 74.865000 ;
        RECT 59.010000 75.070000 59.210000 75.270000 ;
        RECT 59.010000 75.475000 59.210000 75.675000 ;
        RECT 59.010000 75.880000 59.210000 76.080000 ;
        RECT 59.010000 76.285000 59.210000 76.485000 ;
        RECT 59.010000 76.690000 59.210000 76.890000 ;
        RECT 59.010000 77.095000 59.210000 77.295000 ;
        RECT 59.010000 77.500000 59.210000 77.700000 ;
        RECT 59.010000 77.905000 59.210000 78.105000 ;
        RECT 59.010000 78.310000 59.210000 78.510000 ;
        RECT 59.010000 78.715000 59.210000 78.915000 ;
        RECT 59.010000 79.120000 59.210000 79.320000 ;
        RECT 59.010000 79.525000 59.210000 79.725000 ;
        RECT 59.010000 79.930000 59.210000 80.130000 ;
        RECT 59.010000 80.335000 59.210000 80.535000 ;
        RECT 59.010000 80.740000 59.210000 80.940000 ;
        RECT 59.010000 81.145000 59.210000 81.345000 ;
        RECT 59.010000 81.550000 59.210000 81.750000 ;
        RECT 59.010000 81.955000 59.210000 82.155000 ;
        RECT 59.010000 82.360000 59.210000 82.560000 ;
        RECT 59.075000 88.410000 59.275000 88.610000 ;
        RECT 59.075000 88.835000 59.275000 89.035000 ;
        RECT 59.075000 89.265000 59.275000 89.465000 ;
        RECT 59.075000 89.695000 59.275000 89.895000 ;
        RECT 59.075000 90.125000 59.275000 90.325000 ;
        RECT 59.075000 90.555000 59.275000 90.755000 ;
        RECT 59.350000 17.860000 59.550000 18.060000 ;
        RECT 59.350000 18.290000 59.550000 18.490000 ;
        RECT 59.350000 18.720000 59.550000 18.920000 ;
        RECT 59.350000 19.150000 59.550000 19.350000 ;
        RECT 59.350000 19.580000 59.550000 19.780000 ;
        RECT 59.350000 20.010000 59.550000 20.210000 ;
        RECT 59.350000 20.440000 59.550000 20.640000 ;
        RECT 59.350000 20.870000 59.550000 21.070000 ;
        RECT 59.350000 21.300000 59.550000 21.500000 ;
        RECT 59.350000 21.730000 59.550000 21.930000 ;
        RECT 59.350000 22.160000 59.550000 22.360000 ;
        RECT 59.360000 83.055000 59.560000 83.255000 ;
        RECT 59.360000 83.455000 59.560000 83.655000 ;
        RECT 59.360000 83.855000 59.560000 84.055000 ;
        RECT 59.360000 84.255000 59.560000 84.455000 ;
        RECT 59.360000 84.655000 59.560000 84.855000 ;
        RECT 59.360000 85.055000 59.560000 85.255000 ;
        RECT 59.360000 85.455000 59.560000 85.655000 ;
        RECT 59.360000 85.855000 59.560000 86.055000 ;
        RECT 59.360000 86.255000 59.560000 86.455000 ;
        RECT 59.360000 86.660000 59.560000 86.860000 ;
        RECT 59.360000 87.065000 59.560000 87.265000 ;
        RECT 59.360000 87.470000 59.560000 87.670000 ;
        RECT 59.360000 87.875000 59.560000 88.075000 ;
        RECT 59.410000 68.125000 59.610000 68.325000 ;
        RECT 59.410000 68.535000 59.610000 68.735000 ;
        RECT 59.410000 68.945000 59.610000 69.145000 ;
        RECT 59.410000 69.355000 59.610000 69.555000 ;
        RECT 59.410000 69.765000 59.610000 69.965000 ;
        RECT 59.410000 70.175000 59.610000 70.375000 ;
        RECT 59.410000 70.585000 59.610000 70.785000 ;
        RECT 59.410000 70.995000 59.610000 71.195000 ;
        RECT 59.410000 71.405000 59.610000 71.605000 ;
        RECT 59.410000 71.815000 59.610000 72.015000 ;
        RECT 59.410000 72.225000 59.610000 72.425000 ;
        RECT 59.410000 72.635000 59.610000 72.835000 ;
        RECT 59.410000 73.045000 59.610000 73.245000 ;
        RECT 59.410000 73.450000 59.610000 73.650000 ;
        RECT 59.410000 73.855000 59.610000 74.055000 ;
        RECT 59.410000 74.260000 59.610000 74.460000 ;
        RECT 59.410000 74.665000 59.610000 74.865000 ;
        RECT 59.410000 75.070000 59.610000 75.270000 ;
        RECT 59.410000 75.475000 59.610000 75.675000 ;
        RECT 59.410000 75.880000 59.610000 76.080000 ;
        RECT 59.410000 76.285000 59.610000 76.485000 ;
        RECT 59.410000 76.690000 59.610000 76.890000 ;
        RECT 59.410000 77.095000 59.610000 77.295000 ;
        RECT 59.410000 77.500000 59.610000 77.700000 ;
        RECT 59.410000 77.905000 59.610000 78.105000 ;
        RECT 59.410000 78.310000 59.610000 78.510000 ;
        RECT 59.410000 78.715000 59.610000 78.915000 ;
        RECT 59.410000 79.120000 59.610000 79.320000 ;
        RECT 59.410000 79.525000 59.610000 79.725000 ;
        RECT 59.410000 79.930000 59.610000 80.130000 ;
        RECT 59.410000 80.335000 59.610000 80.535000 ;
        RECT 59.410000 80.740000 59.610000 80.940000 ;
        RECT 59.410000 81.145000 59.610000 81.345000 ;
        RECT 59.410000 81.550000 59.610000 81.750000 ;
        RECT 59.410000 81.955000 59.610000 82.155000 ;
        RECT 59.410000 82.360000 59.610000 82.560000 ;
        RECT 59.485000 88.410000 59.685000 88.610000 ;
        RECT 59.485000 88.835000 59.685000 89.035000 ;
        RECT 59.485000 89.265000 59.685000 89.465000 ;
        RECT 59.485000 89.695000 59.685000 89.895000 ;
        RECT 59.485000 90.125000 59.685000 90.325000 ;
        RECT 59.485000 90.555000 59.685000 90.755000 ;
        RECT 59.755000 17.860000 59.955000 18.060000 ;
        RECT 59.755000 18.290000 59.955000 18.490000 ;
        RECT 59.755000 18.720000 59.955000 18.920000 ;
        RECT 59.755000 19.150000 59.955000 19.350000 ;
        RECT 59.755000 19.580000 59.955000 19.780000 ;
        RECT 59.755000 20.010000 59.955000 20.210000 ;
        RECT 59.755000 20.440000 59.955000 20.640000 ;
        RECT 59.755000 20.870000 59.955000 21.070000 ;
        RECT 59.755000 21.300000 59.955000 21.500000 ;
        RECT 59.755000 21.730000 59.955000 21.930000 ;
        RECT 59.755000 22.160000 59.955000 22.360000 ;
        RECT 59.770000 83.055000 59.970000 83.255000 ;
        RECT 59.770000 83.455000 59.970000 83.655000 ;
        RECT 59.770000 83.855000 59.970000 84.055000 ;
        RECT 59.770000 84.255000 59.970000 84.455000 ;
        RECT 59.770000 84.655000 59.970000 84.855000 ;
        RECT 59.770000 85.055000 59.970000 85.255000 ;
        RECT 59.770000 85.455000 59.970000 85.655000 ;
        RECT 59.770000 85.855000 59.970000 86.055000 ;
        RECT 59.770000 86.255000 59.970000 86.455000 ;
        RECT 59.770000 86.660000 59.970000 86.860000 ;
        RECT 59.770000 87.065000 59.970000 87.265000 ;
        RECT 59.770000 87.470000 59.970000 87.670000 ;
        RECT 59.770000 87.875000 59.970000 88.075000 ;
        RECT 59.810000 68.125000 60.010000 68.325000 ;
        RECT 59.810000 68.535000 60.010000 68.735000 ;
        RECT 59.810000 68.945000 60.010000 69.145000 ;
        RECT 59.810000 69.355000 60.010000 69.555000 ;
        RECT 59.810000 69.765000 60.010000 69.965000 ;
        RECT 59.810000 70.175000 60.010000 70.375000 ;
        RECT 59.810000 70.585000 60.010000 70.785000 ;
        RECT 59.810000 70.995000 60.010000 71.195000 ;
        RECT 59.810000 71.405000 60.010000 71.605000 ;
        RECT 59.810000 71.815000 60.010000 72.015000 ;
        RECT 59.810000 72.225000 60.010000 72.425000 ;
        RECT 59.810000 72.635000 60.010000 72.835000 ;
        RECT 59.810000 73.045000 60.010000 73.245000 ;
        RECT 59.810000 73.450000 60.010000 73.650000 ;
        RECT 59.810000 73.855000 60.010000 74.055000 ;
        RECT 59.810000 74.260000 60.010000 74.460000 ;
        RECT 59.810000 74.665000 60.010000 74.865000 ;
        RECT 59.810000 75.070000 60.010000 75.270000 ;
        RECT 59.810000 75.475000 60.010000 75.675000 ;
        RECT 59.810000 75.880000 60.010000 76.080000 ;
        RECT 59.810000 76.285000 60.010000 76.485000 ;
        RECT 59.810000 76.690000 60.010000 76.890000 ;
        RECT 59.810000 77.095000 60.010000 77.295000 ;
        RECT 59.810000 77.500000 60.010000 77.700000 ;
        RECT 59.810000 77.905000 60.010000 78.105000 ;
        RECT 59.810000 78.310000 60.010000 78.510000 ;
        RECT 59.810000 78.715000 60.010000 78.915000 ;
        RECT 59.810000 79.120000 60.010000 79.320000 ;
        RECT 59.810000 79.525000 60.010000 79.725000 ;
        RECT 59.810000 79.930000 60.010000 80.130000 ;
        RECT 59.810000 80.335000 60.010000 80.535000 ;
        RECT 59.810000 80.740000 60.010000 80.940000 ;
        RECT 59.810000 81.145000 60.010000 81.345000 ;
        RECT 59.810000 81.550000 60.010000 81.750000 ;
        RECT 59.810000 81.955000 60.010000 82.155000 ;
        RECT 59.810000 82.360000 60.010000 82.560000 ;
        RECT 59.895000 88.410000 60.095000 88.610000 ;
        RECT 59.895000 88.835000 60.095000 89.035000 ;
        RECT 59.895000 89.265000 60.095000 89.465000 ;
        RECT 59.895000 89.695000 60.095000 89.895000 ;
        RECT 59.895000 90.125000 60.095000 90.325000 ;
        RECT 59.895000 90.555000 60.095000 90.755000 ;
        RECT 59.955000 91.015000 60.155000 91.215000 ;
        RECT 59.955000 91.445000 60.155000 91.645000 ;
        RECT 60.160000 17.860000 60.360000 18.060000 ;
        RECT 60.160000 18.290000 60.360000 18.490000 ;
        RECT 60.160000 18.720000 60.360000 18.920000 ;
        RECT 60.160000 19.150000 60.360000 19.350000 ;
        RECT 60.160000 19.580000 60.360000 19.780000 ;
        RECT 60.160000 20.010000 60.360000 20.210000 ;
        RECT 60.160000 20.440000 60.360000 20.640000 ;
        RECT 60.160000 20.870000 60.360000 21.070000 ;
        RECT 60.160000 21.300000 60.360000 21.500000 ;
        RECT 60.160000 21.730000 60.360000 21.930000 ;
        RECT 60.160000 22.160000 60.360000 22.360000 ;
        RECT 60.180000 83.055000 60.380000 83.255000 ;
        RECT 60.180000 83.455000 60.380000 83.655000 ;
        RECT 60.180000 83.855000 60.380000 84.055000 ;
        RECT 60.180000 84.255000 60.380000 84.455000 ;
        RECT 60.180000 84.655000 60.380000 84.855000 ;
        RECT 60.180000 85.055000 60.380000 85.255000 ;
        RECT 60.180000 85.455000 60.380000 85.655000 ;
        RECT 60.180000 85.855000 60.380000 86.055000 ;
        RECT 60.180000 86.255000 60.380000 86.455000 ;
        RECT 60.180000 86.660000 60.380000 86.860000 ;
        RECT 60.180000 87.065000 60.380000 87.265000 ;
        RECT 60.180000 87.470000 60.380000 87.670000 ;
        RECT 60.180000 87.875000 60.380000 88.075000 ;
        RECT 60.210000 68.125000 60.410000 68.325000 ;
        RECT 60.210000 68.535000 60.410000 68.735000 ;
        RECT 60.210000 68.945000 60.410000 69.145000 ;
        RECT 60.210000 69.355000 60.410000 69.555000 ;
        RECT 60.210000 69.765000 60.410000 69.965000 ;
        RECT 60.210000 70.175000 60.410000 70.375000 ;
        RECT 60.210000 70.585000 60.410000 70.785000 ;
        RECT 60.210000 70.995000 60.410000 71.195000 ;
        RECT 60.210000 71.405000 60.410000 71.605000 ;
        RECT 60.210000 71.815000 60.410000 72.015000 ;
        RECT 60.210000 72.225000 60.410000 72.425000 ;
        RECT 60.210000 72.635000 60.410000 72.835000 ;
        RECT 60.210000 73.045000 60.410000 73.245000 ;
        RECT 60.210000 73.450000 60.410000 73.650000 ;
        RECT 60.210000 73.855000 60.410000 74.055000 ;
        RECT 60.210000 74.260000 60.410000 74.460000 ;
        RECT 60.210000 74.665000 60.410000 74.865000 ;
        RECT 60.210000 75.070000 60.410000 75.270000 ;
        RECT 60.210000 75.475000 60.410000 75.675000 ;
        RECT 60.210000 75.880000 60.410000 76.080000 ;
        RECT 60.210000 76.285000 60.410000 76.485000 ;
        RECT 60.210000 76.690000 60.410000 76.890000 ;
        RECT 60.210000 77.095000 60.410000 77.295000 ;
        RECT 60.210000 77.500000 60.410000 77.700000 ;
        RECT 60.210000 77.905000 60.410000 78.105000 ;
        RECT 60.210000 78.310000 60.410000 78.510000 ;
        RECT 60.210000 78.715000 60.410000 78.915000 ;
        RECT 60.210000 79.120000 60.410000 79.320000 ;
        RECT 60.210000 79.525000 60.410000 79.725000 ;
        RECT 60.210000 79.930000 60.410000 80.130000 ;
        RECT 60.210000 80.335000 60.410000 80.535000 ;
        RECT 60.210000 80.740000 60.410000 80.940000 ;
        RECT 60.210000 81.145000 60.410000 81.345000 ;
        RECT 60.210000 81.550000 60.410000 81.750000 ;
        RECT 60.210000 81.955000 60.410000 82.155000 ;
        RECT 60.210000 82.360000 60.410000 82.560000 ;
        RECT 60.305000 88.410000 60.505000 88.610000 ;
        RECT 60.305000 88.835000 60.505000 89.035000 ;
        RECT 60.305000 89.265000 60.505000 89.465000 ;
        RECT 60.305000 89.695000 60.505000 89.895000 ;
        RECT 60.305000 90.125000 60.505000 90.325000 ;
        RECT 60.305000 90.555000 60.505000 90.755000 ;
        RECT 60.565000 17.860000 60.765000 18.060000 ;
        RECT 60.565000 18.290000 60.765000 18.490000 ;
        RECT 60.565000 18.720000 60.765000 18.920000 ;
        RECT 60.565000 19.150000 60.765000 19.350000 ;
        RECT 60.565000 19.580000 60.765000 19.780000 ;
        RECT 60.565000 20.010000 60.765000 20.210000 ;
        RECT 60.565000 20.440000 60.765000 20.640000 ;
        RECT 60.565000 20.870000 60.765000 21.070000 ;
        RECT 60.565000 21.300000 60.765000 21.500000 ;
        RECT 60.565000 21.730000 60.765000 21.930000 ;
        RECT 60.565000 22.160000 60.765000 22.360000 ;
        RECT 60.590000 83.055000 60.790000 83.255000 ;
        RECT 60.590000 83.455000 60.790000 83.655000 ;
        RECT 60.590000 83.855000 60.790000 84.055000 ;
        RECT 60.590000 84.255000 60.790000 84.455000 ;
        RECT 60.590000 84.655000 60.790000 84.855000 ;
        RECT 60.590000 85.055000 60.790000 85.255000 ;
        RECT 60.590000 85.455000 60.790000 85.655000 ;
        RECT 60.590000 85.855000 60.790000 86.055000 ;
        RECT 60.590000 86.255000 60.790000 86.455000 ;
        RECT 60.590000 86.660000 60.790000 86.860000 ;
        RECT 60.590000 87.065000 60.790000 87.265000 ;
        RECT 60.590000 87.470000 60.790000 87.670000 ;
        RECT 60.590000 87.875000 60.790000 88.075000 ;
        RECT 60.610000 68.125000 60.810000 68.325000 ;
        RECT 60.610000 68.535000 60.810000 68.735000 ;
        RECT 60.610000 68.945000 60.810000 69.145000 ;
        RECT 60.610000 69.355000 60.810000 69.555000 ;
        RECT 60.610000 69.765000 60.810000 69.965000 ;
        RECT 60.610000 70.175000 60.810000 70.375000 ;
        RECT 60.610000 70.585000 60.810000 70.785000 ;
        RECT 60.610000 70.995000 60.810000 71.195000 ;
        RECT 60.610000 71.405000 60.810000 71.605000 ;
        RECT 60.610000 71.815000 60.810000 72.015000 ;
        RECT 60.610000 72.225000 60.810000 72.425000 ;
        RECT 60.610000 72.635000 60.810000 72.835000 ;
        RECT 60.610000 73.045000 60.810000 73.245000 ;
        RECT 60.610000 73.450000 60.810000 73.650000 ;
        RECT 60.610000 73.855000 60.810000 74.055000 ;
        RECT 60.610000 74.260000 60.810000 74.460000 ;
        RECT 60.610000 74.665000 60.810000 74.865000 ;
        RECT 60.610000 75.070000 60.810000 75.270000 ;
        RECT 60.610000 75.475000 60.810000 75.675000 ;
        RECT 60.610000 75.880000 60.810000 76.080000 ;
        RECT 60.610000 76.285000 60.810000 76.485000 ;
        RECT 60.610000 76.690000 60.810000 76.890000 ;
        RECT 60.610000 77.095000 60.810000 77.295000 ;
        RECT 60.610000 77.500000 60.810000 77.700000 ;
        RECT 60.610000 77.905000 60.810000 78.105000 ;
        RECT 60.610000 78.310000 60.810000 78.510000 ;
        RECT 60.610000 78.715000 60.810000 78.915000 ;
        RECT 60.610000 79.120000 60.810000 79.320000 ;
        RECT 60.610000 79.525000 60.810000 79.725000 ;
        RECT 60.610000 79.930000 60.810000 80.130000 ;
        RECT 60.610000 80.335000 60.810000 80.535000 ;
        RECT 60.610000 80.740000 60.810000 80.940000 ;
        RECT 60.610000 81.145000 60.810000 81.345000 ;
        RECT 60.610000 81.550000 60.810000 81.750000 ;
        RECT 60.610000 81.955000 60.810000 82.155000 ;
        RECT 60.610000 82.360000 60.810000 82.560000 ;
        RECT 60.715000 88.410000 60.915000 88.610000 ;
        RECT 60.715000 88.835000 60.915000 89.035000 ;
        RECT 60.715000 89.265000 60.915000 89.465000 ;
        RECT 60.715000 89.695000 60.915000 89.895000 ;
        RECT 60.715000 90.125000 60.915000 90.325000 ;
        RECT 60.715000 90.555000 60.915000 90.755000 ;
        RECT 60.735000 91.015000 60.935000 91.215000 ;
        RECT 60.735000 91.445000 60.935000 91.645000 ;
        RECT 60.970000 17.860000 61.170000 18.060000 ;
        RECT 60.970000 18.290000 61.170000 18.490000 ;
        RECT 60.970000 18.720000 61.170000 18.920000 ;
        RECT 60.970000 19.150000 61.170000 19.350000 ;
        RECT 60.970000 19.580000 61.170000 19.780000 ;
        RECT 60.970000 20.010000 61.170000 20.210000 ;
        RECT 60.970000 20.440000 61.170000 20.640000 ;
        RECT 60.970000 20.870000 61.170000 21.070000 ;
        RECT 60.970000 21.300000 61.170000 21.500000 ;
        RECT 60.970000 21.730000 61.170000 21.930000 ;
        RECT 60.970000 22.160000 61.170000 22.360000 ;
        RECT 61.010000 68.125000 61.210000 68.325000 ;
        RECT 61.010000 68.535000 61.210000 68.735000 ;
        RECT 61.010000 68.945000 61.210000 69.145000 ;
        RECT 61.010000 69.355000 61.210000 69.555000 ;
        RECT 61.010000 69.765000 61.210000 69.965000 ;
        RECT 61.010000 70.175000 61.210000 70.375000 ;
        RECT 61.010000 70.585000 61.210000 70.785000 ;
        RECT 61.010000 70.995000 61.210000 71.195000 ;
        RECT 61.010000 71.405000 61.210000 71.605000 ;
        RECT 61.010000 71.815000 61.210000 72.015000 ;
        RECT 61.010000 72.225000 61.210000 72.425000 ;
        RECT 61.010000 72.635000 61.210000 72.835000 ;
        RECT 61.010000 73.045000 61.210000 73.245000 ;
        RECT 61.010000 73.450000 61.210000 73.650000 ;
        RECT 61.010000 73.855000 61.210000 74.055000 ;
        RECT 61.010000 74.260000 61.210000 74.460000 ;
        RECT 61.010000 74.665000 61.210000 74.865000 ;
        RECT 61.010000 75.070000 61.210000 75.270000 ;
        RECT 61.010000 75.475000 61.210000 75.675000 ;
        RECT 61.010000 75.880000 61.210000 76.080000 ;
        RECT 61.010000 76.285000 61.210000 76.485000 ;
        RECT 61.010000 76.690000 61.210000 76.890000 ;
        RECT 61.010000 77.095000 61.210000 77.295000 ;
        RECT 61.010000 77.500000 61.210000 77.700000 ;
        RECT 61.010000 77.905000 61.210000 78.105000 ;
        RECT 61.010000 78.310000 61.210000 78.510000 ;
        RECT 61.010000 78.715000 61.210000 78.915000 ;
        RECT 61.010000 79.120000 61.210000 79.320000 ;
        RECT 61.010000 79.525000 61.210000 79.725000 ;
        RECT 61.010000 79.930000 61.210000 80.130000 ;
        RECT 61.010000 80.335000 61.210000 80.535000 ;
        RECT 61.010000 80.740000 61.210000 80.940000 ;
        RECT 61.010000 81.145000 61.210000 81.345000 ;
        RECT 61.010000 81.550000 61.210000 81.750000 ;
        RECT 61.010000 81.955000 61.210000 82.155000 ;
        RECT 61.010000 82.360000 61.210000 82.560000 ;
        RECT 61.215000 82.855000 61.415000 83.055000 ;
        RECT 61.215000 83.265000 61.415000 83.465000 ;
        RECT 61.215000 83.675000 61.415000 83.875000 ;
        RECT 61.215000 84.085000 61.415000 84.285000 ;
        RECT 61.215000 84.495000 61.415000 84.695000 ;
        RECT 61.215000 84.905000 61.415000 85.105000 ;
        RECT 61.215000 85.315000 61.415000 85.515000 ;
        RECT 61.215000 85.725000 61.415000 85.925000 ;
        RECT 61.215000 86.135000 61.415000 86.335000 ;
        RECT 61.215000 86.545000 61.415000 86.745000 ;
        RECT 61.215000 86.955000 61.415000 87.155000 ;
        RECT 61.215000 87.365000 61.415000 87.565000 ;
        RECT 61.215000 87.775000 61.415000 87.975000 ;
        RECT 61.215000 88.185000 61.415000 88.385000 ;
        RECT 61.215000 88.595000 61.415000 88.795000 ;
        RECT 61.215000 89.005000 61.415000 89.205000 ;
        RECT 61.215000 89.415000 61.415000 89.615000 ;
        RECT 61.215000 89.825000 61.415000 90.025000 ;
        RECT 61.215000 90.235000 61.415000 90.435000 ;
        RECT 61.215000 90.645000 61.415000 90.845000 ;
        RECT 61.215000 91.055000 61.415000 91.255000 ;
        RECT 61.215000 91.465000 61.415000 91.665000 ;
        RECT 61.215000 91.875000 61.415000 92.075000 ;
        RECT 61.215000 92.285000 61.415000 92.485000 ;
        RECT 61.215000 92.695000 61.415000 92.895000 ;
        RECT 61.375000 17.860000 61.575000 18.060000 ;
        RECT 61.375000 18.290000 61.575000 18.490000 ;
        RECT 61.375000 18.720000 61.575000 18.920000 ;
        RECT 61.375000 19.150000 61.575000 19.350000 ;
        RECT 61.375000 19.580000 61.575000 19.780000 ;
        RECT 61.375000 20.010000 61.575000 20.210000 ;
        RECT 61.375000 20.440000 61.575000 20.640000 ;
        RECT 61.375000 20.870000 61.575000 21.070000 ;
        RECT 61.375000 21.300000 61.575000 21.500000 ;
        RECT 61.375000 21.730000 61.575000 21.930000 ;
        RECT 61.375000 22.160000 61.575000 22.360000 ;
        RECT 61.410000 68.125000 61.610000 68.325000 ;
        RECT 61.410000 68.535000 61.610000 68.735000 ;
        RECT 61.410000 68.945000 61.610000 69.145000 ;
        RECT 61.410000 69.355000 61.610000 69.555000 ;
        RECT 61.410000 69.765000 61.610000 69.965000 ;
        RECT 61.410000 70.175000 61.610000 70.375000 ;
        RECT 61.410000 70.585000 61.610000 70.785000 ;
        RECT 61.410000 70.995000 61.610000 71.195000 ;
        RECT 61.410000 71.405000 61.610000 71.605000 ;
        RECT 61.410000 71.815000 61.610000 72.015000 ;
        RECT 61.410000 72.225000 61.610000 72.425000 ;
        RECT 61.410000 72.635000 61.610000 72.835000 ;
        RECT 61.410000 73.045000 61.610000 73.245000 ;
        RECT 61.410000 73.450000 61.610000 73.650000 ;
        RECT 61.410000 73.855000 61.610000 74.055000 ;
        RECT 61.410000 74.260000 61.610000 74.460000 ;
        RECT 61.410000 74.665000 61.610000 74.865000 ;
        RECT 61.410000 75.070000 61.610000 75.270000 ;
        RECT 61.410000 75.475000 61.610000 75.675000 ;
        RECT 61.410000 75.880000 61.610000 76.080000 ;
        RECT 61.410000 76.285000 61.610000 76.485000 ;
        RECT 61.410000 76.690000 61.610000 76.890000 ;
        RECT 61.410000 77.095000 61.610000 77.295000 ;
        RECT 61.410000 77.500000 61.610000 77.700000 ;
        RECT 61.410000 77.905000 61.610000 78.105000 ;
        RECT 61.410000 78.310000 61.610000 78.510000 ;
        RECT 61.410000 78.715000 61.610000 78.915000 ;
        RECT 61.410000 79.120000 61.610000 79.320000 ;
        RECT 61.410000 79.525000 61.610000 79.725000 ;
        RECT 61.410000 79.930000 61.610000 80.130000 ;
        RECT 61.410000 80.335000 61.610000 80.535000 ;
        RECT 61.410000 80.740000 61.610000 80.940000 ;
        RECT 61.410000 81.145000 61.610000 81.345000 ;
        RECT 61.410000 81.550000 61.610000 81.750000 ;
        RECT 61.410000 81.955000 61.610000 82.155000 ;
        RECT 61.410000 82.360000 61.610000 82.560000 ;
        RECT 61.620000 82.855000 61.820000 83.055000 ;
        RECT 61.620000 83.265000 61.820000 83.465000 ;
        RECT 61.620000 83.675000 61.820000 83.875000 ;
        RECT 61.620000 84.085000 61.820000 84.285000 ;
        RECT 61.620000 84.495000 61.820000 84.695000 ;
        RECT 61.620000 84.905000 61.820000 85.105000 ;
        RECT 61.620000 85.315000 61.820000 85.515000 ;
        RECT 61.620000 85.725000 61.820000 85.925000 ;
        RECT 61.620000 86.135000 61.820000 86.335000 ;
        RECT 61.620000 86.545000 61.820000 86.745000 ;
        RECT 61.620000 86.955000 61.820000 87.155000 ;
        RECT 61.620000 87.365000 61.820000 87.565000 ;
        RECT 61.620000 87.775000 61.820000 87.975000 ;
        RECT 61.620000 88.185000 61.820000 88.385000 ;
        RECT 61.620000 88.595000 61.820000 88.795000 ;
        RECT 61.620000 89.005000 61.820000 89.205000 ;
        RECT 61.620000 89.415000 61.820000 89.615000 ;
        RECT 61.620000 89.825000 61.820000 90.025000 ;
        RECT 61.620000 90.235000 61.820000 90.435000 ;
        RECT 61.620000 90.645000 61.820000 90.845000 ;
        RECT 61.620000 91.055000 61.820000 91.255000 ;
        RECT 61.620000 91.465000 61.820000 91.665000 ;
        RECT 61.620000 91.875000 61.820000 92.075000 ;
        RECT 61.620000 92.285000 61.820000 92.485000 ;
        RECT 61.620000 92.695000 61.820000 92.895000 ;
        RECT 61.780000 17.860000 61.980000 18.060000 ;
        RECT 61.780000 18.290000 61.980000 18.490000 ;
        RECT 61.780000 18.720000 61.980000 18.920000 ;
        RECT 61.780000 19.150000 61.980000 19.350000 ;
        RECT 61.780000 19.580000 61.980000 19.780000 ;
        RECT 61.780000 20.010000 61.980000 20.210000 ;
        RECT 61.780000 20.440000 61.980000 20.640000 ;
        RECT 61.780000 20.870000 61.980000 21.070000 ;
        RECT 61.780000 21.300000 61.980000 21.500000 ;
        RECT 61.780000 21.730000 61.980000 21.930000 ;
        RECT 61.780000 22.160000 61.980000 22.360000 ;
        RECT 61.810000 68.125000 62.010000 68.325000 ;
        RECT 61.810000 68.535000 62.010000 68.735000 ;
        RECT 61.810000 68.945000 62.010000 69.145000 ;
        RECT 61.810000 69.355000 62.010000 69.555000 ;
        RECT 61.810000 69.765000 62.010000 69.965000 ;
        RECT 61.810000 70.175000 62.010000 70.375000 ;
        RECT 61.810000 70.585000 62.010000 70.785000 ;
        RECT 61.810000 70.995000 62.010000 71.195000 ;
        RECT 61.810000 71.405000 62.010000 71.605000 ;
        RECT 61.810000 71.815000 62.010000 72.015000 ;
        RECT 61.810000 72.225000 62.010000 72.425000 ;
        RECT 61.810000 72.635000 62.010000 72.835000 ;
        RECT 61.810000 73.045000 62.010000 73.245000 ;
        RECT 61.810000 73.450000 62.010000 73.650000 ;
        RECT 61.810000 73.855000 62.010000 74.055000 ;
        RECT 61.810000 74.260000 62.010000 74.460000 ;
        RECT 61.810000 74.665000 62.010000 74.865000 ;
        RECT 61.810000 75.070000 62.010000 75.270000 ;
        RECT 61.810000 75.475000 62.010000 75.675000 ;
        RECT 61.810000 75.880000 62.010000 76.080000 ;
        RECT 61.810000 76.285000 62.010000 76.485000 ;
        RECT 61.810000 76.690000 62.010000 76.890000 ;
        RECT 61.810000 77.095000 62.010000 77.295000 ;
        RECT 61.810000 77.500000 62.010000 77.700000 ;
        RECT 61.810000 77.905000 62.010000 78.105000 ;
        RECT 61.810000 78.310000 62.010000 78.510000 ;
        RECT 61.810000 78.715000 62.010000 78.915000 ;
        RECT 61.810000 79.120000 62.010000 79.320000 ;
        RECT 61.810000 79.525000 62.010000 79.725000 ;
        RECT 61.810000 79.930000 62.010000 80.130000 ;
        RECT 61.810000 80.335000 62.010000 80.535000 ;
        RECT 61.810000 80.740000 62.010000 80.940000 ;
        RECT 61.810000 81.145000 62.010000 81.345000 ;
        RECT 61.810000 81.550000 62.010000 81.750000 ;
        RECT 61.810000 81.955000 62.010000 82.155000 ;
        RECT 61.810000 82.360000 62.010000 82.560000 ;
        RECT 62.025000 82.855000 62.225000 83.055000 ;
        RECT 62.025000 83.265000 62.225000 83.465000 ;
        RECT 62.025000 83.675000 62.225000 83.875000 ;
        RECT 62.025000 84.085000 62.225000 84.285000 ;
        RECT 62.025000 84.495000 62.225000 84.695000 ;
        RECT 62.025000 84.905000 62.225000 85.105000 ;
        RECT 62.025000 85.315000 62.225000 85.515000 ;
        RECT 62.025000 85.725000 62.225000 85.925000 ;
        RECT 62.025000 86.135000 62.225000 86.335000 ;
        RECT 62.025000 86.545000 62.225000 86.745000 ;
        RECT 62.025000 86.955000 62.225000 87.155000 ;
        RECT 62.025000 87.365000 62.225000 87.565000 ;
        RECT 62.025000 87.775000 62.225000 87.975000 ;
        RECT 62.025000 88.185000 62.225000 88.385000 ;
        RECT 62.025000 88.595000 62.225000 88.795000 ;
        RECT 62.025000 89.005000 62.225000 89.205000 ;
        RECT 62.025000 89.415000 62.225000 89.615000 ;
        RECT 62.025000 89.825000 62.225000 90.025000 ;
        RECT 62.025000 90.235000 62.225000 90.435000 ;
        RECT 62.025000 90.645000 62.225000 90.845000 ;
        RECT 62.025000 91.055000 62.225000 91.255000 ;
        RECT 62.025000 91.465000 62.225000 91.665000 ;
        RECT 62.025000 91.875000 62.225000 92.075000 ;
        RECT 62.025000 92.285000 62.225000 92.485000 ;
        RECT 62.025000 92.695000 62.225000 92.895000 ;
        RECT 62.185000 17.860000 62.385000 18.060000 ;
        RECT 62.185000 18.290000 62.385000 18.490000 ;
        RECT 62.185000 18.720000 62.385000 18.920000 ;
        RECT 62.185000 19.150000 62.385000 19.350000 ;
        RECT 62.185000 19.580000 62.385000 19.780000 ;
        RECT 62.185000 20.010000 62.385000 20.210000 ;
        RECT 62.185000 20.440000 62.385000 20.640000 ;
        RECT 62.185000 20.870000 62.385000 21.070000 ;
        RECT 62.185000 21.300000 62.385000 21.500000 ;
        RECT 62.185000 21.730000 62.385000 21.930000 ;
        RECT 62.185000 22.160000 62.385000 22.360000 ;
        RECT 62.210000 68.125000 62.410000 68.325000 ;
        RECT 62.210000 68.535000 62.410000 68.735000 ;
        RECT 62.210000 68.945000 62.410000 69.145000 ;
        RECT 62.210000 69.355000 62.410000 69.555000 ;
        RECT 62.210000 69.765000 62.410000 69.965000 ;
        RECT 62.210000 70.175000 62.410000 70.375000 ;
        RECT 62.210000 70.585000 62.410000 70.785000 ;
        RECT 62.210000 70.995000 62.410000 71.195000 ;
        RECT 62.210000 71.405000 62.410000 71.605000 ;
        RECT 62.210000 71.815000 62.410000 72.015000 ;
        RECT 62.210000 72.225000 62.410000 72.425000 ;
        RECT 62.210000 72.635000 62.410000 72.835000 ;
        RECT 62.210000 73.045000 62.410000 73.245000 ;
        RECT 62.210000 73.450000 62.410000 73.650000 ;
        RECT 62.210000 73.855000 62.410000 74.055000 ;
        RECT 62.210000 74.260000 62.410000 74.460000 ;
        RECT 62.210000 74.665000 62.410000 74.865000 ;
        RECT 62.210000 75.070000 62.410000 75.270000 ;
        RECT 62.210000 75.475000 62.410000 75.675000 ;
        RECT 62.210000 75.880000 62.410000 76.080000 ;
        RECT 62.210000 76.285000 62.410000 76.485000 ;
        RECT 62.210000 76.690000 62.410000 76.890000 ;
        RECT 62.210000 77.095000 62.410000 77.295000 ;
        RECT 62.210000 77.500000 62.410000 77.700000 ;
        RECT 62.210000 77.905000 62.410000 78.105000 ;
        RECT 62.210000 78.310000 62.410000 78.510000 ;
        RECT 62.210000 78.715000 62.410000 78.915000 ;
        RECT 62.210000 79.120000 62.410000 79.320000 ;
        RECT 62.210000 79.525000 62.410000 79.725000 ;
        RECT 62.210000 79.930000 62.410000 80.130000 ;
        RECT 62.210000 80.335000 62.410000 80.535000 ;
        RECT 62.210000 80.740000 62.410000 80.940000 ;
        RECT 62.210000 81.145000 62.410000 81.345000 ;
        RECT 62.210000 81.550000 62.410000 81.750000 ;
        RECT 62.210000 81.955000 62.410000 82.155000 ;
        RECT 62.210000 82.360000 62.410000 82.560000 ;
        RECT 62.430000 82.855000 62.630000 83.055000 ;
        RECT 62.430000 83.265000 62.630000 83.465000 ;
        RECT 62.430000 83.675000 62.630000 83.875000 ;
        RECT 62.430000 84.085000 62.630000 84.285000 ;
        RECT 62.430000 84.495000 62.630000 84.695000 ;
        RECT 62.430000 84.905000 62.630000 85.105000 ;
        RECT 62.430000 85.315000 62.630000 85.515000 ;
        RECT 62.430000 85.725000 62.630000 85.925000 ;
        RECT 62.430000 86.135000 62.630000 86.335000 ;
        RECT 62.430000 86.545000 62.630000 86.745000 ;
        RECT 62.430000 86.955000 62.630000 87.155000 ;
        RECT 62.430000 87.365000 62.630000 87.565000 ;
        RECT 62.430000 87.775000 62.630000 87.975000 ;
        RECT 62.430000 88.185000 62.630000 88.385000 ;
        RECT 62.430000 88.595000 62.630000 88.795000 ;
        RECT 62.430000 89.005000 62.630000 89.205000 ;
        RECT 62.430000 89.415000 62.630000 89.615000 ;
        RECT 62.430000 89.825000 62.630000 90.025000 ;
        RECT 62.430000 90.235000 62.630000 90.435000 ;
        RECT 62.430000 90.645000 62.630000 90.845000 ;
        RECT 62.430000 91.055000 62.630000 91.255000 ;
        RECT 62.430000 91.465000 62.630000 91.665000 ;
        RECT 62.430000 91.875000 62.630000 92.075000 ;
        RECT 62.430000 92.285000 62.630000 92.485000 ;
        RECT 62.430000 92.695000 62.630000 92.895000 ;
        RECT 62.590000 17.860000 62.790000 18.060000 ;
        RECT 62.590000 18.290000 62.790000 18.490000 ;
        RECT 62.590000 18.720000 62.790000 18.920000 ;
        RECT 62.590000 19.150000 62.790000 19.350000 ;
        RECT 62.590000 19.580000 62.790000 19.780000 ;
        RECT 62.590000 20.010000 62.790000 20.210000 ;
        RECT 62.590000 20.440000 62.790000 20.640000 ;
        RECT 62.590000 20.870000 62.790000 21.070000 ;
        RECT 62.590000 21.300000 62.790000 21.500000 ;
        RECT 62.590000 21.730000 62.790000 21.930000 ;
        RECT 62.590000 22.160000 62.790000 22.360000 ;
        RECT 62.610000 68.125000 62.810000 68.325000 ;
        RECT 62.610000 68.535000 62.810000 68.735000 ;
        RECT 62.610000 68.945000 62.810000 69.145000 ;
        RECT 62.610000 69.355000 62.810000 69.555000 ;
        RECT 62.610000 69.765000 62.810000 69.965000 ;
        RECT 62.610000 70.175000 62.810000 70.375000 ;
        RECT 62.610000 70.585000 62.810000 70.785000 ;
        RECT 62.610000 70.995000 62.810000 71.195000 ;
        RECT 62.610000 71.405000 62.810000 71.605000 ;
        RECT 62.610000 71.815000 62.810000 72.015000 ;
        RECT 62.610000 72.225000 62.810000 72.425000 ;
        RECT 62.610000 72.635000 62.810000 72.835000 ;
        RECT 62.610000 73.045000 62.810000 73.245000 ;
        RECT 62.610000 73.450000 62.810000 73.650000 ;
        RECT 62.610000 73.855000 62.810000 74.055000 ;
        RECT 62.610000 74.260000 62.810000 74.460000 ;
        RECT 62.610000 74.665000 62.810000 74.865000 ;
        RECT 62.610000 75.070000 62.810000 75.270000 ;
        RECT 62.610000 75.475000 62.810000 75.675000 ;
        RECT 62.610000 75.880000 62.810000 76.080000 ;
        RECT 62.610000 76.285000 62.810000 76.485000 ;
        RECT 62.610000 76.690000 62.810000 76.890000 ;
        RECT 62.610000 77.095000 62.810000 77.295000 ;
        RECT 62.610000 77.500000 62.810000 77.700000 ;
        RECT 62.610000 77.905000 62.810000 78.105000 ;
        RECT 62.610000 78.310000 62.810000 78.510000 ;
        RECT 62.610000 78.715000 62.810000 78.915000 ;
        RECT 62.610000 79.120000 62.810000 79.320000 ;
        RECT 62.610000 79.525000 62.810000 79.725000 ;
        RECT 62.610000 79.930000 62.810000 80.130000 ;
        RECT 62.610000 80.335000 62.810000 80.535000 ;
        RECT 62.610000 80.740000 62.810000 80.940000 ;
        RECT 62.610000 81.145000 62.810000 81.345000 ;
        RECT 62.610000 81.550000 62.810000 81.750000 ;
        RECT 62.610000 81.955000 62.810000 82.155000 ;
        RECT 62.610000 82.360000 62.810000 82.560000 ;
        RECT 62.840000 82.855000 63.040000 83.055000 ;
        RECT 62.840000 83.265000 63.040000 83.465000 ;
        RECT 62.840000 83.675000 63.040000 83.875000 ;
        RECT 62.840000 84.085000 63.040000 84.285000 ;
        RECT 62.840000 84.495000 63.040000 84.695000 ;
        RECT 62.840000 84.905000 63.040000 85.105000 ;
        RECT 62.840000 85.315000 63.040000 85.515000 ;
        RECT 62.840000 85.725000 63.040000 85.925000 ;
        RECT 62.840000 86.135000 63.040000 86.335000 ;
        RECT 62.840000 86.545000 63.040000 86.745000 ;
        RECT 62.840000 86.955000 63.040000 87.155000 ;
        RECT 62.840000 87.365000 63.040000 87.565000 ;
        RECT 62.840000 87.775000 63.040000 87.975000 ;
        RECT 62.840000 88.185000 63.040000 88.385000 ;
        RECT 62.840000 88.595000 63.040000 88.795000 ;
        RECT 62.840000 89.005000 63.040000 89.205000 ;
        RECT 62.840000 89.415000 63.040000 89.615000 ;
        RECT 62.840000 89.825000 63.040000 90.025000 ;
        RECT 62.840000 90.235000 63.040000 90.435000 ;
        RECT 62.840000 90.645000 63.040000 90.845000 ;
        RECT 62.840000 91.055000 63.040000 91.255000 ;
        RECT 62.840000 91.465000 63.040000 91.665000 ;
        RECT 62.840000 91.875000 63.040000 92.075000 ;
        RECT 62.840000 92.285000 63.040000 92.485000 ;
        RECT 62.840000 92.695000 63.040000 92.895000 ;
        RECT 62.995000 17.860000 63.195000 18.060000 ;
        RECT 62.995000 18.290000 63.195000 18.490000 ;
        RECT 62.995000 18.720000 63.195000 18.920000 ;
        RECT 62.995000 19.150000 63.195000 19.350000 ;
        RECT 62.995000 19.580000 63.195000 19.780000 ;
        RECT 62.995000 20.010000 63.195000 20.210000 ;
        RECT 62.995000 20.440000 63.195000 20.640000 ;
        RECT 62.995000 20.870000 63.195000 21.070000 ;
        RECT 62.995000 21.300000 63.195000 21.500000 ;
        RECT 62.995000 21.730000 63.195000 21.930000 ;
        RECT 62.995000 22.160000 63.195000 22.360000 ;
        RECT 63.010000 68.125000 63.210000 68.325000 ;
        RECT 63.010000 68.535000 63.210000 68.735000 ;
        RECT 63.010000 68.945000 63.210000 69.145000 ;
        RECT 63.010000 69.355000 63.210000 69.555000 ;
        RECT 63.010000 69.765000 63.210000 69.965000 ;
        RECT 63.010000 70.175000 63.210000 70.375000 ;
        RECT 63.010000 70.585000 63.210000 70.785000 ;
        RECT 63.010000 70.995000 63.210000 71.195000 ;
        RECT 63.010000 71.405000 63.210000 71.605000 ;
        RECT 63.010000 71.815000 63.210000 72.015000 ;
        RECT 63.010000 72.225000 63.210000 72.425000 ;
        RECT 63.010000 72.635000 63.210000 72.835000 ;
        RECT 63.010000 73.045000 63.210000 73.245000 ;
        RECT 63.010000 73.450000 63.210000 73.650000 ;
        RECT 63.010000 73.855000 63.210000 74.055000 ;
        RECT 63.010000 74.260000 63.210000 74.460000 ;
        RECT 63.010000 74.665000 63.210000 74.865000 ;
        RECT 63.010000 75.070000 63.210000 75.270000 ;
        RECT 63.010000 75.475000 63.210000 75.675000 ;
        RECT 63.010000 75.880000 63.210000 76.080000 ;
        RECT 63.010000 76.285000 63.210000 76.485000 ;
        RECT 63.010000 76.690000 63.210000 76.890000 ;
        RECT 63.010000 77.095000 63.210000 77.295000 ;
        RECT 63.010000 77.500000 63.210000 77.700000 ;
        RECT 63.010000 77.905000 63.210000 78.105000 ;
        RECT 63.010000 78.310000 63.210000 78.510000 ;
        RECT 63.010000 78.715000 63.210000 78.915000 ;
        RECT 63.010000 79.120000 63.210000 79.320000 ;
        RECT 63.010000 79.525000 63.210000 79.725000 ;
        RECT 63.010000 79.930000 63.210000 80.130000 ;
        RECT 63.010000 80.335000 63.210000 80.535000 ;
        RECT 63.010000 80.740000 63.210000 80.940000 ;
        RECT 63.010000 81.145000 63.210000 81.345000 ;
        RECT 63.010000 81.550000 63.210000 81.750000 ;
        RECT 63.010000 81.955000 63.210000 82.155000 ;
        RECT 63.010000 82.360000 63.210000 82.560000 ;
        RECT 63.250000 82.855000 63.450000 83.055000 ;
        RECT 63.250000 83.265000 63.450000 83.465000 ;
        RECT 63.250000 83.675000 63.450000 83.875000 ;
        RECT 63.250000 84.085000 63.450000 84.285000 ;
        RECT 63.250000 84.495000 63.450000 84.695000 ;
        RECT 63.250000 84.905000 63.450000 85.105000 ;
        RECT 63.250000 85.315000 63.450000 85.515000 ;
        RECT 63.250000 85.725000 63.450000 85.925000 ;
        RECT 63.250000 86.135000 63.450000 86.335000 ;
        RECT 63.250000 86.545000 63.450000 86.745000 ;
        RECT 63.250000 86.955000 63.450000 87.155000 ;
        RECT 63.250000 87.365000 63.450000 87.565000 ;
        RECT 63.250000 87.775000 63.450000 87.975000 ;
        RECT 63.250000 88.185000 63.450000 88.385000 ;
        RECT 63.250000 88.595000 63.450000 88.795000 ;
        RECT 63.250000 89.005000 63.450000 89.205000 ;
        RECT 63.250000 89.415000 63.450000 89.615000 ;
        RECT 63.250000 89.825000 63.450000 90.025000 ;
        RECT 63.250000 90.235000 63.450000 90.435000 ;
        RECT 63.250000 90.645000 63.450000 90.845000 ;
        RECT 63.250000 91.055000 63.450000 91.255000 ;
        RECT 63.250000 91.465000 63.450000 91.665000 ;
        RECT 63.250000 91.875000 63.450000 92.075000 ;
        RECT 63.250000 92.285000 63.450000 92.485000 ;
        RECT 63.250000 92.695000 63.450000 92.895000 ;
        RECT 63.400000 17.860000 63.600000 18.060000 ;
        RECT 63.400000 18.290000 63.600000 18.490000 ;
        RECT 63.400000 18.720000 63.600000 18.920000 ;
        RECT 63.400000 19.150000 63.600000 19.350000 ;
        RECT 63.400000 19.580000 63.600000 19.780000 ;
        RECT 63.400000 20.010000 63.600000 20.210000 ;
        RECT 63.400000 20.440000 63.600000 20.640000 ;
        RECT 63.400000 20.870000 63.600000 21.070000 ;
        RECT 63.400000 21.300000 63.600000 21.500000 ;
        RECT 63.400000 21.730000 63.600000 21.930000 ;
        RECT 63.400000 22.160000 63.600000 22.360000 ;
        RECT 63.410000 68.125000 63.610000 68.325000 ;
        RECT 63.410000 68.535000 63.610000 68.735000 ;
        RECT 63.410000 68.945000 63.610000 69.145000 ;
        RECT 63.410000 69.355000 63.610000 69.555000 ;
        RECT 63.410000 69.765000 63.610000 69.965000 ;
        RECT 63.410000 70.175000 63.610000 70.375000 ;
        RECT 63.410000 70.585000 63.610000 70.785000 ;
        RECT 63.410000 70.995000 63.610000 71.195000 ;
        RECT 63.410000 71.405000 63.610000 71.605000 ;
        RECT 63.410000 71.815000 63.610000 72.015000 ;
        RECT 63.410000 72.225000 63.610000 72.425000 ;
        RECT 63.410000 72.635000 63.610000 72.835000 ;
        RECT 63.410000 73.045000 63.610000 73.245000 ;
        RECT 63.410000 73.450000 63.610000 73.650000 ;
        RECT 63.410000 73.855000 63.610000 74.055000 ;
        RECT 63.410000 74.260000 63.610000 74.460000 ;
        RECT 63.410000 74.665000 63.610000 74.865000 ;
        RECT 63.410000 75.070000 63.610000 75.270000 ;
        RECT 63.410000 75.475000 63.610000 75.675000 ;
        RECT 63.410000 75.880000 63.610000 76.080000 ;
        RECT 63.410000 76.285000 63.610000 76.485000 ;
        RECT 63.410000 76.690000 63.610000 76.890000 ;
        RECT 63.410000 77.095000 63.610000 77.295000 ;
        RECT 63.410000 77.500000 63.610000 77.700000 ;
        RECT 63.410000 77.905000 63.610000 78.105000 ;
        RECT 63.410000 78.310000 63.610000 78.510000 ;
        RECT 63.410000 78.715000 63.610000 78.915000 ;
        RECT 63.410000 79.120000 63.610000 79.320000 ;
        RECT 63.410000 79.525000 63.610000 79.725000 ;
        RECT 63.410000 79.930000 63.610000 80.130000 ;
        RECT 63.410000 80.335000 63.610000 80.535000 ;
        RECT 63.410000 80.740000 63.610000 80.940000 ;
        RECT 63.410000 81.145000 63.610000 81.345000 ;
        RECT 63.410000 81.550000 63.610000 81.750000 ;
        RECT 63.410000 81.955000 63.610000 82.155000 ;
        RECT 63.410000 82.360000 63.610000 82.560000 ;
        RECT 63.660000 82.855000 63.860000 83.055000 ;
        RECT 63.660000 83.265000 63.860000 83.465000 ;
        RECT 63.660000 83.675000 63.860000 83.875000 ;
        RECT 63.660000 84.085000 63.860000 84.285000 ;
        RECT 63.660000 84.495000 63.860000 84.695000 ;
        RECT 63.660000 84.905000 63.860000 85.105000 ;
        RECT 63.660000 85.315000 63.860000 85.515000 ;
        RECT 63.660000 85.725000 63.860000 85.925000 ;
        RECT 63.660000 86.135000 63.860000 86.335000 ;
        RECT 63.660000 86.545000 63.860000 86.745000 ;
        RECT 63.660000 86.955000 63.860000 87.155000 ;
        RECT 63.660000 87.365000 63.860000 87.565000 ;
        RECT 63.660000 87.775000 63.860000 87.975000 ;
        RECT 63.660000 88.185000 63.860000 88.385000 ;
        RECT 63.660000 88.595000 63.860000 88.795000 ;
        RECT 63.660000 89.005000 63.860000 89.205000 ;
        RECT 63.660000 89.415000 63.860000 89.615000 ;
        RECT 63.660000 89.825000 63.860000 90.025000 ;
        RECT 63.660000 90.235000 63.860000 90.435000 ;
        RECT 63.660000 90.645000 63.860000 90.845000 ;
        RECT 63.660000 91.055000 63.860000 91.255000 ;
        RECT 63.660000 91.465000 63.860000 91.665000 ;
        RECT 63.660000 91.875000 63.860000 92.075000 ;
        RECT 63.660000 92.285000 63.860000 92.485000 ;
        RECT 63.660000 92.695000 63.860000 92.895000 ;
        RECT 63.805000 17.860000 64.005000 18.060000 ;
        RECT 63.805000 18.290000 64.005000 18.490000 ;
        RECT 63.805000 18.720000 64.005000 18.920000 ;
        RECT 63.805000 19.150000 64.005000 19.350000 ;
        RECT 63.805000 19.580000 64.005000 19.780000 ;
        RECT 63.805000 20.010000 64.005000 20.210000 ;
        RECT 63.805000 20.440000 64.005000 20.640000 ;
        RECT 63.805000 20.870000 64.005000 21.070000 ;
        RECT 63.805000 21.300000 64.005000 21.500000 ;
        RECT 63.805000 21.730000 64.005000 21.930000 ;
        RECT 63.805000 22.160000 64.005000 22.360000 ;
        RECT 63.810000 68.125000 64.010000 68.325000 ;
        RECT 63.810000 68.535000 64.010000 68.735000 ;
        RECT 63.810000 68.945000 64.010000 69.145000 ;
        RECT 63.810000 69.355000 64.010000 69.555000 ;
        RECT 63.810000 69.765000 64.010000 69.965000 ;
        RECT 63.810000 70.175000 64.010000 70.375000 ;
        RECT 63.810000 70.585000 64.010000 70.785000 ;
        RECT 63.810000 70.995000 64.010000 71.195000 ;
        RECT 63.810000 71.405000 64.010000 71.605000 ;
        RECT 63.810000 71.815000 64.010000 72.015000 ;
        RECT 63.810000 72.225000 64.010000 72.425000 ;
        RECT 63.810000 72.635000 64.010000 72.835000 ;
        RECT 63.810000 73.045000 64.010000 73.245000 ;
        RECT 63.810000 73.450000 64.010000 73.650000 ;
        RECT 63.810000 73.855000 64.010000 74.055000 ;
        RECT 63.810000 74.260000 64.010000 74.460000 ;
        RECT 63.810000 74.665000 64.010000 74.865000 ;
        RECT 63.810000 75.070000 64.010000 75.270000 ;
        RECT 63.810000 75.475000 64.010000 75.675000 ;
        RECT 63.810000 75.880000 64.010000 76.080000 ;
        RECT 63.810000 76.285000 64.010000 76.485000 ;
        RECT 63.810000 76.690000 64.010000 76.890000 ;
        RECT 63.810000 77.095000 64.010000 77.295000 ;
        RECT 63.810000 77.500000 64.010000 77.700000 ;
        RECT 63.810000 77.905000 64.010000 78.105000 ;
        RECT 63.810000 78.310000 64.010000 78.510000 ;
        RECT 63.810000 78.715000 64.010000 78.915000 ;
        RECT 63.810000 79.120000 64.010000 79.320000 ;
        RECT 63.810000 79.525000 64.010000 79.725000 ;
        RECT 63.810000 79.930000 64.010000 80.130000 ;
        RECT 63.810000 80.335000 64.010000 80.535000 ;
        RECT 63.810000 80.740000 64.010000 80.940000 ;
        RECT 63.810000 81.145000 64.010000 81.345000 ;
        RECT 63.810000 81.550000 64.010000 81.750000 ;
        RECT 63.810000 81.955000 64.010000 82.155000 ;
        RECT 63.810000 82.360000 64.010000 82.560000 ;
        RECT 64.070000 82.855000 64.270000 83.055000 ;
        RECT 64.070000 83.265000 64.270000 83.465000 ;
        RECT 64.070000 83.675000 64.270000 83.875000 ;
        RECT 64.070000 84.085000 64.270000 84.285000 ;
        RECT 64.070000 84.495000 64.270000 84.695000 ;
        RECT 64.070000 84.905000 64.270000 85.105000 ;
        RECT 64.070000 85.315000 64.270000 85.515000 ;
        RECT 64.070000 85.725000 64.270000 85.925000 ;
        RECT 64.070000 86.135000 64.270000 86.335000 ;
        RECT 64.070000 86.545000 64.270000 86.745000 ;
        RECT 64.070000 86.955000 64.270000 87.155000 ;
        RECT 64.070000 87.365000 64.270000 87.565000 ;
        RECT 64.070000 87.775000 64.270000 87.975000 ;
        RECT 64.070000 88.185000 64.270000 88.385000 ;
        RECT 64.070000 88.595000 64.270000 88.795000 ;
        RECT 64.070000 89.005000 64.270000 89.205000 ;
        RECT 64.070000 89.415000 64.270000 89.615000 ;
        RECT 64.070000 89.825000 64.270000 90.025000 ;
        RECT 64.070000 90.235000 64.270000 90.435000 ;
        RECT 64.070000 90.645000 64.270000 90.845000 ;
        RECT 64.070000 91.055000 64.270000 91.255000 ;
        RECT 64.070000 91.465000 64.270000 91.665000 ;
        RECT 64.070000 91.875000 64.270000 92.075000 ;
        RECT 64.070000 92.285000 64.270000 92.485000 ;
        RECT 64.070000 92.695000 64.270000 92.895000 ;
        RECT 64.210000 17.860000 64.410000 18.060000 ;
        RECT 64.210000 18.290000 64.410000 18.490000 ;
        RECT 64.210000 18.720000 64.410000 18.920000 ;
        RECT 64.210000 19.150000 64.410000 19.350000 ;
        RECT 64.210000 19.580000 64.410000 19.780000 ;
        RECT 64.210000 20.010000 64.410000 20.210000 ;
        RECT 64.210000 20.440000 64.410000 20.640000 ;
        RECT 64.210000 20.870000 64.410000 21.070000 ;
        RECT 64.210000 21.300000 64.410000 21.500000 ;
        RECT 64.210000 21.730000 64.410000 21.930000 ;
        RECT 64.210000 22.160000 64.410000 22.360000 ;
        RECT 64.210000 68.125000 64.410000 68.325000 ;
        RECT 64.210000 68.535000 64.410000 68.735000 ;
        RECT 64.210000 68.945000 64.410000 69.145000 ;
        RECT 64.210000 69.355000 64.410000 69.555000 ;
        RECT 64.210000 69.765000 64.410000 69.965000 ;
        RECT 64.210000 70.175000 64.410000 70.375000 ;
        RECT 64.210000 70.585000 64.410000 70.785000 ;
        RECT 64.210000 70.995000 64.410000 71.195000 ;
        RECT 64.210000 71.405000 64.410000 71.605000 ;
        RECT 64.210000 71.815000 64.410000 72.015000 ;
        RECT 64.210000 72.225000 64.410000 72.425000 ;
        RECT 64.210000 72.635000 64.410000 72.835000 ;
        RECT 64.210000 73.045000 64.410000 73.245000 ;
        RECT 64.210000 73.450000 64.410000 73.650000 ;
        RECT 64.210000 73.855000 64.410000 74.055000 ;
        RECT 64.210000 74.260000 64.410000 74.460000 ;
        RECT 64.210000 74.665000 64.410000 74.865000 ;
        RECT 64.210000 75.070000 64.410000 75.270000 ;
        RECT 64.210000 75.475000 64.410000 75.675000 ;
        RECT 64.210000 75.880000 64.410000 76.080000 ;
        RECT 64.210000 76.285000 64.410000 76.485000 ;
        RECT 64.210000 76.690000 64.410000 76.890000 ;
        RECT 64.210000 77.095000 64.410000 77.295000 ;
        RECT 64.210000 77.500000 64.410000 77.700000 ;
        RECT 64.210000 77.905000 64.410000 78.105000 ;
        RECT 64.210000 78.310000 64.410000 78.510000 ;
        RECT 64.210000 78.715000 64.410000 78.915000 ;
        RECT 64.210000 79.120000 64.410000 79.320000 ;
        RECT 64.210000 79.525000 64.410000 79.725000 ;
        RECT 64.210000 79.930000 64.410000 80.130000 ;
        RECT 64.210000 80.335000 64.410000 80.535000 ;
        RECT 64.210000 80.740000 64.410000 80.940000 ;
        RECT 64.210000 81.145000 64.410000 81.345000 ;
        RECT 64.210000 81.550000 64.410000 81.750000 ;
        RECT 64.210000 81.955000 64.410000 82.155000 ;
        RECT 64.210000 82.360000 64.410000 82.560000 ;
        RECT 64.480000 82.855000 64.680000 83.055000 ;
        RECT 64.480000 83.265000 64.680000 83.465000 ;
        RECT 64.480000 83.675000 64.680000 83.875000 ;
        RECT 64.480000 84.085000 64.680000 84.285000 ;
        RECT 64.480000 84.495000 64.680000 84.695000 ;
        RECT 64.480000 84.905000 64.680000 85.105000 ;
        RECT 64.480000 85.315000 64.680000 85.515000 ;
        RECT 64.480000 85.725000 64.680000 85.925000 ;
        RECT 64.480000 86.135000 64.680000 86.335000 ;
        RECT 64.480000 86.545000 64.680000 86.745000 ;
        RECT 64.480000 86.955000 64.680000 87.155000 ;
        RECT 64.480000 87.365000 64.680000 87.565000 ;
        RECT 64.480000 87.775000 64.680000 87.975000 ;
        RECT 64.480000 88.185000 64.680000 88.385000 ;
        RECT 64.480000 88.595000 64.680000 88.795000 ;
        RECT 64.480000 89.005000 64.680000 89.205000 ;
        RECT 64.480000 89.415000 64.680000 89.615000 ;
        RECT 64.480000 89.825000 64.680000 90.025000 ;
        RECT 64.480000 90.235000 64.680000 90.435000 ;
        RECT 64.480000 90.645000 64.680000 90.845000 ;
        RECT 64.480000 91.055000 64.680000 91.255000 ;
        RECT 64.480000 91.465000 64.680000 91.665000 ;
        RECT 64.480000 91.875000 64.680000 92.075000 ;
        RECT 64.480000 92.285000 64.680000 92.485000 ;
        RECT 64.480000 92.695000 64.680000 92.895000 ;
        RECT 64.610000 68.125000 64.810000 68.325000 ;
        RECT 64.610000 68.535000 64.810000 68.735000 ;
        RECT 64.610000 68.945000 64.810000 69.145000 ;
        RECT 64.610000 69.355000 64.810000 69.555000 ;
        RECT 64.610000 69.765000 64.810000 69.965000 ;
        RECT 64.610000 70.175000 64.810000 70.375000 ;
        RECT 64.610000 70.585000 64.810000 70.785000 ;
        RECT 64.610000 70.995000 64.810000 71.195000 ;
        RECT 64.610000 71.405000 64.810000 71.605000 ;
        RECT 64.610000 71.815000 64.810000 72.015000 ;
        RECT 64.610000 72.225000 64.810000 72.425000 ;
        RECT 64.610000 72.635000 64.810000 72.835000 ;
        RECT 64.610000 73.045000 64.810000 73.245000 ;
        RECT 64.610000 73.450000 64.810000 73.650000 ;
        RECT 64.610000 73.855000 64.810000 74.055000 ;
        RECT 64.610000 74.260000 64.810000 74.460000 ;
        RECT 64.610000 74.665000 64.810000 74.865000 ;
        RECT 64.610000 75.070000 64.810000 75.270000 ;
        RECT 64.610000 75.475000 64.810000 75.675000 ;
        RECT 64.610000 75.880000 64.810000 76.080000 ;
        RECT 64.610000 76.285000 64.810000 76.485000 ;
        RECT 64.610000 76.690000 64.810000 76.890000 ;
        RECT 64.610000 77.095000 64.810000 77.295000 ;
        RECT 64.610000 77.500000 64.810000 77.700000 ;
        RECT 64.610000 77.905000 64.810000 78.105000 ;
        RECT 64.610000 78.310000 64.810000 78.510000 ;
        RECT 64.610000 78.715000 64.810000 78.915000 ;
        RECT 64.610000 79.120000 64.810000 79.320000 ;
        RECT 64.610000 79.525000 64.810000 79.725000 ;
        RECT 64.610000 79.930000 64.810000 80.130000 ;
        RECT 64.610000 80.335000 64.810000 80.535000 ;
        RECT 64.610000 80.740000 64.810000 80.940000 ;
        RECT 64.610000 81.145000 64.810000 81.345000 ;
        RECT 64.610000 81.550000 64.810000 81.750000 ;
        RECT 64.610000 81.955000 64.810000 82.155000 ;
        RECT 64.610000 82.360000 64.810000 82.560000 ;
        RECT 64.615000 17.860000 64.815000 18.060000 ;
        RECT 64.615000 18.290000 64.815000 18.490000 ;
        RECT 64.615000 18.720000 64.815000 18.920000 ;
        RECT 64.615000 19.150000 64.815000 19.350000 ;
        RECT 64.615000 19.580000 64.815000 19.780000 ;
        RECT 64.615000 20.010000 64.815000 20.210000 ;
        RECT 64.615000 20.440000 64.815000 20.640000 ;
        RECT 64.615000 20.870000 64.815000 21.070000 ;
        RECT 64.615000 21.300000 64.815000 21.500000 ;
        RECT 64.615000 21.730000 64.815000 21.930000 ;
        RECT 64.615000 22.160000 64.815000 22.360000 ;
        RECT 64.890000 82.855000 65.090000 83.055000 ;
        RECT 64.890000 83.265000 65.090000 83.465000 ;
        RECT 64.890000 83.675000 65.090000 83.875000 ;
        RECT 64.890000 84.085000 65.090000 84.285000 ;
        RECT 64.890000 84.495000 65.090000 84.695000 ;
        RECT 64.890000 84.905000 65.090000 85.105000 ;
        RECT 64.890000 85.315000 65.090000 85.515000 ;
        RECT 64.890000 85.725000 65.090000 85.925000 ;
        RECT 64.890000 86.135000 65.090000 86.335000 ;
        RECT 64.890000 86.545000 65.090000 86.745000 ;
        RECT 64.890000 86.955000 65.090000 87.155000 ;
        RECT 64.890000 87.365000 65.090000 87.565000 ;
        RECT 64.890000 87.775000 65.090000 87.975000 ;
        RECT 64.890000 88.185000 65.090000 88.385000 ;
        RECT 64.890000 88.595000 65.090000 88.795000 ;
        RECT 64.890000 89.005000 65.090000 89.205000 ;
        RECT 64.890000 89.415000 65.090000 89.615000 ;
        RECT 64.890000 89.825000 65.090000 90.025000 ;
        RECT 64.890000 90.235000 65.090000 90.435000 ;
        RECT 64.890000 90.645000 65.090000 90.845000 ;
        RECT 64.890000 91.055000 65.090000 91.255000 ;
        RECT 64.890000 91.465000 65.090000 91.665000 ;
        RECT 64.890000 91.875000 65.090000 92.075000 ;
        RECT 64.890000 92.285000 65.090000 92.485000 ;
        RECT 64.890000 92.695000 65.090000 92.895000 ;
        RECT 65.010000 68.125000 65.210000 68.325000 ;
        RECT 65.010000 68.535000 65.210000 68.735000 ;
        RECT 65.010000 68.945000 65.210000 69.145000 ;
        RECT 65.010000 69.355000 65.210000 69.555000 ;
        RECT 65.010000 69.765000 65.210000 69.965000 ;
        RECT 65.010000 70.175000 65.210000 70.375000 ;
        RECT 65.010000 70.585000 65.210000 70.785000 ;
        RECT 65.010000 70.995000 65.210000 71.195000 ;
        RECT 65.010000 71.405000 65.210000 71.605000 ;
        RECT 65.010000 71.815000 65.210000 72.015000 ;
        RECT 65.010000 72.225000 65.210000 72.425000 ;
        RECT 65.010000 72.635000 65.210000 72.835000 ;
        RECT 65.010000 73.045000 65.210000 73.245000 ;
        RECT 65.010000 73.450000 65.210000 73.650000 ;
        RECT 65.010000 73.855000 65.210000 74.055000 ;
        RECT 65.010000 74.260000 65.210000 74.460000 ;
        RECT 65.010000 74.665000 65.210000 74.865000 ;
        RECT 65.010000 75.070000 65.210000 75.270000 ;
        RECT 65.010000 75.475000 65.210000 75.675000 ;
        RECT 65.010000 75.880000 65.210000 76.080000 ;
        RECT 65.010000 76.285000 65.210000 76.485000 ;
        RECT 65.010000 76.690000 65.210000 76.890000 ;
        RECT 65.010000 77.095000 65.210000 77.295000 ;
        RECT 65.010000 77.500000 65.210000 77.700000 ;
        RECT 65.010000 77.905000 65.210000 78.105000 ;
        RECT 65.010000 78.310000 65.210000 78.510000 ;
        RECT 65.010000 78.715000 65.210000 78.915000 ;
        RECT 65.010000 79.120000 65.210000 79.320000 ;
        RECT 65.010000 79.525000 65.210000 79.725000 ;
        RECT 65.010000 79.930000 65.210000 80.130000 ;
        RECT 65.010000 80.335000 65.210000 80.535000 ;
        RECT 65.010000 80.740000 65.210000 80.940000 ;
        RECT 65.010000 81.145000 65.210000 81.345000 ;
        RECT 65.010000 81.550000 65.210000 81.750000 ;
        RECT 65.010000 81.955000 65.210000 82.155000 ;
        RECT 65.010000 82.360000 65.210000 82.560000 ;
        RECT 65.020000 17.860000 65.220000 18.060000 ;
        RECT 65.020000 18.290000 65.220000 18.490000 ;
        RECT 65.020000 18.720000 65.220000 18.920000 ;
        RECT 65.020000 19.150000 65.220000 19.350000 ;
        RECT 65.020000 19.580000 65.220000 19.780000 ;
        RECT 65.020000 20.010000 65.220000 20.210000 ;
        RECT 65.020000 20.440000 65.220000 20.640000 ;
        RECT 65.020000 20.870000 65.220000 21.070000 ;
        RECT 65.020000 21.300000 65.220000 21.500000 ;
        RECT 65.020000 21.730000 65.220000 21.930000 ;
        RECT 65.020000 22.160000 65.220000 22.360000 ;
        RECT 65.300000 82.855000 65.500000 83.055000 ;
        RECT 65.300000 83.265000 65.500000 83.465000 ;
        RECT 65.300000 83.675000 65.500000 83.875000 ;
        RECT 65.300000 84.085000 65.500000 84.285000 ;
        RECT 65.300000 84.495000 65.500000 84.695000 ;
        RECT 65.300000 84.905000 65.500000 85.105000 ;
        RECT 65.300000 85.315000 65.500000 85.515000 ;
        RECT 65.300000 85.725000 65.500000 85.925000 ;
        RECT 65.300000 86.135000 65.500000 86.335000 ;
        RECT 65.300000 86.545000 65.500000 86.745000 ;
        RECT 65.300000 86.955000 65.500000 87.155000 ;
        RECT 65.300000 87.365000 65.500000 87.565000 ;
        RECT 65.300000 87.775000 65.500000 87.975000 ;
        RECT 65.300000 88.185000 65.500000 88.385000 ;
        RECT 65.300000 88.595000 65.500000 88.795000 ;
        RECT 65.300000 89.005000 65.500000 89.205000 ;
        RECT 65.300000 89.415000 65.500000 89.615000 ;
        RECT 65.300000 89.825000 65.500000 90.025000 ;
        RECT 65.300000 90.235000 65.500000 90.435000 ;
        RECT 65.300000 90.645000 65.500000 90.845000 ;
        RECT 65.300000 91.055000 65.500000 91.255000 ;
        RECT 65.300000 91.465000 65.500000 91.665000 ;
        RECT 65.300000 91.875000 65.500000 92.075000 ;
        RECT 65.300000 92.285000 65.500000 92.485000 ;
        RECT 65.300000 92.695000 65.500000 92.895000 ;
        RECT 65.410000 68.125000 65.610000 68.325000 ;
        RECT 65.410000 68.535000 65.610000 68.735000 ;
        RECT 65.410000 68.945000 65.610000 69.145000 ;
        RECT 65.410000 69.355000 65.610000 69.555000 ;
        RECT 65.410000 69.765000 65.610000 69.965000 ;
        RECT 65.410000 70.175000 65.610000 70.375000 ;
        RECT 65.410000 70.585000 65.610000 70.785000 ;
        RECT 65.410000 70.995000 65.610000 71.195000 ;
        RECT 65.410000 71.405000 65.610000 71.605000 ;
        RECT 65.410000 71.815000 65.610000 72.015000 ;
        RECT 65.410000 72.225000 65.610000 72.425000 ;
        RECT 65.410000 72.635000 65.610000 72.835000 ;
        RECT 65.410000 73.045000 65.610000 73.245000 ;
        RECT 65.410000 73.450000 65.610000 73.650000 ;
        RECT 65.410000 73.855000 65.610000 74.055000 ;
        RECT 65.410000 74.260000 65.610000 74.460000 ;
        RECT 65.410000 74.665000 65.610000 74.865000 ;
        RECT 65.410000 75.070000 65.610000 75.270000 ;
        RECT 65.410000 75.475000 65.610000 75.675000 ;
        RECT 65.410000 75.880000 65.610000 76.080000 ;
        RECT 65.410000 76.285000 65.610000 76.485000 ;
        RECT 65.410000 76.690000 65.610000 76.890000 ;
        RECT 65.410000 77.095000 65.610000 77.295000 ;
        RECT 65.410000 77.500000 65.610000 77.700000 ;
        RECT 65.410000 77.905000 65.610000 78.105000 ;
        RECT 65.410000 78.310000 65.610000 78.510000 ;
        RECT 65.410000 78.715000 65.610000 78.915000 ;
        RECT 65.410000 79.120000 65.610000 79.320000 ;
        RECT 65.410000 79.525000 65.610000 79.725000 ;
        RECT 65.410000 79.930000 65.610000 80.130000 ;
        RECT 65.410000 80.335000 65.610000 80.535000 ;
        RECT 65.410000 80.740000 65.610000 80.940000 ;
        RECT 65.410000 81.145000 65.610000 81.345000 ;
        RECT 65.410000 81.550000 65.610000 81.750000 ;
        RECT 65.410000 81.955000 65.610000 82.155000 ;
        RECT 65.410000 82.360000 65.610000 82.560000 ;
        RECT 65.425000 17.860000 65.625000 18.060000 ;
        RECT 65.425000 18.290000 65.625000 18.490000 ;
        RECT 65.425000 18.720000 65.625000 18.920000 ;
        RECT 65.425000 19.150000 65.625000 19.350000 ;
        RECT 65.425000 19.580000 65.625000 19.780000 ;
        RECT 65.425000 20.010000 65.625000 20.210000 ;
        RECT 65.425000 20.440000 65.625000 20.640000 ;
        RECT 65.425000 20.870000 65.625000 21.070000 ;
        RECT 65.425000 21.300000 65.625000 21.500000 ;
        RECT 65.425000 21.730000 65.625000 21.930000 ;
        RECT 65.425000 22.160000 65.625000 22.360000 ;
        RECT 65.710000 82.855000 65.910000 83.055000 ;
        RECT 65.710000 83.265000 65.910000 83.465000 ;
        RECT 65.710000 83.675000 65.910000 83.875000 ;
        RECT 65.710000 84.085000 65.910000 84.285000 ;
        RECT 65.710000 84.495000 65.910000 84.695000 ;
        RECT 65.710000 84.905000 65.910000 85.105000 ;
        RECT 65.710000 85.315000 65.910000 85.515000 ;
        RECT 65.710000 85.725000 65.910000 85.925000 ;
        RECT 65.710000 86.135000 65.910000 86.335000 ;
        RECT 65.710000 86.545000 65.910000 86.745000 ;
        RECT 65.710000 86.955000 65.910000 87.155000 ;
        RECT 65.710000 87.365000 65.910000 87.565000 ;
        RECT 65.710000 87.775000 65.910000 87.975000 ;
        RECT 65.710000 88.185000 65.910000 88.385000 ;
        RECT 65.710000 88.595000 65.910000 88.795000 ;
        RECT 65.710000 89.005000 65.910000 89.205000 ;
        RECT 65.710000 89.415000 65.910000 89.615000 ;
        RECT 65.710000 89.825000 65.910000 90.025000 ;
        RECT 65.710000 90.235000 65.910000 90.435000 ;
        RECT 65.710000 90.645000 65.910000 90.845000 ;
        RECT 65.710000 91.055000 65.910000 91.255000 ;
        RECT 65.710000 91.465000 65.910000 91.665000 ;
        RECT 65.710000 91.875000 65.910000 92.075000 ;
        RECT 65.710000 92.285000 65.910000 92.485000 ;
        RECT 65.710000 92.695000 65.910000 92.895000 ;
        RECT 65.810000 68.125000 66.010000 68.325000 ;
        RECT 65.810000 68.535000 66.010000 68.735000 ;
        RECT 65.810000 68.945000 66.010000 69.145000 ;
        RECT 65.810000 69.355000 66.010000 69.555000 ;
        RECT 65.810000 69.765000 66.010000 69.965000 ;
        RECT 65.810000 70.175000 66.010000 70.375000 ;
        RECT 65.810000 70.585000 66.010000 70.785000 ;
        RECT 65.810000 70.995000 66.010000 71.195000 ;
        RECT 65.810000 71.405000 66.010000 71.605000 ;
        RECT 65.810000 71.815000 66.010000 72.015000 ;
        RECT 65.810000 72.225000 66.010000 72.425000 ;
        RECT 65.810000 72.635000 66.010000 72.835000 ;
        RECT 65.810000 73.045000 66.010000 73.245000 ;
        RECT 65.810000 73.450000 66.010000 73.650000 ;
        RECT 65.810000 73.855000 66.010000 74.055000 ;
        RECT 65.810000 74.260000 66.010000 74.460000 ;
        RECT 65.810000 74.665000 66.010000 74.865000 ;
        RECT 65.810000 75.070000 66.010000 75.270000 ;
        RECT 65.810000 75.475000 66.010000 75.675000 ;
        RECT 65.810000 75.880000 66.010000 76.080000 ;
        RECT 65.810000 76.285000 66.010000 76.485000 ;
        RECT 65.810000 76.690000 66.010000 76.890000 ;
        RECT 65.810000 77.095000 66.010000 77.295000 ;
        RECT 65.810000 77.500000 66.010000 77.700000 ;
        RECT 65.810000 77.905000 66.010000 78.105000 ;
        RECT 65.810000 78.310000 66.010000 78.510000 ;
        RECT 65.810000 78.715000 66.010000 78.915000 ;
        RECT 65.810000 79.120000 66.010000 79.320000 ;
        RECT 65.810000 79.525000 66.010000 79.725000 ;
        RECT 65.810000 79.930000 66.010000 80.130000 ;
        RECT 65.810000 80.335000 66.010000 80.535000 ;
        RECT 65.810000 80.740000 66.010000 80.940000 ;
        RECT 65.810000 81.145000 66.010000 81.345000 ;
        RECT 65.810000 81.550000 66.010000 81.750000 ;
        RECT 65.810000 81.955000 66.010000 82.155000 ;
        RECT 65.810000 82.360000 66.010000 82.560000 ;
        RECT 65.830000 17.860000 66.030000 18.060000 ;
        RECT 65.830000 18.290000 66.030000 18.490000 ;
        RECT 65.830000 18.720000 66.030000 18.920000 ;
        RECT 65.830000 19.150000 66.030000 19.350000 ;
        RECT 65.830000 19.580000 66.030000 19.780000 ;
        RECT 65.830000 20.010000 66.030000 20.210000 ;
        RECT 65.830000 20.440000 66.030000 20.640000 ;
        RECT 65.830000 20.870000 66.030000 21.070000 ;
        RECT 65.830000 21.300000 66.030000 21.500000 ;
        RECT 65.830000 21.730000 66.030000 21.930000 ;
        RECT 65.830000 22.160000 66.030000 22.360000 ;
        RECT 66.120000 82.855000 66.320000 83.055000 ;
        RECT 66.120000 83.265000 66.320000 83.465000 ;
        RECT 66.120000 83.675000 66.320000 83.875000 ;
        RECT 66.120000 84.085000 66.320000 84.285000 ;
        RECT 66.120000 84.495000 66.320000 84.695000 ;
        RECT 66.120000 84.905000 66.320000 85.105000 ;
        RECT 66.120000 85.315000 66.320000 85.515000 ;
        RECT 66.120000 85.725000 66.320000 85.925000 ;
        RECT 66.120000 86.135000 66.320000 86.335000 ;
        RECT 66.120000 86.545000 66.320000 86.745000 ;
        RECT 66.120000 86.955000 66.320000 87.155000 ;
        RECT 66.120000 87.365000 66.320000 87.565000 ;
        RECT 66.120000 87.775000 66.320000 87.975000 ;
        RECT 66.120000 88.185000 66.320000 88.385000 ;
        RECT 66.120000 88.595000 66.320000 88.795000 ;
        RECT 66.120000 89.005000 66.320000 89.205000 ;
        RECT 66.120000 89.415000 66.320000 89.615000 ;
        RECT 66.120000 89.825000 66.320000 90.025000 ;
        RECT 66.120000 90.235000 66.320000 90.435000 ;
        RECT 66.120000 90.645000 66.320000 90.845000 ;
        RECT 66.120000 91.055000 66.320000 91.255000 ;
        RECT 66.120000 91.465000 66.320000 91.665000 ;
        RECT 66.120000 91.875000 66.320000 92.075000 ;
        RECT 66.120000 92.285000 66.320000 92.485000 ;
        RECT 66.120000 92.695000 66.320000 92.895000 ;
        RECT 66.210000 68.125000 66.410000 68.325000 ;
        RECT 66.210000 68.535000 66.410000 68.735000 ;
        RECT 66.210000 68.945000 66.410000 69.145000 ;
        RECT 66.210000 69.355000 66.410000 69.555000 ;
        RECT 66.210000 69.765000 66.410000 69.965000 ;
        RECT 66.210000 70.175000 66.410000 70.375000 ;
        RECT 66.210000 70.585000 66.410000 70.785000 ;
        RECT 66.210000 70.995000 66.410000 71.195000 ;
        RECT 66.210000 71.405000 66.410000 71.605000 ;
        RECT 66.210000 71.815000 66.410000 72.015000 ;
        RECT 66.210000 72.225000 66.410000 72.425000 ;
        RECT 66.210000 72.635000 66.410000 72.835000 ;
        RECT 66.210000 73.045000 66.410000 73.245000 ;
        RECT 66.210000 73.450000 66.410000 73.650000 ;
        RECT 66.210000 73.855000 66.410000 74.055000 ;
        RECT 66.210000 74.260000 66.410000 74.460000 ;
        RECT 66.210000 74.665000 66.410000 74.865000 ;
        RECT 66.210000 75.070000 66.410000 75.270000 ;
        RECT 66.210000 75.475000 66.410000 75.675000 ;
        RECT 66.210000 75.880000 66.410000 76.080000 ;
        RECT 66.210000 76.285000 66.410000 76.485000 ;
        RECT 66.210000 76.690000 66.410000 76.890000 ;
        RECT 66.210000 77.095000 66.410000 77.295000 ;
        RECT 66.210000 77.500000 66.410000 77.700000 ;
        RECT 66.210000 77.905000 66.410000 78.105000 ;
        RECT 66.210000 78.310000 66.410000 78.510000 ;
        RECT 66.210000 78.715000 66.410000 78.915000 ;
        RECT 66.210000 79.120000 66.410000 79.320000 ;
        RECT 66.210000 79.525000 66.410000 79.725000 ;
        RECT 66.210000 79.930000 66.410000 80.130000 ;
        RECT 66.210000 80.335000 66.410000 80.535000 ;
        RECT 66.210000 80.740000 66.410000 80.940000 ;
        RECT 66.210000 81.145000 66.410000 81.345000 ;
        RECT 66.210000 81.550000 66.410000 81.750000 ;
        RECT 66.210000 81.955000 66.410000 82.155000 ;
        RECT 66.210000 82.360000 66.410000 82.560000 ;
        RECT 66.235000 17.860000 66.435000 18.060000 ;
        RECT 66.235000 18.290000 66.435000 18.490000 ;
        RECT 66.235000 18.720000 66.435000 18.920000 ;
        RECT 66.235000 19.150000 66.435000 19.350000 ;
        RECT 66.235000 19.580000 66.435000 19.780000 ;
        RECT 66.235000 20.010000 66.435000 20.210000 ;
        RECT 66.235000 20.440000 66.435000 20.640000 ;
        RECT 66.235000 20.870000 66.435000 21.070000 ;
        RECT 66.235000 21.300000 66.435000 21.500000 ;
        RECT 66.235000 21.730000 66.435000 21.930000 ;
        RECT 66.235000 22.160000 66.435000 22.360000 ;
        RECT 66.530000 82.855000 66.730000 83.055000 ;
        RECT 66.530000 83.265000 66.730000 83.465000 ;
        RECT 66.530000 83.675000 66.730000 83.875000 ;
        RECT 66.530000 84.085000 66.730000 84.285000 ;
        RECT 66.530000 84.495000 66.730000 84.695000 ;
        RECT 66.530000 84.905000 66.730000 85.105000 ;
        RECT 66.530000 85.315000 66.730000 85.515000 ;
        RECT 66.530000 85.725000 66.730000 85.925000 ;
        RECT 66.530000 86.135000 66.730000 86.335000 ;
        RECT 66.530000 86.545000 66.730000 86.745000 ;
        RECT 66.530000 86.955000 66.730000 87.155000 ;
        RECT 66.530000 87.365000 66.730000 87.565000 ;
        RECT 66.530000 87.775000 66.730000 87.975000 ;
        RECT 66.530000 88.185000 66.730000 88.385000 ;
        RECT 66.530000 88.595000 66.730000 88.795000 ;
        RECT 66.530000 89.005000 66.730000 89.205000 ;
        RECT 66.530000 89.415000 66.730000 89.615000 ;
        RECT 66.530000 89.825000 66.730000 90.025000 ;
        RECT 66.530000 90.235000 66.730000 90.435000 ;
        RECT 66.530000 90.645000 66.730000 90.845000 ;
        RECT 66.530000 91.055000 66.730000 91.255000 ;
        RECT 66.530000 91.465000 66.730000 91.665000 ;
        RECT 66.530000 91.875000 66.730000 92.075000 ;
        RECT 66.530000 92.285000 66.730000 92.485000 ;
        RECT 66.530000 92.695000 66.730000 92.895000 ;
        RECT 66.610000 68.125000 66.810000 68.325000 ;
        RECT 66.610000 68.535000 66.810000 68.735000 ;
        RECT 66.610000 68.945000 66.810000 69.145000 ;
        RECT 66.610000 69.355000 66.810000 69.555000 ;
        RECT 66.610000 69.765000 66.810000 69.965000 ;
        RECT 66.610000 70.175000 66.810000 70.375000 ;
        RECT 66.610000 70.585000 66.810000 70.785000 ;
        RECT 66.610000 70.995000 66.810000 71.195000 ;
        RECT 66.610000 71.405000 66.810000 71.605000 ;
        RECT 66.610000 71.815000 66.810000 72.015000 ;
        RECT 66.610000 72.225000 66.810000 72.425000 ;
        RECT 66.610000 72.635000 66.810000 72.835000 ;
        RECT 66.610000 73.045000 66.810000 73.245000 ;
        RECT 66.610000 73.450000 66.810000 73.650000 ;
        RECT 66.610000 73.855000 66.810000 74.055000 ;
        RECT 66.610000 74.260000 66.810000 74.460000 ;
        RECT 66.610000 74.665000 66.810000 74.865000 ;
        RECT 66.610000 75.070000 66.810000 75.270000 ;
        RECT 66.610000 75.475000 66.810000 75.675000 ;
        RECT 66.610000 75.880000 66.810000 76.080000 ;
        RECT 66.610000 76.285000 66.810000 76.485000 ;
        RECT 66.610000 76.690000 66.810000 76.890000 ;
        RECT 66.610000 77.095000 66.810000 77.295000 ;
        RECT 66.610000 77.500000 66.810000 77.700000 ;
        RECT 66.610000 77.905000 66.810000 78.105000 ;
        RECT 66.610000 78.310000 66.810000 78.510000 ;
        RECT 66.610000 78.715000 66.810000 78.915000 ;
        RECT 66.610000 79.120000 66.810000 79.320000 ;
        RECT 66.610000 79.525000 66.810000 79.725000 ;
        RECT 66.610000 79.930000 66.810000 80.130000 ;
        RECT 66.610000 80.335000 66.810000 80.535000 ;
        RECT 66.610000 80.740000 66.810000 80.940000 ;
        RECT 66.610000 81.145000 66.810000 81.345000 ;
        RECT 66.610000 81.550000 66.810000 81.750000 ;
        RECT 66.610000 81.955000 66.810000 82.155000 ;
        RECT 66.610000 82.360000 66.810000 82.560000 ;
        RECT 66.640000 17.860000 66.840000 18.060000 ;
        RECT 66.640000 18.290000 66.840000 18.490000 ;
        RECT 66.640000 18.720000 66.840000 18.920000 ;
        RECT 66.640000 19.150000 66.840000 19.350000 ;
        RECT 66.640000 19.580000 66.840000 19.780000 ;
        RECT 66.640000 20.010000 66.840000 20.210000 ;
        RECT 66.640000 20.440000 66.840000 20.640000 ;
        RECT 66.640000 20.870000 66.840000 21.070000 ;
        RECT 66.640000 21.300000 66.840000 21.500000 ;
        RECT 66.640000 21.730000 66.840000 21.930000 ;
        RECT 66.640000 22.160000 66.840000 22.360000 ;
        RECT 66.940000 82.855000 67.140000 83.055000 ;
        RECT 66.940000 83.265000 67.140000 83.465000 ;
        RECT 66.940000 83.675000 67.140000 83.875000 ;
        RECT 66.940000 84.085000 67.140000 84.285000 ;
        RECT 66.940000 84.495000 67.140000 84.695000 ;
        RECT 66.940000 84.905000 67.140000 85.105000 ;
        RECT 66.940000 85.315000 67.140000 85.515000 ;
        RECT 66.940000 85.725000 67.140000 85.925000 ;
        RECT 66.940000 86.135000 67.140000 86.335000 ;
        RECT 66.940000 86.545000 67.140000 86.745000 ;
        RECT 66.940000 86.955000 67.140000 87.155000 ;
        RECT 66.940000 87.365000 67.140000 87.565000 ;
        RECT 66.940000 87.775000 67.140000 87.975000 ;
        RECT 66.940000 88.185000 67.140000 88.385000 ;
        RECT 66.940000 88.595000 67.140000 88.795000 ;
        RECT 66.940000 89.005000 67.140000 89.205000 ;
        RECT 66.940000 89.415000 67.140000 89.615000 ;
        RECT 66.940000 89.825000 67.140000 90.025000 ;
        RECT 66.940000 90.235000 67.140000 90.435000 ;
        RECT 66.940000 90.645000 67.140000 90.845000 ;
        RECT 66.940000 91.055000 67.140000 91.255000 ;
        RECT 66.940000 91.465000 67.140000 91.665000 ;
        RECT 66.940000 91.875000 67.140000 92.075000 ;
        RECT 66.940000 92.285000 67.140000 92.485000 ;
        RECT 66.940000 92.695000 67.140000 92.895000 ;
        RECT 67.010000 68.125000 67.210000 68.325000 ;
        RECT 67.010000 68.535000 67.210000 68.735000 ;
        RECT 67.010000 68.945000 67.210000 69.145000 ;
        RECT 67.010000 69.355000 67.210000 69.555000 ;
        RECT 67.010000 69.765000 67.210000 69.965000 ;
        RECT 67.010000 70.175000 67.210000 70.375000 ;
        RECT 67.010000 70.585000 67.210000 70.785000 ;
        RECT 67.010000 70.995000 67.210000 71.195000 ;
        RECT 67.010000 71.405000 67.210000 71.605000 ;
        RECT 67.010000 71.815000 67.210000 72.015000 ;
        RECT 67.010000 72.225000 67.210000 72.425000 ;
        RECT 67.010000 72.635000 67.210000 72.835000 ;
        RECT 67.010000 73.045000 67.210000 73.245000 ;
        RECT 67.010000 73.450000 67.210000 73.650000 ;
        RECT 67.010000 73.855000 67.210000 74.055000 ;
        RECT 67.010000 74.260000 67.210000 74.460000 ;
        RECT 67.010000 74.665000 67.210000 74.865000 ;
        RECT 67.010000 75.070000 67.210000 75.270000 ;
        RECT 67.010000 75.475000 67.210000 75.675000 ;
        RECT 67.010000 75.880000 67.210000 76.080000 ;
        RECT 67.010000 76.285000 67.210000 76.485000 ;
        RECT 67.010000 76.690000 67.210000 76.890000 ;
        RECT 67.010000 77.095000 67.210000 77.295000 ;
        RECT 67.010000 77.500000 67.210000 77.700000 ;
        RECT 67.010000 77.905000 67.210000 78.105000 ;
        RECT 67.010000 78.310000 67.210000 78.510000 ;
        RECT 67.010000 78.715000 67.210000 78.915000 ;
        RECT 67.010000 79.120000 67.210000 79.320000 ;
        RECT 67.010000 79.525000 67.210000 79.725000 ;
        RECT 67.010000 79.930000 67.210000 80.130000 ;
        RECT 67.010000 80.335000 67.210000 80.535000 ;
        RECT 67.010000 80.740000 67.210000 80.940000 ;
        RECT 67.010000 81.145000 67.210000 81.345000 ;
        RECT 67.010000 81.550000 67.210000 81.750000 ;
        RECT 67.010000 81.955000 67.210000 82.155000 ;
        RECT 67.010000 82.360000 67.210000 82.560000 ;
        RECT 67.045000 17.860000 67.245000 18.060000 ;
        RECT 67.045000 18.290000 67.245000 18.490000 ;
        RECT 67.045000 18.720000 67.245000 18.920000 ;
        RECT 67.045000 19.150000 67.245000 19.350000 ;
        RECT 67.045000 19.580000 67.245000 19.780000 ;
        RECT 67.045000 20.010000 67.245000 20.210000 ;
        RECT 67.045000 20.440000 67.245000 20.640000 ;
        RECT 67.045000 20.870000 67.245000 21.070000 ;
        RECT 67.045000 21.300000 67.245000 21.500000 ;
        RECT 67.045000 21.730000 67.245000 21.930000 ;
        RECT 67.045000 22.160000 67.245000 22.360000 ;
        RECT 67.350000 82.855000 67.550000 83.055000 ;
        RECT 67.350000 83.265000 67.550000 83.465000 ;
        RECT 67.350000 83.675000 67.550000 83.875000 ;
        RECT 67.350000 84.085000 67.550000 84.285000 ;
        RECT 67.350000 84.495000 67.550000 84.695000 ;
        RECT 67.350000 84.905000 67.550000 85.105000 ;
        RECT 67.350000 85.315000 67.550000 85.515000 ;
        RECT 67.350000 85.725000 67.550000 85.925000 ;
        RECT 67.350000 86.135000 67.550000 86.335000 ;
        RECT 67.350000 86.545000 67.550000 86.745000 ;
        RECT 67.350000 86.955000 67.550000 87.155000 ;
        RECT 67.350000 87.365000 67.550000 87.565000 ;
        RECT 67.350000 87.775000 67.550000 87.975000 ;
        RECT 67.350000 88.185000 67.550000 88.385000 ;
        RECT 67.350000 88.595000 67.550000 88.795000 ;
        RECT 67.350000 89.005000 67.550000 89.205000 ;
        RECT 67.350000 89.415000 67.550000 89.615000 ;
        RECT 67.350000 89.825000 67.550000 90.025000 ;
        RECT 67.350000 90.235000 67.550000 90.435000 ;
        RECT 67.350000 90.645000 67.550000 90.845000 ;
        RECT 67.350000 91.055000 67.550000 91.255000 ;
        RECT 67.350000 91.465000 67.550000 91.665000 ;
        RECT 67.350000 91.875000 67.550000 92.075000 ;
        RECT 67.350000 92.285000 67.550000 92.485000 ;
        RECT 67.350000 92.695000 67.550000 92.895000 ;
        RECT 67.410000 68.125000 67.610000 68.325000 ;
        RECT 67.410000 68.535000 67.610000 68.735000 ;
        RECT 67.410000 68.945000 67.610000 69.145000 ;
        RECT 67.410000 69.355000 67.610000 69.555000 ;
        RECT 67.410000 69.765000 67.610000 69.965000 ;
        RECT 67.410000 70.175000 67.610000 70.375000 ;
        RECT 67.410000 70.585000 67.610000 70.785000 ;
        RECT 67.410000 70.995000 67.610000 71.195000 ;
        RECT 67.410000 71.405000 67.610000 71.605000 ;
        RECT 67.410000 71.815000 67.610000 72.015000 ;
        RECT 67.410000 72.225000 67.610000 72.425000 ;
        RECT 67.410000 72.635000 67.610000 72.835000 ;
        RECT 67.410000 73.045000 67.610000 73.245000 ;
        RECT 67.410000 73.450000 67.610000 73.650000 ;
        RECT 67.410000 73.855000 67.610000 74.055000 ;
        RECT 67.410000 74.260000 67.610000 74.460000 ;
        RECT 67.410000 74.665000 67.610000 74.865000 ;
        RECT 67.410000 75.070000 67.610000 75.270000 ;
        RECT 67.410000 75.475000 67.610000 75.675000 ;
        RECT 67.410000 75.880000 67.610000 76.080000 ;
        RECT 67.410000 76.285000 67.610000 76.485000 ;
        RECT 67.410000 76.690000 67.610000 76.890000 ;
        RECT 67.410000 77.095000 67.610000 77.295000 ;
        RECT 67.410000 77.500000 67.610000 77.700000 ;
        RECT 67.410000 77.905000 67.610000 78.105000 ;
        RECT 67.410000 78.310000 67.610000 78.510000 ;
        RECT 67.410000 78.715000 67.610000 78.915000 ;
        RECT 67.410000 79.120000 67.610000 79.320000 ;
        RECT 67.410000 79.525000 67.610000 79.725000 ;
        RECT 67.410000 79.930000 67.610000 80.130000 ;
        RECT 67.410000 80.335000 67.610000 80.535000 ;
        RECT 67.410000 80.740000 67.610000 80.940000 ;
        RECT 67.410000 81.145000 67.610000 81.345000 ;
        RECT 67.410000 81.550000 67.610000 81.750000 ;
        RECT 67.410000 81.955000 67.610000 82.155000 ;
        RECT 67.410000 82.360000 67.610000 82.560000 ;
        RECT 67.450000 17.860000 67.650000 18.060000 ;
        RECT 67.450000 18.290000 67.650000 18.490000 ;
        RECT 67.450000 18.720000 67.650000 18.920000 ;
        RECT 67.450000 19.150000 67.650000 19.350000 ;
        RECT 67.450000 19.580000 67.650000 19.780000 ;
        RECT 67.450000 20.010000 67.650000 20.210000 ;
        RECT 67.450000 20.440000 67.650000 20.640000 ;
        RECT 67.450000 20.870000 67.650000 21.070000 ;
        RECT 67.450000 21.300000 67.650000 21.500000 ;
        RECT 67.450000 21.730000 67.650000 21.930000 ;
        RECT 67.450000 22.160000 67.650000 22.360000 ;
        RECT 67.760000 82.855000 67.960000 83.055000 ;
        RECT 67.760000 83.265000 67.960000 83.465000 ;
        RECT 67.760000 83.675000 67.960000 83.875000 ;
        RECT 67.760000 84.085000 67.960000 84.285000 ;
        RECT 67.760000 84.495000 67.960000 84.695000 ;
        RECT 67.760000 84.905000 67.960000 85.105000 ;
        RECT 67.760000 85.315000 67.960000 85.515000 ;
        RECT 67.760000 85.725000 67.960000 85.925000 ;
        RECT 67.760000 86.135000 67.960000 86.335000 ;
        RECT 67.760000 86.545000 67.960000 86.745000 ;
        RECT 67.760000 86.955000 67.960000 87.155000 ;
        RECT 67.760000 87.365000 67.960000 87.565000 ;
        RECT 67.760000 87.775000 67.960000 87.975000 ;
        RECT 67.760000 88.185000 67.960000 88.385000 ;
        RECT 67.760000 88.595000 67.960000 88.795000 ;
        RECT 67.760000 89.005000 67.960000 89.205000 ;
        RECT 67.760000 89.415000 67.960000 89.615000 ;
        RECT 67.760000 89.825000 67.960000 90.025000 ;
        RECT 67.760000 90.235000 67.960000 90.435000 ;
        RECT 67.760000 90.645000 67.960000 90.845000 ;
        RECT 67.760000 91.055000 67.960000 91.255000 ;
        RECT 67.760000 91.465000 67.960000 91.665000 ;
        RECT 67.760000 91.875000 67.960000 92.075000 ;
        RECT 67.760000 92.285000 67.960000 92.485000 ;
        RECT 67.760000 92.695000 67.960000 92.895000 ;
        RECT 67.810000 68.125000 68.010000 68.325000 ;
        RECT 67.810000 68.535000 68.010000 68.735000 ;
        RECT 67.810000 68.945000 68.010000 69.145000 ;
        RECT 67.810000 69.355000 68.010000 69.555000 ;
        RECT 67.810000 69.765000 68.010000 69.965000 ;
        RECT 67.810000 70.175000 68.010000 70.375000 ;
        RECT 67.810000 70.585000 68.010000 70.785000 ;
        RECT 67.810000 70.995000 68.010000 71.195000 ;
        RECT 67.810000 71.405000 68.010000 71.605000 ;
        RECT 67.810000 71.815000 68.010000 72.015000 ;
        RECT 67.810000 72.225000 68.010000 72.425000 ;
        RECT 67.810000 72.635000 68.010000 72.835000 ;
        RECT 67.810000 73.045000 68.010000 73.245000 ;
        RECT 67.810000 73.450000 68.010000 73.650000 ;
        RECT 67.810000 73.855000 68.010000 74.055000 ;
        RECT 67.810000 74.260000 68.010000 74.460000 ;
        RECT 67.810000 74.665000 68.010000 74.865000 ;
        RECT 67.810000 75.070000 68.010000 75.270000 ;
        RECT 67.810000 75.475000 68.010000 75.675000 ;
        RECT 67.810000 75.880000 68.010000 76.080000 ;
        RECT 67.810000 76.285000 68.010000 76.485000 ;
        RECT 67.810000 76.690000 68.010000 76.890000 ;
        RECT 67.810000 77.095000 68.010000 77.295000 ;
        RECT 67.810000 77.500000 68.010000 77.700000 ;
        RECT 67.810000 77.905000 68.010000 78.105000 ;
        RECT 67.810000 78.310000 68.010000 78.510000 ;
        RECT 67.810000 78.715000 68.010000 78.915000 ;
        RECT 67.810000 79.120000 68.010000 79.320000 ;
        RECT 67.810000 79.525000 68.010000 79.725000 ;
        RECT 67.810000 79.930000 68.010000 80.130000 ;
        RECT 67.810000 80.335000 68.010000 80.535000 ;
        RECT 67.810000 80.740000 68.010000 80.940000 ;
        RECT 67.810000 81.145000 68.010000 81.345000 ;
        RECT 67.810000 81.550000 68.010000 81.750000 ;
        RECT 67.810000 81.955000 68.010000 82.155000 ;
        RECT 67.810000 82.360000 68.010000 82.560000 ;
        RECT 67.855000 17.860000 68.055000 18.060000 ;
        RECT 67.855000 18.290000 68.055000 18.490000 ;
        RECT 67.855000 18.720000 68.055000 18.920000 ;
        RECT 67.855000 19.150000 68.055000 19.350000 ;
        RECT 67.855000 19.580000 68.055000 19.780000 ;
        RECT 67.855000 20.010000 68.055000 20.210000 ;
        RECT 67.855000 20.440000 68.055000 20.640000 ;
        RECT 67.855000 20.870000 68.055000 21.070000 ;
        RECT 67.855000 21.300000 68.055000 21.500000 ;
        RECT 67.855000 21.730000 68.055000 21.930000 ;
        RECT 67.855000 22.160000 68.055000 22.360000 ;
        RECT 68.170000 82.855000 68.370000 83.055000 ;
        RECT 68.170000 83.265000 68.370000 83.465000 ;
        RECT 68.170000 83.675000 68.370000 83.875000 ;
        RECT 68.170000 84.085000 68.370000 84.285000 ;
        RECT 68.170000 84.495000 68.370000 84.695000 ;
        RECT 68.170000 84.905000 68.370000 85.105000 ;
        RECT 68.170000 85.315000 68.370000 85.515000 ;
        RECT 68.170000 85.725000 68.370000 85.925000 ;
        RECT 68.170000 86.135000 68.370000 86.335000 ;
        RECT 68.170000 86.545000 68.370000 86.745000 ;
        RECT 68.170000 86.955000 68.370000 87.155000 ;
        RECT 68.170000 87.365000 68.370000 87.565000 ;
        RECT 68.170000 87.775000 68.370000 87.975000 ;
        RECT 68.170000 88.185000 68.370000 88.385000 ;
        RECT 68.170000 88.595000 68.370000 88.795000 ;
        RECT 68.170000 89.005000 68.370000 89.205000 ;
        RECT 68.170000 89.415000 68.370000 89.615000 ;
        RECT 68.170000 89.825000 68.370000 90.025000 ;
        RECT 68.170000 90.235000 68.370000 90.435000 ;
        RECT 68.170000 90.645000 68.370000 90.845000 ;
        RECT 68.170000 91.055000 68.370000 91.255000 ;
        RECT 68.170000 91.465000 68.370000 91.665000 ;
        RECT 68.170000 91.875000 68.370000 92.075000 ;
        RECT 68.170000 92.285000 68.370000 92.485000 ;
        RECT 68.170000 92.695000 68.370000 92.895000 ;
        RECT 68.210000 68.125000 68.410000 68.325000 ;
        RECT 68.210000 68.535000 68.410000 68.735000 ;
        RECT 68.210000 68.945000 68.410000 69.145000 ;
        RECT 68.210000 69.355000 68.410000 69.555000 ;
        RECT 68.210000 69.765000 68.410000 69.965000 ;
        RECT 68.210000 70.175000 68.410000 70.375000 ;
        RECT 68.210000 70.585000 68.410000 70.785000 ;
        RECT 68.210000 70.995000 68.410000 71.195000 ;
        RECT 68.210000 71.405000 68.410000 71.605000 ;
        RECT 68.210000 71.815000 68.410000 72.015000 ;
        RECT 68.210000 72.225000 68.410000 72.425000 ;
        RECT 68.210000 72.635000 68.410000 72.835000 ;
        RECT 68.210000 73.045000 68.410000 73.245000 ;
        RECT 68.210000 73.450000 68.410000 73.650000 ;
        RECT 68.210000 73.855000 68.410000 74.055000 ;
        RECT 68.210000 74.260000 68.410000 74.460000 ;
        RECT 68.210000 74.665000 68.410000 74.865000 ;
        RECT 68.210000 75.070000 68.410000 75.270000 ;
        RECT 68.210000 75.475000 68.410000 75.675000 ;
        RECT 68.210000 75.880000 68.410000 76.080000 ;
        RECT 68.210000 76.285000 68.410000 76.485000 ;
        RECT 68.210000 76.690000 68.410000 76.890000 ;
        RECT 68.210000 77.095000 68.410000 77.295000 ;
        RECT 68.210000 77.500000 68.410000 77.700000 ;
        RECT 68.210000 77.905000 68.410000 78.105000 ;
        RECT 68.210000 78.310000 68.410000 78.510000 ;
        RECT 68.210000 78.715000 68.410000 78.915000 ;
        RECT 68.210000 79.120000 68.410000 79.320000 ;
        RECT 68.210000 79.525000 68.410000 79.725000 ;
        RECT 68.210000 79.930000 68.410000 80.130000 ;
        RECT 68.210000 80.335000 68.410000 80.535000 ;
        RECT 68.210000 80.740000 68.410000 80.940000 ;
        RECT 68.210000 81.145000 68.410000 81.345000 ;
        RECT 68.210000 81.550000 68.410000 81.750000 ;
        RECT 68.210000 81.955000 68.410000 82.155000 ;
        RECT 68.210000 82.360000 68.410000 82.560000 ;
        RECT 68.260000 17.860000 68.460000 18.060000 ;
        RECT 68.260000 18.290000 68.460000 18.490000 ;
        RECT 68.260000 18.720000 68.460000 18.920000 ;
        RECT 68.260000 19.150000 68.460000 19.350000 ;
        RECT 68.260000 19.580000 68.460000 19.780000 ;
        RECT 68.260000 20.010000 68.460000 20.210000 ;
        RECT 68.260000 20.440000 68.460000 20.640000 ;
        RECT 68.260000 20.870000 68.460000 21.070000 ;
        RECT 68.260000 21.300000 68.460000 21.500000 ;
        RECT 68.260000 21.730000 68.460000 21.930000 ;
        RECT 68.260000 22.160000 68.460000 22.360000 ;
        RECT 68.580000 82.855000 68.780000 83.055000 ;
        RECT 68.580000 83.265000 68.780000 83.465000 ;
        RECT 68.580000 83.675000 68.780000 83.875000 ;
        RECT 68.580000 84.085000 68.780000 84.285000 ;
        RECT 68.580000 84.495000 68.780000 84.695000 ;
        RECT 68.580000 84.905000 68.780000 85.105000 ;
        RECT 68.580000 85.315000 68.780000 85.515000 ;
        RECT 68.580000 85.725000 68.780000 85.925000 ;
        RECT 68.580000 86.135000 68.780000 86.335000 ;
        RECT 68.580000 86.545000 68.780000 86.745000 ;
        RECT 68.580000 86.955000 68.780000 87.155000 ;
        RECT 68.580000 87.365000 68.780000 87.565000 ;
        RECT 68.580000 87.775000 68.780000 87.975000 ;
        RECT 68.580000 88.185000 68.780000 88.385000 ;
        RECT 68.580000 88.595000 68.780000 88.795000 ;
        RECT 68.580000 89.005000 68.780000 89.205000 ;
        RECT 68.580000 89.415000 68.780000 89.615000 ;
        RECT 68.580000 89.825000 68.780000 90.025000 ;
        RECT 68.580000 90.235000 68.780000 90.435000 ;
        RECT 68.580000 90.645000 68.780000 90.845000 ;
        RECT 68.580000 91.055000 68.780000 91.255000 ;
        RECT 68.580000 91.465000 68.780000 91.665000 ;
        RECT 68.580000 91.875000 68.780000 92.075000 ;
        RECT 68.580000 92.285000 68.780000 92.485000 ;
        RECT 68.580000 92.695000 68.780000 92.895000 ;
        RECT 68.610000 68.125000 68.810000 68.325000 ;
        RECT 68.610000 68.535000 68.810000 68.735000 ;
        RECT 68.610000 68.945000 68.810000 69.145000 ;
        RECT 68.610000 69.355000 68.810000 69.555000 ;
        RECT 68.610000 69.765000 68.810000 69.965000 ;
        RECT 68.610000 70.175000 68.810000 70.375000 ;
        RECT 68.610000 70.585000 68.810000 70.785000 ;
        RECT 68.610000 70.995000 68.810000 71.195000 ;
        RECT 68.610000 71.405000 68.810000 71.605000 ;
        RECT 68.610000 71.815000 68.810000 72.015000 ;
        RECT 68.610000 72.225000 68.810000 72.425000 ;
        RECT 68.610000 72.635000 68.810000 72.835000 ;
        RECT 68.610000 73.045000 68.810000 73.245000 ;
        RECT 68.610000 73.450000 68.810000 73.650000 ;
        RECT 68.610000 73.855000 68.810000 74.055000 ;
        RECT 68.610000 74.260000 68.810000 74.460000 ;
        RECT 68.610000 74.665000 68.810000 74.865000 ;
        RECT 68.610000 75.070000 68.810000 75.270000 ;
        RECT 68.610000 75.475000 68.810000 75.675000 ;
        RECT 68.610000 75.880000 68.810000 76.080000 ;
        RECT 68.610000 76.285000 68.810000 76.485000 ;
        RECT 68.610000 76.690000 68.810000 76.890000 ;
        RECT 68.610000 77.095000 68.810000 77.295000 ;
        RECT 68.610000 77.500000 68.810000 77.700000 ;
        RECT 68.610000 77.905000 68.810000 78.105000 ;
        RECT 68.610000 78.310000 68.810000 78.510000 ;
        RECT 68.610000 78.715000 68.810000 78.915000 ;
        RECT 68.610000 79.120000 68.810000 79.320000 ;
        RECT 68.610000 79.525000 68.810000 79.725000 ;
        RECT 68.610000 79.930000 68.810000 80.130000 ;
        RECT 68.610000 80.335000 68.810000 80.535000 ;
        RECT 68.610000 80.740000 68.810000 80.940000 ;
        RECT 68.610000 81.145000 68.810000 81.345000 ;
        RECT 68.610000 81.550000 68.810000 81.750000 ;
        RECT 68.610000 81.955000 68.810000 82.155000 ;
        RECT 68.610000 82.360000 68.810000 82.560000 ;
        RECT 68.665000 17.860000 68.865000 18.060000 ;
        RECT 68.665000 18.290000 68.865000 18.490000 ;
        RECT 68.665000 18.720000 68.865000 18.920000 ;
        RECT 68.665000 19.150000 68.865000 19.350000 ;
        RECT 68.665000 19.580000 68.865000 19.780000 ;
        RECT 68.665000 20.010000 68.865000 20.210000 ;
        RECT 68.665000 20.440000 68.865000 20.640000 ;
        RECT 68.665000 20.870000 68.865000 21.070000 ;
        RECT 68.665000 21.300000 68.865000 21.500000 ;
        RECT 68.665000 21.730000 68.865000 21.930000 ;
        RECT 68.665000 22.160000 68.865000 22.360000 ;
        RECT 68.990000 82.855000 69.190000 83.055000 ;
        RECT 68.990000 83.265000 69.190000 83.465000 ;
        RECT 68.990000 83.675000 69.190000 83.875000 ;
        RECT 68.990000 84.085000 69.190000 84.285000 ;
        RECT 68.990000 84.495000 69.190000 84.695000 ;
        RECT 68.990000 84.905000 69.190000 85.105000 ;
        RECT 68.990000 85.315000 69.190000 85.515000 ;
        RECT 68.990000 85.725000 69.190000 85.925000 ;
        RECT 68.990000 86.135000 69.190000 86.335000 ;
        RECT 68.990000 86.545000 69.190000 86.745000 ;
        RECT 68.990000 86.955000 69.190000 87.155000 ;
        RECT 68.990000 87.365000 69.190000 87.565000 ;
        RECT 68.990000 87.775000 69.190000 87.975000 ;
        RECT 68.990000 88.185000 69.190000 88.385000 ;
        RECT 68.990000 88.595000 69.190000 88.795000 ;
        RECT 68.990000 89.005000 69.190000 89.205000 ;
        RECT 68.990000 89.415000 69.190000 89.615000 ;
        RECT 68.990000 89.825000 69.190000 90.025000 ;
        RECT 68.990000 90.235000 69.190000 90.435000 ;
        RECT 68.990000 90.645000 69.190000 90.845000 ;
        RECT 68.990000 91.055000 69.190000 91.255000 ;
        RECT 68.990000 91.465000 69.190000 91.665000 ;
        RECT 68.990000 91.875000 69.190000 92.075000 ;
        RECT 68.990000 92.285000 69.190000 92.485000 ;
        RECT 68.990000 92.695000 69.190000 92.895000 ;
        RECT 69.010000 68.125000 69.210000 68.325000 ;
        RECT 69.010000 68.535000 69.210000 68.735000 ;
        RECT 69.010000 68.945000 69.210000 69.145000 ;
        RECT 69.010000 69.355000 69.210000 69.555000 ;
        RECT 69.010000 69.765000 69.210000 69.965000 ;
        RECT 69.010000 70.175000 69.210000 70.375000 ;
        RECT 69.010000 70.585000 69.210000 70.785000 ;
        RECT 69.010000 70.995000 69.210000 71.195000 ;
        RECT 69.010000 71.405000 69.210000 71.605000 ;
        RECT 69.010000 71.815000 69.210000 72.015000 ;
        RECT 69.010000 72.225000 69.210000 72.425000 ;
        RECT 69.010000 72.635000 69.210000 72.835000 ;
        RECT 69.010000 73.045000 69.210000 73.245000 ;
        RECT 69.010000 73.450000 69.210000 73.650000 ;
        RECT 69.010000 73.855000 69.210000 74.055000 ;
        RECT 69.010000 74.260000 69.210000 74.460000 ;
        RECT 69.010000 74.665000 69.210000 74.865000 ;
        RECT 69.010000 75.070000 69.210000 75.270000 ;
        RECT 69.010000 75.475000 69.210000 75.675000 ;
        RECT 69.010000 75.880000 69.210000 76.080000 ;
        RECT 69.010000 76.285000 69.210000 76.485000 ;
        RECT 69.010000 76.690000 69.210000 76.890000 ;
        RECT 69.010000 77.095000 69.210000 77.295000 ;
        RECT 69.010000 77.500000 69.210000 77.700000 ;
        RECT 69.010000 77.905000 69.210000 78.105000 ;
        RECT 69.010000 78.310000 69.210000 78.510000 ;
        RECT 69.010000 78.715000 69.210000 78.915000 ;
        RECT 69.010000 79.120000 69.210000 79.320000 ;
        RECT 69.010000 79.525000 69.210000 79.725000 ;
        RECT 69.010000 79.930000 69.210000 80.130000 ;
        RECT 69.010000 80.335000 69.210000 80.535000 ;
        RECT 69.010000 80.740000 69.210000 80.940000 ;
        RECT 69.010000 81.145000 69.210000 81.345000 ;
        RECT 69.010000 81.550000 69.210000 81.750000 ;
        RECT 69.010000 81.955000 69.210000 82.155000 ;
        RECT 69.010000 82.360000 69.210000 82.560000 ;
        RECT 69.070000 17.860000 69.270000 18.060000 ;
        RECT 69.070000 18.290000 69.270000 18.490000 ;
        RECT 69.070000 18.720000 69.270000 18.920000 ;
        RECT 69.070000 19.150000 69.270000 19.350000 ;
        RECT 69.070000 19.580000 69.270000 19.780000 ;
        RECT 69.070000 20.010000 69.270000 20.210000 ;
        RECT 69.070000 20.440000 69.270000 20.640000 ;
        RECT 69.070000 20.870000 69.270000 21.070000 ;
        RECT 69.070000 21.300000 69.270000 21.500000 ;
        RECT 69.070000 21.730000 69.270000 21.930000 ;
        RECT 69.070000 22.160000 69.270000 22.360000 ;
        RECT 69.400000 82.855000 69.600000 83.055000 ;
        RECT 69.400000 83.265000 69.600000 83.465000 ;
        RECT 69.400000 83.675000 69.600000 83.875000 ;
        RECT 69.400000 84.085000 69.600000 84.285000 ;
        RECT 69.400000 84.495000 69.600000 84.695000 ;
        RECT 69.400000 84.905000 69.600000 85.105000 ;
        RECT 69.400000 85.315000 69.600000 85.515000 ;
        RECT 69.400000 85.725000 69.600000 85.925000 ;
        RECT 69.400000 86.135000 69.600000 86.335000 ;
        RECT 69.400000 86.545000 69.600000 86.745000 ;
        RECT 69.400000 86.955000 69.600000 87.155000 ;
        RECT 69.400000 87.365000 69.600000 87.565000 ;
        RECT 69.400000 87.775000 69.600000 87.975000 ;
        RECT 69.400000 88.185000 69.600000 88.385000 ;
        RECT 69.400000 88.595000 69.600000 88.795000 ;
        RECT 69.400000 89.005000 69.600000 89.205000 ;
        RECT 69.400000 89.415000 69.600000 89.615000 ;
        RECT 69.400000 89.825000 69.600000 90.025000 ;
        RECT 69.400000 90.235000 69.600000 90.435000 ;
        RECT 69.400000 90.645000 69.600000 90.845000 ;
        RECT 69.400000 91.055000 69.600000 91.255000 ;
        RECT 69.400000 91.465000 69.600000 91.665000 ;
        RECT 69.400000 91.875000 69.600000 92.075000 ;
        RECT 69.400000 92.285000 69.600000 92.485000 ;
        RECT 69.400000 92.695000 69.600000 92.895000 ;
        RECT 69.410000 68.125000 69.610000 68.325000 ;
        RECT 69.410000 68.535000 69.610000 68.735000 ;
        RECT 69.410000 68.945000 69.610000 69.145000 ;
        RECT 69.410000 69.355000 69.610000 69.555000 ;
        RECT 69.410000 69.765000 69.610000 69.965000 ;
        RECT 69.410000 70.175000 69.610000 70.375000 ;
        RECT 69.410000 70.585000 69.610000 70.785000 ;
        RECT 69.410000 70.995000 69.610000 71.195000 ;
        RECT 69.410000 71.405000 69.610000 71.605000 ;
        RECT 69.410000 71.815000 69.610000 72.015000 ;
        RECT 69.410000 72.225000 69.610000 72.425000 ;
        RECT 69.410000 72.635000 69.610000 72.835000 ;
        RECT 69.410000 73.045000 69.610000 73.245000 ;
        RECT 69.410000 73.450000 69.610000 73.650000 ;
        RECT 69.410000 73.855000 69.610000 74.055000 ;
        RECT 69.410000 74.260000 69.610000 74.460000 ;
        RECT 69.410000 74.665000 69.610000 74.865000 ;
        RECT 69.410000 75.070000 69.610000 75.270000 ;
        RECT 69.410000 75.475000 69.610000 75.675000 ;
        RECT 69.410000 75.880000 69.610000 76.080000 ;
        RECT 69.410000 76.285000 69.610000 76.485000 ;
        RECT 69.410000 76.690000 69.610000 76.890000 ;
        RECT 69.410000 77.095000 69.610000 77.295000 ;
        RECT 69.410000 77.500000 69.610000 77.700000 ;
        RECT 69.410000 77.905000 69.610000 78.105000 ;
        RECT 69.410000 78.310000 69.610000 78.510000 ;
        RECT 69.410000 78.715000 69.610000 78.915000 ;
        RECT 69.410000 79.120000 69.610000 79.320000 ;
        RECT 69.410000 79.525000 69.610000 79.725000 ;
        RECT 69.410000 79.930000 69.610000 80.130000 ;
        RECT 69.410000 80.335000 69.610000 80.535000 ;
        RECT 69.410000 80.740000 69.610000 80.940000 ;
        RECT 69.410000 81.145000 69.610000 81.345000 ;
        RECT 69.410000 81.550000 69.610000 81.750000 ;
        RECT 69.410000 81.955000 69.610000 82.155000 ;
        RECT 69.410000 82.360000 69.610000 82.560000 ;
        RECT 69.475000 17.860000 69.675000 18.060000 ;
        RECT 69.475000 18.290000 69.675000 18.490000 ;
        RECT 69.475000 18.720000 69.675000 18.920000 ;
        RECT 69.475000 19.150000 69.675000 19.350000 ;
        RECT 69.475000 19.580000 69.675000 19.780000 ;
        RECT 69.475000 20.010000 69.675000 20.210000 ;
        RECT 69.475000 20.440000 69.675000 20.640000 ;
        RECT 69.475000 20.870000 69.675000 21.070000 ;
        RECT 69.475000 21.300000 69.675000 21.500000 ;
        RECT 69.475000 21.730000 69.675000 21.930000 ;
        RECT 69.475000 22.160000 69.675000 22.360000 ;
        RECT 69.810000 68.125000 70.010000 68.325000 ;
        RECT 69.810000 68.535000 70.010000 68.735000 ;
        RECT 69.810000 68.945000 70.010000 69.145000 ;
        RECT 69.810000 69.355000 70.010000 69.555000 ;
        RECT 69.810000 69.765000 70.010000 69.965000 ;
        RECT 69.810000 70.175000 70.010000 70.375000 ;
        RECT 69.810000 70.585000 70.010000 70.785000 ;
        RECT 69.810000 70.995000 70.010000 71.195000 ;
        RECT 69.810000 71.405000 70.010000 71.605000 ;
        RECT 69.810000 71.815000 70.010000 72.015000 ;
        RECT 69.810000 72.225000 70.010000 72.425000 ;
        RECT 69.810000 72.635000 70.010000 72.835000 ;
        RECT 69.810000 73.045000 70.010000 73.245000 ;
        RECT 69.810000 73.450000 70.010000 73.650000 ;
        RECT 69.810000 73.855000 70.010000 74.055000 ;
        RECT 69.810000 74.260000 70.010000 74.460000 ;
        RECT 69.810000 74.665000 70.010000 74.865000 ;
        RECT 69.810000 75.070000 70.010000 75.270000 ;
        RECT 69.810000 75.475000 70.010000 75.675000 ;
        RECT 69.810000 75.880000 70.010000 76.080000 ;
        RECT 69.810000 76.285000 70.010000 76.485000 ;
        RECT 69.810000 76.690000 70.010000 76.890000 ;
        RECT 69.810000 77.095000 70.010000 77.295000 ;
        RECT 69.810000 77.500000 70.010000 77.700000 ;
        RECT 69.810000 77.905000 70.010000 78.105000 ;
        RECT 69.810000 78.310000 70.010000 78.510000 ;
        RECT 69.810000 78.715000 70.010000 78.915000 ;
        RECT 69.810000 79.120000 70.010000 79.320000 ;
        RECT 69.810000 79.525000 70.010000 79.725000 ;
        RECT 69.810000 79.930000 70.010000 80.130000 ;
        RECT 69.810000 80.335000 70.010000 80.535000 ;
        RECT 69.810000 80.740000 70.010000 80.940000 ;
        RECT 69.810000 81.145000 70.010000 81.345000 ;
        RECT 69.810000 81.550000 70.010000 81.750000 ;
        RECT 69.810000 81.955000 70.010000 82.155000 ;
        RECT 69.810000 82.360000 70.010000 82.560000 ;
        RECT 69.810000 82.855000 70.010000 83.055000 ;
        RECT 69.810000 83.265000 70.010000 83.465000 ;
        RECT 69.810000 83.675000 70.010000 83.875000 ;
        RECT 69.810000 84.085000 70.010000 84.285000 ;
        RECT 69.810000 84.495000 70.010000 84.695000 ;
        RECT 69.810000 84.905000 70.010000 85.105000 ;
        RECT 69.810000 85.315000 70.010000 85.515000 ;
        RECT 69.810000 85.725000 70.010000 85.925000 ;
        RECT 69.810000 86.135000 70.010000 86.335000 ;
        RECT 69.810000 86.545000 70.010000 86.745000 ;
        RECT 69.810000 86.955000 70.010000 87.155000 ;
        RECT 69.810000 87.365000 70.010000 87.565000 ;
        RECT 69.810000 87.775000 70.010000 87.975000 ;
        RECT 69.810000 88.185000 70.010000 88.385000 ;
        RECT 69.810000 88.595000 70.010000 88.795000 ;
        RECT 69.810000 89.005000 70.010000 89.205000 ;
        RECT 69.810000 89.415000 70.010000 89.615000 ;
        RECT 69.810000 89.825000 70.010000 90.025000 ;
        RECT 69.810000 90.235000 70.010000 90.435000 ;
        RECT 69.810000 90.645000 70.010000 90.845000 ;
        RECT 69.810000 91.055000 70.010000 91.255000 ;
        RECT 69.810000 91.465000 70.010000 91.665000 ;
        RECT 69.810000 91.875000 70.010000 92.075000 ;
        RECT 69.810000 92.285000 70.010000 92.485000 ;
        RECT 69.810000 92.695000 70.010000 92.895000 ;
        RECT 69.880000 17.860000 70.080000 18.060000 ;
        RECT 69.880000 18.290000 70.080000 18.490000 ;
        RECT 69.880000 18.720000 70.080000 18.920000 ;
        RECT 69.880000 19.150000 70.080000 19.350000 ;
        RECT 69.880000 19.580000 70.080000 19.780000 ;
        RECT 69.880000 20.010000 70.080000 20.210000 ;
        RECT 69.880000 20.440000 70.080000 20.640000 ;
        RECT 69.880000 20.870000 70.080000 21.070000 ;
        RECT 69.880000 21.300000 70.080000 21.500000 ;
        RECT 69.880000 21.730000 70.080000 21.930000 ;
        RECT 69.880000 22.160000 70.080000 22.360000 ;
        RECT 70.210000 68.125000 70.410000 68.325000 ;
        RECT 70.210000 68.535000 70.410000 68.735000 ;
        RECT 70.210000 68.945000 70.410000 69.145000 ;
        RECT 70.210000 69.355000 70.410000 69.555000 ;
        RECT 70.210000 69.765000 70.410000 69.965000 ;
        RECT 70.210000 70.175000 70.410000 70.375000 ;
        RECT 70.210000 70.585000 70.410000 70.785000 ;
        RECT 70.210000 70.995000 70.410000 71.195000 ;
        RECT 70.210000 71.405000 70.410000 71.605000 ;
        RECT 70.210000 71.815000 70.410000 72.015000 ;
        RECT 70.210000 72.225000 70.410000 72.425000 ;
        RECT 70.210000 72.635000 70.410000 72.835000 ;
        RECT 70.210000 73.045000 70.410000 73.245000 ;
        RECT 70.210000 73.450000 70.410000 73.650000 ;
        RECT 70.210000 73.855000 70.410000 74.055000 ;
        RECT 70.210000 74.260000 70.410000 74.460000 ;
        RECT 70.210000 74.665000 70.410000 74.865000 ;
        RECT 70.210000 75.070000 70.410000 75.270000 ;
        RECT 70.210000 75.475000 70.410000 75.675000 ;
        RECT 70.210000 75.880000 70.410000 76.080000 ;
        RECT 70.210000 76.285000 70.410000 76.485000 ;
        RECT 70.210000 76.690000 70.410000 76.890000 ;
        RECT 70.210000 77.095000 70.410000 77.295000 ;
        RECT 70.210000 77.500000 70.410000 77.700000 ;
        RECT 70.210000 77.905000 70.410000 78.105000 ;
        RECT 70.210000 78.310000 70.410000 78.510000 ;
        RECT 70.210000 78.715000 70.410000 78.915000 ;
        RECT 70.210000 79.120000 70.410000 79.320000 ;
        RECT 70.210000 79.525000 70.410000 79.725000 ;
        RECT 70.210000 79.930000 70.410000 80.130000 ;
        RECT 70.210000 80.335000 70.410000 80.535000 ;
        RECT 70.210000 80.740000 70.410000 80.940000 ;
        RECT 70.210000 81.145000 70.410000 81.345000 ;
        RECT 70.210000 81.550000 70.410000 81.750000 ;
        RECT 70.210000 81.955000 70.410000 82.155000 ;
        RECT 70.210000 82.360000 70.410000 82.560000 ;
        RECT 70.220000 82.855000 70.420000 83.055000 ;
        RECT 70.220000 83.265000 70.420000 83.465000 ;
        RECT 70.220000 83.675000 70.420000 83.875000 ;
        RECT 70.220000 84.085000 70.420000 84.285000 ;
        RECT 70.220000 84.495000 70.420000 84.695000 ;
        RECT 70.220000 84.905000 70.420000 85.105000 ;
        RECT 70.220000 85.315000 70.420000 85.515000 ;
        RECT 70.220000 85.725000 70.420000 85.925000 ;
        RECT 70.220000 86.135000 70.420000 86.335000 ;
        RECT 70.220000 86.545000 70.420000 86.745000 ;
        RECT 70.220000 86.955000 70.420000 87.155000 ;
        RECT 70.220000 87.365000 70.420000 87.565000 ;
        RECT 70.220000 87.775000 70.420000 87.975000 ;
        RECT 70.220000 88.185000 70.420000 88.385000 ;
        RECT 70.220000 88.595000 70.420000 88.795000 ;
        RECT 70.220000 89.005000 70.420000 89.205000 ;
        RECT 70.220000 89.415000 70.420000 89.615000 ;
        RECT 70.220000 89.825000 70.420000 90.025000 ;
        RECT 70.220000 90.235000 70.420000 90.435000 ;
        RECT 70.220000 90.645000 70.420000 90.845000 ;
        RECT 70.220000 91.055000 70.420000 91.255000 ;
        RECT 70.220000 91.465000 70.420000 91.665000 ;
        RECT 70.220000 91.875000 70.420000 92.075000 ;
        RECT 70.220000 92.285000 70.420000 92.485000 ;
        RECT 70.220000 92.695000 70.420000 92.895000 ;
        RECT 70.285000 17.860000 70.485000 18.060000 ;
        RECT 70.285000 18.290000 70.485000 18.490000 ;
        RECT 70.285000 18.720000 70.485000 18.920000 ;
        RECT 70.285000 19.150000 70.485000 19.350000 ;
        RECT 70.285000 19.580000 70.485000 19.780000 ;
        RECT 70.285000 20.010000 70.485000 20.210000 ;
        RECT 70.285000 20.440000 70.485000 20.640000 ;
        RECT 70.285000 20.870000 70.485000 21.070000 ;
        RECT 70.285000 21.300000 70.485000 21.500000 ;
        RECT 70.285000 21.730000 70.485000 21.930000 ;
        RECT 70.285000 22.160000 70.485000 22.360000 ;
        RECT 70.610000 68.125000 70.810000 68.325000 ;
        RECT 70.610000 68.535000 70.810000 68.735000 ;
        RECT 70.610000 68.945000 70.810000 69.145000 ;
        RECT 70.610000 69.355000 70.810000 69.555000 ;
        RECT 70.610000 69.765000 70.810000 69.965000 ;
        RECT 70.610000 70.175000 70.810000 70.375000 ;
        RECT 70.610000 70.585000 70.810000 70.785000 ;
        RECT 70.610000 70.995000 70.810000 71.195000 ;
        RECT 70.610000 71.405000 70.810000 71.605000 ;
        RECT 70.610000 71.815000 70.810000 72.015000 ;
        RECT 70.610000 72.225000 70.810000 72.425000 ;
        RECT 70.610000 72.635000 70.810000 72.835000 ;
        RECT 70.610000 73.045000 70.810000 73.245000 ;
        RECT 70.610000 73.450000 70.810000 73.650000 ;
        RECT 70.610000 73.855000 70.810000 74.055000 ;
        RECT 70.610000 74.260000 70.810000 74.460000 ;
        RECT 70.610000 74.665000 70.810000 74.865000 ;
        RECT 70.610000 75.070000 70.810000 75.270000 ;
        RECT 70.610000 75.475000 70.810000 75.675000 ;
        RECT 70.610000 75.880000 70.810000 76.080000 ;
        RECT 70.610000 76.285000 70.810000 76.485000 ;
        RECT 70.610000 76.690000 70.810000 76.890000 ;
        RECT 70.610000 77.095000 70.810000 77.295000 ;
        RECT 70.610000 77.500000 70.810000 77.700000 ;
        RECT 70.610000 77.905000 70.810000 78.105000 ;
        RECT 70.610000 78.310000 70.810000 78.510000 ;
        RECT 70.610000 78.715000 70.810000 78.915000 ;
        RECT 70.610000 79.120000 70.810000 79.320000 ;
        RECT 70.610000 79.525000 70.810000 79.725000 ;
        RECT 70.610000 79.930000 70.810000 80.130000 ;
        RECT 70.610000 80.335000 70.810000 80.535000 ;
        RECT 70.610000 80.740000 70.810000 80.940000 ;
        RECT 70.610000 81.145000 70.810000 81.345000 ;
        RECT 70.610000 81.550000 70.810000 81.750000 ;
        RECT 70.610000 81.955000 70.810000 82.155000 ;
        RECT 70.610000 82.360000 70.810000 82.560000 ;
        RECT 70.630000 82.855000 70.830000 83.055000 ;
        RECT 70.630000 83.265000 70.830000 83.465000 ;
        RECT 70.630000 83.675000 70.830000 83.875000 ;
        RECT 70.630000 84.085000 70.830000 84.285000 ;
        RECT 70.630000 84.495000 70.830000 84.695000 ;
        RECT 70.630000 84.905000 70.830000 85.105000 ;
        RECT 70.630000 85.315000 70.830000 85.515000 ;
        RECT 70.630000 85.725000 70.830000 85.925000 ;
        RECT 70.630000 86.135000 70.830000 86.335000 ;
        RECT 70.630000 86.545000 70.830000 86.745000 ;
        RECT 70.630000 86.955000 70.830000 87.155000 ;
        RECT 70.630000 87.365000 70.830000 87.565000 ;
        RECT 70.630000 87.775000 70.830000 87.975000 ;
        RECT 70.630000 88.185000 70.830000 88.385000 ;
        RECT 70.630000 88.595000 70.830000 88.795000 ;
        RECT 70.630000 89.005000 70.830000 89.205000 ;
        RECT 70.630000 89.415000 70.830000 89.615000 ;
        RECT 70.630000 89.825000 70.830000 90.025000 ;
        RECT 70.630000 90.235000 70.830000 90.435000 ;
        RECT 70.630000 90.645000 70.830000 90.845000 ;
        RECT 70.630000 91.055000 70.830000 91.255000 ;
        RECT 70.630000 91.465000 70.830000 91.665000 ;
        RECT 70.630000 91.875000 70.830000 92.075000 ;
        RECT 70.630000 92.285000 70.830000 92.485000 ;
        RECT 70.630000 92.695000 70.830000 92.895000 ;
        RECT 70.690000 17.860000 70.890000 18.060000 ;
        RECT 70.690000 18.290000 70.890000 18.490000 ;
        RECT 70.690000 18.720000 70.890000 18.920000 ;
        RECT 70.690000 19.150000 70.890000 19.350000 ;
        RECT 70.690000 19.580000 70.890000 19.780000 ;
        RECT 70.690000 20.010000 70.890000 20.210000 ;
        RECT 70.690000 20.440000 70.890000 20.640000 ;
        RECT 70.690000 20.870000 70.890000 21.070000 ;
        RECT 70.690000 21.300000 70.890000 21.500000 ;
        RECT 70.690000 21.730000 70.890000 21.930000 ;
        RECT 70.690000 22.160000 70.890000 22.360000 ;
        RECT 71.010000 68.125000 71.210000 68.325000 ;
        RECT 71.010000 68.535000 71.210000 68.735000 ;
        RECT 71.010000 68.945000 71.210000 69.145000 ;
        RECT 71.010000 69.355000 71.210000 69.555000 ;
        RECT 71.010000 69.765000 71.210000 69.965000 ;
        RECT 71.010000 70.175000 71.210000 70.375000 ;
        RECT 71.010000 70.585000 71.210000 70.785000 ;
        RECT 71.010000 70.995000 71.210000 71.195000 ;
        RECT 71.010000 71.405000 71.210000 71.605000 ;
        RECT 71.010000 71.815000 71.210000 72.015000 ;
        RECT 71.010000 72.225000 71.210000 72.425000 ;
        RECT 71.010000 72.635000 71.210000 72.835000 ;
        RECT 71.010000 73.045000 71.210000 73.245000 ;
        RECT 71.010000 73.450000 71.210000 73.650000 ;
        RECT 71.010000 73.855000 71.210000 74.055000 ;
        RECT 71.010000 74.260000 71.210000 74.460000 ;
        RECT 71.010000 74.665000 71.210000 74.865000 ;
        RECT 71.010000 75.070000 71.210000 75.270000 ;
        RECT 71.010000 75.475000 71.210000 75.675000 ;
        RECT 71.010000 75.880000 71.210000 76.080000 ;
        RECT 71.010000 76.285000 71.210000 76.485000 ;
        RECT 71.010000 76.690000 71.210000 76.890000 ;
        RECT 71.010000 77.095000 71.210000 77.295000 ;
        RECT 71.010000 77.500000 71.210000 77.700000 ;
        RECT 71.010000 77.905000 71.210000 78.105000 ;
        RECT 71.010000 78.310000 71.210000 78.510000 ;
        RECT 71.010000 78.715000 71.210000 78.915000 ;
        RECT 71.010000 79.120000 71.210000 79.320000 ;
        RECT 71.010000 79.525000 71.210000 79.725000 ;
        RECT 71.010000 79.930000 71.210000 80.130000 ;
        RECT 71.010000 80.335000 71.210000 80.535000 ;
        RECT 71.010000 80.740000 71.210000 80.940000 ;
        RECT 71.010000 81.145000 71.210000 81.345000 ;
        RECT 71.010000 81.550000 71.210000 81.750000 ;
        RECT 71.010000 81.955000 71.210000 82.155000 ;
        RECT 71.010000 82.360000 71.210000 82.560000 ;
        RECT 71.040000 82.855000 71.240000 83.055000 ;
        RECT 71.040000 83.265000 71.240000 83.465000 ;
        RECT 71.040000 83.675000 71.240000 83.875000 ;
        RECT 71.040000 84.085000 71.240000 84.285000 ;
        RECT 71.040000 84.495000 71.240000 84.695000 ;
        RECT 71.040000 84.905000 71.240000 85.105000 ;
        RECT 71.040000 85.315000 71.240000 85.515000 ;
        RECT 71.040000 85.725000 71.240000 85.925000 ;
        RECT 71.040000 86.135000 71.240000 86.335000 ;
        RECT 71.040000 86.545000 71.240000 86.745000 ;
        RECT 71.040000 86.955000 71.240000 87.155000 ;
        RECT 71.040000 87.365000 71.240000 87.565000 ;
        RECT 71.040000 87.775000 71.240000 87.975000 ;
        RECT 71.040000 88.185000 71.240000 88.385000 ;
        RECT 71.040000 88.595000 71.240000 88.795000 ;
        RECT 71.040000 89.005000 71.240000 89.205000 ;
        RECT 71.040000 89.415000 71.240000 89.615000 ;
        RECT 71.040000 89.825000 71.240000 90.025000 ;
        RECT 71.040000 90.235000 71.240000 90.435000 ;
        RECT 71.040000 90.645000 71.240000 90.845000 ;
        RECT 71.040000 91.055000 71.240000 91.255000 ;
        RECT 71.040000 91.465000 71.240000 91.665000 ;
        RECT 71.040000 91.875000 71.240000 92.075000 ;
        RECT 71.040000 92.285000 71.240000 92.485000 ;
        RECT 71.040000 92.695000 71.240000 92.895000 ;
        RECT 71.095000 17.860000 71.295000 18.060000 ;
        RECT 71.095000 18.290000 71.295000 18.490000 ;
        RECT 71.095000 18.720000 71.295000 18.920000 ;
        RECT 71.095000 19.150000 71.295000 19.350000 ;
        RECT 71.095000 19.580000 71.295000 19.780000 ;
        RECT 71.095000 20.010000 71.295000 20.210000 ;
        RECT 71.095000 20.440000 71.295000 20.640000 ;
        RECT 71.095000 20.870000 71.295000 21.070000 ;
        RECT 71.095000 21.300000 71.295000 21.500000 ;
        RECT 71.095000 21.730000 71.295000 21.930000 ;
        RECT 71.095000 22.160000 71.295000 22.360000 ;
        RECT 71.410000 68.125000 71.610000 68.325000 ;
        RECT 71.410000 68.535000 71.610000 68.735000 ;
        RECT 71.410000 68.945000 71.610000 69.145000 ;
        RECT 71.410000 69.355000 71.610000 69.555000 ;
        RECT 71.410000 69.765000 71.610000 69.965000 ;
        RECT 71.410000 70.175000 71.610000 70.375000 ;
        RECT 71.410000 70.585000 71.610000 70.785000 ;
        RECT 71.410000 70.995000 71.610000 71.195000 ;
        RECT 71.410000 71.405000 71.610000 71.605000 ;
        RECT 71.410000 71.815000 71.610000 72.015000 ;
        RECT 71.410000 72.225000 71.610000 72.425000 ;
        RECT 71.410000 72.635000 71.610000 72.835000 ;
        RECT 71.410000 73.045000 71.610000 73.245000 ;
        RECT 71.410000 73.450000 71.610000 73.650000 ;
        RECT 71.410000 73.855000 71.610000 74.055000 ;
        RECT 71.410000 74.260000 71.610000 74.460000 ;
        RECT 71.410000 74.665000 71.610000 74.865000 ;
        RECT 71.410000 75.070000 71.610000 75.270000 ;
        RECT 71.410000 75.475000 71.610000 75.675000 ;
        RECT 71.410000 75.880000 71.610000 76.080000 ;
        RECT 71.410000 76.285000 71.610000 76.485000 ;
        RECT 71.410000 76.690000 71.610000 76.890000 ;
        RECT 71.410000 77.095000 71.610000 77.295000 ;
        RECT 71.410000 77.500000 71.610000 77.700000 ;
        RECT 71.410000 77.905000 71.610000 78.105000 ;
        RECT 71.410000 78.310000 71.610000 78.510000 ;
        RECT 71.410000 78.715000 71.610000 78.915000 ;
        RECT 71.410000 79.120000 71.610000 79.320000 ;
        RECT 71.410000 79.525000 71.610000 79.725000 ;
        RECT 71.410000 79.930000 71.610000 80.130000 ;
        RECT 71.410000 80.335000 71.610000 80.535000 ;
        RECT 71.410000 80.740000 71.610000 80.940000 ;
        RECT 71.410000 81.145000 71.610000 81.345000 ;
        RECT 71.410000 81.550000 71.610000 81.750000 ;
        RECT 71.410000 81.955000 71.610000 82.155000 ;
        RECT 71.410000 82.360000 71.610000 82.560000 ;
        RECT 71.450000 82.855000 71.650000 83.055000 ;
        RECT 71.450000 83.265000 71.650000 83.465000 ;
        RECT 71.450000 83.675000 71.650000 83.875000 ;
        RECT 71.450000 84.085000 71.650000 84.285000 ;
        RECT 71.450000 84.495000 71.650000 84.695000 ;
        RECT 71.450000 84.905000 71.650000 85.105000 ;
        RECT 71.450000 85.315000 71.650000 85.515000 ;
        RECT 71.450000 85.725000 71.650000 85.925000 ;
        RECT 71.450000 86.135000 71.650000 86.335000 ;
        RECT 71.450000 86.545000 71.650000 86.745000 ;
        RECT 71.450000 86.955000 71.650000 87.155000 ;
        RECT 71.450000 87.365000 71.650000 87.565000 ;
        RECT 71.450000 87.775000 71.650000 87.975000 ;
        RECT 71.450000 88.185000 71.650000 88.385000 ;
        RECT 71.450000 88.595000 71.650000 88.795000 ;
        RECT 71.450000 89.005000 71.650000 89.205000 ;
        RECT 71.450000 89.415000 71.650000 89.615000 ;
        RECT 71.450000 89.825000 71.650000 90.025000 ;
        RECT 71.450000 90.235000 71.650000 90.435000 ;
        RECT 71.450000 90.645000 71.650000 90.845000 ;
        RECT 71.450000 91.055000 71.650000 91.255000 ;
        RECT 71.450000 91.465000 71.650000 91.665000 ;
        RECT 71.450000 91.875000 71.650000 92.075000 ;
        RECT 71.450000 92.285000 71.650000 92.485000 ;
        RECT 71.450000 92.695000 71.650000 92.895000 ;
        RECT 71.500000 17.860000 71.700000 18.060000 ;
        RECT 71.500000 18.290000 71.700000 18.490000 ;
        RECT 71.500000 18.720000 71.700000 18.920000 ;
        RECT 71.500000 19.150000 71.700000 19.350000 ;
        RECT 71.500000 19.580000 71.700000 19.780000 ;
        RECT 71.500000 20.010000 71.700000 20.210000 ;
        RECT 71.500000 20.440000 71.700000 20.640000 ;
        RECT 71.500000 20.870000 71.700000 21.070000 ;
        RECT 71.500000 21.300000 71.700000 21.500000 ;
        RECT 71.500000 21.730000 71.700000 21.930000 ;
        RECT 71.500000 22.160000 71.700000 22.360000 ;
        RECT 71.810000 68.125000 72.010000 68.325000 ;
        RECT 71.810000 68.535000 72.010000 68.735000 ;
        RECT 71.810000 68.945000 72.010000 69.145000 ;
        RECT 71.810000 69.355000 72.010000 69.555000 ;
        RECT 71.810000 69.765000 72.010000 69.965000 ;
        RECT 71.810000 70.175000 72.010000 70.375000 ;
        RECT 71.810000 70.585000 72.010000 70.785000 ;
        RECT 71.810000 70.995000 72.010000 71.195000 ;
        RECT 71.810000 71.405000 72.010000 71.605000 ;
        RECT 71.810000 71.815000 72.010000 72.015000 ;
        RECT 71.810000 72.225000 72.010000 72.425000 ;
        RECT 71.810000 72.635000 72.010000 72.835000 ;
        RECT 71.810000 73.045000 72.010000 73.245000 ;
        RECT 71.810000 73.450000 72.010000 73.650000 ;
        RECT 71.810000 73.855000 72.010000 74.055000 ;
        RECT 71.810000 74.260000 72.010000 74.460000 ;
        RECT 71.810000 74.665000 72.010000 74.865000 ;
        RECT 71.810000 75.070000 72.010000 75.270000 ;
        RECT 71.810000 75.475000 72.010000 75.675000 ;
        RECT 71.810000 75.880000 72.010000 76.080000 ;
        RECT 71.810000 76.285000 72.010000 76.485000 ;
        RECT 71.810000 76.690000 72.010000 76.890000 ;
        RECT 71.810000 77.095000 72.010000 77.295000 ;
        RECT 71.810000 77.500000 72.010000 77.700000 ;
        RECT 71.810000 77.905000 72.010000 78.105000 ;
        RECT 71.810000 78.310000 72.010000 78.510000 ;
        RECT 71.810000 78.715000 72.010000 78.915000 ;
        RECT 71.810000 79.120000 72.010000 79.320000 ;
        RECT 71.810000 79.525000 72.010000 79.725000 ;
        RECT 71.810000 79.930000 72.010000 80.130000 ;
        RECT 71.810000 80.335000 72.010000 80.535000 ;
        RECT 71.810000 80.740000 72.010000 80.940000 ;
        RECT 71.810000 81.145000 72.010000 81.345000 ;
        RECT 71.810000 81.550000 72.010000 81.750000 ;
        RECT 71.810000 81.955000 72.010000 82.155000 ;
        RECT 71.810000 82.360000 72.010000 82.560000 ;
        RECT 71.860000 82.855000 72.060000 83.055000 ;
        RECT 71.860000 83.265000 72.060000 83.465000 ;
        RECT 71.860000 83.675000 72.060000 83.875000 ;
        RECT 71.860000 84.085000 72.060000 84.285000 ;
        RECT 71.860000 84.495000 72.060000 84.695000 ;
        RECT 71.860000 84.905000 72.060000 85.105000 ;
        RECT 71.860000 85.315000 72.060000 85.515000 ;
        RECT 71.860000 85.725000 72.060000 85.925000 ;
        RECT 71.860000 86.135000 72.060000 86.335000 ;
        RECT 71.860000 86.545000 72.060000 86.745000 ;
        RECT 71.860000 86.955000 72.060000 87.155000 ;
        RECT 71.860000 87.365000 72.060000 87.565000 ;
        RECT 71.860000 87.775000 72.060000 87.975000 ;
        RECT 71.860000 88.185000 72.060000 88.385000 ;
        RECT 71.860000 88.595000 72.060000 88.795000 ;
        RECT 71.860000 89.005000 72.060000 89.205000 ;
        RECT 71.860000 89.415000 72.060000 89.615000 ;
        RECT 71.860000 89.825000 72.060000 90.025000 ;
        RECT 71.860000 90.235000 72.060000 90.435000 ;
        RECT 71.860000 90.645000 72.060000 90.845000 ;
        RECT 71.860000 91.055000 72.060000 91.255000 ;
        RECT 71.860000 91.465000 72.060000 91.665000 ;
        RECT 71.860000 91.875000 72.060000 92.075000 ;
        RECT 71.860000 92.285000 72.060000 92.485000 ;
        RECT 71.860000 92.695000 72.060000 92.895000 ;
        RECT 71.905000 17.860000 72.105000 18.060000 ;
        RECT 71.905000 18.290000 72.105000 18.490000 ;
        RECT 71.905000 18.720000 72.105000 18.920000 ;
        RECT 71.905000 19.150000 72.105000 19.350000 ;
        RECT 71.905000 19.580000 72.105000 19.780000 ;
        RECT 71.905000 20.010000 72.105000 20.210000 ;
        RECT 71.905000 20.440000 72.105000 20.640000 ;
        RECT 71.905000 20.870000 72.105000 21.070000 ;
        RECT 71.905000 21.300000 72.105000 21.500000 ;
        RECT 71.905000 21.730000 72.105000 21.930000 ;
        RECT 71.905000 22.160000 72.105000 22.360000 ;
        RECT 72.210000 68.125000 72.410000 68.325000 ;
        RECT 72.210000 68.535000 72.410000 68.735000 ;
        RECT 72.210000 68.945000 72.410000 69.145000 ;
        RECT 72.210000 69.355000 72.410000 69.555000 ;
        RECT 72.210000 69.765000 72.410000 69.965000 ;
        RECT 72.210000 70.175000 72.410000 70.375000 ;
        RECT 72.210000 70.585000 72.410000 70.785000 ;
        RECT 72.210000 70.995000 72.410000 71.195000 ;
        RECT 72.210000 71.405000 72.410000 71.605000 ;
        RECT 72.210000 71.815000 72.410000 72.015000 ;
        RECT 72.210000 72.225000 72.410000 72.425000 ;
        RECT 72.210000 72.635000 72.410000 72.835000 ;
        RECT 72.210000 73.045000 72.410000 73.245000 ;
        RECT 72.210000 73.450000 72.410000 73.650000 ;
        RECT 72.210000 73.855000 72.410000 74.055000 ;
        RECT 72.210000 74.260000 72.410000 74.460000 ;
        RECT 72.210000 74.665000 72.410000 74.865000 ;
        RECT 72.210000 75.070000 72.410000 75.270000 ;
        RECT 72.210000 75.475000 72.410000 75.675000 ;
        RECT 72.210000 75.880000 72.410000 76.080000 ;
        RECT 72.210000 76.285000 72.410000 76.485000 ;
        RECT 72.210000 76.690000 72.410000 76.890000 ;
        RECT 72.210000 77.095000 72.410000 77.295000 ;
        RECT 72.210000 77.500000 72.410000 77.700000 ;
        RECT 72.210000 77.905000 72.410000 78.105000 ;
        RECT 72.210000 78.310000 72.410000 78.510000 ;
        RECT 72.210000 78.715000 72.410000 78.915000 ;
        RECT 72.210000 79.120000 72.410000 79.320000 ;
        RECT 72.210000 79.525000 72.410000 79.725000 ;
        RECT 72.210000 79.930000 72.410000 80.130000 ;
        RECT 72.210000 80.335000 72.410000 80.535000 ;
        RECT 72.210000 80.740000 72.410000 80.940000 ;
        RECT 72.210000 81.145000 72.410000 81.345000 ;
        RECT 72.210000 81.550000 72.410000 81.750000 ;
        RECT 72.210000 81.955000 72.410000 82.155000 ;
        RECT 72.210000 82.360000 72.410000 82.560000 ;
        RECT 72.270000 82.855000 72.470000 83.055000 ;
        RECT 72.270000 83.265000 72.470000 83.465000 ;
        RECT 72.270000 83.675000 72.470000 83.875000 ;
        RECT 72.270000 84.085000 72.470000 84.285000 ;
        RECT 72.270000 84.495000 72.470000 84.695000 ;
        RECT 72.270000 84.905000 72.470000 85.105000 ;
        RECT 72.270000 85.315000 72.470000 85.515000 ;
        RECT 72.270000 85.725000 72.470000 85.925000 ;
        RECT 72.270000 86.135000 72.470000 86.335000 ;
        RECT 72.270000 86.545000 72.470000 86.745000 ;
        RECT 72.270000 86.955000 72.470000 87.155000 ;
        RECT 72.270000 87.365000 72.470000 87.565000 ;
        RECT 72.270000 87.775000 72.470000 87.975000 ;
        RECT 72.270000 88.185000 72.470000 88.385000 ;
        RECT 72.270000 88.595000 72.470000 88.795000 ;
        RECT 72.270000 89.005000 72.470000 89.205000 ;
        RECT 72.270000 89.415000 72.470000 89.615000 ;
        RECT 72.270000 89.825000 72.470000 90.025000 ;
        RECT 72.270000 90.235000 72.470000 90.435000 ;
        RECT 72.270000 90.645000 72.470000 90.845000 ;
        RECT 72.270000 91.055000 72.470000 91.255000 ;
        RECT 72.270000 91.465000 72.470000 91.665000 ;
        RECT 72.270000 91.875000 72.470000 92.075000 ;
        RECT 72.270000 92.285000 72.470000 92.485000 ;
        RECT 72.270000 92.695000 72.470000 92.895000 ;
        RECT 72.315000 17.860000 72.515000 18.060000 ;
        RECT 72.315000 18.290000 72.515000 18.490000 ;
        RECT 72.315000 18.720000 72.515000 18.920000 ;
        RECT 72.315000 19.150000 72.515000 19.350000 ;
        RECT 72.315000 19.580000 72.515000 19.780000 ;
        RECT 72.315000 20.010000 72.515000 20.210000 ;
        RECT 72.315000 20.440000 72.515000 20.640000 ;
        RECT 72.315000 20.870000 72.515000 21.070000 ;
        RECT 72.315000 21.300000 72.515000 21.500000 ;
        RECT 72.315000 21.730000 72.515000 21.930000 ;
        RECT 72.315000 22.160000 72.515000 22.360000 ;
        RECT 72.610000 68.125000 72.810000 68.325000 ;
        RECT 72.610000 68.535000 72.810000 68.735000 ;
        RECT 72.610000 68.945000 72.810000 69.145000 ;
        RECT 72.610000 69.355000 72.810000 69.555000 ;
        RECT 72.610000 69.765000 72.810000 69.965000 ;
        RECT 72.610000 70.175000 72.810000 70.375000 ;
        RECT 72.610000 70.585000 72.810000 70.785000 ;
        RECT 72.610000 70.995000 72.810000 71.195000 ;
        RECT 72.610000 71.405000 72.810000 71.605000 ;
        RECT 72.610000 71.815000 72.810000 72.015000 ;
        RECT 72.610000 72.225000 72.810000 72.425000 ;
        RECT 72.610000 72.635000 72.810000 72.835000 ;
        RECT 72.610000 73.045000 72.810000 73.245000 ;
        RECT 72.610000 73.450000 72.810000 73.650000 ;
        RECT 72.610000 73.855000 72.810000 74.055000 ;
        RECT 72.610000 74.260000 72.810000 74.460000 ;
        RECT 72.610000 74.665000 72.810000 74.865000 ;
        RECT 72.610000 75.070000 72.810000 75.270000 ;
        RECT 72.610000 75.475000 72.810000 75.675000 ;
        RECT 72.610000 75.880000 72.810000 76.080000 ;
        RECT 72.610000 76.285000 72.810000 76.485000 ;
        RECT 72.610000 76.690000 72.810000 76.890000 ;
        RECT 72.610000 77.095000 72.810000 77.295000 ;
        RECT 72.610000 77.500000 72.810000 77.700000 ;
        RECT 72.610000 77.905000 72.810000 78.105000 ;
        RECT 72.610000 78.310000 72.810000 78.510000 ;
        RECT 72.610000 78.715000 72.810000 78.915000 ;
        RECT 72.610000 79.120000 72.810000 79.320000 ;
        RECT 72.610000 79.525000 72.810000 79.725000 ;
        RECT 72.610000 79.930000 72.810000 80.130000 ;
        RECT 72.610000 80.335000 72.810000 80.535000 ;
        RECT 72.610000 80.740000 72.810000 80.940000 ;
        RECT 72.610000 81.145000 72.810000 81.345000 ;
        RECT 72.610000 81.550000 72.810000 81.750000 ;
        RECT 72.610000 81.955000 72.810000 82.155000 ;
        RECT 72.610000 82.360000 72.810000 82.560000 ;
        RECT 72.680000 82.855000 72.880000 83.055000 ;
        RECT 72.680000 83.265000 72.880000 83.465000 ;
        RECT 72.680000 83.675000 72.880000 83.875000 ;
        RECT 72.680000 84.085000 72.880000 84.285000 ;
        RECT 72.680000 84.495000 72.880000 84.695000 ;
        RECT 72.680000 84.905000 72.880000 85.105000 ;
        RECT 72.680000 85.315000 72.880000 85.515000 ;
        RECT 72.680000 85.725000 72.880000 85.925000 ;
        RECT 72.680000 86.135000 72.880000 86.335000 ;
        RECT 72.680000 86.545000 72.880000 86.745000 ;
        RECT 72.680000 86.955000 72.880000 87.155000 ;
        RECT 72.680000 87.365000 72.880000 87.565000 ;
        RECT 72.680000 87.775000 72.880000 87.975000 ;
        RECT 72.680000 88.185000 72.880000 88.385000 ;
        RECT 72.680000 88.595000 72.880000 88.795000 ;
        RECT 72.680000 89.005000 72.880000 89.205000 ;
        RECT 72.680000 89.415000 72.880000 89.615000 ;
        RECT 72.680000 89.825000 72.880000 90.025000 ;
        RECT 72.680000 90.235000 72.880000 90.435000 ;
        RECT 72.680000 90.645000 72.880000 90.845000 ;
        RECT 72.680000 91.055000 72.880000 91.255000 ;
        RECT 72.680000 91.465000 72.880000 91.665000 ;
        RECT 72.680000 91.875000 72.880000 92.075000 ;
        RECT 72.680000 92.285000 72.880000 92.485000 ;
        RECT 72.680000 92.695000 72.880000 92.895000 ;
        RECT 72.725000 17.860000 72.925000 18.060000 ;
        RECT 72.725000 18.290000 72.925000 18.490000 ;
        RECT 72.725000 18.720000 72.925000 18.920000 ;
        RECT 72.725000 19.150000 72.925000 19.350000 ;
        RECT 72.725000 19.580000 72.925000 19.780000 ;
        RECT 72.725000 20.010000 72.925000 20.210000 ;
        RECT 72.725000 20.440000 72.925000 20.640000 ;
        RECT 72.725000 20.870000 72.925000 21.070000 ;
        RECT 72.725000 21.300000 72.925000 21.500000 ;
        RECT 72.725000 21.730000 72.925000 21.930000 ;
        RECT 72.725000 22.160000 72.925000 22.360000 ;
        RECT 73.010000 68.125000 73.210000 68.325000 ;
        RECT 73.010000 68.535000 73.210000 68.735000 ;
        RECT 73.010000 68.945000 73.210000 69.145000 ;
        RECT 73.010000 69.355000 73.210000 69.555000 ;
        RECT 73.010000 69.765000 73.210000 69.965000 ;
        RECT 73.010000 70.175000 73.210000 70.375000 ;
        RECT 73.010000 70.585000 73.210000 70.785000 ;
        RECT 73.010000 70.995000 73.210000 71.195000 ;
        RECT 73.010000 71.405000 73.210000 71.605000 ;
        RECT 73.010000 71.815000 73.210000 72.015000 ;
        RECT 73.010000 72.225000 73.210000 72.425000 ;
        RECT 73.010000 72.635000 73.210000 72.835000 ;
        RECT 73.010000 73.045000 73.210000 73.245000 ;
        RECT 73.010000 73.450000 73.210000 73.650000 ;
        RECT 73.010000 73.855000 73.210000 74.055000 ;
        RECT 73.010000 74.260000 73.210000 74.460000 ;
        RECT 73.010000 74.665000 73.210000 74.865000 ;
        RECT 73.010000 75.070000 73.210000 75.270000 ;
        RECT 73.010000 75.475000 73.210000 75.675000 ;
        RECT 73.010000 75.880000 73.210000 76.080000 ;
        RECT 73.010000 76.285000 73.210000 76.485000 ;
        RECT 73.010000 76.690000 73.210000 76.890000 ;
        RECT 73.010000 77.095000 73.210000 77.295000 ;
        RECT 73.010000 77.500000 73.210000 77.700000 ;
        RECT 73.010000 77.905000 73.210000 78.105000 ;
        RECT 73.010000 78.310000 73.210000 78.510000 ;
        RECT 73.010000 78.715000 73.210000 78.915000 ;
        RECT 73.010000 79.120000 73.210000 79.320000 ;
        RECT 73.010000 79.525000 73.210000 79.725000 ;
        RECT 73.010000 79.930000 73.210000 80.130000 ;
        RECT 73.010000 80.335000 73.210000 80.535000 ;
        RECT 73.010000 80.740000 73.210000 80.940000 ;
        RECT 73.010000 81.145000 73.210000 81.345000 ;
        RECT 73.010000 81.550000 73.210000 81.750000 ;
        RECT 73.010000 81.955000 73.210000 82.155000 ;
        RECT 73.010000 82.360000 73.210000 82.560000 ;
        RECT 73.090000 82.855000 73.290000 83.055000 ;
        RECT 73.090000 83.265000 73.290000 83.465000 ;
        RECT 73.090000 83.675000 73.290000 83.875000 ;
        RECT 73.090000 84.085000 73.290000 84.285000 ;
        RECT 73.090000 84.495000 73.290000 84.695000 ;
        RECT 73.090000 84.905000 73.290000 85.105000 ;
        RECT 73.090000 85.315000 73.290000 85.515000 ;
        RECT 73.090000 85.725000 73.290000 85.925000 ;
        RECT 73.090000 86.135000 73.290000 86.335000 ;
        RECT 73.090000 86.545000 73.290000 86.745000 ;
        RECT 73.090000 86.955000 73.290000 87.155000 ;
        RECT 73.090000 87.365000 73.290000 87.565000 ;
        RECT 73.090000 87.775000 73.290000 87.975000 ;
        RECT 73.090000 88.185000 73.290000 88.385000 ;
        RECT 73.090000 88.595000 73.290000 88.795000 ;
        RECT 73.090000 89.005000 73.290000 89.205000 ;
        RECT 73.090000 89.415000 73.290000 89.615000 ;
        RECT 73.090000 89.825000 73.290000 90.025000 ;
        RECT 73.090000 90.235000 73.290000 90.435000 ;
        RECT 73.090000 90.645000 73.290000 90.845000 ;
        RECT 73.090000 91.055000 73.290000 91.255000 ;
        RECT 73.090000 91.465000 73.290000 91.665000 ;
        RECT 73.090000 91.875000 73.290000 92.075000 ;
        RECT 73.090000 92.285000 73.290000 92.485000 ;
        RECT 73.090000 92.695000 73.290000 92.895000 ;
        RECT 73.135000 17.860000 73.335000 18.060000 ;
        RECT 73.135000 18.290000 73.335000 18.490000 ;
        RECT 73.135000 18.720000 73.335000 18.920000 ;
        RECT 73.135000 19.150000 73.335000 19.350000 ;
        RECT 73.135000 19.580000 73.335000 19.780000 ;
        RECT 73.135000 20.010000 73.335000 20.210000 ;
        RECT 73.135000 20.440000 73.335000 20.640000 ;
        RECT 73.135000 20.870000 73.335000 21.070000 ;
        RECT 73.135000 21.300000 73.335000 21.500000 ;
        RECT 73.135000 21.730000 73.335000 21.930000 ;
        RECT 73.135000 22.160000 73.335000 22.360000 ;
        RECT 73.410000 68.125000 73.610000 68.325000 ;
        RECT 73.410000 68.535000 73.610000 68.735000 ;
        RECT 73.410000 68.945000 73.610000 69.145000 ;
        RECT 73.410000 69.355000 73.610000 69.555000 ;
        RECT 73.410000 69.765000 73.610000 69.965000 ;
        RECT 73.410000 70.175000 73.610000 70.375000 ;
        RECT 73.410000 70.585000 73.610000 70.785000 ;
        RECT 73.410000 70.995000 73.610000 71.195000 ;
        RECT 73.410000 71.405000 73.610000 71.605000 ;
        RECT 73.410000 71.815000 73.610000 72.015000 ;
        RECT 73.410000 72.225000 73.610000 72.425000 ;
        RECT 73.410000 72.635000 73.610000 72.835000 ;
        RECT 73.410000 73.045000 73.610000 73.245000 ;
        RECT 73.410000 73.450000 73.610000 73.650000 ;
        RECT 73.410000 73.855000 73.610000 74.055000 ;
        RECT 73.410000 74.260000 73.610000 74.460000 ;
        RECT 73.410000 74.665000 73.610000 74.865000 ;
        RECT 73.410000 75.070000 73.610000 75.270000 ;
        RECT 73.410000 75.475000 73.610000 75.675000 ;
        RECT 73.410000 75.880000 73.610000 76.080000 ;
        RECT 73.410000 76.285000 73.610000 76.485000 ;
        RECT 73.410000 76.690000 73.610000 76.890000 ;
        RECT 73.410000 77.095000 73.610000 77.295000 ;
        RECT 73.410000 77.500000 73.610000 77.700000 ;
        RECT 73.410000 77.905000 73.610000 78.105000 ;
        RECT 73.410000 78.310000 73.610000 78.510000 ;
        RECT 73.410000 78.715000 73.610000 78.915000 ;
        RECT 73.410000 79.120000 73.610000 79.320000 ;
        RECT 73.410000 79.525000 73.610000 79.725000 ;
        RECT 73.410000 79.930000 73.610000 80.130000 ;
        RECT 73.410000 80.335000 73.610000 80.535000 ;
        RECT 73.410000 80.740000 73.610000 80.940000 ;
        RECT 73.410000 81.145000 73.610000 81.345000 ;
        RECT 73.410000 81.550000 73.610000 81.750000 ;
        RECT 73.410000 81.955000 73.610000 82.155000 ;
        RECT 73.410000 82.360000 73.610000 82.560000 ;
        RECT 73.500000 82.855000 73.700000 83.055000 ;
        RECT 73.500000 83.265000 73.700000 83.465000 ;
        RECT 73.500000 83.675000 73.700000 83.875000 ;
        RECT 73.500000 84.085000 73.700000 84.285000 ;
        RECT 73.500000 84.495000 73.700000 84.695000 ;
        RECT 73.500000 84.905000 73.700000 85.105000 ;
        RECT 73.500000 85.315000 73.700000 85.515000 ;
        RECT 73.500000 85.725000 73.700000 85.925000 ;
        RECT 73.500000 86.135000 73.700000 86.335000 ;
        RECT 73.500000 86.545000 73.700000 86.745000 ;
        RECT 73.500000 86.955000 73.700000 87.155000 ;
        RECT 73.500000 87.365000 73.700000 87.565000 ;
        RECT 73.500000 87.775000 73.700000 87.975000 ;
        RECT 73.500000 88.185000 73.700000 88.385000 ;
        RECT 73.500000 88.595000 73.700000 88.795000 ;
        RECT 73.500000 89.005000 73.700000 89.205000 ;
        RECT 73.500000 89.415000 73.700000 89.615000 ;
        RECT 73.500000 89.825000 73.700000 90.025000 ;
        RECT 73.500000 90.235000 73.700000 90.435000 ;
        RECT 73.500000 90.645000 73.700000 90.845000 ;
        RECT 73.500000 91.055000 73.700000 91.255000 ;
        RECT 73.500000 91.465000 73.700000 91.665000 ;
        RECT 73.500000 91.875000 73.700000 92.075000 ;
        RECT 73.500000 92.285000 73.700000 92.485000 ;
        RECT 73.500000 92.695000 73.700000 92.895000 ;
        RECT 73.545000 17.860000 73.745000 18.060000 ;
        RECT 73.545000 18.290000 73.745000 18.490000 ;
        RECT 73.545000 18.720000 73.745000 18.920000 ;
        RECT 73.545000 19.150000 73.745000 19.350000 ;
        RECT 73.545000 19.580000 73.745000 19.780000 ;
        RECT 73.545000 20.010000 73.745000 20.210000 ;
        RECT 73.545000 20.440000 73.745000 20.640000 ;
        RECT 73.545000 20.870000 73.745000 21.070000 ;
        RECT 73.545000 21.300000 73.745000 21.500000 ;
        RECT 73.545000 21.730000 73.745000 21.930000 ;
        RECT 73.545000 22.160000 73.745000 22.360000 ;
        RECT 73.810000 68.125000 74.010000 68.325000 ;
        RECT 73.810000 68.535000 74.010000 68.735000 ;
        RECT 73.810000 68.945000 74.010000 69.145000 ;
        RECT 73.810000 69.355000 74.010000 69.555000 ;
        RECT 73.810000 69.765000 74.010000 69.965000 ;
        RECT 73.810000 70.175000 74.010000 70.375000 ;
        RECT 73.810000 70.585000 74.010000 70.785000 ;
        RECT 73.810000 70.995000 74.010000 71.195000 ;
        RECT 73.810000 71.405000 74.010000 71.605000 ;
        RECT 73.810000 71.815000 74.010000 72.015000 ;
        RECT 73.810000 72.225000 74.010000 72.425000 ;
        RECT 73.810000 72.635000 74.010000 72.835000 ;
        RECT 73.810000 73.045000 74.010000 73.245000 ;
        RECT 73.810000 73.450000 74.010000 73.650000 ;
        RECT 73.810000 73.855000 74.010000 74.055000 ;
        RECT 73.810000 74.260000 74.010000 74.460000 ;
        RECT 73.810000 74.665000 74.010000 74.865000 ;
        RECT 73.810000 75.070000 74.010000 75.270000 ;
        RECT 73.810000 75.475000 74.010000 75.675000 ;
        RECT 73.810000 75.880000 74.010000 76.080000 ;
        RECT 73.810000 76.285000 74.010000 76.485000 ;
        RECT 73.810000 76.690000 74.010000 76.890000 ;
        RECT 73.810000 77.095000 74.010000 77.295000 ;
        RECT 73.810000 77.500000 74.010000 77.700000 ;
        RECT 73.810000 77.905000 74.010000 78.105000 ;
        RECT 73.810000 78.310000 74.010000 78.510000 ;
        RECT 73.810000 78.715000 74.010000 78.915000 ;
        RECT 73.810000 79.120000 74.010000 79.320000 ;
        RECT 73.810000 79.525000 74.010000 79.725000 ;
        RECT 73.810000 79.930000 74.010000 80.130000 ;
        RECT 73.810000 80.335000 74.010000 80.535000 ;
        RECT 73.810000 80.740000 74.010000 80.940000 ;
        RECT 73.810000 81.145000 74.010000 81.345000 ;
        RECT 73.810000 81.550000 74.010000 81.750000 ;
        RECT 73.810000 81.955000 74.010000 82.155000 ;
        RECT 73.810000 82.360000 74.010000 82.560000 ;
        RECT 73.910000 82.855000 74.110000 83.055000 ;
        RECT 73.910000 83.265000 74.110000 83.465000 ;
        RECT 73.910000 83.675000 74.110000 83.875000 ;
        RECT 73.910000 84.085000 74.110000 84.285000 ;
        RECT 73.910000 84.495000 74.110000 84.695000 ;
        RECT 73.910000 84.905000 74.110000 85.105000 ;
        RECT 73.910000 85.315000 74.110000 85.515000 ;
        RECT 73.910000 85.725000 74.110000 85.925000 ;
        RECT 73.910000 86.135000 74.110000 86.335000 ;
        RECT 73.910000 86.545000 74.110000 86.745000 ;
        RECT 73.910000 86.955000 74.110000 87.155000 ;
        RECT 73.910000 87.365000 74.110000 87.565000 ;
        RECT 73.910000 87.775000 74.110000 87.975000 ;
        RECT 73.910000 88.185000 74.110000 88.385000 ;
        RECT 73.910000 88.595000 74.110000 88.795000 ;
        RECT 73.910000 89.005000 74.110000 89.205000 ;
        RECT 73.910000 89.415000 74.110000 89.615000 ;
        RECT 73.910000 89.825000 74.110000 90.025000 ;
        RECT 73.910000 90.235000 74.110000 90.435000 ;
        RECT 73.910000 90.645000 74.110000 90.845000 ;
        RECT 73.910000 91.055000 74.110000 91.255000 ;
        RECT 73.910000 91.465000 74.110000 91.665000 ;
        RECT 73.910000 91.875000 74.110000 92.075000 ;
        RECT 73.910000 92.285000 74.110000 92.485000 ;
        RECT 73.910000 92.695000 74.110000 92.895000 ;
        RECT 73.955000 17.860000 74.155000 18.060000 ;
        RECT 73.955000 18.290000 74.155000 18.490000 ;
        RECT 73.955000 18.720000 74.155000 18.920000 ;
        RECT 73.955000 19.150000 74.155000 19.350000 ;
        RECT 73.955000 19.580000 74.155000 19.780000 ;
        RECT 73.955000 20.010000 74.155000 20.210000 ;
        RECT 73.955000 20.440000 74.155000 20.640000 ;
        RECT 73.955000 20.870000 74.155000 21.070000 ;
        RECT 73.955000 21.300000 74.155000 21.500000 ;
        RECT 73.955000 21.730000 74.155000 21.930000 ;
        RECT 73.955000 22.160000 74.155000 22.360000 ;
        RECT 74.210000 68.125000 74.410000 68.325000 ;
        RECT 74.210000 68.535000 74.410000 68.735000 ;
        RECT 74.210000 68.945000 74.410000 69.145000 ;
        RECT 74.210000 69.355000 74.410000 69.555000 ;
        RECT 74.210000 69.765000 74.410000 69.965000 ;
        RECT 74.210000 70.175000 74.410000 70.375000 ;
        RECT 74.210000 70.585000 74.410000 70.785000 ;
        RECT 74.210000 70.995000 74.410000 71.195000 ;
        RECT 74.210000 71.405000 74.410000 71.605000 ;
        RECT 74.210000 71.815000 74.410000 72.015000 ;
        RECT 74.210000 72.225000 74.410000 72.425000 ;
        RECT 74.210000 72.635000 74.410000 72.835000 ;
        RECT 74.210000 73.045000 74.410000 73.245000 ;
        RECT 74.210000 73.450000 74.410000 73.650000 ;
        RECT 74.210000 73.855000 74.410000 74.055000 ;
        RECT 74.210000 74.260000 74.410000 74.460000 ;
        RECT 74.210000 74.665000 74.410000 74.865000 ;
        RECT 74.210000 75.070000 74.410000 75.270000 ;
        RECT 74.210000 75.475000 74.410000 75.675000 ;
        RECT 74.210000 75.880000 74.410000 76.080000 ;
        RECT 74.210000 76.285000 74.410000 76.485000 ;
        RECT 74.210000 76.690000 74.410000 76.890000 ;
        RECT 74.210000 77.095000 74.410000 77.295000 ;
        RECT 74.210000 77.500000 74.410000 77.700000 ;
        RECT 74.210000 77.905000 74.410000 78.105000 ;
        RECT 74.210000 78.310000 74.410000 78.510000 ;
        RECT 74.210000 78.715000 74.410000 78.915000 ;
        RECT 74.210000 79.120000 74.410000 79.320000 ;
        RECT 74.210000 79.525000 74.410000 79.725000 ;
        RECT 74.210000 79.930000 74.410000 80.130000 ;
        RECT 74.210000 80.335000 74.410000 80.535000 ;
        RECT 74.210000 80.740000 74.410000 80.940000 ;
        RECT 74.210000 81.145000 74.410000 81.345000 ;
        RECT 74.210000 81.550000 74.410000 81.750000 ;
        RECT 74.210000 81.955000 74.410000 82.155000 ;
        RECT 74.210000 82.360000 74.410000 82.560000 ;
        RECT 74.320000 82.855000 74.520000 83.055000 ;
        RECT 74.320000 83.265000 74.520000 83.465000 ;
        RECT 74.320000 83.675000 74.520000 83.875000 ;
        RECT 74.320000 84.085000 74.520000 84.285000 ;
        RECT 74.320000 84.495000 74.520000 84.695000 ;
        RECT 74.320000 84.905000 74.520000 85.105000 ;
        RECT 74.320000 85.315000 74.520000 85.515000 ;
        RECT 74.320000 85.725000 74.520000 85.925000 ;
        RECT 74.320000 86.135000 74.520000 86.335000 ;
        RECT 74.320000 86.545000 74.520000 86.745000 ;
        RECT 74.320000 86.955000 74.520000 87.155000 ;
        RECT 74.320000 87.365000 74.520000 87.565000 ;
        RECT 74.320000 87.775000 74.520000 87.975000 ;
        RECT 74.320000 88.185000 74.520000 88.385000 ;
        RECT 74.320000 88.595000 74.520000 88.795000 ;
        RECT 74.320000 89.005000 74.520000 89.205000 ;
        RECT 74.320000 89.415000 74.520000 89.615000 ;
        RECT 74.320000 89.825000 74.520000 90.025000 ;
        RECT 74.320000 90.235000 74.520000 90.435000 ;
        RECT 74.320000 90.645000 74.520000 90.845000 ;
        RECT 74.320000 91.055000 74.520000 91.255000 ;
        RECT 74.320000 91.465000 74.520000 91.665000 ;
        RECT 74.320000 91.875000 74.520000 92.075000 ;
        RECT 74.320000 92.285000 74.520000 92.485000 ;
        RECT 74.320000 92.695000 74.520000 92.895000 ;
        RECT 74.365000 17.860000 74.565000 18.060000 ;
        RECT 74.365000 18.290000 74.565000 18.490000 ;
        RECT 74.365000 18.720000 74.565000 18.920000 ;
        RECT 74.365000 19.150000 74.565000 19.350000 ;
        RECT 74.365000 19.580000 74.565000 19.780000 ;
        RECT 74.365000 20.010000 74.565000 20.210000 ;
        RECT 74.365000 20.440000 74.565000 20.640000 ;
        RECT 74.365000 20.870000 74.565000 21.070000 ;
        RECT 74.365000 21.300000 74.565000 21.500000 ;
        RECT 74.365000 21.730000 74.565000 21.930000 ;
        RECT 74.365000 22.160000 74.565000 22.360000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.600000 62.090000 24.500000 66.530000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000 62.090000 74.655000 66.530000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 62.085000 24.475000 66.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.780000 62.085000 75.000000 66.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 62.185000 1.270000 66.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.690000 62.160000  0.890000 62.360000 ;
        RECT  0.690000 62.570000  0.890000 62.770000 ;
        RECT  0.690000 62.980000  0.890000 63.180000 ;
        RECT  0.690000 63.390000  0.890000 63.590000 ;
        RECT  0.690000 63.800000  0.890000 64.000000 ;
        RECT  0.690000 64.210000  0.890000 64.410000 ;
        RECT  0.690000 64.620000  0.890000 64.820000 ;
        RECT  0.690000 65.030000  0.890000 65.230000 ;
        RECT  0.690000 65.440000  0.890000 65.640000 ;
        RECT  0.690000 65.850000  0.890000 66.050000 ;
        RECT  0.690000 66.260000  0.890000 66.460000 ;
        RECT  1.095000 62.160000  1.295000 62.360000 ;
        RECT  1.095000 62.570000  1.295000 62.770000 ;
        RECT  1.095000 62.980000  1.295000 63.180000 ;
        RECT  1.095000 63.390000  1.295000 63.590000 ;
        RECT  1.095000 63.800000  1.295000 64.000000 ;
        RECT  1.095000 64.210000  1.295000 64.410000 ;
        RECT  1.095000 64.620000  1.295000 64.820000 ;
        RECT  1.095000 65.030000  1.295000 65.230000 ;
        RECT  1.095000 65.440000  1.295000 65.640000 ;
        RECT  1.095000 65.850000  1.295000 66.050000 ;
        RECT  1.095000 66.260000  1.295000 66.460000 ;
        RECT  1.500000 62.160000  1.700000 62.360000 ;
        RECT  1.500000 62.570000  1.700000 62.770000 ;
        RECT  1.500000 62.980000  1.700000 63.180000 ;
        RECT  1.500000 63.390000  1.700000 63.590000 ;
        RECT  1.500000 63.800000  1.700000 64.000000 ;
        RECT  1.500000 64.210000  1.700000 64.410000 ;
        RECT  1.500000 64.620000  1.700000 64.820000 ;
        RECT  1.500000 65.030000  1.700000 65.230000 ;
        RECT  1.500000 65.440000  1.700000 65.640000 ;
        RECT  1.500000 65.850000  1.700000 66.050000 ;
        RECT  1.500000 66.260000  1.700000 66.460000 ;
        RECT  1.905000 62.160000  2.105000 62.360000 ;
        RECT  1.905000 62.570000  2.105000 62.770000 ;
        RECT  1.905000 62.980000  2.105000 63.180000 ;
        RECT  1.905000 63.390000  2.105000 63.590000 ;
        RECT  1.905000 63.800000  2.105000 64.000000 ;
        RECT  1.905000 64.210000  2.105000 64.410000 ;
        RECT  1.905000 64.620000  2.105000 64.820000 ;
        RECT  1.905000 65.030000  2.105000 65.230000 ;
        RECT  1.905000 65.440000  2.105000 65.640000 ;
        RECT  1.905000 65.850000  2.105000 66.050000 ;
        RECT  1.905000 66.260000  2.105000 66.460000 ;
        RECT  2.310000 62.160000  2.510000 62.360000 ;
        RECT  2.310000 62.570000  2.510000 62.770000 ;
        RECT  2.310000 62.980000  2.510000 63.180000 ;
        RECT  2.310000 63.390000  2.510000 63.590000 ;
        RECT  2.310000 63.800000  2.510000 64.000000 ;
        RECT  2.310000 64.210000  2.510000 64.410000 ;
        RECT  2.310000 64.620000  2.510000 64.820000 ;
        RECT  2.310000 65.030000  2.510000 65.230000 ;
        RECT  2.310000 65.440000  2.510000 65.640000 ;
        RECT  2.310000 65.850000  2.510000 66.050000 ;
        RECT  2.310000 66.260000  2.510000 66.460000 ;
        RECT  2.715000 62.160000  2.915000 62.360000 ;
        RECT  2.715000 62.570000  2.915000 62.770000 ;
        RECT  2.715000 62.980000  2.915000 63.180000 ;
        RECT  2.715000 63.390000  2.915000 63.590000 ;
        RECT  2.715000 63.800000  2.915000 64.000000 ;
        RECT  2.715000 64.210000  2.915000 64.410000 ;
        RECT  2.715000 64.620000  2.915000 64.820000 ;
        RECT  2.715000 65.030000  2.915000 65.230000 ;
        RECT  2.715000 65.440000  2.915000 65.640000 ;
        RECT  2.715000 65.850000  2.915000 66.050000 ;
        RECT  2.715000 66.260000  2.915000 66.460000 ;
        RECT  3.120000 62.160000  3.320000 62.360000 ;
        RECT  3.120000 62.570000  3.320000 62.770000 ;
        RECT  3.120000 62.980000  3.320000 63.180000 ;
        RECT  3.120000 63.390000  3.320000 63.590000 ;
        RECT  3.120000 63.800000  3.320000 64.000000 ;
        RECT  3.120000 64.210000  3.320000 64.410000 ;
        RECT  3.120000 64.620000  3.320000 64.820000 ;
        RECT  3.120000 65.030000  3.320000 65.230000 ;
        RECT  3.120000 65.440000  3.320000 65.640000 ;
        RECT  3.120000 65.850000  3.320000 66.050000 ;
        RECT  3.120000 66.260000  3.320000 66.460000 ;
        RECT  3.525000 62.160000  3.725000 62.360000 ;
        RECT  3.525000 62.570000  3.725000 62.770000 ;
        RECT  3.525000 62.980000  3.725000 63.180000 ;
        RECT  3.525000 63.390000  3.725000 63.590000 ;
        RECT  3.525000 63.800000  3.725000 64.000000 ;
        RECT  3.525000 64.210000  3.725000 64.410000 ;
        RECT  3.525000 64.620000  3.725000 64.820000 ;
        RECT  3.525000 65.030000  3.725000 65.230000 ;
        RECT  3.525000 65.440000  3.725000 65.640000 ;
        RECT  3.525000 65.850000  3.725000 66.050000 ;
        RECT  3.525000 66.260000  3.725000 66.460000 ;
        RECT  3.930000 62.160000  4.130000 62.360000 ;
        RECT  3.930000 62.570000  4.130000 62.770000 ;
        RECT  3.930000 62.980000  4.130000 63.180000 ;
        RECT  3.930000 63.390000  4.130000 63.590000 ;
        RECT  3.930000 63.800000  4.130000 64.000000 ;
        RECT  3.930000 64.210000  4.130000 64.410000 ;
        RECT  3.930000 64.620000  4.130000 64.820000 ;
        RECT  3.930000 65.030000  4.130000 65.230000 ;
        RECT  3.930000 65.440000  4.130000 65.640000 ;
        RECT  3.930000 65.850000  4.130000 66.050000 ;
        RECT  3.930000 66.260000  4.130000 66.460000 ;
        RECT  4.335000 62.160000  4.535000 62.360000 ;
        RECT  4.335000 62.570000  4.535000 62.770000 ;
        RECT  4.335000 62.980000  4.535000 63.180000 ;
        RECT  4.335000 63.390000  4.535000 63.590000 ;
        RECT  4.335000 63.800000  4.535000 64.000000 ;
        RECT  4.335000 64.210000  4.535000 64.410000 ;
        RECT  4.335000 64.620000  4.535000 64.820000 ;
        RECT  4.335000 65.030000  4.535000 65.230000 ;
        RECT  4.335000 65.440000  4.535000 65.640000 ;
        RECT  4.335000 65.850000  4.535000 66.050000 ;
        RECT  4.335000 66.260000  4.535000 66.460000 ;
        RECT  4.740000 62.160000  4.940000 62.360000 ;
        RECT  4.740000 62.570000  4.940000 62.770000 ;
        RECT  4.740000 62.980000  4.940000 63.180000 ;
        RECT  4.740000 63.390000  4.940000 63.590000 ;
        RECT  4.740000 63.800000  4.940000 64.000000 ;
        RECT  4.740000 64.210000  4.940000 64.410000 ;
        RECT  4.740000 64.620000  4.940000 64.820000 ;
        RECT  4.740000 65.030000  4.940000 65.230000 ;
        RECT  4.740000 65.440000  4.940000 65.640000 ;
        RECT  4.740000 65.850000  4.940000 66.050000 ;
        RECT  4.740000 66.260000  4.940000 66.460000 ;
        RECT  5.145000 62.160000  5.345000 62.360000 ;
        RECT  5.145000 62.570000  5.345000 62.770000 ;
        RECT  5.145000 62.980000  5.345000 63.180000 ;
        RECT  5.145000 63.390000  5.345000 63.590000 ;
        RECT  5.145000 63.800000  5.345000 64.000000 ;
        RECT  5.145000 64.210000  5.345000 64.410000 ;
        RECT  5.145000 64.620000  5.345000 64.820000 ;
        RECT  5.145000 65.030000  5.345000 65.230000 ;
        RECT  5.145000 65.440000  5.345000 65.640000 ;
        RECT  5.145000 65.850000  5.345000 66.050000 ;
        RECT  5.145000 66.260000  5.345000 66.460000 ;
        RECT  5.550000 62.160000  5.750000 62.360000 ;
        RECT  5.550000 62.570000  5.750000 62.770000 ;
        RECT  5.550000 62.980000  5.750000 63.180000 ;
        RECT  5.550000 63.390000  5.750000 63.590000 ;
        RECT  5.550000 63.800000  5.750000 64.000000 ;
        RECT  5.550000 64.210000  5.750000 64.410000 ;
        RECT  5.550000 64.620000  5.750000 64.820000 ;
        RECT  5.550000 65.030000  5.750000 65.230000 ;
        RECT  5.550000 65.440000  5.750000 65.640000 ;
        RECT  5.550000 65.850000  5.750000 66.050000 ;
        RECT  5.550000 66.260000  5.750000 66.460000 ;
        RECT  5.955000 62.160000  6.155000 62.360000 ;
        RECT  5.955000 62.570000  6.155000 62.770000 ;
        RECT  5.955000 62.980000  6.155000 63.180000 ;
        RECT  5.955000 63.390000  6.155000 63.590000 ;
        RECT  5.955000 63.800000  6.155000 64.000000 ;
        RECT  5.955000 64.210000  6.155000 64.410000 ;
        RECT  5.955000 64.620000  6.155000 64.820000 ;
        RECT  5.955000 65.030000  6.155000 65.230000 ;
        RECT  5.955000 65.440000  6.155000 65.640000 ;
        RECT  5.955000 65.850000  6.155000 66.050000 ;
        RECT  5.955000 66.260000  6.155000 66.460000 ;
        RECT  6.360000 62.160000  6.560000 62.360000 ;
        RECT  6.360000 62.570000  6.560000 62.770000 ;
        RECT  6.360000 62.980000  6.560000 63.180000 ;
        RECT  6.360000 63.390000  6.560000 63.590000 ;
        RECT  6.360000 63.800000  6.560000 64.000000 ;
        RECT  6.360000 64.210000  6.560000 64.410000 ;
        RECT  6.360000 64.620000  6.560000 64.820000 ;
        RECT  6.360000 65.030000  6.560000 65.230000 ;
        RECT  6.360000 65.440000  6.560000 65.640000 ;
        RECT  6.360000 65.850000  6.560000 66.050000 ;
        RECT  6.360000 66.260000  6.560000 66.460000 ;
        RECT  6.765000 62.160000  6.965000 62.360000 ;
        RECT  6.765000 62.570000  6.965000 62.770000 ;
        RECT  6.765000 62.980000  6.965000 63.180000 ;
        RECT  6.765000 63.390000  6.965000 63.590000 ;
        RECT  6.765000 63.800000  6.965000 64.000000 ;
        RECT  6.765000 64.210000  6.965000 64.410000 ;
        RECT  6.765000 64.620000  6.965000 64.820000 ;
        RECT  6.765000 65.030000  6.965000 65.230000 ;
        RECT  6.765000 65.440000  6.965000 65.640000 ;
        RECT  6.765000 65.850000  6.965000 66.050000 ;
        RECT  6.765000 66.260000  6.965000 66.460000 ;
        RECT  7.170000 62.160000  7.370000 62.360000 ;
        RECT  7.170000 62.570000  7.370000 62.770000 ;
        RECT  7.170000 62.980000  7.370000 63.180000 ;
        RECT  7.170000 63.390000  7.370000 63.590000 ;
        RECT  7.170000 63.800000  7.370000 64.000000 ;
        RECT  7.170000 64.210000  7.370000 64.410000 ;
        RECT  7.170000 64.620000  7.370000 64.820000 ;
        RECT  7.170000 65.030000  7.370000 65.230000 ;
        RECT  7.170000 65.440000  7.370000 65.640000 ;
        RECT  7.170000 65.850000  7.370000 66.050000 ;
        RECT  7.170000 66.260000  7.370000 66.460000 ;
        RECT  7.575000 62.160000  7.775000 62.360000 ;
        RECT  7.575000 62.570000  7.775000 62.770000 ;
        RECT  7.575000 62.980000  7.775000 63.180000 ;
        RECT  7.575000 63.390000  7.775000 63.590000 ;
        RECT  7.575000 63.800000  7.775000 64.000000 ;
        RECT  7.575000 64.210000  7.775000 64.410000 ;
        RECT  7.575000 64.620000  7.775000 64.820000 ;
        RECT  7.575000 65.030000  7.775000 65.230000 ;
        RECT  7.575000 65.440000  7.775000 65.640000 ;
        RECT  7.575000 65.850000  7.775000 66.050000 ;
        RECT  7.575000 66.260000  7.775000 66.460000 ;
        RECT  7.980000 62.160000  8.180000 62.360000 ;
        RECT  7.980000 62.570000  8.180000 62.770000 ;
        RECT  7.980000 62.980000  8.180000 63.180000 ;
        RECT  7.980000 63.390000  8.180000 63.590000 ;
        RECT  7.980000 63.800000  8.180000 64.000000 ;
        RECT  7.980000 64.210000  8.180000 64.410000 ;
        RECT  7.980000 64.620000  8.180000 64.820000 ;
        RECT  7.980000 65.030000  8.180000 65.230000 ;
        RECT  7.980000 65.440000  8.180000 65.640000 ;
        RECT  7.980000 65.850000  8.180000 66.050000 ;
        RECT  7.980000 66.260000  8.180000 66.460000 ;
        RECT  8.385000 62.160000  8.585000 62.360000 ;
        RECT  8.385000 62.570000  8.585000 62.770000 ;
        RECT  8.385000 62.980000  8.585000 63.180000 ;
        RECT  8.385000 63.390000  8.585000 63.590000 ;
        RECT  8.385000 63.800000  8.585000 64.000000 ;
        RECT  8.385000 64.210000  8.585000 64.410000 ;
        RECT  8.385000 64.620000  8.585000 64.820000 ;
        RECT  8.385000 65.030000  8.585000 65.230000 ;
        RECT  8.385000 65.440000  8.585000 65.640000 ;
        RECT  8.385000 65.850000  8.585000 66.050000 ;
        RECT  8.385000 66.260000  8.585000 66.460000 ;
        RECT  8.790000 62.160000  8.990000 62.360000 ;
        RECT  8.790000 62.570000  8.990000 62.770000 ;
        RECT  8.790000 62.980000  8.990000 63.180000 ;
        RECT  8.790000 63.390000  8.990000 63.590000 ;
        RECT  8.790000 63.800000  8.990000 64.000000 ;
        RECT  8.790000 64.210000  8.990000 64.410000 ;
        RECT  8.790000 64.620000  8.990000 64.820000 ;
        RECT  8.790000 65.030000  8.990000 65.230000 ;
        RECT  8.790000 65.440000  8.990000 65.640000 ;
        RECT  8.790000 65.850000  8.990000 66.050000 ;
        RECT  8.790000 66.260000  8.990000 66.460000 ;
        RECT  9.195000 62.160000  9.395000 62.360000 ;
        RECT  9.195000 62.570000  9.395000 62.770000 ;
        RECT  9.195000 62.980000  9.395000 63.180000 ;
        RECT  9.195000 63.390000  9.395000 63.590000 ;
        RECT  9.195000 63.800000  9.395000 64.000000 ;
        RECT  9.195000 64.210000  9.395000 64.410000 ;
        RECT  9.195000 64.620000  9.395000 64.820000 ;
        RECT  9.195000 65.030000  9.395000 65.230000 ;
        RECT  9.195000 65.440000  9.395000 65.640000 ;
        RECT  9.195000 65.850000  9.395000 66.050000 ;
        RECT  9.195000 66.260000  9.395000 66.460000 ;
        RECT  9.600000 62.160000  9.800000 62.360000 ;
        RECT  9.600000 62.570000  9.800000 62.770000 ;
        RECT  9.600000 62.980000  9.800000 63.180000 ;
        RECT  9.600000 63.390000  9.800000 63.590000 ;
        RECT  9.600000 63.800000  9.800000 64.000000 ;
        RECT  9.600000 64.210000  9.800000 64.410000 ;
        RECT  9.600000 64.620000  9.800000 64.820000 ;
        RECT  9.600000 65.030000  9.800000 65.230000 ;
        RECT  9.600000 65.440000  9.800000 65.640000 ;
        RECT  9.600000 65.850000  9.800000 66.050000 ;
        RECT  9.600000 66.260000  9.800000 66.460000 ;
        RECT 10.005000 62.160000 10.205000 62.360000 ;
        RECT 10.005000 62.570000 10.205000 62.770000 ;
        RECT 10.005000 62.980000 10.205000 63.180000 ;
        RECT 10.005000 63.390000 10.205000 63.590000 ;
        RECT 10.005000 63.800000 10.205000 64.000000 ;
        RECT 10.005000 64.210000 10.205000 64.410000 ;
        RECT 10.005000 64.620000 10.205000 64.820000 ;
        RECT 10.005000 65.030000 10.205000 65.230000 ;
        RECT 10.005000 65.440000 10.205000 65.640000 ;
        RECT 10.005000 65.850000 10.205000 66.050000 ;
        RECT 10.005000 66.260000 10.205000 66.460000 ;
        RECT 10.410000 62.160000 10.610000 62.360000 ;
        RECT 10.410000 62.570000 10.610000 62.770000 ;
        RECT 10.410000 62.980000 10.610000 63.180000 ;
        RECT 10.410000 63.390000 10.610000 63.590000 ;
        RECT 10.410000 63.800000 10.610000 64.000000 ;
        RECT 10.410000 64.210000 10.610000 64.410000 ;
        RECT 10.410000 64.620000 10.610000 64.820000 ;
        RECT 10.410000 65.030000 10.610000 65.230000 ;
        RECT 10.410000 65.440000 10.610000 65.640000 ;
        RECT 10.410000 65.850000 10.610000 66.050000 ;
        RECT 10.410000 66.260000 10.610000 66.460000 ;
        RECT 10.815000 62.160000 11.015000 62.360000 ;
        RECT 10.815000 62.570000 11.015000 62.770000 ;
        RECT 10.815000 62.980000 11.015000 63.180000 ;
        RECT 10.815000 63.390000 11.015000 63.590000 ;
        RECT 10.815000 63.800000 11.015000 64.000000 ;
        RECT 10.815000 64.210000 11.015000 64.410000 ;
        RECT 10.815000 64.620000 11.015000 64.820000 ;
        RECT 10.815000 65.030000 11.015000 65.230000 ;
        RECT 10.815000 65.440000 11.015000 65.640000 ;
        RECT 10.815000 65.850000 11.015000 66.050000 ;
        RECT 10.815000 66.260000 11.015000 66.460000 ;
        RECT 11.220000 62.160000 11.420000 62.360000 ;
        RECT 11.220000 62.570000 11.420000 62.770000 ;
        RECT 11.220000 62.980000 11.420000 63.180000 ;
        RECT 11.220000 63.390000 11.420000 63.590000 ;
        RECT 11.220000 63.800000 11.420000 64.000000 ;
        RECT 11.220000 64.210000 11.420000 64.410000 ;
        RECT 11.220000 64.620000 11.420000 64.820000 ;
        RECT 11.220000 65.030000 11.420000 65.230000 ;
        RECT 11.220000 65.440000 11.420000 65.640000 ;
        RECT 11.220000 65.850000 11.420000 66.050000 ;
        RECT 11.220000 66.260000 11.420000 66.460000 ;
        RECT 11.625000 62.160000 11.825000 62.360000 ;
        RECT 11.625000 62.570000 11.825000 62.770000 ;
        RECT 11.625000 62.980000 11.825000 63.180000 ;
        RECT 11.625000 63.390000 11.825000 63.590000 ;
        RECT 11.625000 63.800000 11.825000 64.000000 ;
        RECT 11.625000 64.210000 11.825000 64.410000 ;
        RECT 11.625000 64.620000 11.825000 64.820000 ;
        RECT 11.625000 65.030000 11.825000 65.230000 ;
        RECT 11.625000 65.440000 11.825000 65.640000 ;
        RECT 11.625000 65.850000 11.825000 66.050000 ;
        RECT 11.625000 66.260000 11.825000 66.460000 ;
        RECT 12.030000 62.160000 12.230000 62.360000 ;
        RECT 12.030000 62.570000 12.230000 62.770000 ;
        RECT 12.030000 62.980000 12.230000 63.180000 ;
        RECT 12.030000 63.390000 12.230000 63.590000 ;
        RECT 12.030000 63.800000 12.230000 64.000000 ;
        RECT 12.030000 64.210000 12.230000 64.410000 ;
        RECT 12.030000 64.620000 12.230000 64.820000 ;
        RECT 12.030000 65.030000 12.230000 65.230000 ;
        RECT 12.030000 65.440000 12.230000 65.640000 ;
        RECT 12.030000 65.850000 12.230000 66.050000 ;
        RECT 12.030000 66.260000 12.230000 66.460000 ;
        RECT 12.435000 62.160000 12.635000 62.360000 ;
        RECT 12.435000 62.570000 12.635000 62.770000 ;
        RECT 12.435000 62.980000 12.635000 63.180000 ;
        RECT 12.435000 63.390000 12.635000 63.590000 ;
        RECT 12.435000 63.800000 12.635000 64.000000 ;
        RECT 12.435000 64.210000 12.635000 64.410000 ;
        RECT 12.435000 64.620000 12.635000 64.820000 ;
        RECT 12.435000 65.030000 12.635000 65.230000 ;
        RECT 12.435000 65.440000 12.635000 65.640000 ;
        RECT 12.435000 65.850000 12.635000 66.050000 ;
        RECT 12.435000 66.260000 12.635000 66.460000 ;
        RECT 12.840000 62.160000 13.040000 62.360000 ;
        RECT 12.840000 62.570000 13.040000 62.770000 ;
        RECT 12.840000 62.980000 13.040000 63.180000 ;
        RECT 12.840000 63.390000 13.040000 63.590000 ;
        RECT 12.840000 63.800000 13.040000 64.000000 ;
        RECT 12.840000 64.210000 13.040000 64.410000 ;
        RECT 12.840000 64.620000 13.040000 64.820000 ;
        RECT 12.840000 65.030000 13.040000 65.230000 ;
        RECT 12.840000 65.440000 13.040000 65.640000 ;
        RECT 12.840000 65.850000 13.040000 66.050000 ;
        RECT 12.840000 66.260000 13.040000 66.460000 ;
        RECT 13.245000 62.160000 13.445000 62.360000 ;
        RECT 13.245000 62.570000 13.445000 62.770000 ;
        RECT 13.245000 62.980000 13.445000 63.180000 ;
        RECT 13.245000 63.390000 13.445000 63.590000 ;
        RECT 13.245000 63.800000 13.445000 64.000000 ;
        RECT 13.245000 64.210000 13.445000 64.410000 ;
        RECT 13.245000 64.620000 13.445000 64.820000 ;
        RECT 13.245000 65.030000 13.445000 65.230000 ;
        RECT 13.245000 65.440000 13.445000 65.640000 ;
        RECT 13.245000 65.850000 13.445000 66.050000 ;
        RECT 13.245000 66.260000 13.445000 66.460000 ;
        RECT 13.650000 62.160000 13.850000 62.360000 ;
        RECT 13.650000 62.570000 13.850000 62.770000 ;
        RECT 13.650000 62.980000 13.850000 63.180000 ;
        RECT 13.650000 63.390000 13.850000 63.590000 ;
        RECT 13.650000 63.800000 13.850000 64.000000 ;
        RECT 13.650000 64.210000 13.850000 64.410000 ;
        RECT 13.650000 64.620000 13.850000 64.820000 ;
        RECT 13.650000 65.030000 13.850000 65.230000 ;
        RECT 13.650000 65.440000 13.850000 65.640000 ;
        RECT 13.650000 65.850000 13.850000 66.050000 ;
        RECT 13.650000 66.260000 13.850000 66.460000 ;
        RECT 14.055000 62.160000 14.255000 62.360000 ;
        RECT 14.055000 62.570000 14.255000 62.770000 ;
        RECT 14.055000 62.980000 14.255000 63.180000 ;
        RECT 14.055000 63.390000 14.255000 63.590000 ;
        RECT 14.055000 63.800000 14.255000 64.000000 ;
        RECT 14.055000 64.210000 14.255000 64.410000 ;
        RECT 14.055000 64.620000 14.255000 64.820000 ;
        RECT 14.055000 65.030000 14.255000 65.230000 ;
        RECT 14.055000 65.440000 14.255000 65.640000 ;
        RECT 14.055000 65.850000 14.255000 66.050000 ;
        RECT 14.055000 66.260000 14.255000 66.460000 ;
        RECT 14.460000 62.160000 14.660000 62.360000 ;
        RECT 14.460000 62.570000 14.660000 62.770000 ;
        RECT 14.460000 62.980000 14.660000 63.180000 ;
        RECT 14.460000 63.390000 14.660000 63.590000 ;
        RECT 14.460000 63.800000 14.660000 64.000000 ;
        RECT 14.460000 64.210000 14.660000 64.410000 ;
        RECT 14.460000 64.620000 14.660000 64.820000 ;
        RECT 14.460000 65.030000 14.660000 65.230000 ;
        RECT 14.460000 65.440000 14.660000 65.640000 ;
        RECT 14.460000 65.850000 14.660000 66.050000 ;
        RECT 14.460000 66.260000 14.660000 66.460000 ;
        RECT 14.865000 62.160000 15.065000 62.360000 ;
        RECT 14.865000 62.570000 15.065000 62.770000 ;
        RECT 14.865000 62.980000 15.065000 63.180000 ;
        RECT 14.865000 63.390000 15.065000 63.590000 ;
        RECT 14.865000 63.800000 15.065000 64.000000 ;
        RECT 14.865000 64.210000 15.065000 64.410000 ;
        RECT 14.865000 64.620000 15.065000 64.820000 ;
        RECT 14.865000 65.030000 15.065000 65.230000 ;
        RECT 14.865000 65.440000 15.065000 65.640000 ;
        RECT 14.865000 65.850000 15.065000 66.050000 ;
        RECT 14.865000 66.260000 15.065000 66.460000 ;
        RECT 15.270000 62.160000 15.470000 62.360000 ;
        RECT 15.270000 62.570000 15.470000 62.770000 ;
        RECT 15.270000 62.980000 15.470000 63.180000 ;
        RECT 15.270000 63.390000 15.470000 63.590000 ;
        RECT 15.270000 63.800000 15.470000 64.000000 ;
        RECT 15.270000 64.210000 15.470000 64.410000 ;
        RECT 15.270000 64.620000 15.470000 64.820000 ;
        RECT 15.270000 65.030000 15.470000 65.230000 ;
        RECT 15.270000 65.440000 15.470000 65.640000 ;
        RECT 15.270000 65.850000 15.470000 66.050000 ;
        RECT 15.270000 66.260000 15.470000 66.460000 ;
        RECT 15.675000 62.160000 15.875000 62.360000 ;
        RECT 15.675000 62.570000 15.875000 62.770000 ;
        RECT 15.675000 62.980000 15.875000 63.180000 ;
        RECT 15.675000 63.390000 15.875000 63.590000 ;
        RECT 15.675000 63.800000 15.875000 64.000000 ;
        RECT 15.675000 64.210000 15.875000 64.410000 ;
        RECT 15.675000 64.620000 15.875000 64.820000 ;
        RECT 15.675000 65.030000 15.875000 65.230000 ;
        RECT 15.675000 65.440000 15.875000 65.640000 ;
        RECT 15.675000 65.850000 15.875000 66.050000 ;
        RECT 15.675000 66.260000 15.875000 66.460000 ;
        RECT 16.080000 62.160000 16.280000 62.360000 ;
        RECT 16.080000 62.570000 16.280000 62.770000 ;
        RECT 16.080000 62.980000 16.280000 63.180000 ;
        RECT 16.080000 63.390000 16.280000 63.590000 ;
        RECT 16.080000 63.800000 16.280000 64.000000 ;
        RECT 16.080000 64.210000 16.280000 64.410000 ;
        RECT 16.080000 64.620000 16.280000 64.820000 ;
        RECT 16.080000 65.030000 16.280000 65.230000 ;
        RECT 16.080000 65.440000 16.280000 65.640000 ;
        RECT 16.080000 65.850000 16.280000 66.050000 ;
        RECT 16.080000 66.260000 16.280000 66.460000 ;
        RECT 16.485000 62.160000 16.685000 62.360000 ;
        RECT 16.485000 62.570000 16.685000 62.770000 ;
        RECT 16.485000 62.980000 16.685000 63.180000 ;
        RECT 16.485000 63.390000 16.685000 63.590000 ;
        RECT 16.485000 63.800000 16.685000 64.000000 ;
        RECT 16.485000 64.210000 16.685000 64.410000 ;
        RECT 16.485000 64.620000 16.685000 64.820000 ;
        RECT 16.485000 65.030000 16.685000 65.230000 ;
        RECT 16.485000 65.440000 16.685000 65.640000 ;
        RECT 16.485000 65.850000 16.685000 66.050000 ;
        RECT 16.485000 66.260000 16.685000 66.460000 ;
        RECT 16.890000 62.160000 17.090000 62.360000 ;
        RECT 16.890000 62.570000 17.090000 62.770000 ;
        RECT 16.890000 62.980000 17.090000 63.180000 ;
        RECT 16.890000 63.390000 17.090000 63.590000 ;
        RECT 16.890000 63.800000 17.090000 64.000000 ;
        RECT 16.890000 64.210000 17.090000 64.410000 ;
        RECT 16.890000 64.620000 17.090000 64.820000 ;
        RECT 16.890000 65.030000 17.090000 65.230000 ;
        RECT 16.890000 65.440000 17.090000 65.640000 ;
        RECT 16.890000 65.850000 17.090000 66.050000 ;
        RECT 16.890000 66.260000 17.090000 66.460000 ;
        RECT 17.295000 62.160000 17.495000 62.360000 ;
        RECT 17.295000 62.570000 17.495000 62.770000 ;
        RECT 17.295000 62.980000 17.495000 63.180000 ;
        RECT 17.295000 63.390000 17.495000 63.590000 ;
        RECT 17.295000 63.800000 17.495000 64.000000 ;
        RECT 17.295000 64.210000 17.495000 64.410000 ;
        RECT 17.295000 64.620000 17.495000 64.820000 ;
        RECT 17.295000 65.030000 17.495000 65.230000 ;
        RECT 17.295000 65.440000 17.495000 65.640000 ;
        RECT 17.295000 65.850000 17.495000 66.050000 ;
        RECT 17.295000 66.260000 17.495000 66.460000 ;
        RECT 17.700000 62.160000 17.900000 62.360000 ;
        RECT 17.700000 62.570000 17.900000 62.770000 ;
        RECT 17.700000 62.980000 17.900000 63.180000 ;
        RECT 17.700000 63.390000 17.900000 63.590000 ;
        RECT 17.700000 63.800000 17.900000 64.000000 ;
        RECT 17.700000 64.210000 17.900000 64.410000 ;
        RECT 17.700000 64.620000 17.900000 64.820000 ;
        RECT 17.700000 65.030000 17.900000 65.230000 ;
        RECT 17.700000 65.440000 17.900000 65.640000 ;
        RECT 17.700000 65.850000 17.900000 66.050000 ;
        RECT 17.700000 66.260000 17.900000 66.460000 ;
        RECT 18.105000 62.160000 18.305000 62.360000 ;
        RECT 18.105000 62.570000 18.305000 62.770000 ;
        RECT 18.105000 62.980000 18.305000 63.180000 ;
        RECT 18.105000 63.390000 18.305000 63.590000 ;
        RECT 18.105000 63.800000 18.305000 64.000000 ;
        RECT 18.105000 64.210000 18.305000 64.410000 ;
        RECT 18.105000 64.620000 18.305000 64.820000 ;
        RECT 18.105000 65.030000 18.305000 65.230000 ;
        RECT 18.105000 65.440000 18.305000 65.640000 ;
        RECT 18.105000 65.850000 18.305000 66.050000 ;
        RECT 18.105000 66.260000 18.305000 66.460000 ;
        RECT 18.510000 62.160000 18.710000 62.360000 ;
        RECT 18.510000 62.570000 18.710000 62.770000 ;
        RECT 18.510000 62.980000 18.710000 63.180000 ;
        RECT 18.510000 63.390000 18.710000 63.590000 ;
        RECT 18.510000 63.800000 18.710000 64.000000 ;
        RECT 18.510000 64.210000 18.710000 64.410000 ;
        RECT 18.510000 64.620000 18.710000 64.820000 ;
        RECT 18.510000 65.030000 18.710000 65.230000 ;
        RECT 18.510000 65.440000 18.710000 65.640000 ;
        RECT 18.510000 65.850000 18.710000 66.050000 ;
        RECT 18.510000 66.260000 18.710000 66.460000 ;
        RECT 18.915000 62.160000 19.115000 62.360000 ;
        RECT 18.915000 62.570000 19.115000 62.770000 ;
        RECT 18.915000 62.980000 19.115000 63.180000 ;
        RECT 18.915000 63.390000 19.115000 63.590000 ;
        RECT 18.915000 63.800000 19.115000 64.000000 ;
        RECT 18.915000 64.210000 19.115000 64.410000 ;
        RECT 18.915000 64.620000 19.115000 64.820000 ;
        RECT 18.915000 65.030000 19.115000 65.230000 ;
        RECT 18.915000 65.440000 19.115000 65.640000 ;
        RECT 18.915000 65.850000 19.115000 66.050000 ;
        RECT 18.915000 66.260000 19.115000 66.460000 ;
        RECT 19.320000 62.160000 19.520000 62.360000 ;
        RECT 19.320000 62.570000 19.520000 62.770000 ;
        RECT 19.320000 62.980000 19.520000 63.180000 ;
        RECT 19.320000 63.390000 19.520000 63.590000 ;
        RECT 19.320000 63.800000 19.520000 64.000000 ;
        RECT 19.320000 64.210000 19.520000 64.410000 ;
        RECT 19.320000 64.620000 19.520000 64.820000 ;
        RECT 19.320000 65.030000 19.520000 65.230000 ;
        RECT 19.320000 65.440000 19.520000 65.640000 ;
        RECT 19.320000 65.850000 19.520000 66.050000 ;
        RECT 19.320000 66.260000 19.520000 66.460000 ;
        RECT 19.725000 62.160000 19.925000 62.360000 ;
        RECT 19.725000 62.570000 19.925000 62.770000 ;
        RECT 19.725000 62.980000 19.925000 63.180000 ;
        RECT 19.725000 63.390000 19.925000 63.590000 ;
        RECT 19.725000 63.800000 19.925000 64.000000 ;
        RECT 19.725000 64.210000 19.925000 64.410000 ;
        RECT 19.725000 64.620000 19.925000 64.820000 ;
        RECT 19.725000 65.030000 19.925000 65.230000 ;
        RECT 19.725000 65.440000 19.925000 65.640000 ;
        RECT 19.725000 65.850000 19.925000 66.050000 ;
        RECT 19.725000 66.260000 19.925000 66.460000 ;
        RECT 20.130000 62.160000 20.330000 62.360000 ;
        RECT 20.130000 62.570000 20.330000 62.770000 ;
        RECT 20.130000 62.980000 20.330000 63.180000 ;
        RECT 20.130000 63.390000 20.330000 63.590000 ;
        RECT 20.130000 63.800000 20.330000 64.000000 ;
        RECT 20.130000 64.210000 20.330000 64.410000 ;
        RECT 20.130000 64.620000 20.330000 64.820000 ;
        RECT 20.130000 65.030000 20.330000 65.230000 ;
        RECT 20.130000 65.440000 20.330000 65.640000 ;
        RECT 20.130000 65.850000 20.330000 66.050000 ;
        RECT 20.130000 66.260000 20.330000 66.460000 ;
        RECT 20.535000 62.160000 20.735000 62.360000 ;
        RECT 20.535000 62.570000 20.735000 62.770000 ;
        RECT 20.535000 62.980000 20.735000 63.180000 ;
        RECT 20.535000 63.390000 20.735000 63.590000 ;
        RECT 20.535000 63.800000 20.735000 64.000000 ;
        RECT 20.535000 64.210000 20.735000 64.410000 ;
        RECT 20.535000 64.620000 20.735000 64.820000 ;
        RECT 20.535000 65.030000 20.735000 65.230000 ;
        RECT 20.535000 65.440000 20.735000 65.640000 ;
        RECT 20.535000 65.850000 20.735000 66.050000 ;
        RECT 20.535000 66.260000 20.735000 66.460000 ;
        RECT 20.940000 62.160000 21.140000 62.360000 ;
        RECT 20.940000 62.570000 21.140000 62.770000 ;
        RECT 20.940000 62.980000 21.140000 63.180000 ;
        RECT 20.940000 63.390000 21.140000 63.590000 ;
        RECT 20.940000 63.800000 21.140000 64.000000 ;
        RECT 20.940000 64.210000 21.140000 64.410000 ;
        RECT 20.940000 64.620000 21.140000 64.820000 ;
        RECT 20.940000 65.030000 21.140000 65.230000 ;
        RECT 20.940000 65.440000 21.140000 65.640000 ;
        RECT 20.940000 65.850000 21.140000 66.050000 ;
        RECT 20.940000 66.260000 21.140000 66.460000 ;
        RECT 21.345000 62.160000 21.545000 62.360000 ;
        RECT 21.345000 62.570000 21.545000 62.770000 ;
        RECT 21.345000 62.980000 21.545000 63.180000 ;
        RECT 21.345000 63.390000 21.545000 63.590000 ;
        RECT 21.345000 63.800000 21.545000 64.000000 ;
        RECT 21.345000 64.210000 21.545000 64.410000 ;
        RECT 21.345000 64.620000 21.545000 64.820000 ;
        RECT 21.345000 65.030000 21.545000 65.230000 ;
        RECT 21.345000 65.440000 21.545000 65.640000 ;
        RECT 21.345000 65.850000 21.545000 66.050000 ;
        RECT 21.345000 66.260000 21.545000 66.460000 ;
        RECT 21.750000 62.160000 21.950000 62.360000 ;
        RECT 21.750000 62.570000 21.950000 62.770000 ;
        RECT 21.750000 62.980000 21.950000 63.180000 ;
        RECT 21.750000 63.390000 21.950000 63.590000 ;
        RECT 21.750000 63.800000 21.950000 64.000000 ;
        RECT 21.750000 64.210000 21.950000 64.410000 ;
        RECT 21.750000 64.620000 21.950000 64.820000 ;
        RECT 21.750000 65.030000 21.950000 65.230000 ;
        RECT 21.750000 65.440000 21.950000 65.640000 ;
        RECT 21.750000 65.850000 21.950000 66.050000 ;
        RECT 21.750000 66.260000 21.950000 66.460000 ;
        RECT 22.160000 62.160000 22.360000 62.360000 ;
        RECT 22.160000 62.570000 22.360000 62.770000 ;
        RECT 22.160000 62.980000 22.360000 63.180000 ;
        RECT 22.160000 63.390000 22.360000 63.590000 ;
        RECT 22.160000 63.800000 22.360000 64.000000 ;
        RECT 22.160000 64.210000 22.360000 64.410000 ;
        RECT 22.160000 64.620000 22.360000 64.820000 ;
        RECT 22.160000 65.030000 22.360000 65.230000 ;
        RECT 22.160000 65.440000 22.360000 65.640000 ;
        RECT 22.160000 65.850000 22.360000 66.050000 ;
        RECT 22.160000 66.260000 22.360000 66.460000 ;
        RECT 22.570000 62.160000 22.770000 62.360000 ;
        RECT 22.570000 62.570000 22.770000 62.770000 ;
        RECT 22.570000 62.980000 22.770000 63.180000 ;
        RECT 22.570000 63.390000 22.770000 63.590000 ;
        RECT 22.570000 63.800000 22.770000 64.000000 ;
        RECT 22.570000 64.210000 22.770000 64.410000 ;
        RECT 22.570000 64.620000 22.770000 64.820000 ;
        RECT 22.570000 65.030000 22.770000 65.230000 ;
        RECT 22.570000 65.440000 22.770000 65.640000 ;
        RECT 22.570000 65.850000 22.770000 66.050000 ;
        RECT 22.570000 66.260000 22.770000 66.460000 ;
        RECT 22.980000 62.160000 23.180000 62.360000 ;
        RECT 22.980000 62.570000 23.180000 62.770000 ;
        RECT 22.980000 62.980000 23.180000 63.180000 ;
        RECT 22.980000 63.390000 23.180000 63.590000 ;
        RECT 22.980000 63.800000 23.180000 64.000000 ;
        RECT 22.980000 64.210000 23.180000 64.410000 ;
        RECT 22.980000 64.620000 23.180000 64.820000 ;
        RECT 22.980000 65.030000 23.180000 65.230000 ;
        RECT 22.980000 65.440000 23.180000 65.640000 ;
        RECT 22.980000 65.850000 23.180000 66.050000 ;
        RECT 22.980000 66.260000 23.180000 66.460000 ;
        RECT 23.390000 62.160000 23.590000 62.360000 ;
        RECT 23.390000 62.570000 23.590000 62.770000 ;
        RECT 23.390000 62.980000 23.590000 63.180000 ;
        RECT 23.390000 63.390000 23.590000 63.590000 ;
        RECT 23.390000 63.800000 23.590000 64.000000 ;
        RECT 23.390000 64.210000 23.590000 64.410000 ;
        RECT 23.390000 64.620000 23.590000 64.820000 ;
        RECT 23.390000 65.030000 23.590000 65.230000 ;
        RECT 23.390000 65.440000 23.590000 65.640000 ;
        RECT 23.390000 65.850000 23.590000 66.050000 ;
        RECT 23.390000 66.260000 23.590000 66.460000 ;
        RECT 23.800000 62.160000 24.000000 62.360000 ;
        RECT 23.800000 62.570000 24.000000 62.770000 ;
        RECT 23.800000 62.980000 24.000000 63.180000 ;
        RECT 23.800000 63.390000 24.000000 63.590000 ;
        RECT 23.800000 63.800000 24.000000 64.000000 ;
        RECT 23.800000 64.210000 24.000000 64.410000 ;
        RECT 23.800000 64.620000 24.000000 64.820000 ;
        RECT 23.800000 65.030000 24.000000 65.230000 ;
        RECT 23.800000 65.440000 24.000000 65.640000 ;
        RECT 23.800000 65.850000 24.000000 66.050000 ;
        RECT 23.800000 66.260000 24.000000 66.460000 ;
        RECT 24.210000 62.160000 24.410000 62.360000 ;
        RECT 24.210000 62.570000 24.410000 62.770000 ;
        RECT 24.210000 62.980000 24.410000 63.180000 ;
        RECT 24.210000 63.390000 24.410000 63.590000 ;
        RECT 24.210000 63.800000 24.410000 64.000000 ;
        RECT 24.210000 64.210000 24.410000 64.410000 ;
        RECT 24.210000 64.620000 24.410000 64.820000 ;
        RECT 24.210000 65.030000 24.410000 65.230000 ;
        RECT 24.210000 65.440000 24.410000 65.640000 ;
        RECT 24.210000 65.850000 24.410000 66.050000 ;
        RECT 24.210000 66.260000 24.410000 66.460000 ;
        RECT 50.845000 62.160000 51.045000 62.360000 ;
        RECT 50.845000 62.570000 51.045000 62.770000 ;
        RECT 50.845000 62.980000 51.045000 63.180000 ;
        RECT 50.845000 63.390000 51.045000 63.590000 ;
        RECT 50.845000 63.800000 51.045000 64.000000 ;
        RECT 50.845000 64.210000 51.045000 64.410000 ;
        RECT 50.845000 64.620000 51.045000 64.820000 ;
        RECT 50.845000 65.030000 51.045000 65.230000 ;
        RECT 50.845000 65.440000 51.045000 65.640000 ;
        RECT 50.845000 65.850000 51.045000 66.050000 ;
        RECT 50.845000 66.260000 51.045000 66.460000 ;
        RECT 51.250000 62.160000 51.450000 62.360000 ;
        RECT 51.250000 62.570000 51.450000 62.770000 ;
        RECT 51.250000 62.980000 51.450000 63.180000 ;
        RECT 51.250000 63.390000 51.450000 63.590000 ;
        RECT 51.250000 63.800000 51.450000 64.000000 ;
        RECT 51.250000 64.210000 51.450000 64.410000 ;
        RECT 51.250000 64.620000 51.450000 64.820000 ;
        RECT 51.250000 65.030000 51.450000 65.230000 ;
        RECT 51.250000 65.440000 51.450000 65.640000 ;
        RECT 51.250000 65.850000 51.450000 66.050000 ;
        RECT 51.250000 66.260000 51.450000 66.460000 ;
        RECT 51.655000 62.160000 51.855000 62.360000 ;
        RECT 51.655000 62.570000 51.855000 62.770000 ;
        RECT 51.655000 62.980000 51.855000 63.180000 ;
        RECT 51.655000 63.390000 51.855000 63.590000 ;
        RECT 51.655000 63.800000 51.855000 64.000000 ;
        RECT 51.655000 64.210000 51.855000 64.410000 ;
        RECT 51.655000 64.620000 51.855000 64.820000 ;
        RECT 51.655000 65.030000 51.855000 65.230000 ;
        RECT 51.655000 65.440000 51.855000 65.640000 ;
        RECT 51.655000 65.850000 51.855000 66.050000 ;
        RECT 51.655000 66.260000 51.855000 66.460000 ;
        RECT 52.060000 62.160000 52.260000 62.360000 ;
        RECT 52.060000 62.570000 52.260000 62.770000 ;
        RECT 52.060000 62.980000 52.260000 63.180000 ;
        RECT 52.060000 63.390000 52.260000 63.590000 ;
        RECT 52.060000 63.800000 52.260000 64.000000 ;
        RECT 52.060000 64.210000 52.260000 64.410000 ;
        RECT 52.060000 64.620000 52.260000 64.820000 ;
        RECT 52.060000 65.030000 52.260000 65.230000 ;
        RECT 52.060000 65.440000 52.260000 65.640000 ;
        RECT 52.060000 65.850000 52.260000 66.050000 ;
        RECT 52.060000 66.260000 52.260000 66.460000 ;
        RECT 52.465000 62.160000 52.665000 62.360000 ;
        RECT 52.465000 62.570000 52.665000 62.770000 ;
        RECT 52.465000 62.980000 52.665000 63.180000 ;
        RECT 52.465000 63.390000 52.665000 63.590000 ;
        RECT 52.465000 63.800000 52.665000 64.000000 ;
        RECT 52.465000 64.210000 52.665000 64.410000 ;
        RECT 52.465000 64.620000 52.665000 64.820000 ;
        RECT 52.465000 65.030000 52.665000 65.230000 ;
        RECT 52.465000 65.440000 52.665000 65.640000 ;
        RECT 52.465000 65.850000 52.665000 66.050000 ;
        RECT 52.465000 66.260000 52.665000 66.460000 ;
        RECT 52.870000 62.160000 53.070000 62.360000 ;
        RECT 52.870000 62.570000 53.070000 62.770000 ;
        RECT 52.870000 62.980000 53.070000 63.180000 ;
        RECT 52.870000 63.390000 53.070000 63.590000 ;
        RECT 52.870000 63.800000 53.070000 64.000000 ;
        RECT 52.870000 64.210000 53.070000 64.410000 ;
        RECT 52.870000 64.620000 53.070000 64.820000 ;
        RECT 52.870000 65.030000 53.070000 65.230000 ;
        RECT 52.870000 65.440000 53.070000 65.640000 ;
        RECT 52.870000 65.850000 53.070000 66.050000 ;
        RECT 52.870000 66.260000 53.070000 66.460000 ;
        RECT 53.275000 62.160000 53.475000 62.360000 ;
        RECT 53.275000 62.570000 53.475000 62.770000 ;
        RECT 53.275000 62.980000 53.475000 63.180000 ;
        RECT 53.275000 63.390000 53.475000 63.590000 ;
        RECT 53.275000 63.800000 53.475000 64.000000 ;
        RECT 53.275000 64.210000 53.475000 64.410000 ;
        RECT 53.275000 64.620000 53.475000 64.820000 ;
        RECT 53.275000 65.030000 53.475000 65.230000 ;
        RECT 53.275000 65.440000 53.475000 65.640000 ;
        RECT 53.275000 65.850000 53.475000 66.050000 ;
        RECT 53.275000 66.260000 53.475000 66.460000 ;
        RECT 53.680000 62.160000 53.880000 62.360000 ;
        RECT 53.680000 62.570000 53.880000 62.770000 ;
        RECT 53.680000 62.980000 53.880000 63.180000 ;
        RECT 53.680000 63.390000 53.880000 63.590000 ;
        RECT 53.680000 63.800000 53.880000 64.000000 ;
        RECT 53.680000 64.210000 53.880000 64.410000 ;
        RECT 53.680000 64.620000 53.880000 64.820000 ;
        RECT 53.680000 65.030000 53.880000 65.230000 ;
        RECT 53.680000 65.440000 53.880000 65.640000 ;
        RECT 53.680000 65.850000 53.880000 66.050000 ;
        RECT 53.680000 66.260000 53.880000 66.460000 ;
        RECT 54.085000 62.160000 54.285000 62.360000 ;
        RECT 54.085000 62.570000 54.285000 62.770000 ;
        RECT 54.085000 62.980000 54.285000 63.180000 ;
        RECT 54.085000 63.390000 54.285000 63.590000 ;
        RECT 54.085000 63.800000 54.285000 64.000000 ;
        RECT 54.085000 64.210000 54.285000 64.410000 ;
        RECT 54.085000 64.620000 54.285000 64.820000 ;
        RECT 54.085000 65.030000 54.285000 65.230000 ;
        RECT 54.085000 65.440000 54.285000 65.640000 ;
        RECT 54.085000 65.850000 54.285000 66.050000 ;
        RECT 54.085000 66.260000 54.285000 66.460000 ;
        RECT 54.490000 62.160000 54.690000 62.360000 ;
        RECT 54.490000 62.570000 54.690000 62.770000 ;
        RECT 54.490000 62.980000 54.690000 63.180000 ;
        RECT 54.490000 63.390000 54.690000 63.590000 ;
        RECT 54.490000 63.800000 54.690000 64.000000 ;
        RECT 54.490000 64.210000 54.690000 64.410000 ;
        RECT 54.490000 64.620000 54.690000 64.820000 ;
        RECT 54.490000 65.030000 54.690000 65.230000 ;
        RECT 54.490000 65.440000 54.690000 65.640000 ;
        RECT 54.490000 65.850000 54.690000 66.050000 ;
        RECT 54.490000 66.260000 54.690000 66.460000 ;
        RECT 54.895000 62.160000 55.095000 62.360000 ;
        RECT 54.895000 62.570000 55.095000 62.770000 ;
        RECT 54.895000 62.980000 55.095000 63.180000 ;
        RECT 54.895000 63.390000 55.095000 63.590000 ;
        RECT 54.895000 63.800000 55.095000 64.000000 ;
        RECT 54.895000 64.210000 55.095000 64.410000 ;
        RECT 54.895000 64.620000 55.095000 64.820000 ;
        RECT 54.895000 65.030000 55.095000 65.230000 ;
        RECT 54.895000 65.440000 55.095000 65.640000 ;
        RECT 54.895000 65.850000 55.095000 66.050000 ;
        RECT 54.895000 66.260000 55.095000 66.460000 ;
        RECT 55.300000 62.160000 55.500000 62.360000 ;
        RECT 55.300000 62.570000 55.500000 62.770000 ;
        RECT 55.300000 62.980000 55.500000 63.180000 ;
        RECT 55.300000 63.390000 55.500000 63.590000 ;
        RECT 55.300000 63.800000 55.500000 64.000000 ;
        RECT 55.300000 64.210000 55.500000 64.410000 ;
        RECT 55.300000 64.620000 55.500000 64.820000 ;
        RECT 55.300000 65.030000 55.500000 65.230000 ;
        RECT 55.300000 65.440000 55.500000 65.640000 ;
        RECT 55.300000 65.850000 55.500000 66.050000 ;
        RECT 55.300000 66.260000 55.500000 66.460000 ;
        RECT 55.705000 62.160000 55.905000 62.360000 ;
        RECT 55.705000 62.570000 55.905000 62.770000 ;
        RECT 55.705000 62.980000 55.905000 63.180000 ;
        RECT 55.705000 63.390000 55.905000 63.590000 ;
        RECT 55.705000 63.800000 55.905000 64.000000 ;
        RECT 55.705000 64.210000 55.905000 64.410000 ;
        RECT 55.705000 64.620000 55.905000 64.820000 ;
        RECT 55.705000 65.030000 55.905000 65.230000 ;
        RECT 55.705000 65.440000 55.905000 65.640000 ;
        RECT 55.705000 65.850000 55.905000 66.050000 ;
        RECT 55.705000 66.260000 55.905000 66.460000 ;
        RECT 56.110000 62.160000 56.310000 62.360000 ;
        RECT 56.110000 62.570000 56.310000 62.770000 ;
        RECT 56.110000 62.980000 56.310000 63.180000 ;
        RECT 56.110000 63.390000 56.310000 63.590000 ;
        RECT 56.110000 63.800000 56.310000 64.000000 ;
        RECT 56.110000 64.210000 56.310000 64.410000 ;
        RECT 56.110000 64.620000 56.310000 64.820000 ;
        RECT 56.110000 65.030000 56.310000 65.230000 ;
        RECT 56.110000 65.440000 56.310000 65.640000 ;
        RECT 56.110000 65.850000 56.310000 66.050000 ;
        RECT 56.110000 66.260000 56.310000 66.460000 ;
        RECT 56.515000 62.160000 56.715000 62.360000 ;
        RECT 56.515000 62.570000 56.715000 62.770000 ;
        RECT 56.515000 62.980000 56.715000 63.180000 ;
        RECT 56.515000 63.390000 56.715000 63.590000 ;
        RECT 56.515000 63.800000 56.715000 64.000000 ;
        RECT 56.515000 64.210000 56.715000 64.410000 ;
        RECT 56.515000 64.620000 56.715000 64.820000 ;
        RECT 56.515000 65.030000 56.715000 65.230000 ;
        RECT 56.515000 65.440000 56.715000 65.640000 ;
        RECT 56.515000 65.850000 56.715000 66.050000 ;
        RECT 56.515000 66.260000 56.715000 66.460000 ;
        RECT 56.920000 62.160000 57.120000 62.360000 ;
        RECT 56.920000 62.570000 57.120000 62.770000 ;
        RECT 56.920000 62.980000 57.120000 63.180000 ;
        RECT 56.920000 63.390000 57.120000 63.590000 ;
        RECT 56.920000 63.800000 57.120000 64.000000 ;
        RECT 56.920000 64.210000 57.120000 64.410000 ;
        RECT 56.920000 64.620000 57.120000 64.820000 ;
        RECT 56.920000 65.030000 57.120000 65.230000 ;
        RECT 56.920000 65.440000 57.120000 65.640000 ;
        RECT 56.920000 65.850000 57.120000 66.050000 ;
        RECT 56.920000 66.260000 57.120000 66.460000 ;
        RECT 57.325000 62.160000 57.525000 62.360000 ;
        RECT 57.325000 62.570000 57.525000 62.770000 ;
        RECT 57.325000 62.980000 57.525000 63.180000 ;
        RECT 57.325000 63.390000 57.525000 63.590000 ;
        RECT 57.325000 63.800000 57.525000 64.000000 ;
        RECT 57.325000 64.210000 57.525000 64.410000 ;
        RECT 57.325000 64.620000 57.525000 64.820000 ;
        RECT 57.325000 65.030000 57.525000 65.230000 ;
        RECT 57.325000 65.440000 57.525000 65.640000 ;
        RECT 57.325000 65.850000 57.525000 66.050000 ;
        RECT 57.325000 66.260000 57.525000 66.460000 ;
        RECT 57.730000 62.160000 57.930000 62.360000 ;
        RECT 57.730000 62.570000 57.930000 62.770000 ;
        RECT 57.730000 62.980000 57.930000 63.180000 ;
        RECT 57.730000 63.390000 57.930000 63.590000 ;
        RECT 57.730000 63.800000 57.930000 64.000000 ;
        RECT 57.730000 64.210000 57.930000 64.410000 ;
        RECT 57.730000 64.620000 57.930000 64.820000 ;
        RECT 57.730000 65.030000 57.930000 65.230000 ;
        RECT 57.730000 65.440000 57.930000 65.640000 ;
        RECT 57.730000 65.850000 57.930000 66.050000 ;
        RECT 57.730000 66.260000 57.930000 66.460000 ;
        RECT 58.135000 62.160000 58.335000 62.360000 ;
        RECT 58.135000 62.570000 58.335000 62.770000 ;
        RECT 58.135000 62.980000 58.335000 63.180000 ;
        RECT 58.135000 63.390000 58.335000 63.590000 ;
        RECT 58.135000 63.800000 58.335000 64.000000 ;
        RECT 58.135000 64.210000 58.335000 64.410000 ;
        RECT 58.135000 64.620000 58.335000 64.820000 ;
        RECT 58.135000 65.030000 58.335000 65.230000 ;
        RECT 58.135000 65.440000 58.335000 65.640000 ;
        RECT 58.135000 65.850000 58.335000 66.050000 ;
        RECT 58.135000 66.260000 58.335000 66.460000 ;
        RECT 58.540000 62.160000 58.740000 62.360000 ;
        RECT 58.540000 62.570000 58.740000 62.770000 ;
        RECT 58.540000 62.980000 58.740000 63.180000 ;
        RECT 58.540000 63.390000 58.740000 63.590000 ;
        RECT 58.540000 63.800000 58.740000 64.000000 ;
        RECT 58.540000 64.210000 58.740000 64.410000 ;
        RECT 58.540000 64.620000 58.740000 64.820000 ;
        RECT 58.540000 65.030000 58.740000 65.230000 ;
        RECT 58.540000 65.440000 58.740000 65.640000 ;
        RECT 58.540000 65.850000 58.740000 66.050000 ;
        RECT 58.540000 66.260000 58.740000 66.460000 ;
        RECT 58.945000 62.160000 59.145000 62.360000 ;
        RECT 58.945000 62.570000 59.145000 62.770000 ;
        RECT 58.945000 62.980000 59.145000 63.180000 ;
        RECT 58.945000 63.390000 59.145000 63.590000 ;
        RECT 58.945000 63.800000 59.145000 64.000000 ;
        RECT 58.945000 64.210000 59.145000 64.410000 ;
        RECT 58.945000 64.620000 59.145000 64.820000 ;
        RECT 58.945000 65.030000 59.145000 65.230000 ;
        RECT 58.945000 65.440000 59.145000 65.640000 ;
        RECT 58.945000 65.850000 59.145000 66.050000 ;
        RECT 58.945000 66.260000 59.145000 66.460000 ;
        RECT 59.350000 62.160000 59.550000 62.360000 ;
        RECT 59.350000 62.570000 59.550000 62.770000 ;
        RECT 59.350000 62.980000 59.550000 63.180000 ;
        RECT 59.350000 63.390000 59.550000 63.590000 ;
        RECT 59.350000 63.800000 59.550000 64.000000 ;
        RECT 59.350000 64.210000 59.550000 64.410000 ;
        RECT 59.350000 64.620000 59.550000 64.820000 ;
        RECT 59.350000 65.030000 59.550000 65.230000 ;
        RECT 59.350000 65.440000 59.550000 65.640000 ;
        RECT 59.350000 65.850000 59.550000 66.050000 ;
        RECT 59.350000 66.260000 59.550000 66.460000 ;
        RECT 59.755000 62.160000 59.955000 62.360000 ;
        RECT 59.755000 62.570000 59.955000 62.770000 ;
        RECT 59.755000 62.980000 59.955000 63.180000 ;
        RECT 59.755000 63.390000 59.955000 63.590000 ;
        RECT 59.755000 63.800000 59.955000 64.000000 ;
        RECT 59.755000 64.210000 59.955000 64.410000 ;
        RECT 59.755000 64.620000 59.955000 64.820000 ;
        RECT 59.755000 65.030000 59.955000 65.230000 ;
        RECT 59.755000 65.440000 59.955000 65.640000 ;
        RECT 59.755000 65.850000 59.955000 66.050000 ;
        RECT 59.755000 66.260000 59.955000 66.460000 ;
        RECT 60.160000 62.160000 60.360000 62.360000 ;
        RECT 60.160000 62.570000 60.360000 62.770000 ;
        RECT 60.160000 62.980000 60.360000 63.180000 ;
        RECT 60.160000 63.390000 60.360000 63.590000 ;
        RECT 60.160000 63.800000 60.360000 64.000000 ;
        RECT 60.160000 64.210000 60.360000 64.410000 ;
        RECT 60.160000 64.620000 60.360000 64.820000 ;
        RECT 60.160000 65.030000 60.360000 65.230000 ;
        RECT 60.160000 65.440000 60.360000 65.640000 ;
        RECT 60.160000 65.850000 60.360000 66.050000 ;
        RECT 60.160000 66.260000 60.360000 66.460000 ;
        RECT 60.565000 62.160000 60.765000 62.360000 ;
        RECT 60.565000 62.570000 60.765000 62.770000 ;
        RECT 60.565000 62.980000 60.765000 63.180000 ;
        RECT 60.565000 63.390000 60.765000 63.590000 ;
        RECT 60.565000 63.800000 60.765000 64.000000 ;
        RECT 60.565000 64.210000 60.765000 64.410000 ;
        RECT 60.565000 64.620000 60.765000 64.820000 ;
        RECT 60.565000 65.030000 60.765000 65.230000 ;
        RECT 60.565000 65.440000 60.765000 65.640000 ;
        RECT 60.565000 65.850000 60.765000 66.050000 ;
        RECT 60.565000 66.260000 60.765000 66.460000 ;
        RECT 60.970000 62.160000 61.170000 62.360000 ;
        RECT 60.970000 62.570000 61.170000 62.770000 ;
        RECT 60.970000 62.980000 61.170000 63.180000 ;
        RECT 60.970000 63.390000 61.170000 63.590000 ;
        RECT 60.970000 63.800000 61.170000 64.000000 ;
        RECT 60.970000 64.210000 61.170000 64.410000 ;
        RECT 60.970000 64.620000 61.170000 64.820000 ;
        RECT 60.970000 65.030000 61.170000 65.230000 ;
        RECT 60.970000 65.440000 61.170000 65.640000 ;
        RECT 60.970000 65.850000 61.170000 66.050000 ;
        RECT 60.970000 66.260000 61.170000 66.460000 ;
        RECT 61.375000 62.160000 61.575000 62.360000 ;
        RECT 61.375000 62.570000 61.575000 62.770000 ;
        RECT 61.375000 62.980000 61.575000 63.180000 ;
        RECT 61.375000 63.390000 61.575000 63.590000 ;
        RECT 61.375000 63.800000 61.575000 64.000000 ;
        RECT 61.375000 64.210000 61.575000 64.410000 ;
        RECT 61.375000 64.620000 61.575000 64.820000 ;
        RECT 61.375000 65.030000 61.575000 65.230000 ;
        RECT 61.375000 65.440000 61.575000 65.640000 ;
        RECT 61.375000 65.850000 61.575000 66.050000 ;
        RECT 61.375000 66.260000 61.575000 66.460000 ;
        RECT 61.780000 62.160000 61.980000 62.360000 ;
        RECT 61.780000 62.570000 61.980000 62.770000 ;
        RECT 61.780000 62.980000 61.980000 63.180000 ;
        RECT 61.780000 63.390000 61.980000 63.590000 ;
        RECT 61.780000 63.800000 61.980000 64.000000 ;
        RECT 61.780000 64.210000 61.980000 64.410000 ;
        RECT 61.780000 64.620000 61.980000 64.820000 ;
        RECT 61.780000 65.030000 61.980000 65.230000 ;
        RECT 61.780000 65.440000 61.980000 65.640000 ;
        RECT 61.780000 65.850000 61.980000 66.050000 ;
        RECT 61.780000 66.260000 61.980000 66.460000 ;
        RECT 62.185000 62.160000 62.385000 62.360000 ;
        RECT 62.185000 62.570000 62.385000 62.770000 ;
        RECT 62.185000 62.980000 62.385000 63.180000 ;
        RECT 62.185000 63.390000 62.385000 63.590000 ;
        RECT 62.185000 63.800000 62.385000 64.000000 ;
        RECT 62.185000 64.210000 62.385000 64.410000 ;
        RECT 62.185000 64.620000 62.385000 64.820000 ;
        RECT 62.185000 65.030000 62.385000 65.230000 ;
        RECT 62.185000 65.440000 62.385000 65.640000 ;
        RECT 62.185000 65.850000 62.385000 66.050000 ;
        RECT 62.185000 66.260000 62.385000 66.460000 ;
        RECT 62.590000 62.160000 62.790000 62.360000 ;
        RECT 62.590000 62.570000 62.790000 62.770000 ;
        RECT 62.590000 62.980000 62.790000 63.180000 ;
        RECT 62.590000 63.390000 62.790000 63.590000 ;
        RECT 62.590000 63.800000 62.790000 64.000000 ;
        RECT 62.590000 64.210000 62.790000 64.410000 ;
        RECT 62.590000 64.620000 62.790000 64.820000 ;
        RECT 62.590000 65.030000 62.790000 65.230000 ;
        RECT 62.590000 65.440000 62.790000 65.640000 ;
        RECT 62.590000 65.850000 62.790000 66.050000 ;
        RECT 62.590000 66.260000 62.790000 66.460000 ;
        RECT 62.995000 62.160000 63.195000 62.360000 ;
        RECT 62.995000 62.570000 63.195000 62.770000 ;
        RECT 62.995000 62.980000 63.195000 63.180000 ;
        RECT 62.995000 63.390000 63.195000 63.590000 ;
        RECT 62.995000 63.800000 63.195000 64.000000 ;
        RECT 62.995000 64.210000 63.195000 64.410000 ;
        RECT 62.995000 64.620000 63.195000 64.820000 ;
        RECT 62.995000 65.030000 63.195000 65.230000 ;
        RECT 62.995000 65.440000 63.195000 65.640000 ;
        RECT 62.995000 65.850000 63.195000 66.050000 ;
        RECT 62.995000 66.260000 63.195000 66.460000 ;
        RECT 63.400000 62.160000 63.600000 62.360000 ;
        RECT 63.400000 62.570000 63.600000 62.770000 ;
        RECT 63.400000 62.980000 63.600000 63.180000 ;
        RECT 63.400000 63.390000 63.600000 63.590000 ;
        RECT 63.400000 63.800000 63.600000 64.000000 ;
        RECT 63.400000 64.210000 63.600000 64.410000 ;
        RECT 63.400000 64.620000 63.600000 64.820000 ;
        RECT 63.400000 65.030000 63.600000 65.230000 ;
        RECT 63.400000 65.440000 63.600000 65.640000 ;
        RECT 63.400000 65.850000 63.600000 66.050000 ;
        RECT 63.400000 66.260000 63.600000 66.460000 ;
        RECT 63.805000 62.160000 64.005000 62.360000 ;
        RECT 63.805000 62.570000 64.005000 62.770000 ;
        RECT 63.805000 62.980000 64.005000 63.180000 ;
        RECT 63.805000 63.390000 64.005000 63.590000 ;
        RECT 63.805000 63.800000 64.005000 64.000000 ;
        RECT 63.805000 64.210000 64.005000 64.410000 ;
        RECT 63.805000 64.620000 64.005000 64.820000 ;
        RECT 63.805000 65.030000 64.005000 65.230000 ;
        RECT 63.805000 65.440000 64.005000 65.640000 ;
        RECT 63.805000 65.850000 64.005000 66.050000 ;
        RECT 63.805000 66.260000 64.005000 66.460000 ;
        RECT 64.210000 62.160000 64.410000 62.360000 ;
        RECT 64.210000 62.570000 64.410000 62.770000 ;
        RECT 64.210000 62.980000 64.410000 63.180000 ;
        RECT 64.210000 63.390000 64.410000 63.590000 ;
        RECT 64.210000 63.800000 64.410000 64.000000 ;
        RECT 64.210000 64.210000 64.410000 64.410000 ;
        RECT 64.210000 64.620000 64.410000 64.820000 ;
        RECT 64.210000 65.030000 64.410000 65.230000 ;
        RECT 64.210000 65.440000 64.410000 65.640000 ;
        RECT 64.210000 65.850000 64.410000 66.050000 ;
        RECT 64.210000 66.260000 64.410000 66.460000 ;
        RECT 64.615000 62.160000 64.815000 62.360000 ;
        RECT 64.615000 62.570000 64.815000 62.770000 ;
        RECT 64.615000 62.980000 64.815000 63.180000 ;
        RECT 64.615000 63.390000 64.815000 63.590000 ;
        RECT 64.615000 63.800000 64.815000 64.000000 ;
        RECT 64.615000 64.210000 64.815000 64.410000 ;
        RECT 64.615000 64.620000 64.815000 64.820000 ;
        RECT 64.615000 65.030000 64.815000 65.230000 ;
        RECT 64.615000 65.440000 64.815000 65.640000 ;
        RECT 64.615000 65.850000 64.815000 66.050000 ;
        RECT 64.615000 66.260000 64.815000 66.460000 ;
        RECT 65.020000 62.160000 65.220000 62.360000 ;
        RECT 65.020000 62.570000 65.220000 62.770000 ;
        RECT 65.020000 62.980000 65.220000 63.180000 ;
        RECT 65.020000 63.390000 65.220000 63.590000 ;
        RECT 65.020000 63.800000 65.220000 64.000000 ;
        RECT 65.020000 64.210000 65.220000 64.410000 ;
        RECT 65.020000 64.620000 65.220000 64.820000 ;
        RECT 65.020000 65.030000 65.220000 65.230000 ;
        RECT 65.020000 65.440000 65.220000 65.640000 ;
        RECT 65.020000 65.850000 65.220000 66.050000 ;
        RECT 65.020000 66.260000 65.220000 66.460000 ;
        RECT 65.425000 62.160000 65.625000 62.360000 ;
        RECT 65.425000 62.570000 65.625000 62.770000 ;
        RECT 65.425000 62.980000 65.625000 63.180000 ;
        RECT 65.425000 63.390000 65.625000 63.590000 ;
        RECT 65.425000 63.800000 65.625000 64.000000 ;
        RECT 65.425000 64.210000 65.625000 64.410000 ;
        RECT 65.425000 64.620000 65.625000 64.820000 ;
        RECT 65.425000 65.030000 65.625000 65.230000 ;
        RECT 65.425000 65.440000 65.625000 65.640000 ;
        RECT 65.425000 65.850000 65.625000 66.050000 ;
        RECT 65.425000 66.260000 65.625000 66.460000 ;
        RECT 65.830000 62.160000 66.030000 62.360000 ;
        RECT 65.830000 62.570000 66.030000 62.770000 ;
        RECT 65.830000 62.980000 66.030000 63.180000 ;
        RECT 65.830000 63.390000 66.030000 63.590000 ;
        RECT 65.830000 63.800000 66.030000 64.000000 ;
        RECT 65.830000 64.210000 66.030000 64.410000 ;
        RECT 65.830000 64.620000 66.030000 64.820000 ;
        RECT 65.830000 65.030000 66.030000 65.230000 ;
        RECT 65.830000 65.440000 66.030000 65.640000 ;
        RECT 65.830000 65.850000 66.030000 66.050000 ;
        RECT 65.830000 66.260000 66.030000 66.460000 ;
        RECT 66.235000 62.160000 66.435000 62.360000 ;
        RECT 66.235000 62.570000 66.435000 62.770000 ;
        RECT 66.235000 62.980000 66.435000 63.180000 ;
        RECT 66.235000 63.390000 66.435000 63.590000 ;
        RECT 66.235000 63.800000 66.435000 64.000000 ;
        RECT 66.235000 64.210000 66.435000 64.410000 ;
        RECT 66.235000 64.620000 66.435000 64.820000 ;
        RECT 66.235000 65.030000 66.435000 65.230000 ;
        RECT 66.235000 65.440000 66.435000 65.640000 ;
        RECT 66.235000 65.850000 66.435000 66.050000 ;
        RECT 66.235000 66.260000 66.435000 66.460000 ;
        RECT 66.640000 62.160000 66.840000 62.360000 ;
        RECT 66.640000 62.570000 66.840000 62.770000 ;
        RECT 66.640000 62.980000 66.840000 63.180000 ;
        RECT 66.640000 63.390000 66.840000 63.590000 ;
        RECT 66.640000 63.800000 66.840000 64.000000 ;
        RECT 66.640000 64.210000 66.840000 64.410000 ;
        RECT 66.640000 64.620000 66.840000 64.820000 ;
        RECT 66.640000 65.030000 66.840000 65.230000 ;
        RECT 66.640000 65.440000 66.840000 65.640000 ;
        RECT 66.640000 65.850000 66.840000 66.050000 ;
        RECT 66.640000 66.260000 66.840000 66.460000 ;
        RECT 67.045000 62.160000 67.245000 62.360000 ;
        RECT 67.045000 62.570000 67.245000 62.770000 ;
        RECT 67.045000 62.980000 67.245000 63.180000 ;
        RECT 67.045000 63.390000 67.245000 63.590000 ;
        RECT 67.045000 63.800000 67.245000 64.000000 ;
        RECT 67.045000 64.210000 67.245000 64.410000 ;
        RECT 67.045000 64.620000 67.245000 64.820000 ;
        RECT 67.045000 65.030000 67.245000 65.230000 ;
        RECT 67.045000 65.440000 67.245000 65.640000 ;
        RECT 67.045000 65.850000 67.245000 66.050000 ;
        RECT 67.045000 66.260000 67.245000 66.460000 ;
        RECT 67.450000 62.160000 67.650000 62.360000 ;
        RECT 67.450000 62.570000 67.650000 62.770000 ;
        RECT 67.450000 62.980000 67.650000 63.180000 ;
        RECT 67.450000 63.390000 67.650000 63.590000 ;
        RECT 67.450000 63.800000 67.650000 64.000000 ;
        RECT 67.450000 64.210000 67.650000 64.410000 ;
        RECT 67.450000 64.620000 67.650000 64.820000 ;
        RECT 67.450000 65.030000 67.650000 65.230000 ;
        RECT 67.450000 65.440000 67.650000 65.640000 ;
        RECT 67.450000 65.850000 67.650000 66.050000 ;
        RECT 67.450000 66.260000 67.650000 66.460000 ;
        RECT 67.855000 62.160000 68.055000 62.360000 ;
        RECT 67.855000 62.570000 68.055000 62.770000 ;
        RECT 67.855000 62.980000 68.055000 63.180000 ;
        RECT 67.855000 63.390000 68.055000 63.590000 ;
        RECT 67.855000 63.800000 68.055000 64.000000 ;
        RECT 67.855000 64.210000 68.055000 64.410000 ;
        RECT 67.855000 64.620000 68.055000 64.820000 ;
        RECT 67.855000 65.030000 68.055000 65.230000 ;
        RECT 67.855000 65.440000 68.055000 65.640000 ;
        RECT 67.855000 65.850000 68.055000 66.050000 ;
        RECT 67.855000 66.260000 68.055000 66.460000 ;
        RECT 68.260000 62.160000 68.460000 62.360000 ;
        RECT 68.260000 62.570000 68.460000 62.770000 ;
        RECT 68.260000 62.980000 68.460000 63.180000 ;
        RECT 68.260000 63.390000 68.460000 63.590000 ;
        RECT 68.260000 63.800000 68.460000 64.000000 ;
        RECT 68.260000 64.210000 68.460000 64.410000 ;
        RECT 68.260000 64.620000 68.460000 64.820000 ;
        RECT 68.260000 65.030000 68.460000 65.230000 ;
        RECT 68.260000 65.440000 68.460000 65.640000 ;
        RECT 68.260000 65.850000 68.460000 66.050000 ;
        RECT 68.260000 66.260000 68.460000 66.460000 ;
        RECT 68.665000 62.160000 68.865000 62.360000 ;
        RECT 68.665000 62.570000 68.865000 62.770000 ;
        RECT 68.665000 62.980000 68.865000 63.180000 ;
        RECT 68.665000 63.390000 68.865000 63.590000 ;
        RECT 68.665000 63.800000 68.865000 64.000000 ;
        RECT 68.665000 64.210000 68.865000 64.410000 ;
        RECT 68.665000 64.620000 68.865000 64.820000 ;
        RECT 68.665000 65.030000 68.865000 65.230000 ;
        RECT 68.665000 65.440000 68.865000 65.640000 ;
        RECT 68.665000 65.850000 68.865000 66.050000 ;
        RECT 68.665000 66.260000 68.865000 66.460000 ;
        RECT 69.070000 62.160000 69.270000 62.360000 ;
        RECT 69.070000 62.570000 69.270000 62.770000 ;
        RECT 69.070000 62.980000 69.270000 63.180000 ;
        RECT 69.070000 63.390000 69.270000 63.590000 ;
        RECT 69.070000 63.800000 69.270000 64.000000 ;
        RECT 69.070000 64.210000 69.270000 64.410000 ;
        RECT 69.070000 64.620000 69.270000 64.820000 ;
        RECT 69.070000 65.030000 69.270000 65.230000 ;
        RECT 69.070000 65.440000 69.270000 65.640000 ;
        RECT 69.070000 65.850000 69.270000 66.050000 ;
        RECT 69.070000 66.260000 69.270000 66.460000 ;
        RECT 69.475000 62.160000 69.675000 62.360000 ;
        RECT 69.475000 62.570000 69.675000 62.770000 ;
        RECT 69.475000 62.980000 69.675000 63.180000 ;
        RECT 69.475000 63.390000 69.675000 63.590000 ;
        RECT 69.475000 63.800000 69.675000 64.000000 ;
        RECT 69.475000 64.210000 69.675000 64.410000 ;
        RECT 69.475000 64.620000 69.675000 64.820000 ;
        RECT 69.475000 65.030000 69.675000 65.230000 ;
        RECT 69.475000 65.440000 69.675000 65.640000 ;
        RECT 69.475000 65.850000 69.675000 66.050000 ;
        RECT 69.475000 66.260000 69.675000 66.460000 ;
        RECT 69.880000 62.160000 70.080000 62.360000 ;
        RECT 69.880000 62.570000 70.080000 62.770000 ;
        RECT 69.880000 62.980000 70.080000 63.180000 ;
        RECT 69.880000 63.390000 70.080000 63.590000 ;
        RECT 69.880000 63.800000 70.080000 64.000000 ;
        RECT 69.880000 64.210000 70.080000 64.410000 ;
        RECT 69.880000 64.620000 70.080000 64.820000 ;
        RECT 69.880000 65.030000 70.080000 65.230000 ;
        RECT 69.880000 65.440000 70.080000 65.640000 ;
        RECT 69.880000 65.850000 70.080000 66.050000 ;
        RECT 69.880000 66.260000 70.080000 66.460000 ;
        RECT 70.285000 62.160000 70.485000 62.360000 ;
        RECT 70.285000 62.570000 70.485000 62.770000 ;
        RECT 70.285000 62.980000 70.485000 63.180000 ;
        RECT 70.285000 63.390000 70.485000 63.590000 ;
        RECT 70.285000 63.800000 70.485000 64.000000 ;
        RECT 70.285000 64.210000 70.485000 64.410000 ;
        RECT 70.285000 64.620000 70.485000 64.820000 ;
        RECT 70.285000 65.030000 70.485000 65.230000 ;
        RECT 70.285000 65.440000 70.485000 65.640000 ;
        RECT 70.285000 65.850000 70.485000 66.050000 ;
        RECT 70.285000 66.260000 70.485000 66.460000 ;
        RECT 70.690000 62.160000 70.890000 62.360000 ;
        RECT 70.690000 62.570000 70.890000 62.770000 ;
        RECT 70.690000 62.980000 70.890000 63.180000 ;
        RECT 70.690000 63.390000 70.890000 63.590000 ;
        RECT 70.690000 63.800000 70.890000 64.000000 ;
        RECT 70.690000 64.210000 70.890000 64.410000 ;
        RECT 70.690000 64.620000 70.890000 64.820000 ;
        RECT 70.690000 65.030000 70.890000 65.230000 ;
        RECT 70.690000 65.440000 70.890000 65.640000 ;
        RECT 70.690000 65.850000 70.890000 66.050000 ;
        RECT 70.690000 66.260000 70.890000 66.460000 ;
        RECT 71.095000 62.160000 71.295000 62.360000 ;
        RECT 71.095000 62.570000 71.295000 62.770000 ;
        RECT 71.095000 62.980000 71.295000 63.180000 ;
        RECT 71.095000 63.390000 71.295000 63.590000 ;
        RECT 71.095000 63.800000 71.295000 64.000000 ;
        RECT 71.095000 64.210000 71.295000 64.410000 ;
        RECT 71.095000 64.620000 71.295000 64.820000 ;
        RECT 71.095000 65.030000 71.295000 65.230000 ;
        RECT 71.095000 65.440000 71.295000 65.640000 ;
        RECT 71.095000 65.850000 71.295000 66.050000 ;
        RECT 71.095000 66.260000 71.295000 66.460000 ;
        RECT 71.500000 62.160000 71.700000 62.360000 ;
        RECT 71.500000 62.570000 71.700000 62.770000 ;
        RECT 71.500000 62.980000 71.700000 63.180000 ;
        RECT 71.500000 63.390000 71.700000 63.590000 ;
        RECT 71.500000 63.800000 71.700000 64.000000 ;
        RECT 71.500000 64.210000 71.700000 64.410000 ;
        RECT 71.500000 64.620000 71.700000 64.820000 ;
        RECT 71.500000 65.030000 71.700000 65.230000 ;
        RECT 71.500000 65.440000 71.700000 65.640000 ;
        RECT 71.500000 65.850000 71.700000 66.050000 ;
        RECT 71.500000 66.260000 71.700000 66.460000 ;
        RECT 71.905000 62.160000 72.105000 62.360000 ;
        RECT 71.905000 62.570000 72.105000 62.770000 ;
        RECT 71.905000 62.980000 72.105000 63.180000 ;
        RECT 71.905000 63.390000 72.105000 63.590000 ;
        RECT 71.905000 63.800000 72.105000 64.000000 ;
        RECT 71.905000 64.210000 72.105000 64.410000 ;
        RECT 71.905000 64.620000 72.105000 64.820000 ;
        RECT 71.905000 65.030000 72.105000 65.230000 ;
        RECT 71.905000 65.440000 72.105000 65.640000 ;
        RECT 71.905000 65.850000 72.105000 66.050000 ;
        RECT 71.905000 66.260000 72.105000 66.460000 ;
        RECT 72.315000 62.160000 72.515000 62.360000 ;
        RECT 72.315000 62.570000 72.515000 62.770000 ;
        RECT 72.315000 62.980000 72.515000 63.180000 ;
        RECT 72.315000 63.390000 72.515000 63.590000 ;
        RECT 72.315000 63.800000 72.515000 64.000000 ;
        RECT 72.315000 64.210000 72.515000 64.410000 ;
        RECT 72.315000 64.620000 72.515000 64.820000 ;
        RECT 72.315000 65.030000 72.515000 65.230000 ;
        RECT 72.315000 65.440000 72.515000 65.640000 ;
        RECT 72.315000 65.850000 72.515000 66.050000 ;
        RECT 72.315000 66.260000 72.515000 66.460000 ;
        RECT 72.725000 62.160000 72.925000 62.360000 ;
        RECT 72.725000 62.570000 72.925000 62.770000 ;
        RECT 72.725000 62.980000 72.925000 63.180000 ;
        RECT 72.725000 63.390000 72.925000 63.590000 ;
        RECT 72.725000 63.800000 72.925000 64.000000 ;
        RECT 72.725000 64.210000 72.925000 64.410000 ;
        RECT 72.725000 64.620000 72.925000 64.820000 ;
        RECT 72.725000 65.030000 72.925000 65.230000 ;
        RECT 72.725000 65.440000 72.925000 65.640000 ;
        RECT 72.725000 65.850000 72.925000 66.050000 ;
        RECT 72.725000 66.260000 72.925000 66.460000 ;
        RECT 73.135000 62.160000 73.335000 62.360000 ;
        RECT 73.135000 62.570000 73.335000 62.770000 ;
        RECT 73.135000 62.980000 73.335000 63.180000 ;
        RECT 73.135000 63.390000 73.335000 63.590000 ;
        RECT 73.135000 63.800000 73.335000 64.000000 ;
        RECT 73.135000 64.210000 73.335000 64.410000 ;
        RECT 73.135000 64.620000 73.335000 64.820000 ;
        RECT 73.135000 65.030000 73.335000 65.230000 ;
        RECT 73.135000 65.440000 73.335000 65.640000 ;
        RECT 73.135000 65.850000 73.335000 66.050000 ;
        RECT 73.135000 66.260000 73.335000 66.460000 ;
        RECT 73.545000 62.160000 73.745000 62.360000 ;
        RECT 73.545000 62.570000 73.745000 62.770000 ;
        RECT 73.545000 62.980000 73.745000 63.180000 ;
        RECT 73.545000 63.390000 73.745000 63.590000 ;
        RECT 73.545000 63.800000 73.745000 64.000000 ;
        RECT 73.545000 64.210000 73.745000 64.410000 ;
        RECT 73.545000 64.620000 73.745000 64.820000 ;
        RECT 73.545000 65.030000 73.745000 65.230000 ;
        RECT 73.545000 65.440000 73.745000 65.640000 ;
        RECT 73.545000 65.850000 73.745000 66.050000 ;
        RECT 73.545000 66.260000 73.745000 66.460000 ;
        RECT 73.955000 62.160000 74.155000 62.360000 ;
        RECT 73.955000 62.570000 74.155000 62.770000 ;
        RECT 73.955000 62.980000 74.155000 63.180000 ;
        RECT 73.955000 63.390000 74.155000 63.590000 ;
        RECT 73.955000 63.800000 74.155000 64.000000 ;
        RECT 73.955000 64.210000 74.155000 64.410000 ;
        RECT 73.955000 64.620000 74.155000 64.820000 ;
        RECT 73.955000 65.030000 74.155000 65.230000 ;
        RECT 73.955000 65.440000 74.155000 65.640000 ;
        RECT 73.955000 65.850000 74.155000 66.050000 ;
        RECT 73.955000 66.260000 74.155000 66.460000 ;
        RECT 74.365000 62.160000 74.565000 62.360000 ;
        RECT 74.365000 62.570000 74.565000 62.770000 ;
        RECT 74.365000 62.980000 74.565000 63.180000 ;
        RECT 74.365000 63.390000 74.565000 63.590000 ;
        RECT 74.365000 63.800000 74.565000 64.000000 ;
        RECT 74.365000 64.210000 74.565000 64.410000 ;
        RECT 74.365000 64.620000 74.565000 64.820000 ;
        RECT 74.365000 65.030000 74.565000 65.230000 ;
        RECT 74.365000 65.440000 74.565000 65.640000 ;
        RECT 74.365000 65.850000 74.565000 66.050000 ;
        RECT 74.365000 66.260000 74.565000 66.460000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 34.735000 1.270000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 45.735000 1.270000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 49.645000 1.270000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 54.405000 1.270000 54.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 34.735000 75.000000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 45.735000 75.000000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 49.645000 75.000000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 54.405000 75.000000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 34.840000 1.270000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 45.735000 1.270000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 34.840000 75.000000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 39.585000 1.270000 44.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 39.585000 75.000000 44.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 39.685000 1.270000 44.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 23.835000 1.270000 28.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 23.835000 75.000000 28.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 23.935000 1.270000 28.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 56.235000 1.270000 60.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.235000 75.000000 60.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 56.335000 1.270000 60.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 29.885000 1.270000 33.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 29.885000 75.000000 33.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 29.985000 1.270000 33.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 198.000000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 75.000000 198.000000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000 24.900000   3.005000 ;
      RECT  0.000000   3.005000  3.005000  14.385000 ;
      RECT  0.000000  14.385000 24.900000  17.390000 ;
      RECT  0.000000  22.830000 24.900000  25.835000 ;
      RECT  0.000000  25.835000  3.005000  58.685000 ;
      RECT  0.000000  58.685000 24.900000  61.690000 ;
      RECT  0.000000  66.930000 24.895000  67.635000 ;
      RECT  0.000000  93.355000 60.885000  93.360000 ;
      RECT  0.000000  93.360000 18.610000  96.365000 ;
      RECT  0.000000  96.365000  3.005000 194.995000 ;
      RECT  0.000000 194.995000 24.895000 198.000000 ;
      RECT  3.000000   3.002000 72.000000  14.390000 ;
      RECT  3.000000  25.830000 72.000000  58.690000 ;
      RECT  3.000000  96.355000 59.640000  96.360000 ;
      RECT  3.000000  96.355000 59.640000  96.360000 ;
      RECT  3.000000  96.360000 72.000000 195.000000 ;
      RECT 14.395000  93.330000 60.860000  93.355000 ;
      RECT 14.545000  93.180000 60.710000  93.330000 ;
      RECT 14.695000  93.030000 60.560000  93.180000 ;
      RECT 14.845000  92.880000 60.410000  93.030000 ;
      RECT 14.995000  92.730000 60.260000  92.880000 ;
      RECT 15.145000  92.580000 60.110000  92.730000 ;
      RECT 15.295000  92.430000 59.960000  92.580000 ;
      RECT 15.445000  92.280000 59.810000  92.430000 ;
      RECT 15.595000  92.130000 59.660000  92.280000 ;
      RECT 15.745000  91.980000 59.510000  92.130000 ;
      RECT 15.745000  96.225000 59.510000  96.355000 ;
      RECT 15.745000  96.225000 59.510000  96.355000 ;
      RECT 15.895000  91.830000 59.360000  91.980000 ;
      RECT 15.895000  96.075000 59.360000  96.225000 ;
      RECT 15.895000  96.075000 59.360000  96.225000 ;
      RECT 16.045000  91.680000 59.210000  91.830000 ;
      RECT 16.045000  95.925000 59.210000  96.075000 ;
      RECT 16.045000  95.925000 59.210000  96.075000 ;
      RECT 16.195000  91.530000 59.060000  91.680000 ;
      RECT 16.195000  95.775000 59.060000  95.925000 ;
      RECT 16.195000  95.775000 59.060000  95.925000 ;
      RECT 16.345000  91.380000 58.910000  91.530000 ;
      RECT 16.345000  95.625000 58.910000  95.775000 ;
      RECT 16.345000  95.625000 58.910000  95.775000 ;
      RECT 16.495000  91.230000 58.760000  91.380000 ;
      RECT 16.495000  95.475000 58.760000  95.625000 ;
      RECT 16.495000  95.475000 58.760000  95.625000 ;
      RECT 16.645000  91.080000 58.610000  91.230000 ;
      RECT 16.645000  95.325000 58.610000  95.475000 ;
      RECT 16.645000  95.325000 58.610000  95.475000 ;
      RECT 16.795000  90.930000 58.460000  91.080000 ;
      RECT 16.795000  95.175000 58.460000  95.325000 ;
      RECT 16.795000  95.175000 58.460000  95.325000 ;
      RECT 16.945000  90.780000 58.310000  90.930000 ;
      RECT 16.945000  95.025000 58.310000  95.175000 ;
      RECT 16.945000  95.025000 58.310000  95.175000 ;
      RECT 17.095000  90.630000 58.160000  90.780000 ;
      RECT 17.095000  94.875000 58.160000  95.025000 ;
      RECT 17.095000  94.875000 58.160000  95.025000 ;
      RECT 17.245000  90.480000 58.010000  90.630000 ;
      RECT 17.245000  94.725000 58.010000  94.875000 ;
      RECT 17.245000  94.725000 58.010000  94.875000 ;
      RECT 17.395000  90.330000 57.860000  90.480000 ;
      RECT 17.395000  94.575000 57.860000  94.725000 ;
      RECT 17.395000  94.575000 57.860000  94.725000 ;
      RECT 17.545000  90.180000 57.710000  90.330000 ;
      RECT 17.545000  94.425000 57.710000  94.575000 ;
      RECT 17.545000  94.425000 57.710000  94.575000 ;
      RECT 17.695000  90.030000 57.560000  90.180000 ;
      RECT 17.695000  94.275000 57.560000  94.425000 ;
      RECT 17.695000  94.275000 57.560000  94.425000 ;
      RECT 17.845000  89.880000 57.410000  90.030000 ;
      RECT 17.845000  94.125000 57.410000  94.275000 ;
      RECT 17.845000  94.125000 57.410000  94.275000 ;
      RECT 17.995000  89.730000 57.260000  89.880000 ;
      RECT 17.995000  93.975000 57.260000  94.125000 ;
      RECT 17.995000  93.975000 57.260000  94.125000 ;
      RECT 18.145000  89.580000 57.110000  89.730000 ;
      RECT 18.145000  93.825000 57.110000  93.975000 ;
      RECT 18.145000  93.825000 57.110000  93.975000 ;
      RECT 18.295000  89.430000 56.960000  89.580000 ;
      RECT 18.295000  93.675000 56.960000  93.825000 ;
      RECT 18.295000  93.675000 56.960000  93.825000 ;
      RECT 18.445000  89.280000 56.810000  89.430000 ;
      RECT 18.445000  93.525000 56.810000  93.675000 ;
      RECT 18.445000  93.525000 56.810000  93.675000 ;
      RECT 18.595000  89.130000 56.660000  89.280000 ;
      RECT 18.595000  93.375000 56.660000  93.525000 ;
      RECT 18.595000  93.375000 56.660000  93.525000 ;
      RECT 18.745000  88.980000 56.510000  89.130000 ;
      RECT 18.745000  93.225000 56.510000  93.375000 ;
      RECT 18.745000  93.225000 56.510000  93.375000 ;
      RECT 18.895000  88.830000 56.360000  88.980000 ;
      RECT 18.895000  93.075000 56.360000  93.225000 ;
      RECT 18.895000  93.075000 56.360000  93.225000 ;
      RECT 19.045000  88.680000 56.210000  88.830000 ;
      RECT 19.045000  92.925000 56.210000  93.075000 ;
      RECT 19.045000  92.925000 56.210000  93.075000 ;
      RECT 19.195000  88.530000 56.060000  88.680000 ;
      RECT 19.195000  92.775000 56.060000  92.925000 ;
      RECT 19.195000  92.775000 56.060000  92.925000 ;
      RECT 19.345000  88.380000 55.910000  88.530000 ;
      RECT 19.345000  92.625000 55.910000  92.775000 ;
      RECT 19.345000  92.625000 55.910000  92.775000 ;
      RECT 19.495000  88.230000 55.760000  88.380000 ;
      RECT 19.495000  92.475000 55.760000  92.625000 ;
      RECT 19.495000  92.475000 55.760000  92.625000 ;
      RECT 19.645000  88.080000 55.610000  88.230000 ;
      RECT 19.645000  92.325000 55.610000  92.475000 ;
      RECT 19.645000  92.325000 55.610000  92.475000 ;
      RECT 19.795000  87.930000 55.460000  88.080000 ;
      RECT 19.795000  92.175000 55.460000  92.325000 ;
      RECT 19.795000  92.175000 55.460000  92.325000 ;
      RECT 19.945000  87.780000 55.310000  87.930000 ;
      RECT 19.945000  92.025000 55.310000  92.175000 ;
      RECT 19.945000  92.025000 55.310000  92.175000 ;
      RECT 20.095000  87.630000 55.160000  87.780000 ;
      RECT 20.095000  91.875000 55.160000  92.025000 ;
      RECT 20.095000  91.875000 55.160000  92.025000 ;
      RECT 20.245000  87.480000 55.010000  87.630000 ;
      RECT 20.245000  91.725000 55.010000  91.875000 ;
      RECT 20.245000  91.725000 55.010000  91.875000 ;
      RECT 20.395000  87.330000 54.860000  87.480000 ;
      RECT 20.395000  91.575000 54.860000  91.725000 ;
      RECT 20.395000  91.575000 54.860000  91.725000 ;
      RECT 20.545000  87.180000 54.710000  87.330000 ;
      RECT 20.545000  91.425000 54.710000  91.575000 ;
      RECT 20.545000  91.425000 54.710000  91.575000 ;
      RECT 20.695000  87.030000 54.560000  87.180000 ;
      RECT 20.695000  91.275000 54.560000  91.425000 ;
      RECT 20.695000  91.275000 54.560000  91.425000 ;
      RECT 20.845000  86.880000 54.410000  87.030000 ;
      RECT 20.845000  91.125000 54.410000  91.275000 ;
      RECT 20.845000  91.125000 54.410000  91.275000 ;
      RECT 20.995000  86.730000 54.260000  86.880000 ;
      RECT 20.995000  90.975000 54.260000  91.125000 ;
      RECT 20.995000  90.975000 54.260000  91.125000 ;
      RECT 21.145000  86.580000 54.110000  86.730000 ;
      RECT 21.145000  90.825000 54.110000  90.975000 ;
      RECT 21.145000  90.825000 54.110000  90.975000 ;
      RECT 21.295000  86.430000 53.960000  86.580000 ;
      RECT 21.295000  90.675000 53.960000  90.825000 ;
      RECT 21.295000  90.675000 53.960000  90.825000 ;
      RECT 21.445000  86.280000 53.810000  86.430000 ;
      RECT 21.445000  90.525000 53.810000  90.675000 ;
      RECT 21.445000  90.525000 53.810000  90.675000 ;
      RECT 21.595000  86.130000 53.660000  86.280000 ;
      RECT 21.595000  90.375000 53.660000  90.525000 ;
      RECT 21.595000  90.375000 53.660000  90.525000 ;
      RECT 21.745000  85.980000 53.510000  86.130000 ;
      RECT 21.745000  90.225000 53.510000  90.375000 ;
      RECT 21.745000  90.225000 53.510000  90.375000 ;
      RECT 21.895000  85.830000 53.360000  85.980000 ;
      RECT 21.895000  90.075000 53.360000  90.225000 ;
      RECT 21.895000  90.075000 53.360000  90.225000 ;
      RECT 22.045000  85.680000 53.210000  85.830000 ;
      RECT 22.045000  89.925000 53.210000  90.075000 ;
      RECT 22.045000  89.925000 53.210000  90.075000 ;
      RECT 22.195000  85.530000 53.060000  85.680000 ;
      RECT 22.195000  89.775000 53.060000  89.925000 ;
      RECT 22.195000  89.775000 53.060000  89.925000 ;
      RECT 22.345000  85.380000 52.910000  85.530000 ;
      RECT 22.345000  89.625000 52.910000  89.775000 ;
      RECT 22.345000  89.625000 52.910000  89.775000 ;
      RECT 22.495000  85.230000 52.760000  85.380000 ;
      RECT 22.495000  89.475000 52.760000  89.625000 ;
      RECT 22.495000  89.475000 52.760000  89.625000 ;
      RECT 22.645000  85.080000 52.610000  85.230000 ;
      RECT 22.645000  89.325000 52.610000  89.475000 ;
      RECT 22.645000  89.325000 52.610000  89.475000 ;
      RECT 22.795000  84.930000 52.460000  85.080000 ;
      RECT 22.795000  89.175000 52.460000  89.325000 ;
      RECT 22.795000  89.175000 52.460000  89.325000 ;
      RECT 22.945000  84.780000 52.310000  84.930000 ;
      RECT 22.945000  89.025000 52.310000  89.175000 ;
      RECT 22.945000  89.025000 52.310000  89.175000 ;
      RECT 23.095000  84.630000 52.160000  84.780000 ;
      RECT 23.095000  88.875000 52.160000  89.025000 ;
      RECT 23.095000  88.875000 52.160000  89.025000 ;
      RECT 23.245000  84.480000 52.010000  84.630000 ;
      RECT 23.245000  88.725000 52.010000  88.875000 ;
      RECT 23.245000  88.725000 52.010000  88.875000 ;
      RECT 23.395000  84.330000 51.860000  84.480000 ;
      RECT 23.395000  88.575000 51.860000  88.725000 ;
      RECT 23.395000  88.575000 51.860000  88.725000 ;
      RECT 23.545000  84.180000 51.710000  84.330000 ;
      RECT 23.545000  88.425000 51.710000  88.575000 ;
      RECT 23.545000  88.425000 51.710000  88.575000 ;
      RECT 23.695000  84.030000 51.560000  84.180000 ;
      RECT 23.695000  88.275000 51.560000  88.425000 ;
      RECT 23.695000  88.275000 51.560000  88.425000 ;
      RECT 23.845000  83.880000 51.410000  84.030000 ;
      RECT 23.845000  88.125000 51.410000  88.275000 ;
      RECT 23.845000  88.125000 51.410000  88.275000 ;
      RECT 23.995000  83.730000 51.260000  83.880000 ;
      RECT 23.995000  87.975000 51.260000  88.125000 ;
      RECT 23.995000  87.975000 51.260000  88.125000 ;
      RECT 24.145000  83.580000 51.110000  83.730000 ;
      RECT 24.145000  87.825000 51.110000  87.975000 ;
      RECT 24.145000  87.825000 51.110000  87.975000 ;
      RECT 24.295000  83.430000 50.960000  83.580000 ;
      RECT 24.295000  87.675000 50.960000  87.825000 ;
      RECT 24.295000  87.675000 50.960000  87.825000 ;
      RECT 24.445000  83.280000 50.810000  83.430000 ;
      RECT 24.445000  87.525000 50.810000  87.675000 ;
      RECT 24.445000  87.525000 50.810000  87.675000 ;
      RECT 24.595000  83.130000 50.660000  83.280000 ;
      RECT 24.595000  87.375000 50.660000  87.525000 ;
      RECT 24.595000  87.375000 50.660000  87.525000 ;
      RECT 24.745000  82.980000 50.510000  83.130000 ;
      RECT 24.745000  87.225000 50.510000  87.375000 ;
      RECT 24.745000  87.225000 50.510000  87.375000 ;
      RECT 24.895000  66.930000 50.360000 198.000000 ;
      RECT 24.895000  82.830000 50.360000  82.980000 ;
      RECT 24.895000  87.075000 50.360000  87.225000 ;
      RECT 24.895000  87.075000 50.360000  87.225000 ;
      RECT 24.900000   0.000000 50.355000 198.000000 ;
      RECT 24.900000   0.000000 50.355000 198.000000 ;
      RECT 25.045000  86.925000 50.210000  87.075000 ;
      RECT 25.045000  86.925000 50.210000  87.075000 ;
      RECT 25.195000  86.775000 50.060000  86.925000 ;
      RECT 25.195000  86.775000 50.060000  86.925000 ;
      RECT 25.345000  86.625000 49.910000  86.775000 ;
      RECT 25.345000  86.625000 49.910000  86.775000 ;
      RECT 25.495000  86.475000 49.760000  86.625000 ;
      RECT 25.495000  86.475000 49.760000  86.625000 ;
      RECT 25.645000  86.325000 49.610000  86.475000 ;
      RECT 25.645000  86.325000 49.610000  86.475000 ;
      RECT 25.795000  86.175000 49.460000  86.325000 ;
      RECT 25.795000  86.175000 49.460000  86.325000 ;
      RECT 25.945000  86.025000 49.310000  86.175000 ;
      RECT 25.945000  86.025000 49.310000  86.175000 ;
      RECT 26.095000  85.875000 49.160000  86.025000 ;
      RECT 26.095000  85.875000 49.160000  86.025000 ;
      RECT 26.245000  85.725000 49.010000  85.875000 ;
      RECT 26.245000  85.725000 49.010000  85.875000 ;
      RECT 26.395000  85.575000 48.860000  85.725000 ;
      RECT 26.395000  85.575000 48.860000  85.725000 ;
      RECT 26.545000  85.425000 48.710000  85.575000 ;
      RECT 26.545000  85.425000 48.710000  85.575000 ;
      RECT 26.695000  85.275000 48.560000  85.425000 ;
      RECT 26.695000  85.275000 48.560000  85.425000 ;
      RECT 26.845000  85.125000 48.410000  85.275000 ;
      RECT 26.845000  85.125000 48.410000  85.275000 ;
      RECT 26.995000  84.975000 48.260000  85.125000 ;
      RECT 26.995000  84.975000 48.260000  85.125000 ;
      RECT 27.145000  84.825000 48.110000  84.975000 ;
      RECT 27.145000  84.825000 48.110000  84.975000 ;
      RECT 27.295000  84.675000 47.960000  84.825000 ;
      RECT 27.295000  84.675000 47.960000  84.825000 ;
      RECT 27.445000  84.525000 47.810000  84.675000 ;
      RECT 27.445000  84.525000 47.810000  84.675000 ;
      RECT 27.595000  84.375000 47.660000  84.525000 ;
      RECT 27.595000  84.375000 47.660000  84.525000 ;
      RECT 27.745000  84.225000 47.510000  84.375000 ;
      RECT 27.745000  84.225000 47.510000  84.375000 ;
      RECT 27.895000  69.930000 47.360000  84.075000 ;
      RECT 27.895000  84.075000 47.360000  84.225000 ;
      RECT 27.895000  84.075000 47.360000  84.225000 ;
      RECT 27.900000  14.390000 47.355000  25.830000 ;
      RECT 27.900000  58.690000 47.355000  69.930000 ;
      RECT 50.355000   0.000000 75.000000   3.005000 ;
      RECT 50.355000  14.385000 75.000000  17.390000 ;
      RECT 50.355000  22.830000 75.000000  25.835000 ;
      RECT 50.355000  58.685000 75.000000  61.690000 ;
      RECT 50.360000  66.930000 75.000000  67.635000 ;
      RECT 50.360000 194.995000 75.000000 198.000000 ;
      RECT 56.645000  93.360000 75.000000  96.365000 ;
      RECT 71.995000   3.005000 75.000000  14.385000 ;
      RECT 71.995000  25.835000 75.000000  58.685000 ;
      RECT 71.995000  96.365000 75.000000 194.995000 ;
    LAYER met4 ;
      RECT  0.000000   5.885000 75.000000   6.485000 ;
      RECT  0.000000  11.935000  1.365000  12.535000 ;
      RECT  0.000000  16.785000  1.365000  17.385000 ;
      RECT  0.000000  22.835000  1.670000  23.435000 ;
      RECT  0.000000  28.885000  1.670000  29.485000 ;
      RECT  0.000000  33.735000  1.670000  34.335000 ;
      RECT  0.000000  38.585000  1.670000  39.185000 ;
      RECT  0.000000  44.635000  1.670000  45.335000 ;
      RECT  0.000000  55.135000  1.670000  55.835000 ;
      RECT  0.000000  61.085000  1.670000  61.685000 ;
      RECT  0.000000  66.935000 75.000000  67.635000 ;
      RECT  0.000000  93.400000 75.000000 173.385000 ;
      RECT  1.365000  11.935000 73.635000  17.385000 ;
      RECT  1.670000   0.000000 73.330000   5.885000 ;
      RECT  1.670000   6.485000 73.330000  11.935000 ;
      RECT  1.670000  22.835000 73.330000  61.685000 ;
      RECT  1.670000  67.635000 73.330000  67.660000 ;
      RECT  1.670000  93.360000 60.750000  93.365000 ;
      RECT  1.670000  93.360000 60.750000 173.385000 ;
      RECT  1.670000  93.360000 60.750000 173.385000 ;
      RECT  1.670000  93.360000 60.750000 173.385000 ;
      RECT  1.670000  93.360000 60.750000 173.385000 ;
      RECT  1.670000  93.360000 60.750000 173.385000 ;
      RECT  1.670000  93.365000 73.330000  93.400000 ;
      RECT  1.670000  93.365000 73.330000 173.385000 ;
      RECT  1.670000  93.365000 73.330000 173.385000 ;
      RECT  1.670000  93.365000 73.330000 173.385000 ;
      RECT  1.670000  93.365000 73.330000 173.385000 ;
      RECT  1.670000  93.365000 73.330000 173.385000 ;
      RECT  1.670000 173.385000 73.330000 198.000000 ;
      RECT 14.505000  92.110000 60.750000  93.360000 ;
      RECT 14.505000  92.110000 60.750000 173.385000 ;
      RECT 14.505000  92.110000 60.750000 173.385000 ;
      RECT 14.505000  92.110000 60.750000 173.385000 ;
      RECT 14.505000  92.110000 60.750000 173.385000 ;
      RECT 14.505000  92.110000 60.750000 173.385000 ;
      RECT 15.765000  91.220000 59.490000  92.110000 ;
      RECT 16.650000  89.930000 58.605000  91.220000 ;
      RECT 17.925000  88.540000 57.330000  89.930000 ;
      RECT 19.255000  87.415000 56.000000  88.540000 ;
      RECT 20.465000  85.990000 54.790000  87.415000 ;
      RECT 21.850000  84.685000 53.405000  85.990000 ;
      RECT 21.850000  84.685000 53.405000  88.540000 ;
      RECT 23.170000  83.025000 52.085000  84.685000 ;
      RECT 23.170000  83.025000 52.085000  87.415000 ;
      RECT 24.875000  17.385000 50.380000  22.835000 ;
      RECT 24.875000  61.685000 50.380000  66.935000 ;
      RECT 24.900000  67.660000 50.355000  85.990000 ;
      RECT 24.900000  67.660000 50.355000  85.990000 ;
      RECT 24.900000  67.660000 50.355000  85.990000 ;
      RECT 73.330000  22.835000 75.000000  23.435000 ;
      RECT 73.330000  28.885000 75.000000  29.485000 ;
      RECT 73.330000  33.735000 75.000000  34.335000 ;
      RECT 73.330000  38.585000 75.000000  39.185000 ;
      RECT 73.330000  44.635000 75.000000  45.335000 ;
      RECT 73.330000  55.135000 75.000000  55.835000 ;
      RECT 73.330000  61.085000 75.000000  61.685000 ;
      RECT 73.635000  11.935000 75.000000  12.535000 ;
      RECT 73.635000  16.785000 75.000000  17.385000 ;
    LAYER met5 ;
      RECT 0.000000  93.785000 75.000000 172.985000 ;
      RECT 1.765000  12.235000 73.235000  17.085000 ;
      RECT 2.070000   0.000000 72.930000  12.235000 ;
      RECT 2.070000  17.085000 72.930000  93.785000 ;
      RECT 2.070000 172.985000 72.930000 198.000000 ;
  END
END sky130_fd_io__overlay_vddio_lvc
END LIBRARY
