# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__overlay_vssd_hvc
  CLASS BLOCK ;
  FOREIGN sky130_fd_io__overlay_vssd_hvc ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  75.00000 BY  200.0000 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 1.000000 41.600000 1.320000 41.920000 ;
      LAYER met4 ;
        RECT 1.000000 41.600000 1.320000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000000 42.030000 1.320000 42.350000 ;
      LAYER met4 ;
        RECT 1.000000 42.030000 1.320000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000000 42.460000 1.320000 42.780000 ;
      LAYER met4 ;
        RECT 1.000000 42.460000 1.320000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000000 42.890000 1.320000 43.210000 ;
      LAYER met4 ;
        RECT 1.000000 42.890000 1.320000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000000 43.320000 1.320000 43.640000 ;
      LAYER met4 ;
        RECT 1.000000 43.320000 1.320000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000000 43.750000 1.320000 44.070000 ;
      LAYER met4 ;
        RECT 1.000000 43.750000 1.320000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000000 44.180000 1.320000 44.500000 ;
      LAYER met4 ;
        RECT 1.000000 44.180000 1.320000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000000 44.610000 1.320000 44.930000 ;
      LAYER met4 ;
        RECT 1.000000 44.610000 1.320000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000000 45.040000 1.320000 45.360000 ;
      LAYER met4 ;
        RECT 1.000000 45.040000 1.320000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000000 45.470000 1.320000 45.790000 ;
      LAYER met4 ;
        RECT 1.000000 45.470000 1.320000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000000 45.900000 1.320000 46.220000 ;
      LAYER met4 ;
        RECT 1.000000 45.900000 1.320000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405000 41.600000 1.725000 41.920000 ;
      LAYER met4 ;
        RECT 1.405000 41.600000 1.725000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405000 42.030000 1.725000 42.350000 ;
      LAYER met4 ;
        RECT 1.405000 42.030000 1.725000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405000 42.460000 1.725000 42.780000 ;
      LAYER met4 ;
        RECT 1.405000 42.460000 1.725000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405000 42.890000 1.725000 43.210000 ;
      LAYER met4 ;
        RECT 1.405000 42.890000 1.725000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405000 43.320000 1.725000 43.640000 ;
      LAYER met4 ;
        RECT 1.405000 43.320000 1.725000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405000 43.750000 1.725000 44.070000 ;
      LAYER met4 ;
        RECT 1.405000 43.750000 1.725000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405000 44.180000 1.725000 44.500000 ;
      LAYER met4 ;
        RECT 1.405000 44.180000 1.725000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405000 44.610000 1.725000 44.930000 ;
      LAYER met4 ;
        RECT 1.405000 44.610000 1.725000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405000 45.040000 1.725000 45.360000 ;
      LAYER met4 ;
        RECT 1.405000 45.040000 1.725000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405000 45.470000 1.725000 45.790000 ;
      LAYER met4 ;
        RECT 1.405000 45.470000 1.725000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405000 45.900000 1.725000 46.220000 ;
      LAYER met4 ;
        RECT 1.405000 45.900000 1.725000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810000 41.600000 2.130000 41.920000 ;
      LAYER met4 ;
        RECT 1.810000 41.600000 2.130000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810000 42.030000 2.130000 42.350000 ;
      LAYER met4 ;
        RECT 1.810000 42.030000 2.130000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810000 42.460000 2.130000 42.780000 ;
      LAYER met4 ;
        RECT 1.810000 42.460000 2.130000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810000 42.890000 2.130000 43.210000 ;
      LAYER met4 ;
        RECT 1.810000 42.890000 2.130000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810000 43.320000 2.130000 43.640000 ;
      LAYER met4 ;
        RECT 1.810000 43.320000 2.130000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810000 43.750000 2.130000 44.070000 ;
      LAYER met4 ;
        RECT 1.810000 43.750000 2.130000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810000 44.180000 2.130000 44.500000 ;
      LAYER met4 ;
        RECT 1.810000 44.180000 2.130000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810000 44.610000 2.130000 44.930000 ;
      LAYER met4 ;
        RECT 1.810000 44.610000 2.130000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810000 45.040000 2.130000 45.360000 ;
      LAYER met4 ;
        RECT 1.810000 45.040000 2.130000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810000 45.470000 2.130000 45.790000 ;
      LAYER met4 ;
        RECT 1.810000 45.470000 2.130000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810000 45.900000 2.130000 46.220000 ;
      LAYER met4 ;
        RECT 1.810000 45.900000 2.130000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315000 41.600000 10.635000 41.920000 ;
      LAYER met4 ;
        RECT 10.315000 41.600000 10.635000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315000 42.030000 10.635000 42.350000 ;
      LAYER met4 ;
        RECT 10.315000 42.030000 10.635000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315000 42.460000 10.635000 42.780000 ;
      LAYER met4 ;
        RECT 10.315000 42.460000 10.635000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315000 42.890000 10.635000 43.210000 ;
      LAYER met4 ;
        RECT 10.315000 42.890000 10.635000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315000 43.320000 10.635000 43.640000 ;
      LAYER met4 ;
        RECT 10.315000 43.320000 10.635000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315000 43.750000 10.635000 44.070000 ;
      LAYER met4 ;
        RECT 10.315000 43.750000 10.635000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315000 44.180000 10.635000 44.500000 ;
      LAYER met4 ;
        RECT 10.315000 44.180000 10.635000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315000 44.610000 10.635000 44.930000 ;
      LAYER met4 ;
        RECT 10.315000 44.610000 10.635000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315000 45.040000 10.635000 45.360000 ;
      LAYER met4 ;
        RECT 10.315000 45.040000 10.635000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315000 45.470000 10.635000 45.790000 ;
      LAYER met4 ;
        RECT 10.315000 45.470000 10.635000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315000 45.900000 10.635000 46.220000 ;
      LAYER met4 ;
        RECT 10.315000 45.900000 10.635000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720000 41.600000 11.040000 41.920000 ;
      LAYER met4 ;
        RECT 10.720000 41.600000 11.040000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720000 42.030000 11.040000 42.350000 ;
      LAYER met4 ;
        RECT 10.720000 42.030000 11.040000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720000 42.460000 11.040000 42.780000 ;
      LAYER met4 ;
        RECT 10.720000 42.460000 11.040000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720000 42.890000 11.040000 43.210000 ;
      LAYER met4 ;
        RECT 10.720000 42.890000 11.040000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720000 43.320000 11.040000 43.640000 ;
      LAYER met4 ;
        RECT 10.720000 43.320000 11.040000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720000 43.750000 11.040000 44.070000 ;
      LAYER met4 ;
        RECT 10.720000 43.750000 11.040000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720000 44.180000 11.040000 44.500000 ;
      LAYER met4 ;
        RECT 10.720000 44.180000 11.040000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720000 44.610000 11.040000 44.930000 ;
      LAYER met4 ;
        RECT 10.720000 44.610000 11.040000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720000 45.040000 11.040000 45.360000 ;
      LAYER met4 ;
        RECT 10.720000 45.040000 11.040000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720000 45.470000 11.040000 45.790000 ;
      LAYER met4 ;
        RECT 10.720000 45.470000 11.040000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720000 45.900000 11.040000 46.220000 ;
      LAYER met4 ;
        RECT 10.720000 45.900000 11.040000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125000 41.600000 11.445000 41.920000 ;
      LAYER met4 ;
        RECT 11.125000 41.600000 11.445000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125000 42.030000 11.445000 42.350000 ;
      LAYER met4 ;
        RECT 11.125000 42.030000 11.445000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125000 42.460000 11.445000 42.780000 ;
      LAYER met4 ;
        RECT 11.125000 42.460000 11.445000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125000 42.890000 11.445000 43.210000 ;
      LAYER met4 ;
        RECT 11.125000 42.890000 11.445000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125000 43.320000 11.445000 43.640000 ;
      LAYER met4 ;
        RECT 11.125000 43.320000 11.445000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125000 43.750000 11.445000 44.070000 ;
      LAYER met4 ;
        RECT 11.125000 43.750000 11.445000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125000 44.180000 11.445000 44.500000 ;
      LAYER met4 ;
        RECT 11.125000 44.180000 11.445000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125000 44.610000 11.445000 44.930000 ;
      LAYER met4 ;
        RECT 11.125000 44.610000 11.445000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125000 45.040000 11.445000 45.360000 ;
      LAYER met4 ;
        RECT 11.125000 45.040000 11.445000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125000 45.470000 11.445000 45.790000 ;
      LAYER met4 ;
        RECT 11.125000 45.470000 11.445000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125000 45.900000 11.445000 46.220000 ;
      LAYER met4 ;
        RECT 11.125000 45.900000 11.445000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530000 41.600000 11.850000 41.920000 ;
      LAYER met4 ;
        RECT 11.530000 41.600000 11.850000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530000 42.030000 11.850000 42.350000 ;
      LAYER met4 ;
        RECT 11.530000 42.030000 11.850000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530000 42.460000 11.850000 42.780000 ;
      LAYER met4 ;
        RECT 11.530000 42.460000 11.850000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530000 42.890000 11.850000 43.210000 ;
      LAYER met4 ;
        RECT 11.530000 42.890000 11.850000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530000 43.320000 11.850000 43.640000 ;
      LAYER met4 ;
        RECT 11.530000 43.320000 11.850000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530000 43.750000 11.850000 44.070000 ;
      LAYER met4 ;
        RECT 11.530000 43.750000 11.850000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530000 44.180000 11.850000 44.500000 ;
      LAYER met4 ;
        RECT 11.530000 44.180000 11.850000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530000 44.610000 11.850000 44.930000 ;
      LAYER met4 ;
        RECT 11.530000 44.610000 11.850000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530000 45.040000 11.850000 45.360000 ;
      LAYER met4 ;
        RECT 11.530000 45.040000 11.850000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530000 45.470000 11.850000 45.790000 ;
      LAYER met4 ;
        RECT 11.530000 45.470000 11.850000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530000 45.900000 11.850000 46.220000 ;
      LAYER met4 ;
        RECT 11.530000 45.900000 11.850000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935000 41.600000 12.255000 41.920000 ;
      LAYER met4 ;
        RECT 11.935000 41.600000 12.255000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935000 42.030000 12.255000 42.350000 ;
      LAYER met4 ;
        RECT 11.935000 42.030000 12.255000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935000 42.460000 12.255000 42.780000 ;
      LAYER met4 ;
        RECT 11.935000 42.460000 12.255000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935000 42.890000 12.255000 43.210000 ;
      LAYER met4 ;
        RECT 11.935000 42.890000 12.255000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935000 43.320000 12.255000 43.640000 ;
      LAYER met4 ;
        RECT 11.935000 43.320000 12.255000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935000 43.750000 12.255000 44.070000 ;
      LAYER met4 ;
        RECT 11.935000 43.750000 12.255000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935000 44.180000 12.255000 44.500000 ;
      LAYER met4 ;
        RECT 11.935000 44.180000 12.255000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935000 44.610000 12.255000 44.930000 ;
      LAYER met4 ;
        RECT 11.935000 44.610000 12.255000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935000 45.040000 12.255000 45.360000 ;
      LAYER met4 ;
        RECT 11.935000 45.040000 12.255000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935000 45.470000 12.255000 45.790000 ;
      LAYER met4 ;
        RECT 11.935000 45.470000 12.255000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935000 45.900000 12.255000 46.220000 ;
      LAYER met4 ;
        RECT 11.935000 45.900000 12.255000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340000 41.600000 12.660000 41.920000 ;
      LAYER met4 ;
        RECT 12.340000 41.600000 12.660000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340000 42.030000 12.660000 42.350000 ;
      LAYER met4 ;
        RECT 12.340000 42.030000 12.660000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340000 42.460000 12.660000 42.780000 ;
      LAYER met4 ;
        RECT 12.340000 42.460000 12.660000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340000 42.890000 12.660000 43.210000 ;
      LAYER met4 ;
        RECT 12.340000 42.890000 12.660000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340000 43.320000 12.660000 43.640000 ;
      LAYER met4 ;
        RECT 12.340000 43.320000 12.660000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340000 43.750000 12.660000 44.070000 ;
      LAYER met4 ;
        RECT 12.340000 43.750000 12.660000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340000 44.180000 12.660000 44.500000 ;
      LAYER met4 ;
        RECT 12.340000 44.180000 12.660000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340000 44.610000 12.660000 44.930000 ;
      LAYER met4 ;
        RECT 12.340000 44.610000 12.660000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340000 45.040000 12.660000 45.360000 ;
      LAYER met4 ;
        RECT 12.340000 45.040000 12.660000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340000 45.470000 12.660000 45.790000 ;
      LAYER met4 ;
        RECT 12.340000 45.470000 12.660000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340000 45.900000 12.660000 46.220000 ;
      LAYER met4 ;
        RECT 12.340000 45.900000 12.660000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745000 41.600000 13.065000 41.920000 ;
      LAYER met4 ;
        RECT 12.745000 41.600000 13.065000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745000 42.030000 13.065000 42.350000 ;
      LAYER met4 ;
        RECT 12.745000 42.030000 13.065000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745000 42.460000 13.065000 42.780000 ;
      LAYER met4 ;
        RECT 12.745000 42.460000 13.065000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745000 42.890000 13.065000 43.210000 ;
      LAYER met4 ;
        RECT 12.745000 42.890000 13.065000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745000 43.320000 13.065000 43.640000 ;
      LAYER met4 ;
        RECT 12.745000 43.320000 13.065000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745000 43.750000 13.065000 44.070000 ;
      LAYER met4 ;
        RECT 12.745000 43.750000 13.065000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745000 44.180000 13.065000 44.500000 ;
      LAYER met4 ;
        RECT 12.745000 44.180000 13.065000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745000 44.610000 13.065000 44.930000 ;
      LAYER met4 ;
        RECT 12.745000 44.610000 13.065000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745000 45.040000 13.065000 45.360000 ;
      LAYER met4 ;
        RECT 12.745000 45.040000 13.065000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745000 45.470000 13.065000 45.790000 ;
      LAYER met4 ;
        RECT 12.745000 45.470000 13.065000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745000 45.900000 13.065000 46.220000 ;
      LAYER met4 ;
        RECT 12.745000 45.900000 13.065000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150000 41.600000 13.470000 41.920000 ;
      LAYER met4 ;
        RECT 13.150000 41.600000 13.470000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150000 42.030000 13.470000 42.350000 ;
      LAYER met4 ;
        RECT 13.150000 42.030000 13.470000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150000 42.460000 13.470000 42.780000 ;
      LAYER met4 ;
        RECT 13.150000 42.460000 13.470000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150000 42.890000 13.470000 43.210000 ;
      LAYER met4 ;
        RECT 13.150000 42.890000 13.470000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150000 43.320000 13.470000 43.640000 ;
      LAYER met4 ;
        RECT 13.150000 43.320000 13.470000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150000 43.750000 13.470000 44.070000 ;
      LAYER met4 ;
        RECT 13.150000 43.750000 13.470000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150000 44.180000 13.470000 44.500000 ;
      LAYER met4 ;
        RECT 13.150000 44.180000 13.470000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150000 44.610000 13.470000 44.930000 ;
      LAYER met4 ;
        RECT 13.150000 44.610000 13.470000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150000 45.040000 13.470000 45.360000 ;
      LAYER met4 ;
        RECT 13.150000 45.040000 13.470000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150000 45.470000 13.470000 45.790000 ;
      LAYER met4 ;
        RECT 13.150000 45.470000 13.470000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150000 45.900000 13.470000 46.220000 ;
      LAYER met4 ;
        RECT 13.150000 45.900000 13.470000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555000 41.600000 13.875000 41.920000 ;
      LAYER met4 ;
        RECT 13.555000 41.600000 13.875000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555000 42.030000 13.875000 42.350000 ;
      LAYER met4 ;
        RECT 13.555000 42.030000 13.875000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555000 42.460000 13.875000 42.780000 ;
      LAYER met4 ;
        RECT 13.555000 42.460000 13.875000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555000 42.890000 13.875000 43.210000 ;
      LAYER met4 ;
        RECT 13.555000 42.890000 13.875000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555000 43.320000 13.875000 43.640000 ;
      LAYER met4 ;
        RECT 13.555000 43.320000 13.875000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555000 43.750000 13.875000 44.070000 ;
      LAYER met4 ;
        RECT 13.555000 43.750000 13.875000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555000 44.180000 13.875000 44.500000 ;
      LAYER met4 ;
        RECT 13.555000 44.180000 13.875000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555000 44.610000 13.875000 44.930000 ;
      LAYER met4 ;
        RECT 13.555000 44.610000 13.875000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555000 45.040000 13.875000 45.360000 ;
      LAYER met4 ;
        RECT 13.555000 45.040000 13.875000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555000 45.470000 13.875000 45.790000 ;
      LAYER met4 ;
        RECT 13.555000 45.470000 13.875000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555000 45.900000 13.875000 46.220000 ;
      LAYER met4 ;
        RECT 13.555000 45.900000 13.875000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960000 41.600000 14.280000 41.920000 ;
      LAYER met4 ;
        RECT 13.960000 41.600000 14.280000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960000 42.030000 14.280000 42.350000 ;
      LAYER met4 ;
        RECT 13.960000 42.030000 14.280000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960000 42.460000 14.280000 42.780000 ;
      LAYER met4 ;
        RECT 13.960000 42.460000 14.280000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960000 42.890000 14.280000 43.210000 ;
      LAYER met4 ;
        RECT 13.960000 42.890000 14.280000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960000 43.320000 14.280000 43.640000 ;
      LAYER met4 ;
        RECT 13.960000 43.320000 14.280000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960000 43.750000 14.280000 44.070000 ;
      LAYER met4 ;
        RECT 13.960000 43.750000 14.280000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960000 44.180000 14.280000 44.500000 ;
      LAYER met4 ;
        RECT 13.960000 44.180000 14.280000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960000 44.610000 14.280000 44.930000 ;
      LAYER met4 ;
        RECT 13.960000 44.610000 14.280000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960000 45.040000 14.280000 45.360000 ;
      LAYER met4 ;
        RECT 13.960000 45.040000 14.280000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960000 45.470000 14.280000 45.790000 ;
      LAYER met4 ;
        RECT 13.960000 45.470000 14.280000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960000 45.900000 14.280000 46.220000 ;
      LAYER met4 ;
        RECT 13.960000 45.900000 14.280000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365000 41.600000 14.685000 41.920000 ;
      LAYER met4 ;
        RECT 14.365000 41.600000 14.685000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365000 42.030000 14.685000 42.350000 ;
      LAYER met4 ;
        RECT 14.365000 42.030000 14.685000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365000 42.460000 14.685000 42.780000 ;
      LAYER met4 ;
        RECT 14.365000 42.460000 14.685000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365000 42.890000 14.685000 43.210000 ;
      LAYER met4 ;
        RECT 14.365000 42.890000 14.685000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365000 43.320000 14.685000 43.640000 ;
      LAYER met4 ;
        RECT 14.365000 43.320000 14.685000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365000 43.750000 14.685000 44.070000 ;
      LAYER met4 ;
        RECT 14.365000 43.750000 14.685000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365000 44.180000 14.685000 44.500000 ;
      LAYER met4 ;
        RECT 14.365000 44.180000 14.685000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365000 44.610000 14.685000 44.930000 ;
      LAYER met4 ;
        RECT 14.365000 44.610000 14.685000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365000 45.040000 14.685000 45.360000 ;
      LAYER met4 ;
        RECT 14.365000 45.040000 14.685000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365000 45.470000 14.685000 45.790000 ;
      LAYER met4 ;
        RECT 14.365000 45.470000 14.685000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365000 45.900000 14.685000 46.220000 ;
      LAYER met4 ;
        RECT 14.365000 45.900000 14.685000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770000 41.600000 15.090000 41.920000 ;
      LAYER met4 ;
        RECT 14.770000 41.600000 15.090000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770000 42.030000 15.090000 42.350000 ;
      LAYER met4 ;
        RECT 14.770000 42.030000 15.090000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770000 42.460000 15.090000 42.780000 ;
      LAYER met4 ;
        RECT 14.770000 42.460000 15.090000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770000 42.890000 15.090000 43.210000 ;
      LAYER met4 ;
        RECT 14.770000 42.890000 15.090000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770000 43.320000 15.090000 43.640000 ;
      LAYER met4 ;
        RECT 14.770000 43.320000 15.090000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770000 43.750000 15.090000 44.070000 ;
      LAYER met4 ;
        RECT 14.770000 43.750000 15.090000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770000 44.180000 15.090000 44.500000 ;
      LAYER met4 ;
        RECT 14.770000 44.180000 15.090000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770000 44.610000 15.090000 44.930000 ;
      LAYER met4 ;
        RECT 14.770000 44.610000 15.090000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770000 45.040000 15.090000 45.360000 ;
      LAYER met4 ;
        RECT 14.770000 45.040000 15.090000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770000 45.470000 15.090000 45.790000 ;
      LAYER met4 ;
        RECT 14.770000 45.470000 15.090000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770000 45.900000 15.090000 46.220000 ;
      LAYER met4 ;
        RECT 14.770000 45.900000 15.090000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175000 41.600000 15.495000 41.920000 ;
      LAYER met4 ;
        RECT 15.175000 41.600000 15.495000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175000 42.030000 15.495000 42.350000 ;
      LAYER met4 ;
        RECT 15.175000 42.030000 15.495000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175000 42.460000 15.495000 42.780000 ;
      LAYER met4 ;
        RECT 15.175000 42.460000 15.495000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175000 42.890000 15.495000 43.210000 ;
      LAYER met4 ;
        RECT 15.175000 42.890000 15.495000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175000 43.320000 15.495000 43.640000 ;
      LAYER met4 ;
        RECT 15.175000 43.320000 15.495000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175000 43.750000 15.495000 44.070000 ;
      LAYER met4 ;
        RECT 15.175000 43.750000 15.495000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175000 44.180000 15.495000 44.500000 ;
      LAYER met4 ;
        RECT 15.175000 44.180000 15.495000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175000 44.610000 15.495000 44.930000 ;
      LAYER met4 ;
        RECT 15.175000 44.610000 15.495000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175000 45.040000 15.495000 45.360000 ;
      LAYER met4 ;
        RECT 15.175000 45.040000 15.495000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175000 45.470000 15.495000 45.790000 ;
      LAYER met4 ;
        RECT 15.175000 45.470000 15.495000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175000 45.900000 15.495000 46.220000 ;
      LAYER met4 ;
        RECT 15.175000 45.900000 15.495000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580000 41.600000 15.900000 41.920000 ;
      LAYER met4 ;
        RECT 15.580000 41.600000 15.900000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580000 42.030000 15.900000 42.350000 ;
      LAYER met4 ;
        RECT 15.580000 42.030000 15.900000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580000 42.460000 15.900000 42.780000 ;
      LAYER met4 ;
        RECT 15.580000 42.460000 15.900000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580000 42.890000 15.900000 43.210000 ;
      LAYER met4 ;
        RECT 15.580000 42.890000 15.900000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580000 43.320000 15.900000 43.640000 ;
      LAYER met4 ;
        RECT 15.580000 43.320000 15.900000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580000 43.750000 15.900000 44.070000 ;
      LAYER met4 ;
        RECT 15.580000 43.750000 15.900000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580000 44.180000 15.900000 44.500000 ;
      LAYER met4 ;
        RECT 15.580000 44.180000 15.900000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580000 44.610000 15.900000 44.930000 ;
      LAYER met4 ;
        RECT 15.580000 44.610000 15.900000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580000 45.040000 15.900000 45.360000 ;
      LAYER met4 ;
        RECT 15.580000 45.040000 15.900000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580000 45.470000 15.900000 45.790000 ;
      LAYER met4 ;
        RECT 15.580000 45.470000 15.900000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580000 45.900000 15.900000 46.220000 ;
      LAYER met4 ;
        RECT 15.580000 45.900000 15.900000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 41.600000 16.305000 41.920000 ;
      LAYER met4 ;
        RECT 15.985000 41.600000 16.305000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 42.030000 16.305000 42.350000 ;
      LAYER met4 ;
        RECT 15.985000 42.030000 16.305000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 42.460000 16.305000 42.780000 ;
      LAYER met4 ;
        RECT 15.985000 42.460000 16.305000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 42.890000 16.305000 43.210000 ;
      LAYER met4 ;
        RECT 15.985000 42.890000 16.305000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 43.320000 16.305000 43.640000 ;
      LAYER met4 ;
        RECT 15.985000 43.320000 16.305000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 43.750000 16.305000 44.070000 ;
      LAYER met4 ;
        RECT 15.985000 43.750000 16.305000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 44.180000 16.305000 44.500000 ;
      LAYER met4 ;
        RECT 15.985000 44.180000 16.305000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 44.610000 16.305000 44.930000 ;
      LAYER met4 ;
        RECT 15.985000 44.610000 16.305000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 45.040000 16.305000 45.360000 ;
      LAYER met4 ;
        RECT 15.985000 45.040000 16.305000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 45.470000 16.305000 45.790000 ;
      LAYER met4 ;
        RECT 15.985000 45.470000 16.305000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 45.900000 16.305000 46.220000 ;
      LAYER met4 ;
        RECT 15.985000 45.900000 16.305000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390000 41.600000 16.710000 41.920000 ;
      LAYER met4 ;
        RECT 16.390000 41.600000 16.710000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390000 42.030000 16.710000 42.350000 ;
      LAYER met4 ;
        RECT 16.390000 42.030000 16.710000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390000 42.460000 16.710000 42.780000 ;
      LAYER met4 ;
        RECT 16.390000 42.460000 16.710000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390000 42.890000 16.710000 43.210000 ;
      LAYER met4 ;
        RECT 16.390000 42.890000 16.710000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390000 43.320000 16.710000 43.640000 ;
      LAYER met4 ;
        RECT 16.390000 43.320000 16.710000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390000 43.750000 16.710000 44.070000 ;
      LAYER met4 ;
        RECT 16.390000 43.750000 16.710000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390000 44.180000 16.710000 44.500000 ;
      LAYER met4 ;
        RECT 16.390000 44.180000 16.710000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390000 44.610000 16.710000 44.930000 ;
      LAYER met4 ;
        RECT 16.390000 44.610000 16.710000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390000 45.040000 16.710000 45.360000 ;
      LAYER met4 ;
        RECT 16.390000 45.040000 16.710000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390000 45.470000 16.710000 45.790000 ;
      LAYER met4 ;
        RECT 16.390000 45.470000 16.710000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390000 45.900000 16.710000 46.220000 ;
      LAYER met4 ;
        RECT 16.390000 45.900000 16.710000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795000 41.600000 17.115000 41.920000 ;
      LAYER met4 ;
        RECT 16.795000 41.600000 17.115000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795000 42.030000 17.115000 42.350000 ;
      LAYER met4 ;
        RECT 16.795000 42.030000 17.115000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795000 42.460000 17.115000 42.780000 ;
      LAYER met4 ;
        RECT 16.795000 42.460000 17.115000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795000 42.890000 17.115000 43.210000 ;
      LAYER met4 ;
        RECT 16.795000 42.890000 17.115000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795000 43.320000 17.115000 43.640000 ;
      LAYER met4 ;
        RECT 16.795000 43.320000 17.115000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795000 43.750000 17.115000 44.070000 ;
      LAYER met4 ;
        RECT 16.795000 43.750000 17.115000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795000 44.180000 17.115000 44.500000 ;
      LAYER met4 ;
        RECT 16.795000 44.180000 17.115000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795000 44.610000 17.115000 44.930000 ;
      LAYER met4 ;
        RECT 16.795000 44.610000 17.115000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795000 45.040000 17.115000 45.360000 ;
      LAYER met4 ;
        RECT 16.795000 45.040000 17.115000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795000 45.470000 17.115000 45.790000 ;
      LAYER met4 ;
        RECT 16.795000 45.470000 17.115000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795000 45.900000 17.115000 46.220000 ;
      LAYER met4 ;
        RECT 16.795000 45.900000 17.115000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200000 41.600000 17.520000 41.920000 ;
      LAYER met4 ;
        RECT 17.200000 41.600000 17.520000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200000 42.030000 17.520000 42.350000 ;
      LAYER met4 ;
        RECT 17.200000 42.030000 17.520000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200000 42.460000 17.520000 42.780000 ;
      LAYER met4 ;
        RECT 17.200000 42.460000 17.520000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200000 42.890000 17.520000 43.210000 ;
      LAYER met4 ;
        RECT 17.200000 42.890000 17.520000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200000 43.320000 17.520000 43.640000 ;
      LAYER met4 ;
        RECT 17.200000 43.320000 17.520000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200000 43.750000 17.520000 44.070000 ;
      LAYER met4 ;
        RECT 17.200000 43.750000 17.520000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200000 44.180000 17.520000 44.500000 ;
      LAYER met4 ;
        RECT 17.200000 44.180000 17.520000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200000 44.610000 17.520000 44.930000 ;
      LAYER met4 ;
        RECT 17.200000 44.610000 17.520000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200000 45.040000 17.520000 45.360000 ;
      LAYER met4 ;
        RECT 17.200000 45.040000 17.520000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200000 45.470000 17.520000 45.790000 ;
      LAYER met4 ;
        RECT 17.200000 45.470000 17.520000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200000 45.900000 17.520000 46.220000 ;
      LAYER met4 ;
        RECT 17.200000 45.900000 17.520000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605000 41.600000 17.925000 41.920000 ;
      LAYER met4 ;
        RECT 17.605000 41.600000 17.925000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605000 42.030000 17.925000 42.350000 ;
      LAYER met4 ;
        RECT 17.605000 42.030000 17.925000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605000 42.460000 17.925000 42.780000 ;
      LAYER met4 ;
        RECT 17.605000 42.460000 17.925000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605000 42.890000 17.925000 43.210000 ;
      LAYER met4 ;
        RECT 17.605000 42.890000 17.925000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605000 43.320000 17.925000 43.640000 ;
      LAYER met4 ;
        RECT 17.605000 43.320000 17.925000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605000 43.750000 17.925000 44.070000 ;
      LAYER met4 ;
        RECT 17.605000 43.750000 17.925000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605000 44.180000 17.925000 44.500000 ;
      LAYER met4 ;
        RECT 17.605000 44.180000 17.925000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605000 44.610000 17.925000 44.930000 ;
      LAYER met4 ;
        RECT 17.605000 44.610000 17.925000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605000 45.040000 17.925000 45.360000 ;
      LAYER met4 ;
        RECT 17.605000 45.040000 17.925000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605000 45.470000 17.925000 45.790000 ;
      LAYER met4 ;
        RECT 17.605000 45.470000 17.925000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605000 45.900000 17.925000 46.220000 ;
      LAYER met4 ;
        RECT 17.605000 45.900000 17.925000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010000 41.600000 18.330000 41.920000 ;
      LAYER met4 ;
        RECT 18.010000 41.600000 18.330000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010000 42.030000 18.330000 42.350000 ;
      LAYER met4 ;
        RECT 18.010000 42.030000 18.330000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010000 42.460000 18.330000 42.780000 ;
      LAYER met4 ;
        RECT 18.010000 42.460000 18.330000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010000 42.890000 18.330000 43.210000 ;
      LAYER met4 ;
        RECT 18.010000 42.890000 18.330000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010000 43.320000 18.330000 43.640000 ;
      LAYER met4 ;
        RECT 18.010000 43.320000 18.330000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010000 43.750000 18.330000 44.070000 ;
      LAYER met4 ;
        RECT 18.010000 43.750000 18.330000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010000 44.180000 18.330000 44.500000 ;
      LAYER met4 ;
        RECT 18.010000 44.180000 18.330000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010000 44.610000 18.330000 44.930000 ;
      LAYER met4 ;
        RECT 18.010000 44.610000 18.330000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010000 45.040000 18.330000 45.360000 ;
      LAYER met4 ;
        RECT 18.010000 45.040000 18.330000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010000 45.470000 18.330000 45.790000 ;
      LAYER met4 ;
        RECT 18.010000 45.470000 18.330000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010000 45.900000 18.330000 46.220000 ;
      LAYER met4 ;
        RECT 18.010000 45.900000 18.330000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415000 41.600000 18.735000 41.920000 ;
      LAYER met4 ;
        RECT 18.415000 41.600000 18.735000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415000 42.030000 18.735000 42.350000 ;
      LAYER met4 ;
        RECT 18.415000 42.030000 18.735000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415000 42.460000 18.735000 42.780000 ;
      LAYER met4 ;
        RECT 18.415000 42.460000 18.735000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415000 42.890000 18.735000 43.210000 ;
      LAYER met4 ;
        RECT 18.415000 42.890000 18.735000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415000 43.320000 18.735000 43.640000 ;
      LAYER met4 ;
        RECT 18.415000 43.320000 18.735000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415000 43.750000 18.735000 44.070000 ;
      LAYER met4 ;
        RECT 18.415000 43.750000 18.735000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415000 44.180000 18.735000 44.500000 ;
      LAYER met4 ;
        RECT 18.415000 44.180000 18.735000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415000 44.610000 18.735000 44.930000 ;
      LAYER met4 ;
        RECT 18.415000 44.610000 18.735000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415000 45.040000 18.735000 45.360000 ;
      LAYER met4 ;
        RECT 18.415000 45.040000 18.735000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415000 45.470000 18.735000 45.790000 ;
      LAYER met4 ;
        RECT 18.415000 45.470000 18.735000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415000 45.900000 18.735000 46.220000 ;
      LAYER met4 ;
        RECT 18.415000 45.900000 18.735000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820000 41.600000 19.140000 41.920000 ;
      LAYER met4 ;
        RECT 18.820000 41.600000 19.140000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820000 42.030000 19.140000 42.350000 ;
      LAYER met4 ;
        RECT 18.820000 42.030000 19.140000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820000 42.460000 19.140000 42.780000 ;
      LAYER met4 ;
        RECT 18.820000 42.460000 19.140000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820000 42.890000 19.140000 43.210000 ;
      LAYER met4 ;
        RECT 18.820000 42.890000 19.140000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820000 43.320000 19.140000 43.640000 ;
      LAYER met4 ;
        RECT 18.820000 43.320000 19.140000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820000 43.750000 19.140000 44.070000 ;
      LAYER met4 ;
        RECT 18.820000 43.750000 19.140000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820000 44.180000 19.140000 44.500000 ;
      LAYER met4 ;
        RECT 18.820000 44.180000 19.140000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820000 44.610000 19.140000 44.930000 ;
      LAYER met4 ;
        RECT 18.820000 44.610000 19.140000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820000 45.040000 19.140000 45.360000 ;
      LAYER met4 ;
        RECT 18.820000 45.040000 19.140000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820000 45.470000 19.140000 45.790000 ;
      LAYER met4 ;
        RECT 18.820000 45.470000 19.140000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820000 45.900000 19.140000 46.220000 ;
      LAYER met4 ;
        RECT 18.820000 45.900000 19.140000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225000 41.600000 19.545000 41.920000 ;
      LAYER met4 ;
        RECT 19.225000 41.600000 19.545000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225000 42.030000 19.545000 42.350000 ;
      LAYER met4 ;
        RECT 19.225000 42.030000 19.545000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225000 42.460000 19.545000 42.780000 ;
      LAYER met4 ;
        RECT 19.225000 42.460000 19.545000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225000 42.890000 19.545000 43.210000 ;
      LAYER met4 ;
        RECT 19.225000 42.890000 19.545000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225000 43.320000 19.545000 43.640000 ;
      LAYER met4 ;
        RECT 19.225000 43.320000 19.545000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225000 43.750000 19.545000 44.070000 ;
      LAYER met4 ;
        RECT 19.225000 43.750000 19.545000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225000 44.180000 19.545000 44.500000 ;
      LAYER met4 ;
        RECT 19.225000 44.180000 19.545000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225000 44.610000 19.545000 44.930000 ;
      LAYER met4 ;
        RECT 19.225000 44.610000 19.545000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225000 45.040000 19.545000 45.360000 ;
      LAYER met4 ;
        RECT 19.225000 45.040000 19.545000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225000 45.470000 19.545000 45.790000 ;
      LAYER met4 ;
        RECT 19.225000 45.470000 19.545000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225000 45.900000 19.545000 46.220000 ;
      LAYER met4 ;
        RECT 19.225000 45.900000 19.545000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630000 41.600000 19.950000 41.920000 ;
      LAYER met4 ;
        RECT 19.630000 41.600000 19.950000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630000 42.030000 19.950000 42.350000 ;
      LAYER met4 ;
        RECT 19.630000 42.030000 19.950000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630000 42.460000 19.950000 42.780000 ;
      LAYER met4 ;
        RECT 19.630000 42.460000 19.950000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630000 42.890000 19.950000 43.210000 ;
      LAYER met4 ;
        RECT 19.630000 42.890000 19.950000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630000 43.320000 19.950000 43.640000 ;
      LAYER met4 ;
        RECT 19.630000 43.320000 19.950000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630000 43.750000 19.950000 44.070000 ;
      LAYER met4 ;
        RECT 19.630000 43.750000 19.950000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630000 44.180000 19.950000 44.500000 ;
      LAYER met4 ;
        RECT 19.630000 44.180000 19.950000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630000 44.610000 19.950000 44.930000 ;
      LAYER met4 ;
        RECT 19.630000 44.610000 19.950000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630000 45.040000 19.950000 45.360000 ;
      LAYER met4 ;
        RECT 19.630000 45.040000 19.950000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630000 45.470000 19.950000 45.790000 ;
      LAYER met4 ;
        RECT 19.630000 45.470000 19.950000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630000 45.900000 19.950000 46.220000 ;
      LAYER met4 ;
        RECT 19.630000 45.900000 19.950000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 41.600000 2.535000 41.920000 ;
      LAYER met4 ;
        RECT 2.215000 41.600000 2.535000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 42.030000 2.535000 42.350000 ;
      LAYER met4 ;
        RECT 2.215000 42.030000 2.535000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 42.460000 2.535000 42.780000 ;
      LAYER met4 ;
        RECT 2.215000 42.460000 2.535000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 42.890000 2.535000 43.210000 ;
      LAYER met4 ;
        RECT 2.215000 42.890000 2.535000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 43.320000 2.535000 43.640000 ;
      LAYER met4 ;
        RECT 2.215000 43.320000 2.535000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 43.750000 2.535000 44.070000 ;
      LAYER met4 ;
        RECT 2.215000 43.750000 2.535000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 44.180000 2.535000 44.500000 ;
      LAYER met4 ;
        RECT 2.215000 44.180000 2.535000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 44.610000 2.535000 44.930000 ;
      LAYER met4 ;
        RECT 2.215000 44.610000 2.535000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 45.040000 2.535000 45.360000 ;
      LAYER met4 ;
        RECT 2.215000 45.040000 2.535000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 45.470000 2.535000 45.790000 ;
      LAYER met4 ;
        RECT 2.215000 45.470000 2.535000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 45.900000 2.535000 46.220000 ;
      LAYER met4 ;
        RECT 2.215000 45.900000 2.535000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620000 41.600000 2.940000 41.920000 ;
      LAYER met4 ;
        RECT 2.620000 41.600000 2.940000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620000 42.030000 2.940000 42.350000 ;
      LAYER met4 ;
        RECT 2.620000 42.030000 2.940000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620000 42.460000 2.940000 42.780000 ;
      LAYER met4 ;
        RECT 2.620000 42.460000 2.940000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620000 42.890000 2.940000 43.210000 ;
      LAYER met4 ;
        RECT 2.620000 42.890000 2.940000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620000 43.320000 2.940000 43.640000 ;
      LAYER met4 ;
        RECT 2.620000 43.320000 2.940000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620000 43.750000 2.940000 44.070000 ;
      LAYER met4 ;
        RECT 2.620000 43.750000 2.940000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620000 44.180000 2.940000 44.500000 ;
      LAYER met4 ;
        RECT 2.620000 44.180000 2.940000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620000 44.610000 2.940000 44.930000 ;
      LAYER met4 ;
        RECT 2.620000 44.610000 2.940000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620000 45.040000 2.940000 45.360000 ;
      LAYER met4 ;
        RECT 2.620000 45.040000 2.940000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620000 45.470000 2.940000 45.790000 ;
      LAYER met4 ;
        RECT 2.620000 45.470000 2.940000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620000 45.900000 2.940000 46.220000 ;
      LAYER met4 ;
        RECT 2.620000 45.900000 2.940000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035000 41.600000 20.355000 41.920000 ;
      LAYER met4 ;
        RECT 20.035000 41.600000 20.355000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035000 42.030000 20.355000 42.350000 ;
      LAYER met4 ;
        RECT 20.035000 42.030000 20.355000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035000 42.460000 20.355000 42.780000 ;
      LAYER met4 ;
        RECT 20.035000 42.460000 20.355000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035000 42.890000 20.355000 43.210000 ;
      LAYER met4 ;
        RECT 20.035000 42.890000 20.355000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035000 43.320000 20.355000 43.640000 ;
      LAYER met4 ;
        RECT 20.035000 43.320000 20.355000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035000 43.750000 20.355000 44.070000 ;
      LAYER met4 ;
        RECT 20.035000 43.750000 20.355000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035000 44.180000 20.355000 44.500000 ;
      LAYER met4 ;
        RECT 20.035000 44.180000 20.355000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035000 44.610000 20.355000 44.930000 ;
      LAYER met4 ;
        RECT 20.035000 44.610000 20.355000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035000 45.040000 20.355000 45.360000 ;
      LAYER met4 ;
        RECT 20.035000 45.040000 20.355000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035000 45.470000 20.355000 45.790000 ;
      LAYER met4 ;
        RECT 20.035000 45.470000 20.355000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035000 45.900000 20.355000 46.220000 ;
      LAYER met4 ;
        RECT 20.035000 45.900000 20.355000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440000 41.600000 20.760000 41.920000 ;
      LAYER met4 ;
        RECT 20.440000 41.600000 20.760000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440000 42.030000 20.760000 42.350000 ;
      LAYER met4 ;
        RECT 20.440000 42.030000 20.760000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440000 42.460000 20.760000 42.780000 ;
      LAYER met4 ;
        RECT 20.440000 42.460000 20.760000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440000 42.890000 20.760000 43.210000 ;
      LAYER met4 ;
        RECT 20.440000 42.890000 20.760000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440000 43.320000 20.760000 43.640000 ;
      LAYER met4 ;
        RECT 20.440000 43.320000 20.760000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440000 43.750000 20.760000 44.070000 ;
      LAYER met4 ;
        RECT 20.440000 43.750000 20.760000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440000 44.180000 20.760000 44.500000 ;
      LAYER met4 ;
        RECT 20.440000 44.180000 20.760000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440000 44.610000 20.760000 44.930000 ;
      LAYER met4 ;
        RECT 20.440000 44.610000 20.760000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440000 45.040000 20.760000 45.360000 ;
      LAYER met4 ;
        RECT 20.440000 45.040000 20.760000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440000 45.470000 20.760000 45.790000 ;
      LAYER met4 ;
        RECT 20.440000 45.470000 20.760000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440000 45.900000 20.760000 46.220000 ;
      LAYER met4 ;
        RECT 20.440000 45.900000 20.760000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845000 41.600000 21.165000 41.920000 ;
      LAYER met4 ;
        RECT 20.845000 41.600000 21.165000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845000 42.030000 21.165000 42.350000 ;
      LAYER met4 ;
        RECT 20.845000 42.030000 21.165000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845000 42.460000 21.165000 42.780000 ;
      LAYER met4 ;
        RECT 20.845000 42.460000 21.165000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845000 42.890000 21.165000 43.210000 ;
      LAYER met4 ;
        RECT 20.845000 42.890000 21.165000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845000 43.320000 21.165000 43.640000 ;
      LAYER met4 ;
        RECT 20.845000 43.320000 21.165000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845000 43.750000 21.165000 44.070000 ;
      LAYER met4 ;
        RECT 20.845000 43.750000 21.165000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845000 44.180000 21.165000 44.500000 ;
      LAYER met4 ;
        RECT 20.845000 44.180000 21.165000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845000 44.610000 21.165000 44.930000 ;
      LAYER met4 ;
        RECT 20.845000 44.610000 21.165000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845000 45.040000 21.165000 45.360000 ;
      LAYER met4 ;
        RECT 20.845000 45.040000 21.165000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845000 45.470000 21.165000 45.790000 ;
      LAYER met4 ;
        RECT 20.845000 45.470000 21.165000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845000 45.900000 21.165000 46.220000 ;
      LAYER met4 ;
        RECT 20.845000 45.900000 21.165000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245000 41.600000 21.565000 41.920000 ;
      LAYER met4 ;
        RECT 21.245000 41.600000 21.565000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245000 42.030000 21.565000 42.350000 ;
      LAYER met4 ;
        RECT 21.245000 42.030000 21.565000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245000 42.460000 21.565000 42.780000 ;
      LAYER met4 ;
        RECT 21.245000 42.460000 21.565000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245000 42.890000 21.565000 43.210000 ;
      LAYER met4 ;
        RECT 21.245000 42.890000 21.565000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245000 43.320000 21.565000 43.640000 ;
      LAYER met4 ;
        RECT 21.245000 43.320000 21.565000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245000 43.750000 21.565000 44.070000 ;
      LAYER met4 ;
        RECT 21.245000 43.750000 21.565000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245000 44.180000 21.565000 44.500000 ;
      LAYER met4 ;
        RECT 21.245000 44.180000 21.565000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245000 44.610000 21.565000 44.930000 ;
      LAYER met4 ;
        RECT 21.245000 44.610000 21.565000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245000 45.040000 21.565000 45.360000 ;
      LAYER met4 ;
        RECT 21.245000 45.040000 21.565000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245000 45.470000 21.565000 45.790000 ;
      LAYER met4 ;
        RECT 21.245000 45.470000 21.565000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245000 45.900000 21.565000 46.220000 ;
      LAYER met4 ;
        RECT 21.245000 45.900000 21.565000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645000 41.600000 21.965000 41.920000 ;
      LAYER met4 ;
        RECT 21.645000 41.600000 21.965000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645000 42.030000 21.965000 42.350000 ;
      LAYER met4 ;
        RECT 21.645000 42.030000 21.965000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645000 42.460000 21.965000 42.780000 ;
      LAYER met4 ;
        RECT 21.645000 42.460000 21.965000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645000 42.890000 21.965000 43.210000 ;
      LAYER met4 ;
        RECT 21.645000 42.890000 21.965000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645000 43.320000 21.965000 43.640000 ;
      LAYER met4 ;
        RECT 21.645000 43.320000 21.965000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645000 43.750000 21.965000 44.070000 ;
      LAYER met4 ;
        RECT 21.645000 43.750000 21.965000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645000 44.180000 21.965000 44.500000 ;
      LAYER met4 ;
        RECT 21.645000 44.180000 21.965000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645000 44.610000 21.965000 44.930000 ;
      LAYER met4 ;
        RECT 21.645000 44.610000 21.965000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645000 45.040000 21.965000 45.360000 ;
      LAYER met4 ;
        RECT 21.645000 45.040000 21.965000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645000 45.470000 21.965000 45.790000 ;
      LAYER met4 ;
        RECT 21.645000 45.470000 21.965000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645000 45.900000 21.965000 46.220000 ;
      LAYER met4 ;
        RECT 21.645000 45.900000 21.965000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045000 41.600000 22.365000 41.920000 ;
      LAYER met4 ;
        RECT 22.045000 41.600000 22.365000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045000 42.030000 22.365000 42.350000 ;
      LAYER met4 ;
        RECT 22.045000 42.030000 22.365000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045000 42.460000 22.365000 42.780000 ;
      LAYER met4 ;
        RECT 22.045000 42.460000 22.365000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045000 42.890000 22.365000 43.210000 ;
      LAYER met4 ;
        RECT 22.045000 42.890000 22.365000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045000 43.320000 22.365000 43.640000 ;
      LAYER met4 ;
        RECT 22.045000 43.320000 22.365000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045000 43.750000 22.365000 44.070000 ;
      LAYER met4 ;
        RECT 22.045000 43.750000 22.365000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045000 44.180000 22.365000 44.500000 ;
      LAYER met4 ;
        RECT 22.045000 44.180000 22.365000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045000 44.610000 22.365000 44.930000 ;
      LAYER met4 ;
        RECT 22.045000 44.610000 22.365000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045000 45.040000 22.365000 45.360000 ;
      LAYER met4 ;
        RECT 22.045000 45.040000 22.365000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045000 45.470000 22.365000 45.790000 ;
      LAYER met4 ;
        RECT 22.045000 45.470000 22.365000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045000 45.900000 22.365000 46.220000 ;
      LAYER met4 ;
        RECT 22.045000 45.900000 22.365000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445000 41.600000 22.765000 41.920000 ;
      LAYER met4 ;
        RECT 22.445000 41.600000 22.765000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445000 42.030000 22.765000 42.350000 ;
      LAYER met4 ;
        RECT 22.445000 42.030000 22.765000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445000 42.460000 22.765000 42.780000 ;
      LAYER met4 ;
        RECT 22.445000 42.460000 22.765000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445000 42.890000 22.765000 43.210000 ;
      LAYER met4 ;
        RECT 22.445000 42.890000 22.765000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445000 43.320000 22.765000 43.640000 ;
      LAYER met4 ;
        RECT 22.445000 43.320000 22.765000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445000 43.750000 22.765000 44.070000 ;
      LAYER met4 ;
        RECT 22.445000 43.750000 22.765000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445000 44.180000 22.765000 44.500000 ;
      LAYER met4 ;
        RECT 22.445000 44.180000 22.765000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445000 44.610000 22.765000 44.930000 ;
      LAYER met4 ;
        RECT 22.445000 44.610000 22.765000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445000 45.040000 22.765000 45.360000 ;
      LAYER met4 ;
        RECT 22.445000 45.040000 22.765000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445000 45.470000 22.765000 45.790000 ;
      LAYER met4 ;
        RECT 22.445000 45.470000 22.765000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445000 45.900000 22.765000 46.220000 ;
      LAYER met4 ;
        RECT 22.445000 45.900000 22.765000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845000 41.600000 23.165000 41.920000 ;
      LAYER met4 ;
        RECT 22.845000 41.600000 23.165000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845000 42.030000 23.165000 42.350000 ;
      LAYER met4 ;
        RECT 22.845000 42.030000 23.165000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845000 42.460000 23.165000 42.780000 ;
      LAYER met4 ;
        RECT 22.845000 42.460000 23.165000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845000 42.890000 23.165000 43.210000 ;
      LAYER met4 ;
        RECT 22.845000 42.890000 23.165000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845000 43.320000 23.165000 43.640000 ;
      LAYER met4 ;
        RECT 22.845000 43.320000 23.165000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845000 43.750000 23.165000 44.070000 ;
      LAYER met4 ;
        RECT 22.845000 43.750000 23.165000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845000 44.180000 23.165000 44.500000 ;
      LAYER met4 ;
        RECT 22.845000 44.180000 23.165000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845000 44.610000 23.165000 44.930000 ;
      LAYER met4 ;
        RECT 22.845000 44.610000 23.165000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845000 45.040000 23.165000 45.360000 ;
      LAYER met4 ;
        RECT 22.845000 45.040000 23.165000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845000 45.470000 23.165000 45.790000 ;
      LAYER met4 ;
        RECT 22.845000 45.470000 23.165000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845000 45.900000 23.165000 46.220000 ;
      LAYER met4 ;
        RECT 22.845000 45.900000 23.165000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245000 41.600000 23.565000 41.920000 ;
      LAYER met4 ;
        RECT 23.245000 41.600000 23.565000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245000 42.030000 23.565000 42.350000 ;
      LAYER met4 ;
        RECT 23.245000 42.030000 23.565000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245000 42.460000 23.565000 42.780000 ;
      LAYER met4 ;
        RECT 23.245000 42.460000 23.565000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245000 42.890000 23.565000 43.210000 ;
      LAYER met4 ;
        RECT 23.245000 42.890000 23.565000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245000 43.320000 23.565000 43.640000 ;
      LAYER met4 ;
        RECT 23.245000 43.320000 23.565000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245000 43.750000 23.565000 44.070000 ;
      LAYER met4 ;
        RECT 23.245000 43.750000 23.565000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245000 44.180000 23.565000 44.500000 ;
      LAYER met4 ;
        RECT 23.245000 44.180000 23.565000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245000 44.610000 23.565000 44.930000 ;
      LAYER met4 ;
        RECT 23.245000 44.610000 23.565000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245000 45.040000 23.565000 45.360000 ;
      LAYER met4 ;
        RECT 23.245000 45.040000 23.565000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245000 45.470000 23.565000 45.790000 ;
      LAYER met4 ;
        RECT 23.245000 45.470000 23.565000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245000 45.900000 23.565000 46.220000 ;
      LAYER met4 ;
        RECT 23.245000 45.900000 23.565000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 41.600000 23.965000 41.920000 ;
      LAYER met4 ;
        RECT 23.645000 41.600000 23.965000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 42.030000 23.965000 42.350000 ;
      LAYER met4 ;
        RECT 23.645000 42.030000 23.965000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 42.460000 23.965000 42.780000 ;
      LAYER met4 ;
        RECT 23.645000 42.460000 23.965000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 42.890000 23.965000 43.210000 ;
      LAYER met4 ;
        RECT 23.645000 42.890000 23.965000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 43.320000 23.965000 43.640000 ;
      LAYER met4 ;
        RECT 23.645000 43.320000 23.965000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 43.750000 23.965000 44.070000 ;
      LAYER met4 ;
        RECT 23.645000 43.750000 23.965000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 44.180000 23.965000 44.500000 ;
      LAYER met4 ;
        RECT 23.645000 44.180000 23.965000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 44.610000 23.965000 44.930000 ;
      LAYER met4 ;
        RECT 23.645000 44.610000 23.965000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 45.040000 23.965000 45.360000 ;
      LAYER met4 ;
        RECT 23.645000 45.040000 23.965000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 45.470000 23.965000 45.790000 ;
      LAYER met4 ;
        RECT 23.645000 45.470000 23.965000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 45.900000 23.965000 46.220000 ;
      LAYER met4 ;
        RECT 23.645000 45.900000 23.965000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 41.600000 24.365000 41.920000 ;
      LAYER met4 ;
        RECT 24.045000 41.600000 24.365000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 42.030000 24.365000 42.350000 ;
      LAYER met4 ;
        RECT 24.045000 42.030000 24.365000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 42.460000 24.365000 42.780000 ;
      LAYER met4 ;
        RECT 24.045000 42.460000 24.365000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 42.890000 24.365000 43.210000 ;
      LAYER met4 ;
        RECT 24.045000 42.890000 24.365000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 43.320000 24.365000 43.640000 ;
      LAYER met4 ;
        RECT 24.045000 43.320000 24.365000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 43.750000 24.365000 44.070000 ;
      LAYER met4 ;
        RECT 24.045000 43.750000 24.365000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 44.180000 24.365000 44.500000 ;
      LAYER met4 ;
        RECT 24.045000 44.180000 24.365000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 44.610000 24.365000 44.930000 ;
      LAYER met4 ;
        RECT 24.045000 44.610000 24.365000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 45.040000 24.365000 45.360000 ;
      LAYER met4 ;
        RECT 24.045000 45.040000 24.365000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 45.470000 24.365000 45.790000 ;
      LAYER met4 ;
        RECT 24.045000 45.470000 24.365000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 45.900000 24.365000 46.220000 ;
      LAYER met4 ;
        RECT 24.045000 45.900000 24.365000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 41.600000 3.345000 41.920000 ;
      LAYER met4 ;
        RECT 3.025000 41.600000 3.345000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 42.030000 3.345000 42.350000 ;
      LAYER met4 ;
        RECT 3.025000 42.030000 3.345000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 42.460000 3.345000 42.780000 ;
      LAYER met4 ;
        RECT 3.025000 42.460000 3.345000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 42.890000 3.345000 43.210000 ;
      LAYER met4 ;
        RECT 3.025000 42.890000 3.345000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 43.320000 3.345000 43.640000 ;
      LAYER met4 ;
        RECT 3.025000 43.320000 3.345000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 43.750000 3.345000 44.070000 ;
      LAYER met4 ;
        RECT 3.025000 43.750000 3.345000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 44.180000 3.345000 44.500000 ;
      LAYER met4 ;
        RECT 3.025000 44.180000 3.345000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 44.610000 3.345000 44.930000 ;
      LAYER met4 ;
        RECT 3.025000 44.610000 3.345000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 45.040000 3.345000 45.360000 ;
      LAYER met4 ;
        RECT 3.025000 45.040000 3.345000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 45.470000 3.345000 45.790000 ;
      LAYER met4 ;
        RECT 3.025000 45.470000 3.345000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 45.900000 3.345000 46.220000 ;
      LAYER met4 ;
        RECT 3.025000 45.900000 3.345000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430000 41.600000 3.750000 41.920000 ;
      LAYER met4 ;
        RECT 3.430000 41.600000 3.750000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430000 42.030000 3.750000 42.350000 ;
      LAYER met4 ;
        RECT 3.430000 42.030000 3.750000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430000 42.460000 3.750000 42.780000 ;
      LAYER met4 ;
        RECT 3.430000 42.460000 3.750000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430000 42.890000 3.750000 43.210000 ;
      LAYER met4 ;
        RECT 3.430000 42.890000 3.750000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430000 43.320000 3.750000 43.640000 ;
      LAYER met4 ;
        RECT 3.430000 43.320000 3.750000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430000 43.750000 3.750000 44.070000 ;
      LAYER met4 ;
        RECT 3.430000 43.750000 3.750000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430000 44.180000 3.750000 44.500000 ;
      LAYER met4 ;
        RECT 3.430000 44.180000 3.750000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430000 44.610000 3.750000 44.930000 ;
      LAYER met4 ;
        RECT 3.430000 44.610000 3.750000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430000 45.040000 3.750000 45.360000 ;
      LAYER met4 ;
        RECT 3.430000 45.040000 3.750000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430000 45.470000 3.750000 45.790000 ;
      LAYER met4 ;
        RECT 3.430000 45.470000 3.750000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430000 45.900000 3.750000 46.220000 ;
      LAYER met4 ;
        RECT 3.430000 45.900000 3.750000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835000 41.600000 4.155000 41.920000 ;
      LAYER met4 ;
        RECT 3.835000 41.600000 4.155000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835000 42.030000 4.155000 42.350000 ;
      LAYER met4 ;
        RECT 3.835000 42.030000 4.155000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835000 42.460000 4.155000 42.780000 ;
      LAYER met4 ;
        RECT 3.835000 42.460000 4.155000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835000 42.890000 4.155000 43.210000 ;
      LAYER met4 ;
        RECT 3.835000 42.890000 4.155000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835000 43.320000 4.155000 43.640000 ;
      LAYER met4 ;
        RECT 3.835000 43.320000 4.155000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835000 43.750000 4.155000 44.070000 ;
      LAYER met4 ;
        RECT 3.835000 43.750000 4.155000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835000 44.180000 4.155000 44.500000 ;
      LAYER met4 ;
        RECT 3.835000 44.180000 4.155000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835000 44.610000 4.155000 44.930000 ;
      LAYER met4 ;
        RECT 3.835000 44.610000 4.155000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835000 45.040000 4.155000 45.360000 ;
      LAYER met4 ;
        RECT 3.835000 45.040000 4.155000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835000 45.470000 4.155000 45.790000 ;
      LAYER met4 ;
        RECT 3.835000 45.470000 4.155000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835000 45.900000 4.155000 46.220000 ;
      LAYER met4 ;
        RECT 3.835000 45.900000 4.155000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240000 41.600000 4.560000 41.920000 ;
      LAYER met4 ;
        RECT 4.240000 41.600000 4.560000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240000 42.030000 4.560000 42.350000 ;
      LAYER met4 ;
        RECT 4.240000 42.030000 4.560000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240000 42.460000 4.560000 42.780000 ;
      LAYER met4 ;
        RECT 4.240000 42.460000 4.560000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240000 42.890000 4.560000 43.210000 ;
      LAYER met4 ;
        RECT 4.240000 42.890000 4.560000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240000 43.320000 4.560000 43.640000 ;
      LAYER met4 ;
        RECT 4.240000 43.320000 4.560000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240000 43.750000 4.560000 44.070000 ;
      LAYER met4 ;
        RECT 4.240000 43.750000 4.560000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240000 44.180000 4.560000 44.500000 ;
      LAYER met4 ;
        RECT 4.240000 44.180000 4.560000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240000 44.610000 4.560000 44.930000 ;
      LAYER met4 ;
        RECT 4.240000 44.610000 4.560000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240000 45.040000 4.560000 45.360000 ;
      LAYER met4 ;
        RECT 4.240000 45.040000 4.560000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240000 45.470000 4.560000 45.790000 ;
      LAYER met4 ;
        RECT 4.240000 45.470000 4.560000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240000 45.900000 4.560000 46.220000 ;
      LAYER met4 ;
        RECT 4.240000 45.900000 4.560000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645000 41.600000 4.965000 41.920000 ;
      LAYER met4 ;
        RECT 4.645000 41.600000 4.965000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645000 42.030000 4.965000 42.350000 ;
      LAYER met4 ;
        RECT 4.645000 42.030000 4.965000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645000 42.460000 4.965000 42.780000 ;
      LAYER met4 ;
        RECT 4.645000 42.460000 4.965000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645000 42.890000 4.965000 43.210000 ;
      LAYER met4 ;
        RECT 4.645000 42.890000 4.965000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645000 43.320000 4.965000 43.640000 ;
      LAYER met4 ;
        RECT 4.645000 43.320000 4.965000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645000 43.750000 4.965000 44.070000 ;
      LAYER met4 ;
        RECT 4.645000 43.750000 4.965000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645000 44.180000 4.965000 44.500000 ;
      LAYER met4 ;
        RECT 4.645000 44.180000 4.965000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645000 44.610000 4.965000 44.930000 ;
      LAYER met4 ;
        RECT 4.645000 44.610000 4.965000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645000 45.040000 4.965000 45.360000 ;
      LAYER met4 ;
        RECT 4.645000 45.040000 4.965000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645000 45.470000 4.965000 45.790000 ;
      LAYER met4 ;
        RECT 4.645000 45.470000 4.965000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645000 45.900000 4.965000 46.220000 ;
      LAYER met4 ;
        RECT 4.645000 45.900000 4.965000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050000 41.600000 5.370000 41.920000 ;
      LAYER met4 ;
        RECT 5.050000 41.600000 5.370000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050000 42.030000 5.370000 42.350000 ;
      LAYER met4 ;
        RECT 5.050000 42.030000 5.370000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050000 42.460000 5.370000 42.780000 ;
      LAYER met4 ;
        RECT 5.050000 42.460000 5.370000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050000 42.890000 5.370000 43.210000 ;
      LAYER met4 ;
        RECT 5.050000 42.890000 5.370000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050000 43.320000 5.370000 43.640000 ;
      LAYER met4 ;
        RECT 5.050000 43.320000 5.370000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050000 43.750000 5.370000 44.070000 ;
      LAYER met4 ;
        RECT 5.050000 43.750000 5.370000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050000 44.180000 5.370000 44.500000 ;
      LAYER met4 ;
        RECT 5.050000 44.180000 5.370000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050000 44.610000 5.370000 44.930000 ;
      LAYER met4 ;
        RECT 5.050000 44.610000 5.370000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050000 45.040000 5.370000 45.360000 ;
      LAYER met4 ;
        RECT 5.050000 45.040000 5.370000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050000 45.470000 5.370000 45.790000 ;
      LAYER met4 ;
        RECT 5.050000 45.470000 5.370000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050000 45.900000 5.370000 46.220000 ;
      LAYER met4 ;
        RECT 5.050000 45.900000 5.370000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455000 41.600000 5.775000 41.920000 ;
      LAYER met4 ;
        RECT 5.455000 41.600000 5.775000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455000 42.030000 5.775000 42.350000 ;
      LAYER met4 ;
        RECT 5.455000 42.030000 5.775000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455000 42.460000 5.775000 42.780000 ;
      LAYER met4 ;
        RECT 5.455000 42.460000 5.775000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455000 42.890000 5.775000 43.210000 ;
      LAYER met4 ;
        RECT 5.455000 42.890000 5.775000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455000 43.320000 5.775000 43.640000 ;
      LAYER met4 ;
        RECT 5.455000 43.320000 5.775000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455000 43.750000 5.775000 44.070000 ;
      LAYER met4 ;
        RECT 5.455000 43.750000 5.775000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455000 44.180000 5.775000 44.500000 ;
      LAYER met4 ;
        RECT 5.455000 44.180000 5.775000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455000 44.610000 5.775000 44.930000 ;
      LAYER met4 ;
        RECT 5.455000 44.610000 5.775000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455000 45.040000 5.775000 45.360000 ;
      LAYER met4 ;
        RECT 5.455000 45.040000 5.775000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455000 45.470000 5.775000 45.790000 ;
      LAYER met4 ;
        RECT 5.455000 45.470000 5.775000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455000 45.900000 5.775000 46.220000 ;
      LAYER met4 ;
        RECT 5.455000 45.900000 5.775000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860000 41.600000 6.180000 41.920000 ;
      LAYER met4 ;
        RECT 5.860000 41.600000 6.180000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860000 42.030000 6.180000 42.350000 ;
      LAYER met4 ;
        RECT 5.860000 42.030000 6.180000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860000 42.460000 6.180000 42.780000 ;
      LAYER met4 ;
        RECT 5.860000 42.460000 6.180000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860000 42.890000 6.180000 43.210000 ;
      LAYER met4 ;
        RECT 5.860000 42.890000 6.180000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860000 43.320000 6.180000 43.640000 ;
      LAYER met4 ;
        RECT 5.860000 43.320000 6.180000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860000 43.750000 6.180000 44.070000 ;
      LAYER met4 ;
        RECT 5.860000 43.750000 6.180000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860000 44.180000 6.180000 44.500000 ;
      LAYER met4 ;
        RECT 5.860000 44.180000 6.180000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860000 44.610000 6.180000 44.930000 ;
      LAYER met4 ;
        RECT 5.860000 44.610000 6.180000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860000 45.040000 6.180000 45.360000 ;
      LAYER met4 ;
        RECT 5.860000 45.040000 6.180000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860000 45.470000 6.180000 45.790000 ;
      LAYER met4 ;
        RECT 5.860000 45.470000 6.180000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860000 45.900000 6.180000 46.220000 ;
      LAYER met4 ;
        RECT 5.860000 45.900000 6.180000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 41.600000 50.740000 41.920000 ;
      LAYER met4 ;
        RECT 50.420000 41.600000 50.740000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 42.030000 50.740000 42.350000 ;
      LAYER met4 ;
        RECT 50.420000 42.030000 50.740000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 42.460000 50.740000 42.780000 ;
      LAYER met4 ;
        RECT 50.420000 42.460000 50.740000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 42.890000 50.740000 43.210000 ;
      LAYER met4 ;
        RECT 50.420000 42.890000 50.740000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 43.320000 50.740000 43.640000 ;
      LAYER met4 ;
        RECT 50.420000 43.320000 50.740000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 43.750000 50.740000 44.070000 ;
      LAYER met4 ;
        RECT 50.420000 43.750000 50.740000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 44.180000 50.740000 44.500000 ;
      LAYER met4 ;
        RECT 50.420000 44.180000 50.740000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 44.610000 50.740000 44.930000 ;
      LAYER met4 ;
        RECT 50.420000 44.610000 50.740000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 45.040000 50.740000 45.360000 ;
      LAYER met4 ;
        RECT 50.420000 45.040000 50.740000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 45.470000 50.740000 45.790000 ;
      LAYER met4 ;
        RECT 50.420000 45.470000 50.740000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 45.900000 50.740000 46.220000 ;
      LAYER met4 ;
        RECT 50.420000 45.900000 50.740000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 41.600000 51.150000 41.920000 ;
      LAYER met4 ;
        RECT 50.830000 41.600000 51.150000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 42.030000 51.150000 42.350000 ;
      LAYER met4 ;
        RECT 50.830000 42.030000 51.150000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 42.460000 51.150000 42.780000 ;
      LAYER met4 ;
        RECT 50.830000 42.460000 51.150000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 42.890000 51.150000 43.210000 ;
      LAYER met4 ;
        RECT 50.830000 42.890000 51.150000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 43.320000 51.150000 43.640000 ;
      LAYER met4 ;
        RECT 50.830000 43.320000 51.150000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 43.750000 51.150000 44.070000 ;
      LAYER met4 ;
        RECT 50.830000 43.750000 51.150000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 44.180000 51.150000 44.500000 ;
      LAYER met4 ;
        RECT 50.830000 44.180000 51.150000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 44.610000 51.150000 44.930000 ;
      LAYER met4 ;
        RECT 50.830000 44.610000 51.150000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 45.040000 51.150000 45.360000 ;
      LAYER met4 ;
        RECT 50.830000 45.040000 51.150000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 45.470000 51.150000 45.790000 ;
      LAYER met4 ;
        RECT 50.830000 45.470000 51.150000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 45.900000 51.150000 46.220000 ;
      LAYER met4 ;
        RECT 50.830000 45.900000 51.150000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 41.600000 51.560000 41.920000 ;
      LAYER met4 ;
        RECT 51.240000 41.600000 51.560000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 42.030000 51.560000 42.350000 ;
      LAYER met4 ;
        RECT 51.240000 42.030000 51.560000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 42.460000 51.560000 42.780000 ;
      LAYER met4 ;
        RECT 51.240000 42.460000 51.560000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 42.890000 51.560000 43.210000 ;
      LAYER met4 ;
        RECT 51.240000 42.890000 51.560000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 43.320000 51.560000 43.640000 ;
      LAYER met4 ;
        RECT 51.240000 43.320000 51.560000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 43.750000 51.560000 44.070000 ;
      LAYER met4 ;
        RECT 51.240000 43.750000 51.560000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 44.180000 51.560000 44.500000 ;
      LAYER met4 ;
        RECT 51.240000 44.180000 51.560000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 44.610000 51.560000 44.930000 ;
      LAYER met4 ;
        RECT 51.240000 44.610000 51.560000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 45.040000 51.560000 45.360000 ;
      LAYER met4 ;
        RECT 51.240000 45.040000 51.560000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 45.470000 51.560000 45.790000 ;
      LAYER met4 ;
        RECT 51.240000 45.470000 51.560000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 45.900000 51.560000 46.220000 ;
      LAYER met4 ;
        RECT 51.240000 45.900000 51.560000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 41.600000 51.970000 41.920000 ;
      LAYER met4 ;
        RECT 51.650000 41.600000 51.970000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 42.030000 51.970000 42.350000 ;
      LAYER met4 ;
        RECT 51.650000 42.030000 51.970000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 42.460000 51.970000 42.780000 ;
      LAYER met4 ;
        RECT 51.650000 42.460000 51.970000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 42.890000 51.970000 43.210000 ;
      LAYER met4 ;
        RECT 51.650000 42.890000 51.970000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 43.320000 51.970000 43.640000 ;
      LAYER met4 ;
        RECT 51.650000 43.320000 51.970000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 43.750000 51.970000 44.070000 ;
      LAYER met4 ;
        RECT 51.650000 43.750000 51.970000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 44.180000 51.970000 44.500000 ;
      LAYER met4 ;
        RECT 51.650000 44.180000 51.970000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 44.610000 51.970000 44.930000 ;
      LAYER met4 ;
        RECT 51.650000 44.610000 51.970000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 45.040000 51.970000 45.360000 ;
      LAYER met4 ;
        RECT 51.650000 45.040000 51.970000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 45.470000 51.970000 45.790000 ;
      LAYER met4 ;
        RECT 51.650000 45.470000 51.970000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 45.900000 51.970000 46.220000 ;
      LAYER met4 ;
        RECT 51.650000 45.900000 51.970000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 41.600000 52.380000 41.920000 ;
      LAYER met4 ;
        RECT 52.060000 41.600000 52.380000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 42.030000 52.380000 42.350000 ;
      LAYER met4 ;
        RECT 52.060000 42.030000 52.380000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 42.460000 52.380000 42.780000 ;
      LAYER met4 ;
        RECT 52.060000 42.460000 52.380000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 42.890000 52.380000 43.210000 ;
      LAYER met4 ;
        RECT 52.060000 42.890000 52.380000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 43.320000 52.380000 43.640000 ;
      LAYER met4 ;
        RECT 52.060000 43.320000 52.380000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 43.750000 52.380000 44.070000 ;
      LAYER met4 ;
        RECT 52.060000 43.750000 52.380000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 44.180000 52.380000 44.500000 ;
      LAYER met4 ;
        RECT 52.060000 44.180000 52.380000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 44.610000 52.380000 44.930000 ;
      LAYER met4 ;
        RECT 52.060000 44.610000 52.380000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 45.040000 52.380000 45.360000 ;
      LAYER met4 ;
        RECT 52.060000 45.040000 52.380000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 45.470000 52.380000 45.790000 ;
      LAYER met4 ;
        RECT 52.060000 45.470000 52.380000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 45.900000 52.380000 46.220000 ;
      LAYER met4 ;
        RECT 52.060000 45.900000 52.380000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 41.600000 52.790000 41.920000 ;
      LAYER met4 ;
        RECT 52.470000 41.600000 52.790000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 42.030000 52.790000 42.350000 ;
      LAYER met4 ;
        RECT 52.470000 42.030000 52.790000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 42.460000 52.790000 42.780000 ;
      LAYER met4 ;
        RECT 52.470000 42.460000 52.790000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 42.890000 52.790000 43.210000 ;
      LAYER met4 ;
        RECT 52.470000 42.890000 52.790000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 43.320000 52.790000 43.640000 ;
      LAYER met4 ;
        RECT 52.470000 43.320000 52.790000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 43.750000 52.790000 44.070000 ;
      LAYER met4 ;
        RECT 52.470000 43.750000 52.790000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 44.180000 52.790000 44.500000 ;
      LAYER met4 ;
        RECT 52.470000 44.180000 52.790000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 44.610000 52.790000 44.930000 ;
      LAYER met4 ;
        RECT 52.470000 44.610000 52.790000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 45.040000 52.790000 45.360000 ;
      LAYER met4 ;
        RECT 52.470000 45.040000 52.790000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 45.470000 52.790000 45.790000 ;
      LAYER met4 ;
        RECT 52.470000 45.470000 52.790000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 45.900000 52.790000 46.220000 ;
      LAYER met4 ;
        RECT 52.470000 45.900000 52.790000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 41.600000 53.200000 41.920000 ;
      LAYER met4 ;
        RECT 52.880000 41.600000 53.200000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 42.030000 53.200000 42.350000 ;
      LAYER met4 ;
        RECT 52.880000 42.030000 53.200000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 42.460000 53.200000 42.780000 ;
      LAYER met4 ;
        RECT 52.880000 42.460000 53.200000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 42.890000 53.200000 43.210000 ;
      LAYER met4 ;
        RECT 52.880000 42.890000 53.200000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 43.320000 53.200000 43.640000 ;
      LAYER met4 ;
        RECT 52.880000 43.320000 53.200000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 43.750000 53.200000 44.070000 ;
      LAYER met4 ;
        RECT 52.880000 43.750000 53.200000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 44.180000 53.200000 44.500000 ;
      LAYER met4 ;
        RECT 52.880000 44.180000 53.200000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 44.610000 53.200000 44.930000 ;
      LAYER met4 ;
        RECT 52.880000 44.610000 53.200000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 45.040000 53.200000 45.360000 ;
      LAYER met4 ;
        RECT 52.880000 45.040000 53.200000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 45.470000 53.200000 45.790000 ;
      LAYER met4 ;
        RECT 52.880000 45.470000 53.200000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 45.900000 53.200000 46.220000 ;
      LAYER met4 ;
        RECT 52.880000 45.900000 53.200000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 41.600000 53.605000 41.920000 ;
      LAYER met4 ;
        RECT 53.285000 41.600000 53.605000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 42.030000 53.605000 42.350000 ;
      LAYER met4 ;
        RECT 53.285000 42.030000 53.605000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 42.460000 53.605000 42.780000 ;
      LAYER met4 ;
        RECT 53.285000 42.460000 53.605000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 42.890000 53.605000 43.210000 ;
      LAYER met4 ;
        RECT 53.285000 42.890000 53.605000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 43.320000 53.605000 43.640000 ;
      LAYER met4 ;
        RECT 53.285000 43.320000 53.605000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 43.750000 53.605000 44.070000 ;
      LAYER met4 ;
        RECT 53.285000 43.750000 53.605000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 44.180000 53.605000 44.500000 ;
      LAYER met4 ;
        RECT 53.285000 44.180000 53.605000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 44.610000 53.605000 44.930000 ;
      LAYER met4 ;
        RECT 53.285000 44.610000 53.605000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 45.040000 53.605000 45.360000 ;
      LAYER met4 ;
        RECT 53.285000 45.040000 53.605000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 45.470000 53.605000 45.790000 ;
      LAYER met4 ;
        RECT 53.285000 45.470000 53.605000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 45.900000 53.605000 46.220000 ;
      LAYER met4 ;
        RECT 53.285000 45.900000 53.605000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 41.600000 54.010000 41.920000 ;
      LAYER met4 ;
        RECT 53.690000 41.600000 54.010000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 42.030000 54.010000 42.350000 ;
      LAYER met4 ;
        RECT 53.690000 42.030000 54.010000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 42.460000 54.010000 42.780000 ;
      LAYER met4 ;
        RECT 53.690000 42.460000 54.010000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 42.890000 54.010000 43.210000 ;
      LAYER met4 ;
        RECT 53.690000 42.890000 54.010000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 43.320000 54.010000 43.640000 ;
      LAYER met4 ;
        RECT 53.690000 43.320000 54.010000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 43.750000 54.010000 44.070000 ;
      LAYER met4 ;
        RECT 53.690000 43.750000 54.010000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 44.180000 54.010000 44.500000 ;
      LAYER met4 ;
        RECT 53.690000 44.180000 54.010000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 44.610000 54.010000 44.930000 ;
      LAYER met4 ;
        RECT 53.690000 44.610000 54.010000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 45.040000 54.010000 45.360000 ;
      LAYER met4 ;
        RECT 53.690000 45.040000 54.010000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 45.470000 54.010000 45.790000 ;
      LAYER met4 ;
        RECT 53.690000 45.470000 54.010000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 45.900000 54.010000 46.220000 ;
      LAYER met4 ;
        RECT 53.690000 45.900000 54.010000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 41.600000 54.415000 41.920000 ;
      LAYER met4 ;
        RECT 54.095000 41.600000 54.415000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 42.030000 54.415000 42.350000 ;
      LAYER met4 ;
        RECT 54.095000 42.030000 54.415000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 42.460000 54.415000 42.780000 ;
      LAYER met4 ;
        RECT 54.095000 42.460000 54.415000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 42.890000 54.415000 43.210000 ;
      LAYER met4 ;
        RECT 54.095000 42.890000 54.415000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 43.320000 54.415000 43.640000 ;
      LAYER met4 ;
        RECT 54.095000 43.320000 54.415000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 43.750000 54.415000 44.070000 ;
      LAYER met4 ;
        RECT 54.095000 43.750000 54.415000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 44.180000 54.415000 44.500000 ;
      LAYER met4 ;
        RECT 54.095000 44.180000 54.415000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 44.610000 54.415000 44.930000 ;
      LAYER met4 ;
        RECT 54.095000 44.610000 54.415000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 45.040000 54.415000 45.360000 ;
      LAYER met4 ;
        RECT 54.095000 45.040000 54.415000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 45.470000 54.415000 45.790000 ;
      LAYER met4 ;
        RECT 54.095000 45.470000 54.415000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 45.900000 54.415000 46.220000 ;
      LAYER met4 ;
        RECT 54.095000 45.900000 54.415000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 41.600000 54.820000 41.920000 ;
      LAYER met4 ;
        RECT 54.500000 41.600000 54.820000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 42.030000 54.820000 42.350000 ;
      LAYER met4 ;
        RECT 54.500000 42.030000 54.820000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 42.460000 54.820000 42.780000 ;
      LAYER met4 ;
        RECT 54.500000 42.460000 54.820000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 42.890000 54.820000 43.210000 ;
      LAYER met4 ;
        RECT 54.500000 42.890000 54.820000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 43.320000 54.820000 43.640000 ;
      LAYER met4 ;
        RECT 54.500000 43.320000 54.820000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 43.750000 54.820000 44.070000 ;
      LAYER met4 ;
        RECT 54.500000 43.750000 54.820000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 44.180000 54.820000 44.500000 ;
      LAYER met4 ;
        RECT 54.500000 44.180000 54.820000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 44.610000 54.820000 44.930000 ;
      LAYER met4 ;
        RECT 54.500000 44.610000 54.820000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 45.040000 54.820000 45.360000 ;
      LAYER met4 ;
        RECT 54.500000 45.040000 54.820000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 45.470000 54.820000 45.790000 ;
      LAYER met4 ;
        RECT 54.500000 45.470000 54.820000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 45.900000 54.820000 46.220000 ;
      LAYER met4 ;
        RECT 54.500000 45.900000 54.820000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 41.600000 55.225000 41.920000 ;
      LAYER met4 ;
        RECT 54.905000 41.600000 55.225000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 42.030000 55.225000 42.350000 ;
      LAYER met4 ;
        RECT 54.905000 42.030000 55.225000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 42.460000 55.225000 42.780000 ;
      LAYER met4 ;
        RECT 54.905000 42.460000 55.225000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 42.890000 55.225000 43.210000 ;
      LAYER met4 ;
        RECT 54.905000 42.890000 55.225000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 43.320000 55.225000 43.640000 ;
      LAYER met4 ;
        RECT 54.905000 43.320000 55.225000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 43.750000 55.225000 44.070000 ;
      LAYER met4 ;
        RECT 54.905000 43.750000 55.225000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 44.180000 55.225000 44.500000 ;
      LAYER met4 ;
        RECT 54.905000 44.180000 55.225000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 44.610000 55.225000 44.930000 ;
      LAYER met4 ;
        RECT 54.905000 44.610000 55.225000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 45.040000 55.225000 45.360000 ;
      LAYER met4 ;
        RECT 54.905000 45.040000 55.225000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 45.470000 55.225000 45.790000 ;
      LAYER met4 ;
        RECT 54.905000 45.470000 55.225000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 45.900000 55.225000 46.220000 ;
      LAYER met4 ;
        RECT 54.905000 45.900000 55.225000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 41.600000 55.630000 41.920000 ;
      LAYER met4 ;
        RECT 55.310000 41.600000 55.630000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 42.030000 55.630000 42.350000 ;
      LAYER met4 ;
        RECT 55.310000 42.030000 55.630000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 42.460000 55.630000 42.780000 ;
      LAYER met4 ;
        RECT 55.310000 42.460000 55.630000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 42.890000 55.630000 43.210000 ;
      LAYER met4 ;
        RECT 55.310000 42.890000 55.630000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 43.320000 55.630000 43.640000 ;
      LAYER met4 ;
        RECT 55.310000 43.320000 55.630000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 43.750000 55.630000 44.070000 ;
      LAYER met4 ;
        RECT 55.310000 43.750000 55.630000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 44.180000 55.630000 44.500000 ;
      LAYER met4 ;
        RECT 55.310000 44.180000 55.630000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 44.610000 55.630000 44.930000 ;
      LAYER met4 ;
        RECT 55.310000 44.610000 55.630000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 45.040000 55.630000 45.360000 ;
      LAYER met4 ;
        RECT 55.310000 45.040000 55.630000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 45.470000 55.630000 45.790000 ;
      LAYER met4 ;
        RECT 55.310000 45.470000 55.630000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 45.900000 55.630000 46.220000 ;
      LAYER met4 ;
        RECT 55.310000 45.900000 55.630000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 41.600000 56.035000 41.920000 ;
      LAYER met4 ;
        RECT 55.715000 41.600000 56.035000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 42.030000 56.035000 42.350000 ;
      LAYER met4 ;
        RECT 55.715000 42.030000 56.035000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 42.460000 56.035000 42.780000 ;
      LAYER met4 ;
        RECT 55.715000 42.460000 56.035000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 42.890000 56.035000 43.210000 ;
      LAYER met4 ;
        RECT 55.715000 42.890000 56.035000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 43.320000 56.035000 43.640000 ;
      LAYER met4 ;
        RECT 55.715000 43.320000 56.035000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 43.750000 56.035000 44.070000 ;
      LAYER met4 ;
        RECT 55.715000 43.750000 56.035000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 44.180000 56.035000 44.500000 ;
      LAYER met4 ;
        RECT 55.715000 44.180000 56.035000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 44.610000 56.035000 44.930000 ;
      LAYER met4 ;
        RECT 55.715000 44.610000 56.035000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 45.040000 56.035000 45.360000 ;
      LAYER met4 ;
        RECT 55.715000 45.040000 56.035000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 45.470000 56.035000 45.790000 ;
      LAYER met4 ;
        RECT 55.715000 45.470000 56.035000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 45.900000 56.035000 46.220000 ;
      LAYER met4 ;
        RECT 55.715000 45.900000 56.035000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 41.600000 56.440000 41.920000 ;
      LAYER met4 ;
        RECT 56.120000 41.600000 56.440000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 42.030000 56.440000 42.350000 ;
      LAYER met4 ;
        RECT 56.120000 42.030000 56.440000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 42.460000 56.440000 42.780000 ;
      LAYER met4 ;
        RECT 56.120000 42.460000 56.440000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 42.890000 56.440000 43.210000 ;
      LAYER met4 ;
        RECT 56.120000 42.890000 56.440000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 43.320000 56.440000 43.640000 ;
      LAYER met4 ;
        RECT 56.120000 43.320000 56.440000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 43.750000 56.440000 44.070000 ;
      LAYER met4 ;
        RECT 56.120000 43.750000 56.440000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 44.180000 56.440000 44.500000 ;
      LAYER met4 ;
        RECT 56.120000 44.180000 56.440000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 44.610000 56.440000 44.930000 ;
      LAYER met4 ;
        RECT 56.120000 44.610000 56.440000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 45.040000 56.440000 45.360000 ;
      LAYER met4 ;
        RECT 56.120000 45.040000 56.440000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 45.470000 56.440000 45.790000 ;
      LAYER met4 ;
        RECT 56.120000 45.470000 56.440000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 45.900000 56.440000 46.220000 ;
      LAYER met4 ;
        RECT 56.120000 45.900000 56.440000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 41.600000 56.845000 41.920000 ;
      LAYER met4 ;
        RECT 56.525000 41.600000 56.845000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 42.030000 56.845000 42.350000 ;
      LAYER met4 ;
        RECT 56.525000 42.030000 56.845000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 42.460000 56.845000 42.780000 ;
      LAYER met4 ;
        RECT 56.525000 42.460000 56.845000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 42.890000 56.845000 43.210000 ;
      LAYER met4 ;
        RECT 56.525000 42.890000 56.845000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 43.320000 56.845000 43.640000 ;
      LAYER met4 ;
        RECT 56.525000 43.320000 56.845000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 43.750000 56.845000 44.070000 ;
      LAYER met4 ;
        RECT 56.525000 43.750000 56.845000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 44.180000 56.845000 44.500000 ;
      LAYER met4 ;
        RECT 56.525000 44.180000 56.845000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 44.610000 56.845000 44.930000 ;
      LAYER met4 ;
        RECT 56.525000 44.610000 56.845000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 45.040000 56.845000 45.360000 ;
      LAYER met4 ;
        RECT 56.525000 45.040000 56.845000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 45.470000 56.845000 45.790000 ;
      LAYER met4 ;
        RECT 56.525000 45.470000 56.845000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 45.900000 56.845000 46.220000 ;
      LAYER met4 ;
        RECT 56.525000 45.900000 56.845000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 41.600000 57.250000 41.920000 ;
      LAYER met4 ;
        RECT 56.930000 41.600000 57.250000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 42.030000 57.250000 42.350000 ;
      LAYER met4 ;
        RECT 56.930000 42.030000 57.250000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 42.460000 57.250000 42.780000 ;
      LAYER met4 ;
        RECT 56.930000 42.460000 57.250000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 42.890000 57.250000 43.210000 ;
      LAYER met4 ;
        RECT 56.930000 42.890000 57.250000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 43.320000 57.250000 43.640000 ;
      LAYER met4 ;
        RECT 56.930000 43.320000 57.250000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 43.750000 57.250000 44.070000 ;
      LAYER met4 ;
        RECT 56.930000 43.750000 57.250000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 44.180000 57.250000 44.500000 ;
      LAYER met4 ;
        RECT 56.930000 44.180000 57.250000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 44.610000 57.250000 44.930000 ;
      LAYER met4 ;
        RECT 56.930000 44.610000 57.250000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 45.040000 57.250000 45.360000 ;
      LAYER met4 ;
        RECT 56.930000 45.040000 57.250000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 45.470000 57.250000 45.790000 ;
      LAYER met4 ;
        RECT 56.930000 45.470000 57.250000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 45.900000 57.250000 46.220000 ;
      LAYER met4 ;
        RECT 56.930000 45.900000 57.250000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 41.600000 57.655000 41.920000 ;
      LAYER met4 ;
        RECT 57.335000 41.600000 57.655000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 42.030000 57.655000 42.350000 ;
      LAYER met4 ;
        RECT 57.335000 42.030000 57.655000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 42.460000 57.655000 42.780000 ;
      LAYER met4 ;
        RECT 57.335000 42.460000 57.655000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 42.890000 57.655000 43.210000 ;
      LAYER met4 ;
        RECT 57.335000 42.890000 57.655000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 43.320000 57.655000 43.640000 ;
      LAYER met4 ;
        RECT 57.335000 43.320000 57.655000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 43.750000 57.655000 44.070000 ;
      LAYER met4 ;
        RECT 57.335000 43.750000 57.655000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 44.180000 57.655000 44.500000 ;
      LAYER met4 ;
        RECT 57.335000 44.180000 57.655000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 44.610000 57.655000 44.930000 ;
      LAYER met4 ;
        RECT 57.335000 44.610000 57.655000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 45.040000 57.655000 45.360000 ;
      LAYER met4 ;
        RECT 57.335000 45.040000 57.655000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 45.470000 57.655000 45.790000 ;
      LAYER met4 ;
        RECT 57.335000 45.470000 57.655000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 45.900000 57.655000 46.220000 ;
      LAYER met4 ;
        RECT 57.335000 45.900000 57.655000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 41.600000 58.060000 41.920000 ;
      LAYER met4 ;
        RECT 57.740000 41.600000 58.060000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 42.030000 58.060000 42.350000 ;
      LAYER met4 ;
        RECT 57.740000 42.030000 58.060000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 42.460000 58.060000 42.780000 ;
      LAYER met4 ;
        RECT 57.740000 42.460000 58.060000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 42.890000 58.060000 43.210000 ;
      LAYER met4 ;
        RECT 57.740000 42.890000 58.060000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 43.320000 58.060000 43.640000 ;
      LAYER met4 ;
        RECT 57.740000 43.320000 58.060000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 43.750000 58.060000 44.070000 ;
      LAYER met4 ;
        RECT 57.740000 43.750000 58.060000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 44.180000 58.060000 44.500000 ;
      LAYER met4 ;
        RECT 57.740000 44.180000 58.060000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 44.610000 58.060000 44.930000 ;
      LAYER met4 ;
        RECT 57.740000 44.610000 58.060000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 45.040000 58.060000 45.360000 ;
      LAYER met4 ;
        RECT 57.740000 45.040000 58.060000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 45.470000 58.060000 45.790000 ;
      LAYER met4 ;
        RECT 57.740000 45.470000 58.060000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 45.900000 58.060000 46.220000 ;
      LAYER met4 ;
        RECT 57.740000 45.900000 58.060000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 41.600000 58.465000 41.920000 ;
      LAYER met4 ;
        RECT 58.145000 41.600000 58.465000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 42.030000 58.465000 42.350000 ;
      LAYER met4 ;
        RECT 58.145000 42.030000 58.465000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 42.460000 58.465000 42.780000 ;
      LAYER met4 ;
        RECT 58.145000 42.460000 58.465000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 42.890000 58.465000 43.210000 ;
      LAYER met4 ;
        RECT 58.145000 42.890000 58.465000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 43.320000 58.465000 43.640000 ;
      LAYER met4 ;
        RECT 58.145000 43.320000 58.465000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 43.750000 58.465000 44.070000 ;
      LAYER met4 ;
        RECT 58.145000 43.750000 58.465000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 44.180000 58.465000 44.500000 ;
      LAYER met4 ;
        RECT 58.145000 44.180000 58.465000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 44.610000 58.465000 44.930000 ;
      LAYER met4 ;
        RECT 58.145000 44.610000 58.465000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 45.040000 58.465000 45.360000 ;
      LAYER met4 ;
        RECT 58.145000 45.040000 58.465000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 45.470000 58.465000 45.790000 ;
      LAYER met4 ;
        RECT 58.145000 45.470000 58.465000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 45.900000 58.465000 46.220000 ;
      LAYER met4 ;
        RECT 58.145000 45.900000 58.465000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 41.600000 58.870000 41.920000 ;
      LAYER met4 ;
        RECT 58.550000 41.600000 58.870000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 42.030000 58.870000 42.350000 ;
      LAYER met4 ;
        RECT 58.550000 42.030000 58.870000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 42.460000 58.870000 42.780000 ;
      LAYER met4 ;
        RECT 58.550000 42.460000 58.870000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 42.890000 58.870000 43.210000 ;
      LAYER met4 ;
        RECT 58.550000 42.890000 58.870000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 43.320000 58.870000 43.640000 ;
      LAYER met4 ;
        RECT 58.550000 43.320000 58.870000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 43.750000 58.870000 44.070000 ;
      LAYER met4 ;
        RECT 58.550000 43.750000 58.870000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 44.180000 58.870000 44.500000 ;
      LAYER met4 ;
        RECT 58.550000 44.180000 58.870000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 44.610000 58.870000 44.930000 ;
      LAYER met4 ;
        RECT 58.550000 44.610000 58.870000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 45.040000 58.870000 45.360000 ;
      LAYER met4 ;
        RECT 58.550000 45.040000 58.870000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 45.470000 58.870000 45.790000 ;
      LAYER met4 ;
        RECT 58.550000 45.470000 58.870000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 45.900000 58.870000 46.220000 ;
      LAYER met4 ;
        RECT 58.550000 45.900000 58.870000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 41.600000 59.275000 41.920000 ;
      LAYER met4 ;
        RECT 58.955000 41.600000 59.275000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 42.030000 59.275000 42.350000 ;
      LAYER met4 ;
        RECT 58.955000 42.030000 59.275000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 42.460000 59.275000 42.780000 ;
      LAYER met4 ;
        RECT 58.955000 42.460000 59.275000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 42.890000 59.275000 43.210000 ;
      LAYER met4 ;
        RECT 58.955000 42.890000 59.275000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 43.320000 59.275000 43.640000 ;
      LAYER met4 ;
        RECT 58.955000 43.320000 59.275000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 43.750000 59.275000 44.070000 ;
      LAYER met4 ;
        RECT 58.955000 43.750000 59.275000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 44.180000 59.275000 44.500000 ;
      LAYER met4 ;
        RECT 58.955000 44.180000 59.275000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 44.610000 59.275000 44.930000 ;
      LAYER met4 ;
        RECT 58.955000 44.610000 59.275000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 45.040000 59.275000 45.360000 ;
      LAYER met4 ;
        RECT 58.955000 45.040000 59.275000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 45.470000 59.275000 45.790000 ;
      LAYER met4 ;
        RECT 58.955000 45.470000 59.275000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 45.900000 59.275000 46.220000 ;
      LAYER met4 ;
        RECT 58.955000 45.900000 59.275000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 41.600000 59.680000 41.920000 ;
      LAYER met4 ;
        RECT 59.360000 41.600000 59.680000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 42.030000 59.680000 42.350000 ;
      LAYER met4 ;
        RECT 59.360000 42.030000 59.680000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 42.460000 59.680000 42.780000 ;
      LAYER met4 ;
        RECT 59.360000 42.460000 59.680000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 42.890000 59.680000 43.210000 ;
      LAYER met4 ;
        RECT 59.360000 42.890000 59.680000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 43.320000 59.680000 43.640000 ;
      LAYER met4 ;
        RECT 59.360000 43.320000 59.680000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 43.750000 59.680000 44.070000 ;
      LAYER met4 ;
        RECT 59.360000 43.750000 59.680000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 44.180000 59.680000 44.500000 ;
      LAYER met4 ;
        RECT 59.360000 44.180000 59.680000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 44.610000 59.680000 44.930000 ;
      LAYER met4 ;
        RECT 59.360000 44.610000 59.680000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 45.040000 59.680000 45.360000 ;
      LAYER met4 ;
        RECT 59.360000 45.040000 59.680000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 45.470000 59.680000 45.790000 ;
      LAYER met4 ;
        RECT 59.360000 45.470000 59.680000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 45.900000 59.680000 46.220000 ;
      LAYER met4 ;
        RECT 59.360000 45.900000 59.680000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 41.600000 60.085000 41.920000 ;
      LAYER met4 ;
        RECT 59.765000 41.600000 60.085000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 42.030000 60.085000 42.350000 ;
      LAYER met4 ;
        RECT 59.765000 42.030000 60.085000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 42.460000 60.085000 42.780000 ;
      LAYER met4 ;
        RECT 59.765000 42.460000 60.085000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 42.890000 60.085000 43.210000 ;
      LAYER met4 ;
        RECT 59.765000 42.890000 60.085000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 43.320000 60.085000 43.640000 ;
      LAYER met4 ;
        RECT 59.765000 43.320000 60.085000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 43.750000 60.085000 44.070000 ;
      LAYER met4 ;
        RECT 59.765000 43.750000 60.085000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 44.180000 60.085000 44.500000 ;
      LAYER met4 ;
        RECT 59.765000 44.180000 60.085000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 44.610000 60.085000 44.930000 ;
      LAYER met4 ;
        RECT 59.765000 44.610000 60.085000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 45.040000 60.085000 45.360000 ;
      LAYER met4 ;
        RECT 59.765000 45.040000 60.085000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 45.470000 60.085000 45.790000 ;
      LAYER met4 ;
        RECT 59.765000 45.470000 60.085000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 45.900000 60.085000 46.220000 ;
      LAYER met4 ;
        RECT 59.765000 45.900000 60.085000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265000 41.600000 6.585000 41.920000 ;
      LAYER met4 ;
        RECT 6.265000 41.600000 6.585000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265000 42.030000 6.585000 42.350000 ;
      LAYER met4 ;
        RECT 6.265000 42.030000 6.585000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265000 42.460000 6.585000 42.780000 ;
      LAYER met4 ;
        RECT 6.265000 42.460000 6.585000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265000 42.890000 6.585000 43.210000 ;
      LAYER met4 ;
        RECT 6.265000 42.890000 6.585000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265000 43.320000 6.585000 43.640000 ;
      LAYER met4 ;
        RECT 6.265000 43.320000 6.585000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265000 43.750000 6.585000 44.070000 ;
      LAYER met4 ;
        RECT 6.265000 43.750000 6.585000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265000 44.180000 6.585000 44.500000 ;
      LAYER met4 ;
        RECT 6.265000 44.180000 6.585000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265000 44.610000 6.585000 44.930000 ;
      LAYER met4 ;
        RECT 6.265000 44.610000 6.585000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265000 45.040000 6.585000 45.360000 ;
      LAYER met4 ;
        RECT 6.265000 45.040000 6.585000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265000 45.470000 6.585000 45.790000 ;
      LAYER met4 ;
        RECT 6.265000 45.470000 6.585000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265000 45.900000 6.585000 46.220000 ;
      LAYER met4 ;
        RECT 6.265000 45.900000 6.585000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670000 41.600000 6.990000 41.920000 ;
      LAYER met4 ;
        RECT 6.670000 41.600000 6.990000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670000 42.030000 6.990000 42.350000 ;
      LAYER met4 ;
        RECT 6.670000 42.030000 6.990000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670000 42.460000 6.990000 42.780000 ;
      LAYER met4 ;
        RECT 6.670000 42.460000 6.990000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670000 42.890000 6.990000 43.210000 ;
      LAYER met4 ;
        RECT 6.670000 42.890000 6.990000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670000 43.320000 6.990000 43.640000 ;
      LAYER met4 ;
        RECT 6.670000 43.320000 6.990000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670000 43.750000 6.990000 44.070000 ;
      LAYER met4 ;
        RECT 6.670000 43.750000 6.990000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670000 44.180000 6.990000 44.500000 ;
      LAYER met4 ;
        RECT 6.670000 44.180000 6.990000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670000 44.610000 6.990000 44.930000 ;
      LAYER met4 ;
        RECT 6.670000 44.610000 6.990000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670000 45.040000 6.990000 45.360000 ;
      LAYER met4 ;
        RECT 6.670000 45.040000 6.990000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670000 45.470000 6.990000 45.790000 ;
      LAYER met4 ;
        RECT 6.670000 45.470000 6.990000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670000 45.900000 6.990000 46.220000 ;
      LAYER met4 ;
        RECT 6.670000 45.900000 6.990000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 41.600000 60.490000 41.920000 ;
      LAYER met4 ;
        RECT 60.170000 41.600000 60.490000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 42.030000 60.490000 42.350000 ;
      LAYER met4 ;
        RECT 60.170000 42.030000 60.490000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 42.460000 60.490000 42.780000 ;
      LAYER met4 ;
        RECT 60.170000 42.460000 60.490000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 42.890000 60.490000 43.210000 ;
      LAYER met4 ;
        RECT 60.170000 42.890000 60.490000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 43.320000 60.490000 43.640000 ;
      LAYER met4 ;
        RECT 60.170000 43.320000 60.490000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 43.750000 60.490000 44.070000 ;
      LAYER met4 ;
        RECT 60.170000 43.750000 60.490000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 44.180000 60.490000 44.500000 ;
      LAYER met4 ;
        RECT 60.170000 44.180000 60.490000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 44.610000 60.490000 44.930000 ;
      LAYER met4 ;
        RECT 60.170000 44.610000 60.490000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 45.040000 60.490000 45.360000 ;
      LAYER met4 ;
        RECT 60.170000 45.040000 60.490000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 45.470000 60.490000 45.790000 ;
      LAYER met4 ;
        RECT 60.170000 45.470000 60.490000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 45.900000 60.490000 46.220000 ;
      LAYER met4 ;
        RECT 60.170000 45.900000 60.490000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 41.600000 60.895000 41.920000 ;
      LAYER met4 ;
        RECT 60.575000 41.600000 60.895000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 42.030000 60.895000 42.350000 ;
      LAYER met4 ;
        RECT 60.575000 42.030000 60.895000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 42.460000 60.895000 42.780000 ;
      LAYER met4 ;
        RECT 60.575000 42.460000 60.895000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 42.890000 60.895000 43.210000 ;
      LAYER met4 ;
        RECT 60.575000 42.890000 60.895000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 43.320000 60.895000 43.640000 ;
      LAYER met4 ;
        RECT 60.575000 43.320000 60.895000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 43.750000 60.895000 44.070000 ;
      LAYER met4 ;
        RECT 60.575000 43.750000 60.895000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 44.180000 60.895000 44.500000 ;
      LAYER met4 ;
        RECT 60.575000 44.180000 60.895000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 44.610000 60.895000 44.930000 ;
      LAYER met4 ;
        RECT 60.575000 44.610000 60.895000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 45.040000 60.895000 45.360000 ;
      LAYER met4 ;
        RECT 60.575000 45.040000 60.895000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 45.470000 60.895000 45.790000 ;
      LAYER met4 ;
        RECT 60.575000 45.470000 60.895000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 45.900000 60.895000 46.220000 ;
      LAYER met4 ;
        RECT 60.575000 45.900000 60.895000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 41.600000 61.300000 41.920000 ;
      LAYER met4 ;
        RECT 60.980000 41.600000 61.300000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 42.030000 61.300000 42.350000 ;
      LAYER met4 ;
        RECT 60.980000 42.030000 61.300000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 42.460000 61.300000 42.780000 ;
      LAYER met4 ;
        RECT 60.980000 42.460000 61.300000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 42.890000 61.300000 43.210000 ;
      LAYER met4 ;
        RECT 60.980000 42.890000 61.300000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 43.320000 61.300000 43.640000 ;
      LAYER met4 ;
        RECT 60.980000 43.320000 61.300000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 43.750000 61.300000 44.070000 ;
      LAYER met4 ;
        RECT 60.980000 43.750000 61.300000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 44.180000 61.300000 44.500000 ;
      LAYER met4 ;
        RECT 60.980000 44.180000 61.300000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 44.610000 61.300000 44.930000 ;
      LAYER met4 ;
        RECT 60.980000 44.610000 61.300000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 45.040000 61.300000 45.360000 ;
      LAYER met4 ;
        RECT 60.980000 45.040000 61.300000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 45.470000 61.300000 45.790000 ;
      LAYER met4 ;
        RECT 60.980000 45.470000 61.300000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 45.900000 61.300000 46.220000 ;
      LAYER met4 ;
        RECT 60.980000 45.900000 61.300000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 41.600000 61.705000 41.920000 ;
      LAYER met4 ;
        RECT 61.385000 41.600000 61.705000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 42.030000 61.705000 42.350000 ;
      LAYER met4 ;
        RECT 61.385000 42.030000 61.705000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 42.460000 61.705000 42.780000 ;
      LAYER met4 ;
        RECT 61.385000 42.460000 61.705000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 42.890000 61.705000 43.210000 ;
      LAYER met4 ;
        RECT 61.385000 42.890000 61.705000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 43.320000 61.705000 43.640000 ;
      LAYER met4 ;
        RECT 61.385000 43.320000 61.705000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 43.750000 61.705000 44.070000 ;
      LAYER met4 ;
        RECT 61.385000 43.750000 61.705000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 44.180000 61.705000 44.500000 ;
      LAYER met4 ;
        RECT 61.385000 44.180000 61.705000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 44.610000 61.705000 44.930000 ;
      LAYER met4 ;
        RECT 61.385000 44.610000 61.705000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 45.040000 61.705000 45.360000 ;
      LAYER met4 ;
        RECT 61.385000 45.040000 61.705000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 45.470000 61.705000 45.790000 ;
      LAYER met4 ;
        RECT 61.385000 45.470000 61.705000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 45.900000 61.705000 46.220000 ;
      LAYER met4 ;
        RECT 61.385000 45.900000 61.705000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 41.600000 62.110000 41.920000 ;
      LAYER met4 ;
        RECT 61.790000 41.600000 62.110000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 42.030000 62.110000 42.350000 ;
      LAYER met4 ;
        RECT 61.790000 42.030000 62.110000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 42.460000 62.110000 42.780000 ;
      LAYER met4 ;
        RECT 61.790000 42.460000 62.110000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 42.890000 62.110000 43.210000 ;
      LAYER met4 ;
        RECT 61.790000 42.890000 62.110000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 43.320000 62.110000 43.640000 ;
      LAYER met4 ;
        RECT 61.790000 43.320000 62.110000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 43.750000 62.110000 44.070000 ;
      LAYER met4 ;
        RECT 61.790000 43.750000 62.110000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 44.180000 62.110000 44.500000 ;
      LAYER met4 ;
        RECT 61.790000 44.180000 62.110000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 44.610000 62.110000 44.930000 ;
      LAYER met4 ;
        RECT 61.790000 44.610000 62.110000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 45.040000 62.110000 45.360000 ;
      LAYER met4 ;
        RECT 61.790000 45.040000 62.110000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 45.470000 62.110000 45.790000 ;
      LAYER met4 ;
        RECT 61.790000 45.470000 62.110000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 45.900000 62.110000 46.220000 ;
      LAYER met4 ;
        RECT 61.790000 45.900000 62.110000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 41.600000 62.515000 41.920000 ;
      LAYER met4 ;
        RECT 62.195000 41.600000 62.515000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 42.030000 62.515000 42.350000 ;
      LAYER met4 ;
        RECT 62.195000 42.030000 62.515000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 42.460000 62.515000 42.780000 ;
      LAYER met4 ;
        RECT 62.195000 42.460000 62.515000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 42.890000 62.515000 43.210000 ;
      LAYER met4 ;
        RECT 62.195000 42.890000 62.515000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 43.320000 62.515000 43.640000 ;
      LAYER met4 ;
        RECT 62.195000 43.320000 62.515000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 43.750000 62.515000 44.070000 ;
      LAYER met4 ;
        RECT 62.195000 43.750000 62.515000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 44.180000 62.515000 44.500000 ;
      LAYER met4 ;
        RECT 62.195000 44.180000 62.515000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 44.610000 62.515000 44.930000 ;
      LAYER met4 ;
        RECT 62.195000 44.610000 62.515000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 45.040000 62.515000 45.360000 ;
      LAYER met4 ;
        RECT 62.195000 45.040000 62.515000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 45.470000 62.515000 45.790000 ;
      LAYER met4 ;
        RECT 62.195000 45.470000 62.515000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 45.900000 62.515000 46.220000 ;
      LAYER met4 ;
        RECT 62.195000 45.900000 62.515000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 41.600000 62.920000 41.920000 ;
      LAYER met4 ;
        RECT 62.600000 41.600000 62.920000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 42.030000 62.920000 42.350000 ;
      LAYER met4 ;
        RECT 62.600000 42.030000 62.920000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 42.460000 62.920000 42.780000 ;
      LAYER met4 ;
        RECT 62.600000 42.460000 62.920000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 42.890000 62.920000 43.210000 ;
      LAYER met4 ;
        RECT 62.600000 42.890000 62.920000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 43.320000 62.920000 43.640000 ;
      LAYER met4 ;
        RECT 62.600000 43.320000 62.920000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 43.750000 62.920000 44.070000 ;
      LAYER met4 ;
        RECT 62.600000 43.750000 62.920000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 44.180000 62.920000 44.500000 ;
      LAYER met4 ;
        RECT 62.600000 44.180000 62.920000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 44.610000 62.920000 44.930000 ;
      LAYER met4 ;
        RECT 62.600000 44.610000 62.920000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 45.040000 62.920000 45.360000 ;
      LAYER met4 ;
        RECT 62.600000 45.040000 62.920000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 45.470000 62.920000 45.790000 ;
      LAYER met4 ;
        RECT 62.600000 45.470000 62.920000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 45.900000 62.920000 46.220000 ;
      LAYER met4 ;
        RECT 62.600000 45.900000 62.920000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 41.600000 63.325000 41.920000 ;
      LAYER met4 ;
        RECT 63.005000 41.600000 63.325000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 42.030000 63.325000 42.350000 ;
      LAYER met4 ;
        RECT 63.005000 42.030000 63.325000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 42.460000 63.325000 42.780000 ;
      LAYER met4 ;
        RECT 63.005000 42.460000 63.325000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 42.890000 63.325000 43.210000 ;
      LAYER met4 ;
        RECT 63.005000 42.890000 63.325000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 43.320000 63.325000 43.640000 ;
      LAYER met4 ;
        RECT 63.005000 43.320000 63.325000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 43.750000 63.325000 44.070000 ;
      LAYER met4 ;
        RECT 63.005000 43.750000 63.325000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 44.180000 63.325000 44.500000 ;
      LAYER met4 ;
        RECT 63.005000 44.180000 63.325000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 44.610000 63.325000 44.930000 ;
      LAYER met4 ;
        RECT 63.005000 44.610000 63.325000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 45.040000 63.325000 45.360000 ;
      LAYER met4 ;
        RECT 63.005000 45.040000 63.325000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 45.470000 63.325000 45.790000 ;
      LAYER met4 ;
        RECT 63.005000 45.470000 63.325000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 45.900000 63.325000 46.220000 ;
      LAYER met4 ;
        RECT 63.005000 45.900000 63.325000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 41.600000 63.730000 41.920000 ;
      LAYER met4 ;
        RECT 63.410000 41.600000 63.730000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 42.030000 63.730000 42.350000 ;
      LAYER met4 ;
        RECT 63.410000 42.030000 63.730000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 42.460000 63.730000 42.780000 ;
      LAYER met4 ;
        RECT 63.410000 42.460000 63.730000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 42.890000 63.730000 43.210000 ;
      LAYER met4 ;
        RECT 63.410000 42.890000 63.730000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 43.320000 63.730000 43.640000 ;
      LAYER met4 ;
        RECT 63.410000 43.320000 63.730000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 43.750000 63.730000 44.070000 ;
      LAYER met4 ;
        RECT 63.410000 43.750000 63.730000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 44.180000 63.730000 44.500000 ;
      LAYER met4 ;
        RECT 63.410000 44.180000 63.730000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 44.610000 63.730000 44.930000 ;
      LAYER met4 ;
        RECT 63.410000 44.610000 63.730000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 45.040000 63.730000 45.360000 ;
      LAYER met4 ;
        RECT 63.410000 45.040000 63.730000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 45.470000 63.730000 45.790000 ;
      LAYER met4 ;
        RECT 63.410000 45.470000 63.730000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 45.900000 63.730000 46.220000 ;
      LAYER met4 ;
        RECT 63.410000 45.900000 63.730000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 41.600000 64.135000 41.920000 ;
      LAYER met4 ;
        RECT 63.815000 41.600000 64.135000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 42.030000 64.135000 42.350000 ;
      LAYER met4 ;
        RECT 63.815000 42.030000 64.135000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 42.460000 64.135000 42.780000 ;
      LAYER met4 ;
        RECT 63.815000 42.460000 64.135000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 42.890000 64.135000 43.210000 ;
      LAYER met4 ;
        RECT 63.815000 42.890000 64.135000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 43.320000 64.135000 43.640000 ;
      LAYER met4 ;
        RECT 63.815000 43.320000 64.135000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 43.750000 64.135000 44.070000 ;
      LAYER met4 ;
        RECT 63.815000 43.750000 64.135000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 44.180000 64.135000 44.500000 ;
      LAYER met4 ;
        RECT 63.815000 44.180000 64.135000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 44.610000 64.135000 44.930000 ;
      LAYER met4 ;
        RECT 63.815000 44.610000 64.135000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 45.040000 64.135000 45.360000 ;
      LAYER met4 ;
        RECT 63.815000 45.040000 64.135000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 45.470000 64.135000 45.790000 ;
      LAYER met4 ;
        RECT 63.815000 45.470000 64.135000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 45.900000 64.135000 46.220000 ;
      LAYER met4 ;
        RECT 63.815000 45.900000 64.135000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 41.600000 64.540000 41.920000 ;
      LAYER met4 ;
        RECT 64.220000 41.600000 64.540000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 42.030000 64.540000 42.350000 ;
      LAYER met4 ;
        RECT 64.220000 42.030000 64.540000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 42.460000 64.540000 42.780000 ;
      LAYER met4 ;
        RECT 64.220000 42.460000 64.540000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 42.890000 64.540000 43.210000 ;
      LAYER met4 ;
        RECT 64.220000 42.890000 64.540000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 43.320000 64.540000 43.640000 ;
      LAYER met4 ;
        RECT 64.220000 43.320000 64.540000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 43.750000 64.540000 44.070000 ;
      LAYER met4 ;
        RECT 64.220000 43.750000 64.540000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 44.180000 64.540000 44.500000 ;
      LAYER met4 ;
        RECT 64.220000 44.180000 64.540000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 44.610000 64.540000 44.930000 ;
      LAYER met4 ;
        RECT 64.220000 44.610000 64.540000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 45.040000 64.540000 45.360000 ;
      LAYER met4 ;
        RECT 64.220000 45.040000 64.540000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 45.470000 64.540000 45.790000 ;
      LAYER met4 ;
        RECT 64.220000 45.470000 64.540000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 45.900000 64.540000 46.220000 ;
      LAYER met4 ;
        RECT 64.220000 45.900000 64.540000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 41.600000 64.945000 41.920000 ;
      LAYER met4 ;
        RECT 64.625000 41.600000 64.945000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 42.030000 64.945000 42.350000 ;
      LAYER met4 ;
        RECT 64.625000 42.030000 64.945000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 42.460000 64.945000 42.780000 ;
      LAYER met4 ;
        RECT 64.625000 42.460000 64.945000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 42.890000 64.945000 43.210000 ;
      LAYER met4 ;
        RECT 64.625000 42.890000 64.945000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 43.320000 64.945000 43.640000 ;
      LAYER met4 ;
        RECT 64.625000 43.320000 64.945000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 43.750000 64.945000 44.070000 ;
      LAYER met4 ;
        RECT 64.625000 43.750000 64.945000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 44.180000 64.945000 44.500000 ;
      LAYER met4 ;
        RECT 64.625000 44.180000 64.945000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 44.610000 64.945000 44.930000 ;
      LAYER met4 ;
        RECT 64.625000 44.610000 64.945000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 45.040000 64.945000 45.360000 ;
      LAYER met4 ;
        RECT 64.625000 45.040000 64.945000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 45.470000 64.945000 45.790000 ;
      LAYER met4 ;
        RECT 64.625000 45.470000 64.945000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 45.900000 64.945000 46.220000 ;
      LAYER met4 ;
        RECT 64.625000 45.900000 64.945000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 41.600000 65.350000 41.920000 ;
      LAYER met4 ;
        RECT 65.030000 41.600000 65.350000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 42.030000 65.350000 42.350000 ;
      LAYER met4 ;
        RECT 65.030000 42.030000 65.350000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 42.460000 65.350000 42.780000 ;
      LAYER met4 ;
        RECT 65.030000 42.460000 65.350000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 42.890000 65.350000 43.210000 ;
      LAYER met4 ;
        RECT 65.030000 42.890000 65.350000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 43.320000 65.350000 43.640000 ;
      LAYER met4 ;
        RECT 65.030000 43.320000 65.350000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 43.750000 65.350000 44.070000 ;
      LAYER met4 ;
        RECT 65.030000 43.750000 65.350000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 44.180000 65.350000 44.500000 ;
      LAYER met4 ;
        RECT 65.030000 44.180000 65.350000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 44.610000 65.350000 44.930000 ;
      LAYER met4 ;
        RECT 65.030000 44.610000 65.350000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 45.040000 65.350000 45.360000 ;
      LAYER met4 ;
        RECT 65.030000 45.040000 65.350000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 45.470000 65.350000 45.790000 ;
      LAYER met4 ;
        RECT 65.030000 45.470000 65.350000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 45.900000 65.350000 46.220000 ;
      LAYER met4 ;
        RECT 65.030000 45.900000 65.350000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 41.600000 65.755000 41.920000 ;
      LAYER met4 ;
        RECT 65.435000 41.600000 65.755000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 42.030000 65.755000 42.350000 ;
      LAYER met4 ;
        RECT 65.435000 42.030000 65.755000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 42.460000 65.755000 42.780000 ;
      LAYER met4 ;
        RECT 65.435000 42.460000 65.755000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 42.890000 65.755000 43.210000 ;
      LAYER met4 ;
        RECT 65.435000 42.890000 65.755000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 43.320000 65.755000 43.640000 ;
      LAYER met4 ;
        RECT 65.435000 43.320000 65.755000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 43.750000 65.755000 44.070000 ;
      LAYER met4 ;
        RECT 65.435000 43.750000 65.755000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 44.180000 65.755000 44.500000 ;
      LAYER met4 ;
        RECT 65.435000 44.180000 65.755000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 44.610000 65.755000 44.930000 ;
      LAYER met4 ;
        RECT 65.435000 44.610000 65.755000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 45.040000 65.755000 45.360000 ;
      LAYER met4 ;
        RECT 65.435000 45.040000 65.755000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 45.470000 65.755000 45.790000 ;
      LAYER met4 ;
        RECT 65.435000 45.470000 65.755000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 45.900000 65.755000 46.220000 ;
      LAYER met4 ;
        RECT 65.435000 45.900000 65.755000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 41.600000 66.160000 41.920000 ;
      LAYER met4 ;
        RECT 65.840000 41.600000 66.160000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 42.030000 66.160000 42.350000 ;
      LAYER met4 ;
        RECT 65.840000 42.030000 66.160000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 42.460000 66.160000 42.780000 ;
      LAYER met4 ;
        RECT 65.840000 42.460000 66.160000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 42.890000 66.160000 43.210000 ;
      LAYER met4 ;
        RECT 65.840000 42.890000 66.160000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 43.320000 66.160000 43.640000 ;
      LAYER met4 ;
        RECT 65.840000 43.320000 66.160000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 43.750000 66.160000 44.070000 ;
      LAYER met4 ;
        RECT 65.840000 43.750000 66.160000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 44.180000 66.160000 44.500000 ;
      LAYER met4 ;
        RECT 65.840000 44.180000 66.160000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 44.610000 66.160000 44.930000 ;
      LAYER met4 ;
        RECT 65.840000 44.610000 66.160000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 45.040000 66.160000 45.360000 ;
      LAYER met4 ;
        RECT 65.840000 45.040000 66.160000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 45.470000 66.160000 45.790000 ;
      LAYER met4 ;
        RECT 65.840000 45.470000 66.160000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 45.900000 66.160000 46.220000 ;
      LAYER met4 ;
        RECT 65.840000 45.900000 66.160000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 41.600000 66.565000 41.920000 ;
      LAYER met4 ;
        RECT 66.245000 41.600000 66.565000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 42.030000 66.565000 42.350000 ;
      LAYER met4 ;
        RECT 66.245000 42.030000 66.565000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 42.460000 66.565000 42.780000 ;
      LAYER met4 ;
        RECT 66.245000 42.460000 66.565000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 42.890000 66.565000 43.210000 ;
      LAYER met4 ;
        RECT 66.245000 42.890000 66.565000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 43.320000 66.565000 43.640000 ;
      LAYER met4 ;
        RECT 66.245000 43.320000 66.565000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 43.750000 66.565000 44.070000 ;
      LAYER met4 ;
        RECT 66.245000 43.750000 66.565000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 44.180000 66.565000 44.500000 ;
      LAYER met4 ;
        RECT 66.245000 44.180000 66.565000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 44.610000 66.565000 44.930000 ;
      LAYER met4 ;
        RECT 66.245000 44.610000 66.565000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 45.040000 66.565000 45.360000 ;
      LAYER met4 ;
        RECT 66.245000 45.040000 66.565000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 45.470000 66.565000 45.790000 ;
      LAYER met4 ;
        RECT 66.245000 45.470000 66.565000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 45.900000 66.565000 46.220000 ;
      LAYER met4 ;
        RECT 66.245000 45.900000 66.565000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 41.600000 66.970000 41.920000 ;
      LAYER met4 ;
        RECT 66.650000 41.600000 66.970000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 42.030000 66.970000 42.350000 ;
      LAYER met4 ;
        RECT 66.650000 42.030000 66.970000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 42.460000 66.970000 42.780000 ;
      LAYER met4 ;
        RECT 66.650000 42.460000 66.970000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 42.890000 66.970000 43.210000 ;
      LAYER met4 ;
        RECT 66.650000 42.890000 66.970000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 43.320000 66.970000 43.640000 ;
      LAYER met4 ;
        RECT 66.650000 43.320000 66.970000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 43.750000 66.970000 44.070000 ;
      LAYER met4 ;
        RECT 66.650000 43.750000 66.970000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 44.180000 66.970000 44.500000 ;
      LAYER met4 ;
        RECT 66.650000 44.180000 66.970000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 44.610000 66.970000 44.930000 ;
      LAYER met4 ;
        RECT 66.650000 44.610000 66.970000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 45.040000 66.970000 45.360000 ;
      LAYER met4 ;
        RECT 66.650000 45.040000 66.970000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 45.470000 66.970000 45.790000 ;
      LAYER met4 ;
        RECT 66.650000 45.470000 66.970000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 45.900000 66.970000 46.220000 ;
      LAYER met4 ;
        RECT 66.650000 45.900000 66.970000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 41.600000 67.375000 41.920000 ;
      LAYER met4 ;
        RECT 67.055000 41.600000 67.375000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 42.030000 67.375000 42.350000 ;
      LAYER met4 ;
        RECT 67.055000 42.030000 67.375000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 42.460000 67.375000 42.780000 ;
      LAYER met4 ;
        RECT 67.055000 42.460000 67.375000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 42.890000 67.375000 43.210000 ;
      LAYER met4 ;
        RECT 67.055000 42.890000 67.375000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 43.320000 67.375000 43.640000 ;
      LAYER met4 ;
        RECT 67.055000 43.320000 67.375000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 43.750000 67.375000 44.070000 ;
      LAYER met4 ;
        RECT 67.055000 43.750000 67.375000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 44.180000 67.375000 44.500000 ;
      LAYER met4 ;
        RECT 67.055000 44.180000 67.375000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 44.610000 67.375000 44.930000 ;
      LAYER met4 ;
        RECT 67.055000 44.610000 67.375000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 45.040000 67.375000 45.360000 ;
      LAYER met4 ;
        RECT 67.055000 45.040000 67.375000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 45.470000 67.375000 45.790000 ;
      LAYER met4 ;
        RECT 67.055000 45.470000 67.375000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 45.900000 67.375000 46.220000 ;
      LAYER met4 ;
        RECT 67.055000 45.900000 67.375000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 41.600000 67.780000 41.920000 ;
      LAYER met4 ;
        RECT 67.460000 41.600000 67.780000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 42.030000 67.780000 42.350000 ;
      LAYER met4 ;
        RECT 67.460000 42.030000 67.780000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 42.460000 67.780000 42.780000 ;
      LAYER met4 ;
        RECT 67.460000 42.460000 67.780000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 42.890000 67.780000 43.210000 ;
      LAYER met4 ;
        RECT 67.460000 42.890000 67.780000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 43.320000 67.780000 43.640000 ;
      LAYER met4 ;
        RECT 67.460000 43.320000 67.780000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 43.750000 67.780000 44.070000 ;
      LAYER met4 ;
        RECT 67.460000 43.750000 67.780000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 44.180000 67.780000 44.500000 ;
      LAYER met4 ;
        RECT 67.460000 44.180000 67.780000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 44.610000 67.780000 44.930000 ;
      LAYER met4 ;
        RECT 67.460000 44.610000 67.780000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 45.040000 67.780000 45.360000 ;
      LAYER met4 ;
        RECT 67.460000 45.040000 67.780000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 45.470000 67.780000 45.790000 ;
      LAYER met4 ;
        RECT 67.460000 45.470000 67.780000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 45.900000 67.780000 46.220000 ;
      LAYER met4 ;
        RECT 67.460000 45.900000 67.780000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 41.600000 68.185000 41.920000 ;
      LAYER met4 ;
        RECT 67.865000 41.600000 68.185000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 42.030000 68.185000 42.350000 ;
      LAYER met4 ;
        RECT 67.865000 42.030000 68.185000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 42.460000 68.185000 42.780000 ;
      LAYER met4 ;
        RECT 67.865000 42.460000 68.185000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 42.890000 68.185000 43.210000 ;
      LAYER met4 ;
        RECT 67.865000 42.890000 68.185000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 43.320000 68.185000 43.640000 ;
      LAYER met4 ;
        RECT 67.865000 43.320000 68.185000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 43.750000 68.185000 44.070000 ;
      LAYER met4 ;
        RECT 67.865000 43.750000 68.185000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 44.180000 68.185000 44.500000 ;
      LAYER met4 ;
        RECT 67.865000 44.180000 68.185000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 44.610000 68.185000 44.930000 ;
      LAYER met4 ;
        RECT 67.865000 44.610000 68.185000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 45.040000 68.185000 45.360000 ;
      LAYER met4 ;
        RECT 67.865000 45.040000 68.185000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 45.470000 68.185000 45.790000 ;
      LAYER met4 ;
        RECT 67.865000 45.470000 68.185000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 45.900000 68.185000 46.220000 ;
      LAYER met4 ;
        RECT 67.865000 45.900000 68.185000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 41.600000 68.590000 41.920000 ;
      LAYER met4 ;
        RECT 68.270000 41.600000 68.590000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 42.030000 68.590000 42.350000 ;
      LAYER met4 ;
        RECT 68.270000 42.030000 68.590000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 42.460000 68.590000 42.780000 ;
      LAYER met4 ;
        RECT 68.270000 42.460000 68.590000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 42.890000 68.590000 43.210000 ;
      LAYER met4 ;
        RECT 68.270000 42.890000 68.590000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 43.320000 68.590000 43.640000 ;
      LAYER met4 ;
        RECT 68.270000 43.320000 68.590000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 43.750000 68.590000 44.070000 ;
      LAYER met4 ;
        RECT 68.270000 43.750000 68.590000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 44.180000 68.590000 44.500000 ;
      LAYER met4 ;
        RECT 68.270000 44.180000 68.590000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 44.610000 68.590000 44.930000 ;
      LAYER met4 ;
        RECT 68.270000 44.610000 68.590000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 45.040000 68.590000 45.360000 ;
      LAYER met4 ;
        RECT 68.270000 45.040000 68.590000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 45.470000 68.590000 45.790000 ;
      LAYER met4 ;
        RECT 68.270000 45.470000 68.590000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 45.900000 68.590000 46.220000 ;
      LAYER met4 ;
        RECT 68.270000 45.900000 68.590000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 41.600000 68.995000 41.920000 ;
      LAYER met4 ;
        RECT 68.675000 41.600000 68.995000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 42.030000 68.995000 42.350000 ;
      LAYER met4 ;
        RECT 68.675000 42.030000 68.995000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 42.460000 68.995000 42.780000 ;
      LAYER met4 ;
        RECT 68.675000 42.460000 68.995000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 42.890000 68.995000 43.210000 ;
      LAYER met4 ;
        RECT 68.675000 42.890000 68.995000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 43.320000 68.995000 43.640000 ;
      LAYER met4 ;
        RECT 68.675000 43.320000 68.995000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 43.750000 68.995000 44.070000 ;
      LAYER met4 ;
        RECT 68.675000 43.750000 68.995000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 44.180000 68.995000 44.500000 ;
      LAYER met4 ;
        RECT 68.675000 44.180000 68.995000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 44.610000 68.995000 44.930000 ;
      LAYER met4 ;
        RECT 68.675000 44.610000 68.995000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 45.040000 68.995000 45.360000 ;
      LAYER met4 ;
        RECT 68.675000 45.040000 68.995000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 45.470000 68.995000 45.790000 ;
      LAYER met4 ;
        RECT 68.675000 45.470000 68.995000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 45.900000 68.995000 46.220000 ;
      LAYER met4 ;
        RECT 68.675000 45.900000 68.995000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 41.600000 69.400000 41.920000 ;
      LAYER met4 ;
        RECT 69.080000 41.600000 69.400000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 42.030000 69.400000 42.350000 ;
      LAYER met4 ;
        RECT 69.080000 42.030000 69.400000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 42.460000 69.400000 42.780000 ;
      LAYER met4 ;
        RECT 69.080000 42.460000 69.400000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 42.890000 69.400000 43.210000 ;
      LAYER met4 ;
        RECT 69.080000 42.890000 69.400000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 43.320000 69.400000 43.640000 ;
      LAYER met4 ;
        RECT 69.080000 43.320000 69.400000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 43.750000 69.400000 44.070000 ;
      LAYER met4 ;
        RECT 69.080000 43.750000 69.400000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 44.180000 69.400000 44.500000 ;
      LAYER met4 ;
        RECT 69.080000 44.180000 69.400000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 44.610000 69.400000 44.930000 ;
      LAYER met4 ;
        RECT 69.080000 44.610000 69.400000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 45.040000 69.400000 45.360000 ;
      LAYER met4 ;
        RECT 69.080000 45.040000 69.400000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 45.470000 69.400000 45.790000 ;
      LAYER met4 ;
        RECT 69.080000 45.470000 69.400000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 45.900000 69.400000 46.220000 ;
      LAYER met4 ;
        RECT 69.080000 45.900000 69.400000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 41.600000 69.805000 41.920000 ;
      LAYER met4 ;
        RECT 69.485000 41.600000 69.805000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 42.030000 69.805000 42.350000 ;
      LAYER met4 ;
        RECT 69.485000 42.030000 69.805000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 42.460000 69.805000 42.780000 ;
      LAYER met4 ;
        RECT 69.485000 42.460000 69.805000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 42.890000 69.805000 43.210000 ;
      LAYER met4 ;
        RECT 69.485000 42.890000 69.805000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 43.320000 69.805000 43.640000 ;
      LAYER met4 ;
        RECT 69.485000 43.320000 69.805000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 43.750000 69.805000 44.070000 ;
      LAYER met4 ;
        RECT 69.485000 43.750000 69.805000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 44.180000 69.805000 44.500000 ;
      LAYER met4 ;
        RECT 69.485000 44.180000 69.805000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 44.610000 69.805000 44.930000 ;
      LAYER met4 ;
        RECT 69.485000 44.610000 69.805000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 45.040000 69.805000 45.360000 ;
      LAYER met4 ;
        RECT 69.485000 45.040000 69.805000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 45.470000 69.805000 45.790000 ;
      LAYER met4 ;
        RECT 69.485000 45.470000 69.805000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 45.900000 69.805000 46.220000 ;
      LAYER met4 ;
        RECT 69.485000 45.900000 69.805000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 41.600000 70.210000 41.920000 ;
      LAYER met4 ;
        RECT 69.890000 41.600000 70.210000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 42.030000 70.210000 42.350000 ;
      LAYER met4 ;
        RECT 69.890000 42.030000 70.210000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 42.460000 70.210000 42.780000 ;
      LAYER met4 ;
        RECT 69.890000 42.460000 70.210000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 42.890000 70.210000 43.210000 ;
      LAYER met4 ;
        RECT 69.890000 42.890000 70.210000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 43.320000 70.210000 43.640000 ;
      LAYER met4 ;
        RECT 69.890000 43.320000 70.210000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 43.750000 70.210000 44.070000 ;
      LAYER met4 ;
        RECT 69.890000 43.750000 70.210000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 44.180000 70.210000 44.500000 ;
      LAYER met4 ;
        RECT 69.890000 44.180000 70.210000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 44.610000 70.210000 44.930000 ;
      LAYER met4 ;
        RECT 69.890000 44.610000 70.210000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 45.040000 70.210000 45.360000 ;
      LAYER met4 ;
        RECT 69.890000 45.040000 70.210000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 45.470000 70.210000 45.790000 ;
      LAYER met4 ;
        RECT 69.890000 45.470000 70.210000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 45.900000 70.210000 46.220000 ;
      LAYER met4 ;
        RECT 69.890000 45.900000 70.210000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075000 41.600000 7.395000 41.920000 ;
      LAYER met4 ;
        RECT 7.075000 41.600000 7.395000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075000 42.030000 7.395000 42.350000 ;
      LAYER met4 ;
        RECT 7.075000 42.030000 7.395000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075000 42.460000 7.395000 42.780000 ;
      LAYER met4 ;
        RECT 7.075000 42.460000 7.395000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075000 42.890000 7.395000 43.210000 ;
      LAYER met4 ;
        RECT 7.075000 42.890000 7.395000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075000 43.320000 7.395000 43.640000 ;
      LAYER met4 ;
        RECT 7.075000 43.320000 7.395000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075000 43.750000 7.395000 44.070000 ;
      LAYER met4 ;
        RECT 7.075000 43.750000 7.395000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075000 44.180000 7.395000 44.500000 ;
      LAYER met4 ;
        RECT 7.075000 44.180000 7.395000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075000 44.610000 7.395000 44.930000 ;
      LAYER met4 ;
        RECT 7.075000 44.610000 7.395000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075000 45.040000 7.395000 45.360000 ;
      LAYER met4 ;
        RECT 7.075000 45.040000 7.395000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075000 45.470000 7.395000 45.790000 ;
      LAYER met4 ;
        RECT 7.075000 45.470000 7.395000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075000 45.900000 7.395000 46.220000 ;
      LAYER met4 ;
        RECT 7.075000 45.900000 7.395000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480000 41.600000 7.800000 41.920000 ;
      LAYER met4 ;
        RECT 7.480000 41.600000 7.800000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480000 42.030000 7.800000 42.350000 ;
      LAYER met4 ;
        RECT 7.480000 42.030000 7.800000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480000 42.460000 7.800000 42.780000 ;
      LAYER met4 ;
        RECT 7.480000 42.460000 7.800000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480000 42.890000 7.800000 43.210000 ;
      LAYER met4 ;
        RECT 7.480000 42.890000 7.800000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480000 43.320000 7.800000 43.640000 ;
      LAYER met4 ;
        RECT 7.480000 43.320000 7.800000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480000 43.750000 7.800000 44.070000 ;
      LAYER met4 ;
        RECT 7.480000 43.750000 7.800000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480000 44.180000 7.800000 44.500000 ;
      LAYER met4 ;
        RECT 7.480000 44.180000 7.800000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480000 44.610000 7.800000 44.930000 ;
      LAYER met4 ;
        RECT 7.480000 44.610000 7.800000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480000 45.040000 7.800000 45.360000 ;
      LAYER met4 ;
        RECT 7.480000 45.040000 7.800000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480000 45.470000 7.800000 45.790000 ;
      LAYER met4 ;
        RECT 7.480000 45.470000 7.800000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480000 45.900000 7.800000 46.220000 ;
      LAYER met4 ;
        RECT 7.480000 45.900000 7.800000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 41.600000 8.205000 41.920000 ;
      LAYER met4 ;
        RECT 7.885000 41.600000 8.205000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 42.030000 8.205000 42.350000 ;
      LAYER met4 ;
        RECT 7.885000 42.030000 8.205000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 42.460000 8.205000 42.780000 ;
      LAYER met4 ;
        RECT 7.885000 42.460000 8.205000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 42.890000 8.205000 43.210000 ;
      LAYER met4 ;
        RECT 7.885000 42.890000 8.205000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 43.320000 8.205000 43.640000 ;
      LAYER met4 ;
        RECT 7.885000 43.320000 8.205000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 43.750000 8.205000 44.070000 ;
      LAYER met4 ;
        RECT 7.885000 43.750000 8.205000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 44.180000 8.205000 44.500000 ;
      LAYER met4 ;
        RECT 7.885000 44.180000 8.205000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 44.610000 8.205000 44.930000 ;
      LAYER met4 ;
        RECT 7.885000 44.610000 8.205000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 45.040000 8.205000 45.360000 ;
      LAYER met4 ;
        RECT 7.885000 45.040000 8.205000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 45.470000 8.205000 45.790000 ;
      LAYER met4 ;
        RECT 7.885000 45.470000 8.205000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 45.900000 8.205000 46.220000 ;
      LAYER met4 ;
        RECT 7.885000 45.900000 8.205000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 41.600000 70.615000 41.920000 ;
      LAYER met4 ;
        RECT 70.295000 41.600000 70.615000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 42.030000 70.615000 42.350000 ;
      LAYER met4 ;
        RECT 70.295000 42.030000 70.615000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 42.460000 70.615000 42.780000 ;
      LAYER met4 ;
        RECT 70.295000 42.460000 70.615000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 42.890000 70.615000 43.210000 ;
      LAYER met4 ;
        RECT 70.295000 42.890000 70.615000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 43.320000 70.615000 43.640000 ;
      LAYER met4 ;
        RECT 70.295000 43.320000 70.615000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 43.750000 70.615000 44.070000 ;
      LAYER met4 ;
        RECT 70.295000 43.750000 70.615000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 44.180000 70.615000 44.500000 ;
      LAYER met4 ;
        RECT 70.295000 44.180000 70.615000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 44.610000 70.615000 44.930000 ;
      LAYER met4 ;
        RECT 70.295000 44.610000 70.615000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 45.040000 70.615000 45.360000 ;
      LAYER met4 ;
        RECT 70.295000 45.040000 70.615000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 45.470000 70.615000 45.790000 ;
      LAYER met4 ;
        RECT 70.295000 45.470000 70.615000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 45.900000 70.615000 46.220000 ;
      LAYER met4 ;
        RECT 70.295000 45.900000 70.615000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 41.600000 71.020000 41.920000 ;
      LAYER met4 ;
        RECT 70.700000 41.600000 71.020000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 42.030000 71.020000 42.350000 ;
      LAYER met4 ;
        RECT 70.700000 42.030000 71.020000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 42.460000 71.020000 42.780000 ;
      LAYER met4 ;
        RECT 70.700000 42.460000 71.020000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 42.890000 71.020000 43.210000 ;
      LAYER met4 ;
        RECT 70.700000 42.890000 71.020000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 43.320000 71.020000 43.640000 ;
      LAYER met4 ;
        RECT 70.700000 43.320000 71.020000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 43.750000 71.020000 44.070000 ;
      LAYER met4 ;
        RECT 70.700000 43.750000 71.020000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 44.180000 71.020000 44.500000 ;
      LAYER met4 ;
        RECT 70.700000 44.180000 71.020000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 44.610000 71.020000 44.930000 ;
      LAYER met4 ;
        RECT 70.700000 44.610000 71.020000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 45.040000 71.020000 45.360000 ;
      LAYER met4 ;
        RECT 70.700000 45.040000 71.020000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 45.470000 71.020000 45.790000 ;
      LAYER met4 ;
        RECT 70.700000 45.470000 71.020000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 45.900000 71.020000 46.220000 ;
      LAYER met4 ;
        RECT 70.700000 45.900000 71.020000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 41.600000 71.425000 41.920000 ;
      LAYER met4 ;
        RECT 71.105000 41.600000 71.425000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 42.030000 71.425000 42.350000 ;
      LAYER met4 ;
        RECT 71.105000 42.030000 71.425000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 42.460000 71.425000 42.780000 ;
      LAYER met4 ;
        RECT 71.105000 42.460000 71.425000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 42.890000 71.425000 43.210000 ;
      LAYER met4 ;
        RECT 71.105000 42.890000 71.425000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 43.320000 71.425000 43.640000 ;
      LAYER met4 ;
        RECT 71.105000 43.320000 71.425000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 43.750000 71.425000 44.070000 ;
      LAYER met4 ;
        RECT 71.105000 43.750000 71.425000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 44.180000 71.425000 44.500000 ;
      LAYER met4 ;
        RECT 71.105000 44.180000 71.425000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 44.610000 71.425000 44.930000 ;
      LAYER met4 ;
        RECT 71.105000 44.610000 71.425000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 45.040000 71.425000 45.360000 ;
      LAYER met4 ;
        RECT 71.105000 45.040000 71.425000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 45.470000 71.425000 45.790000 ;
      LAYER met4 ;
        RECT 71.105000 45.470000 71.425000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 45.900000 71.425000 46.220000 ;
      LAYER met4 ;
        RECT 71.105000 45.900000 71.425000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 41.600000 71.830000 41.920000 ;
      LAYER met4 ;
        RECT 71.510000 41.600000 71.830000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 42.030000 71.830000 42.350000 ;
      LAYER met4 ;
        RECT 71.510000 42.030000 71.830000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 42.460000 71.830000 42.780000 ;
      LAYER met4 ;
        RECT 71.510000 42.460000 71.830000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 42.890000 71.830000 43.210000 ;
      LAYER met4 ;
        RECT 71.510000 42.890000 71.830000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 43.320000 71.830000 43.640000 ;
      LAYER met4 ;
        RECT 71.510000 43.320000 71.830000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 43.750000 71.830000 44.070000 ;
      LAYER met4 ;
        RECT 71.510000 43.750000 71.830000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 44.180000 71.830000 44.500000 ;
      LAYER met4 ;
        RECT 71.510000 44.180000 71.830000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 44.610000 71.830000 44.930000 ;
      LAYER met4 ;
        RECT 71.510000 44.610000 71.830000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 45.040000 71.830000 45.360000 ;
      LAYER met4 ;
        RECT 71.510000 45.040000 71.830000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 45.470000 71.830000 45.790000 ;
      LAYER met4 ;
        RECT 71.510000 45.470000 71.830000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 45.900000 71.830000 46.220000 ;
      LAYER met4 ;
        RECT 71.510000 45.900000 71.830000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 41.600000 72.235000 41.920000 ;
      LAYER met4 ;
        RECT 71.915000 41.600000 72.235000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 42.030000 72.235000 42.350000 ;
      LAYER met4 ;
        RECT 71.915000 42.030000 72.235000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 42.460000 72.235000 42.780000 ;
      LAYER met4 ;
        RECT 71.915000 42.460000 72.235000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 42.890000 72.235000 43.210000 ;
      LAYER met4 ;
        RECT 71.915000 42.890000 72.235000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 43.320000 72.235000 43.640000 ;
      LAYER met4 ;
        RECT 71.915000 43.320000 72.235000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 43.750000 72.235000 44.070000 ;
      LAYER met4 ;
        RECT 71.915000 43.750000 72.235000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 44.180000 72.235000 44.500000 ;
      LAYER met4 ;
        RECT 71.915000 44.180000 72.235000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 44.610000 72.235000 44.930000 ;
      LAYER met4 ;
        RECT 71.915000 44.610000 72.235000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 45.040000 72.235000 45.360000 ;
      LAYER met4 ;
        RECT 71.915000 45.040000 72.235000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 45.470000 72.235000 45.790000 ;
      LAYER met4 ;
        RECT 71.915000 45.470000 72.235000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 45.900000 72.235000 46.220000 ;
      LAYER met4 ;
        RECT 71.915000 45.900000 72.235000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 41.600000 72.640000 41.920000 ;
      LAYER met4 ;
        RECT 72.320000 41.600000 72.640000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 42.030000 72.640000 42.350000 ;
      LAYER met4 ;
        RECT 72.320000 42.030000 72.640000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 42.460000 72.640000 42.780000 ;
      LAYER met4 ;
        RECT 72.320000 42.460000 72.640000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 42.890000 72.640000 43.210000 ;
      LAYER met4 ;
        RECT 72.320000 42.890000 72.640000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 43.320000 72.640000 43.640000 ;
      LAYER met4 ;
        RECT 72.320000 43.320000 72.640000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 43.750000 72.640000 44.070000 ;
      LAYER met4 ;
        RECT 72.320000 43.750000 72.640000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 44.180000 72.640000 44.500000 ;
      LAYER met4 ;
        RECT 72.320000 44.180000 72.640000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 44.610000 72.640000 44.930000 ;
      LAYER met4 ;
        RECT 72.320000 44.610000 72.640000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 45.040000 72.640000 45.360000 ;
      LAYER met4 ;
        RECT 72.320000 45.040000 72.640000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 45.470000 72.640000 45.790000 ;
      LAYER met4 ;
        RECT 72.320000 45.470000 72.640000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 45.900000 72.640000 46.220000 ;
      LAYER met4 ;
        RECT 72.320000 45.900000 72.640000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 41.600000 73.045000 41.920000 ;
      LAYER met4 ;
        RECT 72.725000 41.600000 73.045000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 42.030000 73.045000 42.350000 ;
      LAYER met4 ;
        RECT 72.725000 42.030000 73.045000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 42.460000 73.045000 42.780000 ;
      LAYER met4 ;
        RECT 72.725000 42.460000 73.045000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 42.890000 73.045000 43.210000 ;
      LAYER met4 ;
        RECT 72.725000 42.890000 73.045000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 43.320000 73.045000 43.640000 ;
      LAYER met4 ;
        RECT 72.725000 43.320000 73.045000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 43.750000 73.045000 44.070000 ;
      LAYER met4 ;
        RECT 72.725000 43.750000 73.045000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 44.180000 73.045000 44.500000 ;
      LAYER met4 ;
        RECT 72.725000 44.180000 73.045000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 44.610000 73.045000 44.930000 ;
      LAYER met4 ;
        RECT 72.725000 44.610000 73.045000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 45.040000 73.045000 45.360000 ;
      LAYER met4 ;
        RECT 72.725000 45.040000 73.045000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 45.470000 73.045000 45.790000 ;
      LAYER met4 ;
        RECT 72.725000 45.470000 73.045000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 45.900000 73.045000 46.220000 ;
      LAYER met4 ;
        RECT 72.725000 45.900000 73.045000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 41.600000 73.450000 41.920000 ;
      LAYER met4 ;
        RECT 73.130000 41.600000 73.450000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 42.030000 73.450000 42.350000 ;
      LAYER met4 ;
        RECT 73.130000 42.030000 73.450000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 42.460000 73.450000 42.780000 ;
      LAYER met4 ;
        RECT 73.130000 42.460000 73.450000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 42.890000 73.450000 43.210000 ;
      LAYER met4 ;
        RECT 73.130000 42.890000 73.450000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 43.320000 73.450000 43.640000 ;
      LAYER met4 ;
        RECT 73.130000 43.320000 73.450000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 43.750000 73.450000 44.070000 ;
      LAYER met4 ;
        RECT 73.130000 43.750000 73.450000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 44.180000 73.450000 44.500000 ;
      LAYER met4 ;
        RECT 73.130000 44.180000 73.450000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 44.610000 73.450000 44.930000 ;
      LAYER met4 ;
        RECT 73.130000 44.610000 73.450000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 45.040000 73.450000 45.360000 ;
      LAYER met4 ;
        RECT 73.130000 45.040000 73.450000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 45.470000 73.450000 45.790000 ;
      LAYER met4 ;
        RECT 73.130000 45.470000 73.450000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 45.900000 73.450000 46.220000 ;
      LAYER met4 ;
        RECT 73.130000 45.900000 73.450000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 41.600000 73.855000 41.920000 ;
      LAYER met4 ;
        RECT 73.535000 41.600000 73.855000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 42.030000 73.855000 42.350000 ;
      LAYER met4 ;
        RECT 73.535000 42.030000 73.855000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 42.460000 73.855000 42.780000 ;
      LAYER met4 ;
        RECT 73.535000 42.460000 73.855000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 42.890000 73.855000 43.210000 ;
      LAYER met4 ;
        RECT 73.535000 42.890000 73.855000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 43.320000 73.855000 43.640000 ;
      LAYER met4 ;
        RECT 73.535000 43.320000 73.855000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 43.750000 73.855000 44.070000 ;
      LAYER met4 ;
        RECT 73.535000 43.750000 73.855000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 44.180000 73.855000 44.500000 ;
      LAYER met4 ;
        RECT 73.535000 44.180000 73.855000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 44.610000 73.855000 44.930000 ;
      LAYER met4 ;
        RECT 73.535000 44.610000 73.855000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 45.040000 73.855000 45.360000 ;
      LAYER met4 ;
        RECT 73.535000 45.040000 73.855000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 45.470000 73.855000 45.790000 ;
      LAYER met4 ;
        RECT 73.535000 45.470000 73.855000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 45.900000 73.855000 46.220000 ;
      LAYER met4 ;
        RECT 73.535000 45.900000 73.855000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 41.600000 74.260000 41.920000 ;
      LAYER met4 ;
        RECT 73.940000 41.600000 74.260000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 42.030000 74.260000 42.350000 ;
      LAYER met4 ;
        RECT 73.940000 42.030000 74.260000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 42.460000 74.260000 42.780000 ;
      LAYER met4 ;
        RECT 73.940000 42.460000 74.260000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 42.890000 74.260000 43.210000 ;
      LAYER met4 ;
        RECT 73.940000 42.890000 74.260000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 43.320000 74.260000 43.640000 ;
      LAYER met4 ;
        RECT 73.940000 43.320000 74.260000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 43.750000 74.260000 44.070000 ;
      LAYER met4 ;
        RECT 73.940000 43.750000 74.260000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 44.180000 74.260000 44.500000 ;
      LAYER met4 ;
        RECT 73.940000 44.180000 74.260000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 44.610000 74.260000 44.930000 ;
      LAYER met4 ;
        RECT 73.940000 44.610000 74.260000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 45.040000 74.260000 45.360000 ;
      LAYER met4 ;
        RECT 73.940000 45.040000 74.260000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 45.470000 74.260000 45.790000 ;
      LAYER met4 ;
        RECT 73.940000 45.470000 74.260000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 45.900000 74.260000 46.220000 ;
      LAYER met4 ;
        RECT 73.940000 45.900000 74.260000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290000 41.600000 8.610000 41.920000 ;
      LAYER met4 ;
        RECT 8.290000 41.600000 8.610000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290000 42.030000 8.610000 42.350000 ;
      LAYER met4 ;
        RECT 8.290000 42.030000 8.610000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290000 42.460000 8.610000 42.780000 ;
      LAYER met4 ;
        RECT 8.290000 42.460000 8.610000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290000 42.890000 8.610000 43.210000 ;
      LAYER met4 ;
        RECT 8.290000 42.890000 8.610000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290000 43.320000 8.610000 43.640000 ;
      LAYER met4 ;
        RECT 8.290000 43.320000 8.610000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290000 43.750000 8.610000 44.070000 ;
      LAYER met4 ;
        RECT 8.290000 43.750000 8.610000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290000 44.180000 8.610000 44.500000 ;
      LAYER met4 ;
        RECT 8.290000 44.180000 8.610000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290000 44.610000 8.610000 44.930000 ;
      LAYER met4 ;
        RECT 8.290000 44.610000 8.610000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290000 45.040000 8.610000 45.360000 ;
      LAYER met4 ;
        RECT 8.290000 45.040000 8.610000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290000 45.470000 8.610000 45.790000 ;
      LAYER met4 ;
        RECT 8.290000 45.470000 8.610000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290000 45.900000 8.610000 46.220000 ;
      LAYER met4 ;
        RECT 8.290000 45.900000 8.610000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695000 41.600000 9.015000 41.920000 ;
      LAYER met4 ;
        RECT 8.695000 41.600000 9.015000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695000 42.030000 9.015000 42.350000 ;
      LAYER met4 ;
        RECT 8.695000 42.030000 9.015000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695000 42.460000 9.015000 42.780000 ;
      LAYER met4 ;
        RECT 8.695000 42.460000 9.015000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695000 42.890000 9.015000 43.210000 ;
      LAYER met4 ;
        RECT 8.695000 42.890000 9.015000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695000 43.320000 9.015000 43.640000 ;
      LAYER met4 ;
        RECT 8.695000 43.320000 9.015000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695000 43.750000 9.015000 44.070000 ;
      LAYER met4 ;
        RECT 8.695000 43.750000 9.015000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695000 44.180000 9.015000 44.500000 ;
      LAYER met4 ;
        RECT 8.695000 44.180000 9.015000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695000 44.610000 9.015000 44.930000 ;
      LAYER met4 ;
        RECT 8.695000 44.610000 9.015000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695000 45.040000 9.015000 45.360000 ;
      LAYER met4 ;
        RECT 8.695000 45.040000 9.015000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695000 45.470000 9.015000 45.790000 ;
      LAYER met4 ;
        RECT 8.695000 45.470000 9.015000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695000 45.900000 9.015000 46.220000 ;
      LAYER met4 ;
        RECT 8.695000 45.900000 9.015000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100000 41.600000 9.420000 41.920000 ;
      LAYER met4 ;
        RECT 9.100000 41.600000 9.420000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100000 42.030000 9.420000 42.350000 ;
      LAYER met4 ;
        RECT 9.100000 42.030000 9.420000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100000 42.460000 9.420000 42.780000 ;
      LAYER met4 ;
        RECT 9.100000 42.460000 9.420000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100000 42.890000 9.420000 43.210000 ;
      LAYER met4 ;
        RECT 9.100000 42.890000 9.420000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100000 43.320000 9.420000 43.640000 ;
      LAYER met4 ;
        RECT 9.100000 43.320000 9.420000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100000 43.750000 9.420000 44.070000 ;
      LAYER met4 ;
        RECT 9.100000 43.750000 9.420000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100000 44.180000 9.420000 44.500000 ;
      LAYER met4 ;
        RECT 9.100000 44.180000 9.420000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100000 44.610000 9.420000 44.930000 ;
      LAYER met4 ;
        RECT 9.100000 44.610000 9.420000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100000 45.040000 9.420000 45.360000 ;
      LAYER met4 ;
        RECT 9.100000 45.040000 9.420000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100000 45.470000 9.420000 45.790000 ;
      LAYER met4 ;
        RECT 9.100000 45.470000 9.420000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100000 45.900000 9.420000 46.220000 ;
      LAYER met4 ;
        RECT 9.100000 45.900000 9.420000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505000 41.600000 9.825000 41.920000 ;
      LAYER met4 ;
        RECT 9.505000 41.600000 9.825000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505000 42.030000 9.825000 42.350000 ;
      LAYER met4 ;
        RECT 9.505000 42.030000 9.825000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505000 42.460000 9.825000 42.780000 ;
      LAYER met4 ;
        RECT 9.505000 42.460000 9.825000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505000 42.890000 9.825000 43.210000 ;
      LAYER met4 ;
        RECT 9.505000 42.890000 9.825000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505000 43.320000 9.825000 43.640000 ;
      LAYER met4 ;
        RECT 9.505000 43.320000 9.825000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505000 43.750000 9.825000 44.070000 ;
      LAYER met4 ;
        RECT 9.505000 43.750000 9.825000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505000 44.180000 9.825000 44.500000 ;
      LAYER met4 ;
        RECT 9.505000 44.180000 9.825000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505000 44.610000 9.825000 44.930000 ;
      LAYER met4 ;
        RECT 9.505000 44.610000 9.825000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505000 45.040000 9.825000 45.360000 ;
      LAYER met4 ;
        RECT 9.505000 45.040000 9.825000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505000 45.470000 9.825000 45.790000 ;
      LAYER met4 ;
        RECT 9.505000 45.470000 9.825000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505000 45.900000 9.825000 46.220000 ;
      LAYER met4 ;
        RECT 9.505000 45.900000 9.825000 46.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910000 41.600000 10.230000 41.920000 ;
      LAYER met4 ;
        RECT 9.910000 41.600000 10.230000 41.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910000 42.030000 10.230000 42.350000 ;
      LAYER met4 ;
        RECT 9.910000 42.030000 10.230000 42.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910000 42.460000 10.230000 42.780000 ;
      LAYER met4 ;
        RECT 9.910000 42.460000 10.230000 42.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910000 42.890000 10.230000 43.210000 ;
      LAYER met4 ;
        RECT 9.910000 42.890000 10.230000 43.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910000 43.320000 10.230000 43.640000 ;
      LAYER met4 ;
        RECT 9.910000 43.320000 10.230000 43.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910000 43.750000 10.230000 44.070000 ;
      LAYER met4 ;
        RECT 9.910000 43.750000 10.230000 44.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910000 44.180000 10.230000 44.500000 ;
      LAYER met4 ;
        RECT 9.910000 44.180000 10.230000 44.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910000 44.610000 10.230000 44.930000 ;
      LAYER met4 ;
        RECT 9.910000 44.610000 10.230000 44.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910000 45.040000 10.230000 45.360000 ;
      LAYER met4 ;
        RECT 9.910000 45.040000 10.230000 45.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910000 45.470000 10.230000 45.790000 ;
      LAYER met4 ;
        RECT 9.910000 45.470000 10.230000 45.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910000 45.900000 10.230000 46.220000 ;
      LAYER met4 ;
        RECT 9.910000 45.900000 10.230000 46.220000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met3 ;
      RECT 0.970000 41.590000 74.290000 46.230000 ;
    LAYER met4 ;
      RECT 0.000000  2.035000 75.000000  47.965000 ;
      RECT 0.000000 51.745000 75.000000  52.725000 ;
      RECT 0.000000 56.505000 75.000000 200.000000 ;
    LAYER met5 ;
      RECT 0.000000  2.135000 72.130000  15.035000 ;
      RECT 0.000000 15.035000 72.435000  19.885000 ;
      RECT 0.000000 19.885000 75.000000  24.335000 ;
      RECT 0.000000 24.335000 72.130000  36.835000 ;
      RECT 0.000000 36.835000 75.000000  46.135000 ;
      RECT 0.000000 46.135000 72.130000  96.585000 ;
      RECT 0.000000 96.585000 75.000000 200.000000 ;
  END
END sky130_fd_io__overlay_vssd_hvc
END LIBRARY
