/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_IO__TOP_XRES4V2_BLACKBOX_V
`define SKY130_FD_IO__TOP_XRES4V2_BLACKBOX_V

/**
 * top_xres4v2: XRES (Input buffer with Glitch filter).
 *
 * Verilog stub definition (black box without power pins).
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_io__top_xres4v2 (
           XRES_H_N        ,
           AMUXBUS_A       ,
           AMUXBUS_B       ,
           PAD             ,
           DISABLE_PULLUP_H,
           ENABLE_H        ,
           EN_VDDIO_SIG_H  ,
           INP_SEL_H       ,
           FILT_IN_H       ,
           PULLUP_H        ,
           ENABLE_VDDIO    ,
           PAD_A_ESD_H     ,
           TIE_HI_ESD      ,
           TIE_LO_ESD      ,
           TIE_WEAK_HI_H
       );

output XRES_H_N        ;
inout  AMUXBUS_A       ;
inout  AMUXBUS_B       ;
inout  PAD             ;
input  DISABLE_PULLUP_H;
input  ENABLE_H        ;
input  EN_VDDIO_SIG_H  ;
input  INP_SEL_H       ;
input  FILT_IN_H       ;
inout  PULLUP_H        ;
input  ENABLE_VDDIO    ;
inout  PAD_A_ESD_H     ;
output TIE_HI_ESD      ;
output TIE_LO_ESD      ;
inout  TIE_WEAK_HI_H   ;

// Voltage supply signals
supply1 VCCD   ;
supply1 VCCHIB ;
supply1 VDDA   ;
supply1 VDDIO  ;
supply1 VDDIO_Q;
supply0 VSSA   ;
supply0 VSSD   ;
supply0 VSSIO  ;
supply0 VSSIO_Q;
supply1 VSWITCH;

endmodule

`default_nettype wire
`endif  // SKY130_FD_IO__TOP_XRES4V2_BLACKBOX_V
