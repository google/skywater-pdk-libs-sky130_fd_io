# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__top_sio
  CLASS BLOCK ;
  FOREIGN sky130_fd_io__top_sio ;
  ORIGIN  16.58000  0.000000 ;
  SIZE  184.8400 BY  254.8600 ;
  PIN DM[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.350000 0.000000 19.610000 28.955000 ;
    END
  END DM[0]
  PIN DM[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.750000 0.000000 20.010000 33.225000 ;
    END
  END DM[1]
  PIN DM[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.920000 0.000000 22.180000 42.095000 ;
    END
  END DM[2]
  PIN DM_H[0]
    PORT
      LAYER met2 ;
        RECT 7.495000 42.730000 7.755000 54.975000 ;
    END
  END DM_H[0]
  PIN DM_H[1]
    PORT
      LAYER met2 ;
        RECT 13.035000 43.665000 13.295000 51.025000 ;
    END
  END DM_H[1]
  PIN DM_H[2]
    PORT
      LAYER met2 ;
        RECT 28.700000 45.680000 28.710000 45.690000 ;
    END
  END DM_H[2]
  PIN DM_H_N[0]
    PORT
      LAYER met2 ;
        RECT 4.905000 37.535000 5.165000 62.945000 ;
    END
  END DM_H_N[0]
  PIN DM_H_N[1]
    PORT
      LAYER met2 ;
        RECT 11.855000 41.150000 12.115000 67.085000 ;
    END
  END DM_H_N[1]
  PIN DM_H_N[2]
    PORT
      LAYER met2 ;
        RECT 29.695000 41.150000 29.955000 70.675000 ;
    END
  END DM_H_N[2]
  PIN ENABLE_H
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.320000 0.000000 22.580000 28.955000 ;
    END
  END ENABLE_H
  PIN HLD_H_N
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.155000 0.000000 40.415000 36.690000 ;
    END
  END HLD_H_N
  PIN HLD_I_H_N
    PORT
      LAYER met2 ;
        RECT 24.375000 48.815000 24.605000 52.135000 ;
    END
  END HLD_I_H_N
  PIN HLD_OVR
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.445000 0.000000 34.790000 2.085000 ;
    END
  END HLD_OVR
  PIN IBUF_SEL
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.555000 0.000000 40.815000 28.950000 ;
    END
  END IBUF_SEL
  PIN IBUF_SEL_H
    PORT
      LAYER met2 ;
        RECT 33.255000 19.050000 33.515000 42.405000 ;
    END
  END IBUF_SEL_H
  PIN IBUF_SEL_H_N
    PORT
      LAYER met2 ;
        RECT 33.655000 19.050000 33.915000 40.570000 ;
    END
  END IBUF_SEL_H_N
  PIN IN
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 33.725000 0.000000 33.985000 6.970000 ;
    END
  END IN
  PIN INP_DIS
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.020000 0.000000 69.280000 1.350000 ;
    END
  END INP_DIS
  PIN IN_H
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 33.325000 0.000000 33.585000 9.980000 ;
    END
  END IN_H
  PIN OE_N
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.515000 0.000000 28.775000 26.920000 ;
    END
  END OE_N
  PIN OUT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.275000 0.000000 54.535000 46.020000 ;
    END
  END OUT
  PIN PAD
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT 6.100000 131.985000 68.800000 194.600000 ;
    END
  END PAD
  PIN PAD_A_ESD_0_H
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 89.885000 0.000000 90.730000 29.615000 ;
    END
  END PAD_A_ESD_0_H
  PIN PAD_A_ESD_1_H
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT -3.000000 0.000000 -1.000000 23.820000 ;
    END
  END PAD_A_ESD_1_H
  PIN PAD_A_NOESD_H
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 88.895000 0.000000 89.745000 30.555000 ;
    END
  END PAD_A_NOESD_H
  PIN REFLEAK_BIAS
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 158.575000 199.485000 161.505000 199.715000 ;
    END
  END REFLEAK_BIAS
  PIN SIO_DIFF_HYST_EN_H
    PORT
      LAYER met1 ;
        RECT 78.355000 34.300000 81.140000 34.440000 ;
    END
  END SIO_DIFF_HYST_EN_H
  PIN SIO_DIFF_HYST_EN_H_N
    PORT
      LAYER met1 ;
        RECT 54.605000 40.680000 54.615000 40.690000 ;
    END
  END SIO_DIFF_HYST_EN_H_N
  PIN SLOW
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.115000 0.000000 28.375000 45.525000 ;
    END
  END SLOW
  PIN TIE_LO_ESD
    DIRECTION OUTPUT ;
    PORT
      LAYER met2 ;
        RECT 65.640000 0.000000 65.900000 17.465000 ;
    END
  END TIE_LO_ESD
  PIN TRIP_SEL_H
    PORT
      LAYER met2 ;
        RECT 49.440000 17.645000 49.700000 40.610000 ;
    END
  END TRIP_SEL_H
  PIN TRIP_SEL_H_N
    PORT
      LAYER met2 ;
        RECT 50.715000 28.065000 50.975000 40.570000 ;
    END
  END TRIP_SEL_H_N
  PIN VCCD
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000000 46.015000 5.385000 52.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 52.805000 5.360000 58.995000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000000 11.670000 43.885000 17.860000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 5.830000 41.010000 11.070000 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000000 66.385000 1.395000 72.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.560000 96.120000 0.710000 96.270000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000000 25.250000 6.240000 31.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 39.225000 31.465000 45.415000 ;
    END
  END VDDIO_Q
  PIN VINREF
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 163.520000 28.495000 163.905000 28.750000 ;
    END
  END VINREF
  PIN VOUTREF
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 157.645000 200.680000 161.505000 200.940000 ;
    END
    PORT
      LAYER met1 ;
        RECT 161.350000 200.805000 161.360000 200.815000 ;
    END
  END VOUTREF
  PIN VREG_EN
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.925000 0.000000 26.185000 28.250000 ;
    END
  END VREG_EN
  PIN VSSD
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000000 59.595000 3.105000 65.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.490000 32.040000 7.675000 38.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.625000 20.920000 3.775000 21.070000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -11.015000 75.975000 4.580000 90.145000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.560000 111.810000 0.710000 111.960000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 138.290000 111.950000 148.040000 116.400000 ;
    END
  END VSSIO_Q
  PIN VTRIP_SEL
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.605000 0.000000 47.865000 10.175000 ;
    END
  END VTRIP_SEL
  OBS
    LAYER li1 ;
      RECT -14.845000 0.710000 168.210000 253.385000 ;
    LAYER met1 ;
      RECT -16.580000   0.250000 168.210000  28.215000 ;
      RECT -16.580000  28.215000 163.240000  29.030000 ;
      RECT -16.580000  29.030000 168.210000  34.020000 ;
      RECT -16.580000  34.020000  78.075000  34.720000 ;
      RECT -16.580000  34.720000 168.210000  40.400000 ;
      RECT -16.580000  40.400000  54.325000  40.970000 ;
      RECT -16.580000  40.970000 168.210000 199.205000 ;
      RECT -16.580000 199.205000 158.295000 199.995000 ;
      RECT -16.580000 199.995000 168.210000 200.400000 ;
      RECT -16.580000 200.400000 157.365000 201.220000 ;
      RECT -16.580000 201.220000 168.210000 253.410000 ;
      RECT  54.895000  40.400000 168.210000  40.970000 ;
      RECT  81.420000  34.020000 168.210000  34.720000 ;
      RECT 161.785000 199.205000 168.210000 199.995000 ;
      RECT 161.785000 200.400000 168.210000 201.220000 ;
      RECT 164.185000  28.215000 168.210000  29.030000 ;
    LAYER met2 ;
      RECT -16.580000  0.000000  -3.280000  24.100000 ;
      RECT -16.580000 24.100000  19.070000  29.235000 ;
      RECT -16.580000 29.235000  19.470000  33.505000 ;
      RECT -16.580000 33.505000  21.640000  37.255000 ;
      RECT -16.580000 37.255000   4.625000  63.225000 ;
      RECT -16.580000 63.225000  11.575000  67.365000 ;
      RECT -16.580000 67.365000  29.415000  70.955000 ;
      RECT -16.580000 70.955000 164.345000 239.150000 ;
      RECT  -0.720000  0.000000  19.070000  24.100000 ;
      RECT   5.445000 37.255000  21.640000  40.870000 ;
      RECT   5.445000 40.870000  11.575000  42.450000 ;
      RECT   5.445000 42.450000   7.215000  55.255000 ;
      RECT   5.445000 55.255000  11.575000  63.225000 ;
      RECT   8.035000 42.450000  11.575000  55.255000 ;
      RECT  12.395000 40.870000  21.640000  42.375000 ;
      RECT  12.395000 42.375000  27.835000  43.385000 ;
      RECT  12.395000 43.385000  12.755000  51.305000 ;
      RECT  12.395000 51.305000  24.095000  52.415000 ;
      RECT  12.395000 52.415000  29.415000  67.365000 ;
      RECT  13.575000 43.385000  27.835000  45.805000 ;
      RECT  13.575000 45.805000  28.420000  45.970000 ;
      RECT  13.575000 45.970000  29.415000  48.535000 ;
      RECT  13.575000 48.535000  24.095000  51.305000 ;
      RECT  20.290000  0.000000  21.640000  33.505000 ;
      RECT  22.460000 29.235000  27.835000  42.375000 ;
      RECT  22.860000  0.000000  25.645000  28.530000 ;
      RECT  22.860000 28.530000  27.835000  29.235000 ;
      RECT  24.885000 48.535000  29.415000  52.415000 ;
      RECT  26.465000  0.000000  27.835000  28.530000 ;
      RECT  28.655000 27.200000  32.975000  40.870000 ;
      RECT  28.655000 40.870000  29.415000  45.400000 ;
      RECT  28.990000 45.400000  29.415000  45.970000 ;
      RECT  29.055000  0.000000  33.045000  10.260000 ;
      RECT  29.055000 10.260000  39.875000  18.770000 ;
      RECT  29.055000 18.770000  32.975000  27.200000 ;
      RECT  30.235000 40.870000  32.975000  42.685000 ;
      RECT  30.235000 42.685000  53.995000  46.300000 ;
      RECT  30.235000 46.300000 164.345000  70.955000 ;
      RECT  33.795000 40.850000  49.160000  40.890000 ;
      RECT  33.795000 40.890000  53.995000  42.685000 ;
      RECT  33.865000  7.250000  39.875000  10.260000 ;
      RECT  34.195000 18.770000  39.875000  36.970000 ;
      RECT  34.195000 36.970000  49.160000  40.850000 ;
      RECT  34.265000  2.365000  39.875000   7.250000 ;
      RECT  35.070000  0.000000  39.875000   2.365000 ;
      RECT  40.695000 29.230000  49.160000  36.970000 ;
      RECT  41.095000  0.000000  47.325000  10.455000 ;
      RECT  41.095000 10.455000  53.995000  17.365000 ;
      RECT  41.095000 17.365000  49.160000  29.230000 ;
      RECT  48.145000  0.000000  53.995000  10.455000 ;
      RECT  49.980000 17.365000  53.995000  27.785000 ;
      RECT  49.980000 27.785000  50.435000  40.850000 ;
      RECT  49.980000 40.850000  53.995000  40.890000 ;
      RECT  51.255000 27.785000  53.995000  40.850000 ;
      RECT  54.815000  0.000000  65.360000  17.745000 ;
      RECT  54.815000 17.745000  88.615000  30.835000 ;
      RECT  54.815000 30.835000 164.345000  46.300000 ;
      RECT  66.180000  0.000000  68.740000   1.630000 ;
      RECT  66.180000  1.630000  88.615000  17.745000 ;
      RECT  69.560000  0.000000  88.615000   1.630000 ;
      RECT  90.025000 29.895000 164.345000  30.835000 ;
      RECT  91.010000  0.000000 164.345000  29.895000 ;
    LAYER met3 ;
      RECT -10.350000   5.830000  -0.400000  18.260000 ;
      RECT -10.350000  18.260000 163.650000  20.520000 ;
      RECT -10.350000  20.520000   3.225000  21.470000 ;
      RECT -10.350000  21.470000 163.650000  24.850000 ;
      RECT -10.350000  24.850000  -0.400000  31.840000 ;
      RECT -10.350000  31.840000   3.090000  38.825000 ;
      RECT -10.350000  38.825000  -0.400000  72.975000 ;
      RECT -10.350000  72.975000 163.650000  75.575000 ;
      RECT -10.350000  90.545000 163.650000  95.720000 ;
      RECT -10.350000  95.720000   0.160000  96.670000 ;
      RECT -10.350000  96.670000 163.650000 111.410000 ;
      RECT -10.350000 111.410000   0.160000 112.360000 ;
      RECT -10.350000 112.360000 163.650000 211.070000 ;
      RECT   1.110000  95.720000 163.650000  96.670000 ;
      RECT   1.110000 111.410000 163.650000 112.360000 ;
      RECT   1.795000  66.185000 163.650000  72.975000 ;
      RECT   3.505000  59.395000 163.650000  66.185000 ;
      RECT   4.175000  20.520000 163.650000  21.470000 ;
      RECT   4.980000  75.575000 163.650000  90.545000 ;
      RECT   5.760000  52.605000 163.650000  59.395000 ;
      RECT   5.785000  45.815000 163.650000  52.605000 ;
      RECT   6.640000  24.850000 163.650000  31.640000 ;
      RECT   8.075000  31.640000 163.650000  38.825000 ;
      RECT  31.865000  38.825000 163.650000  45.815000 ;
      RECT  41.410000   5.830000 163.650000  11.270000 ;
      RECT  44.285000  11.270000 163.650000  18.260000 ;
    LAYER met4 ;
      RECT -5.840000 125.675000 162.170000 203.240000 ;
    LAYER met5 ;
      RECT  4.800000 125.675000 162.290000 130.385000 ;
      RECT  4.800000 196.200000 162.290000 202.060000 ;
      RECT 70.400000 130.385000 162.290000 196.200000 ;
  END
END sky130_fd_io__top_sio
END LIBRARY
