# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sky130_fd_io__top_pwrdetv2
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 56 BY 200 ;
  SYMMETRY R90 ;

  PIN tie_lo_esd
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.415 0 12.805 0.82 ;
    END
    PORT
      LAYER met1 ;
        RECT 12.415 0 12.805 0.82 ;
    END
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 3.92015 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 219.312 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2 ;
  END tie_lo_esd

  PIN vddio_present_vddd_hv
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.88 0 41.14 0.64 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.88 3.96 42.2 4.22 ;
        RECT 40.88 3.79 41.14 3.86 ;
        RECT 40.88 3.86 41.21 3.93 ;
        RECT 40.88 3.93 41.28 3.96 ;
        RECT 40.88 0 41.14 3.79 ;
        RECT 41.94 4.39 42.2 5.475 ;
        RECT 41.84 4.22 42.2 4.29 ;
        RECT 41.91 4.29 42.2 4.36 ;
        RECT 41.94 4.36 42.2 4.39 ;
    END
    ANTENNADIFFAREA 1.26 LAYER met1 ;
    ANTENNADIFFAREA 1.26 LAYER met2 ;
    ANTENNADIFFAREA 1.26 LAYER met3 ;
    ANTENNADIFFAREA 1.26 LAYER met4 ;
    ANTENNADIFFAREA 1.26 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.05679 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 23.3739 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 78.7443 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.09 LAYER via ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2 ;
  END vddio_present_vddd_hv

  PIN in1_vddio_hv
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.92 0 49.18 0.64 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.26 1.455 49.18 1.715 ;
        RECT 48.92 1.285 49.18 1.355 ;
        RECT 48.85 1.355 49.18 1.425 ;
        RECT 48.78 1.425 49.18 1.455 ;
        RECT 48.92 0 49.18 1.285 ;
        RECT 48.26 1.715 48.62 1.785 ;
        RECT 48.26 1.785 48.55 1.855 ;
        RECT 48.26 1.855 48.52 1.885 ;
        RECT 48.26 1.885 48.52 61.34 ;
    END
    ANTENNAGATEAREA 0.75 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 42.8823 LAYER met1 ;
    ANTENNAGATEAREA 0.75 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 38.5878 LAYER met2 ;
    ANTENNAGATEAREA 0.75 LAYER met3 ;
    ANTENNAGATEAREA 0.75 LAYER met4 ;
    ANTENNAGATEAREA 0.75 LAYER met5 ;
    ANTENNAPARTIALCUTAREA 0.225 LAYER via ;
  END in1_vddio_hv

  PIN out1_vddd_hv
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.145 0 50.425 0.77 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.155 0 50.415 0.64 ;
    END
    ANTENNADIFFAREA 4.2 LAYER met1 ;
    ANTENNADIFFAREA 4.2 LAYER met2 ;
    ANTENNADIFFAREA 4.2 LAYER met3 ;
    ANTENNADIFFAREA 4.2 LAYER met4 ;
    ANTENNADIFFAREA 4.2 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7695 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 131.937 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2 ;
  END out1_vddd_hv

  PIN in2_vddd_hv
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.86 0 48.12 0.64 ;
    END
    PORT
      LAYER met1 ;
        RECT 47.86 0 48.12 5.43 ;
    END
    ANTENNAGATEAREA 0.75 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 3.355 LAYER met1 ;
    ANTENNAGATEAREA 0.75 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 28.5119 LAYER met2 ;
    ANTENNAGATEAREA 0.75 LAYER met3 ;
    ANTENNAGATEAREA 0.75 LAYER met4 ;
    ANTENNAGATEAREA 0.75 LAYER met5 ;
    ANTENNAPARTIALCUTAREA 0.315 LAYER via ;
  END in2_vddd_hv

  PIN out2_vddio_hv
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.305 0 51.585 0.77 ;
    END
    PORT
      LAYER met1 ;
        RECT 51.315 0 51.575 0.64 ;
    END
    ANTENNADIFFAREA 4.2 LAYER met1 ;
    ANTENNADIFFAREA 4.2 LAYER met2 ;
    ANTENNADIFFAREA 4.2 LAYER met3 ;
    ANTENNADIFFAREA 4.2 LAYER met4 ;
    ANTENNADIFFAREA 4.2 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 22.1213 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 85.112 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via ;
    ANTENNAPARTIALCUTAREA 0.24 LAYER via2 ;
  END out2_vddio_hv

  PIN in1_vddd_hv
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.16 0 46.42 0.64 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.16 1.5 47.72 1.76 ;
        RECT 46.16 1.33 46.42 1.4 ;
        RECT 46.16 1.4 46.49 1.47 ;
        RECT 46.16 1.47 46.56 1.5 ;
        RECT 46.16 0 46.42 1.33 ;
        RECT 47.36 1.76 47.72 1.83 ;
        RECT 47.43 1.83 47.72 1.9 ;
        RECT 47.46 1.9 47.72 1.93 ;
        RECT 47.46 1.93 47.72 4.76 ;
    END
    ANTENNAGATEAREA 0.75 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 3.72429 LAYER met1 ;
    ANTENNAGATEAREA 0.75 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 22.4286 LAYER met2 ;
    ANTENNAGATEAREA 0.75 LAYER met3 ;
    ANTENNAGATEAREA 0.75 LAYER met4 ;
    ANTENNAGATEAREA 0.75 LAYER met5 ;
    ANTENNAPARTIALCUTAREA 0.36 LAYER via ;
  END in1_vddd_hv

  PIN out1_vddio_hv
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.58 0 44.86 0.77 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.59 0 44.85 0.64 ;
    END
    ANTENNADIFFAREA 4.2 LAYER met1 ;
    ANTENNADIFFAREA 4.2 LAYER met2 ;
    ANTENNADIFFAREA 4.2 LAYER met3 ;
    ANTENNADIFFAREA 4.2 LAYER met4 ;
    ANTENNADIFFAREA 4.2 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 13.699 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 81.816 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via ;
    ANTENNAPARTIALCUTAREA 0.24 LAYER via2 ;
  END out1_vddio_hv

  PIN out3_vddio_hv
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.2 0 34.48 0.77 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.215 0 34.475 0.64 ;
    END
    ANTENNADIFFAREA 4.2 LAYER met1 ;
    ANTENNADIFFAREA 4.2 LAYER met2 ;
    ANTENNADIFFAREA 4.2 LAYER met3 ;
    ANTENNADIFFAREA 4.2 LAYER met4 ;
    ANTENNADIFFAREA 4.2 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.85765 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 90.08 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via ;
    ANTENNAPARTIALCUTAREA 0.24 LAYER via2 ;
  END out3_vddio_hv

  PIN in3_vddd_hv
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.815 0 11.075 0.64 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.435 10.825 11.075 11.085 ;
        RECT 9.065 9.98 11.075 10.24 ;
        RECT 10.815 0 11.075 9.81 ;
        RECT 10.815 9.81 11.075 9.88 ;
        RECT 10.745 9.88 11.075 9.95 ;
        RECT 10.675 9.95 11.075 9.98 ;
        RECT 10.715 10.24 11.075 10.31 ;
        RECT 10.785 10.31 11.075 10.38 ;
        RECT 10.815 10.38 11.075 10.41 ;
        RECT 10.815 10.41 11.075 10.655 ;
        RECT 10.815 10.655 11.075 10.725 ;
        RECT 10.745 10.725 11.075 10.795 ;
        RECT 10.675 10.795 11.075 10.825 ;
        RECT 9.065 10.41 9.325 51.79 ;
        RECT 9.065 10.24 9.425 10.31 ;
        RECT 9.065 10.31 9.355 10.38 ;
        RECT 9.065 10.38 9.325 10.41 ;
    END
    ANTENNAGATEAREA 0.75 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 37.7481 LAYER met1 ;
    ANTENNAGATEAREA 0.75 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.8439 LAYER met2 ;
    ANTENNAGATEAREA 0.75 LAYER met3 ;
    ANTENNAGATEAREA 0.75 LAYER met4 ;
    ANTENNAGATEAREA 0.75 LAYER met5 ;
    ANTENNAPARTIALCUTAREA 0.225 LAYER via ;
  END in3_vddd_hv

  PIN vddd_present_vddio_hv
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.545 0 9.805 0.64 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.665 9.07 9.805 9.33 ;
        RECT 9.545 0 9.805 8.9 ;
        RECT 9.545 8.9 9.805 8.97 ;
        RECT 9.475 8.97 9.805 9.04 ;
        RECT 9.405 9.04 9.805 9.07 ;
        RECT 8.665 9.33 9.025 9.4 ;
        RECT 8.665 9.4 8.955 9.47 ;
        RECT 8.665 9.47 8.925 9.5 ;
        RECT 8.665 9.5 8.925 55.215 ;
    END
    ANTENNADIFFAREA 1.26 LAYER met1 ;
    ANTENNADIFFAREA 1.26 LAYER met2 ;
    ANTENNADIFFAREA 1.26 LAYER met3 ;
    ANTENNADIFFAREA 1.26 LAYER met4 ;
    ANTENNADIFFAREA 1.26 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 38.7488 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 20.3983 LAYER met2 ;
    ANTENNAPARTIALCUTAREA 0.315 LAYER via ;
  END vddd_present_vddio_hv

  PIN in2_vddio_hv
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.26 0 8.52 0.64 ;
    END
    PORT
      LAYER met1 ;
        RECT 7.88 10.425 8.52 10.685 ;
        RECT 7.88 57.2 9.435 57.34 ;
        RECT 9.295 64.175 9.935 64.435 ;
        RECT 8.26 0 8.52 10.255 ;
        RECT 8.26 10.255 8.52 10.325 ;
        RECT 8.19 10.325 8.52 10.395 ;
        RECT 8.12 10.395 8.52 10.425 ;
        RECT 7.88 10.685 8.12 10.755 ;
        RECT 7.88 10.755 8.05 10.825 ;
        RECT 7.88 10.825 8.02 10.855 ;
        RECT 7.88 10.855 8.02 57.03 ;
        RECT 7.88 57.03 8.02 57.1 ;
        RECT 7.88 57.1 8.09 57.17 ;
        RECT 7.88 57.17 8.16 57.2 ;
        RECT 9.195 57.34 9.435 57.41 ;
        RECT 9.265 57.41 9.435 57.48 ;
        RECT 9.295 57.48 9.435 57.51 ;
        RECT 9.295 57.51 9.435 64.005 ;
        RECT 9.295 64.005 9.435 64.075 ;
        RECT 9.295 64.075 9.505 64.145 ;
        RECT 9.295 64.145 9.575 64.175 ;
    END
    ANTENNAGATEAREA 0.75 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 46.0887 LAYER met1 ;
    ANTENNAGATEAREA 0.75 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.0516 LAYER met2 ;
    ANTENNAGATEAREA 0.75 LAYER met3 ;
    ANTENNAGATEAREA 0.75 LAYER met4 ;
    ANTENNAGATEAREA 0.75 LAYER met5 ;
    ANTENNAPARTIALCUTAREA 0.225 LAYER via ;
  END in2_vddio_hv

  PIN in3_vddio_hv
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.075 0 7.335 0.64 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.48 59.46 8.035 59.6 ;
        RECT 7.895 68.975 8.535 69.235 ;
        RECT 6.48 6 7.335 6.26 ;
        RECT 7.075 0 7.335 5.83 ;
        RECT 7.075 5.83 7.335 5.9 ;
        RECT 7.005 5.9 7.335 5.97 ;
        RECT 6.935 5.97 7.335 6 ;
        RECT 6.48 6.26 6.72 6.33 ;
        RECT 6.48 6.33 6.65 6.4 ;
        RECT 6.48 6.4 6.62 6.43 ;
        RECT 6.48 6.43 6.62 59.29 ;
        RECT 6.48 59.29 6.62 59.36 ;
        RECT 6.48 59.36 6.69 59.43 ;
        RECT 6.48 59.43 6.76 59.46 ;
        RECT 7.795 59.6 8.035 59.67 ;
        RECT 7.865 59.67 8.035 59.74 ;
        RECT 7.895 59.74 8.035 59.77 ;
        RECT 7.895 59.77 8.035 68.805 ;
        RECT 7.895 68.805 8.035 68.875 ;
        RECT 7.895 68.875 8.105 68.945 ;
        RECT 7.895 68.945 8.175 68.975 ;
    END
    ANTENNAGATEAREA 0.75 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 49.5992 LAYER met1 ;
    ANTENNAGATEAREA 0.75 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.9556 LAYER met2 ;
    ANTENNAGATEAREA 0.75 LAYER met3 ;
    ANTENNAGATEAREA 0.75 LAYER met4 ;
    ANTENNAGATEAREA 0.75 LAYER met5 ;
    ANTENNAPARTIALCUTAREA 0.225 LAYER via ;
  END in3_vddio_hv

  PIN out2_vddd_hv
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.5 0 43.78 0.77 ;
    END
    PORT
      LAYER met1 ;
        RECT 43.505 0 43.765 0.64 ;
    END
    ANTENNADIFFAREA 4.2 LAYER met1 ;
    ANTENNADIFFAREA 4.2 LAYER met2 ;
    ANTENNADIFFAREA 4.2 LAYER met3 ;
    ANTENNADIFFAREA 4.2 LAYER met4 ;
    ANTENNADIFFAREA 4.2 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 25.4138 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 86.585 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2 ;
  END out2_vddd_hv

  PIN out3_vddd_hv
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.335 0 42.615 0.77 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.345 0 42.605 0.64 ;
    END
    ANTENNADIFFAREA 4.2 LAYER met1 ;
    ANTENNADIFFAREA 4.2 LAYER met2 ;
    ANTENNADIFFAREA 4.2 LAYER met3 ;
    ANTENNADIFFAREA 4.2 LAYER met4 ;
    ANTENNADIFFAREA 4.2 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 17.5841 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 84.0403 LAYER met3 ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via ;
    ANTENNAPARTIALCUTAREA 0.16 LAYER via2 ;
  END out3_vddd_hv

  PIN rst_por_hv_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.41 0 1.67 0.64 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.41 0 1.67 113.775 ;
    END
    ANTENNAGATEAREA 13 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 79.1945 LAYER met1 ;
    ANTENNAGATEAREA 13 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 52.6894 LAYER met2 ;
    ANTENNAGATEAREA 13 LAYER met3 ;
    ANTENNAGATEAREA 13 LAYER met4 ;
    ANTENNAGATEAREA 13 LAYER met5 ;
    ANTENNAPARTIALCUTAREA 0.4275 LAYER via ;
  END rst_por_hv_n

  PIN vssio_q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 1.41 0 7.115 3.155 ;
    END
  END vssio_q

  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 13.305 0 17.715 200 ;
    END
  END vssd

  PIN vddd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 18.515 0 22.515 200 ;
    END
  END vddd1

  PIN vddd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 33.665 64.965 39.54 200 ;
        RECT 35 49.635 39.59 58.11 ;
        RECT 35 0 39.59 46.715 ;
        RECT 35 63.63 39.54 63.78 ;
        RECT 34.85 63.78 39.54 63.93 ;
        RECT 34.7 63.93 39.54 64.08 ;
        RECT 34.55 64.08 39.54 64.23 ;
        RECT 34.4 64.23 39.54 64.38 ;
        RECT 34.25 64.38 39.54 64.53 ;
        RECT 34.1 64.53 39.54 64.68 ;
        RECT 33.95 64.68 39.54 64.83 ;
        RECT 33.8 64.83 39.54 64.965 ;
        RECT 35 60.055 39.54 63.63 ;
        RECT 35 59.645 39.13 59.795 ;
        RECT 35 59.795 39.28 59.945 ;
        RECT 35 59.945 39.43 60.055 ;
        RECT 35 58.57 39.13 59.645 ;
        RECT 35 58.11 39.44 58.26 ;
        RECT 35 58.26 39.29 58.41 ;
        RECT 35 58.41 39.14 58.56 ;
        RECT 35 58.56 39.13 58.57 ;
        RECT 35 49.235 39.19 49.385 ;
        RECT 35 49.385 39.34 49.535 ;
        RECT 35 49.535 39.49 49.635 ;
        RECT 35 47.115 39.19 49.235 ;
        RECT 35 46.715 39.44 46.865 ;
        RECT 35 46.865 39.29 47.015 ;
        RECT 35 47.015 39.19 47.115 ;
    END
  END vddd2

  PIN vssa
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 23.315 0 28.315 200 ;
    END
  END vssa

  PIN vddio_q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 29.115 0 33.625 33.58 ;
        RECT 29.115 33.58 33.475 33.73 ;
        RECT 29.115 33.73 33.325 33.88 ;
        RECT 29.115 33.88 33.175 34.03 ;
        RECT 29.115 34.03 33.115 34.09 ;
        RECT 29.115 34.09 33.115 200 ;
    END
  END vddio_q

  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 7.915 137.425 12.505 200 ;
        RECT 7.915 136.835 11.915 136.985 ;
        RECT 7.915 136.985 12.065 137.135 ;
        RECT 7.915 137.135 12.215 137.285 ;
        RECT 7.915 137.285 12.365 137.425 ;
        RECT 7.915 0 11.915 136.835 ;
    END
  END vccd
  OBS
    LAYER met2 ;
      RECT 42.755 0 43.36 0.91 ;
      RECT 43.92 0 44.44 0.91 ;
      RECT 45 0.78 50.005 0.91 ;
      RECT 45 0 46.02 0.78 ;
      RECT 46.56 0 47.72 0.78 ;
      RECT 48.26 0 48.78 0.78 ;
      RECT 49.32 0 50.005 0.78 ;
      RECT 50.565 0 51.165 0.91 ;
      RECT 51.725 0 56 0.91 ;
      RECT 0 0 1.27 0.78 ;
      RECT 0 0.78 12.275 0.96 ;
      RECT 0 0.96 56 200 ;
      RECT 1.81 0 6.935 0.78 ;
      RECT 7.475 0 8.12 0.78 ;
      RECT 8.66 0 9.405 0.78 ;
      RECT 9.945 0 10.675 0.78 ;
      RECT 11.215 0 12.275 0.78 ;
      RECT 12.945 0 34.06 0.91 ;
      RECT 12.945 0.91 56 0.96 ;
      RECT 34.62 0 40.74 0.78 ;
      RECT 34.62 0.78 42.195 0.91 ;
      RECT 41.28 0 42.195 0.78 ;
      RECT 0 0 1.13 0.92 ;
      RECT 7.615 0 7.98 0.92 ;
      RECT 8.8 0 9.265 0.92 ;
      RECT 10.085 0 10.535 0.92 ;
      RECT 11.355 0 12.135 0.92 ;
      RECT 41.42 0 42.055 0.92 ;
      RECT 42.895 0 43.22 1.05 ;
      RECT 44.06 0 44.3 1.05 ;
      RECT 45.14 0 45.88 0.92 ;
      RECT 46.7 0 47.58 0.92 ;
      RECT 48.4 0 48.64 0.92 ;
      RECT 49.46 0 49.865 0.92 ;
      RECT 50.705 0 51.025 1.05 ;
      RECT 51.865 0 56 4.055 ;
      RECT 45.14 0.92 49.865 4.055 ;
      RECT 13.085 0 33.92 4.055 ;
      RECT 0 0.92 12.135 4.105 ;
      RECT 1.95 0 6.795 3.925 ;
      RECT 0 1.1 56 200 ;
      RECT 13.085 1.05 56 4.105 ;
      RECT 34.76 0.92 42.055 4.055 ;
      RECT 34.76 0 40.6 3.925 ;
    LAYER met1 ;
      RECT 0 113.915 56 200 ;
      RECT 1.81 69.375 56 113.915 ;
      RECT 8.675 68.835 56 69.375 ;
      RECT 8.175 68.745 56 68.835 ;
      RECT 8.175 64.575 56 68.745 ;
      RECT 10.075 64.035 56 64.575 ;
      RECT 9.575 63.945 56 64.035 ;
      RECT 9.575 61.48 56 63.945 ;
      RECT 1.81 59.83 7.755 69.375 ;
      RECT 1.81 59.74 7.755 59.83 ;
      RECT 8.175 59.32 9.155 64.575 ;
      RECT 6.76 59.23 9.155 59.32 ;
      RECT 6.76 57.57 9.155 59.23 ;
      RECT 6.76 57.48 9.155 57.57 ;
      RECT 9.575 57.06 48.12 61.48 ;
      RECT 8.16 56.97 48.12 57.06 ;
      RECT 8.16 55.355 48.12 56.97 ;
      RECT 9.065 51.93 48.12 55.355 ;
      RECT 9.465 11.225 48.12 51.93 ;
      RECT 8.16 10.915 8.525 55.355 ;
      RECT 8.25 10.825 8.525 10.915 ;
      RECT 9.465 10.685 10.295 11.225 ;
      RECT 9.465 10.595 10.585 10.685 ;
      RECT 9.465 10.47 10.675 10.595 ;
      RECT 9.555 10.38 10.675 10.47 ;
      RECT 6.76 10.285 7.74 57.48 ;
      RECT 6.76 10.195 8.03 10.285 ;
      RECT 9.065 9.75 10.585 9.84 ;
      RECT 9.065 9.56 10.675 9.75 ;
      RECT 9.155 9.47 10.675 9.56 ;
      RECT 8.66 8.84 9.315 8.93 ;
      RECT 6.76 6.49 8.12 10.195 ;
      RECT 6.85 6.4 8.12 6.49 ;
      RECT 1.81 5.86 6.34 59.74 ;
      RECT 1.81 5.77 6.845 5.86 ;
      RECT 11.215 5.615 48.12 11.225 ;
      RECT 42.34 5.57 48.12 5.615 ;
      RECT 42.34 4.9 47.72 5.57 ;
      RECT 11.215 4.45 41.8 5.615 ;
      RECT 11.215 4.36 41.8 4.45 ;
      RECT 42.34 3.82 47.32 4.9 ;
      RECT 41.28 3.73 47.32 3.82 ;
      RECT 41.28 1.99 47.32 3.73 ;
      RECT 48.66 1.945 56 61.48 ;
      RECT 41.28 1.9 47.32 1.99 ;
      RECT 48.75 1.855 56 1.945 ;
      RECT 46.56 1.27 47.72 1.36 ;
      RECT 48.26 1.225 48.69 1.315 ;
      RECT 11.215 0.96 40.74 4.36 ;
      RECT 12.945 0.78 40.74 0.96 ;
      RECT 12.945 0 34.075 0.78 ;
      RECT 41.28 0.78 46.02 1.9 ;
      RECT 49.32 0.78 56 1.855 ;
      RECT 46.56 0 47.72 1.27 ;
      RECT 48.26 0 48.78 1.225 ;
      RECT 34.615 0 40.74 0.78 ;
      RECT 41.28 0 42.205 0.78 ;
      RECT 42.745 0 43.365 0.78 ;
      RECT 43.905 0 44.45 0.78 ;
      RECT 44.99 0 46.02 0.78 ;
      RECT 49.32 0 50.015 0.78 ;
      RECT 50.555 0 51.175 0.78 ;
      RECT 51.715 0 56 0.78 ;
      RECT 0 0 1.27 113.915 ;
      RECT 9.945 0 10.675 9.47 ;
      RECT 8.66 0 9.405 8.84 ;
      RECT 7.475 0 8.12 6.4 ;
      RECT 1.81 0 6.935 5.77 ;
      RECT 11.215 0 12.275 0.96 ;
      RECT 9.715 61.62 56 63.895 ;
      RECT 10.215 61.62 56 68.695 ;
      RECT 10.215 61.62 56 68.695 ;
      RECT 48.8 1.995 56 68.695 ;
      RECT 48.8 1.995 56 68.695 ;
      RECT 48.8 1.995 56 61.62 ;
      RECT 51.855 0 56 61.62 ;
      RECT 51.855 0 56 61.62 ;
      RECT 51.855 0 56 0.92 ;
      RECT 10.085 0 10.535 9.7 ;
      RECT 8.8 0 9.265 8.79 ;
      RECT 46.7 0 47.58 1.22 ;
      RECT 48.4 0 48.64 1.175 ;
      RECT 9.605 10.52 10.155 11.365 ;
      RECT 11.355 0 12.135 1.1 ;
      RECT 41.42 0 42.065 0.92 ;
      RECT 42.885 0 43.225 0.92 ;
      RECT 44.045 0 44.31 0.92 ;
      RECT 45.13 0 45.88 0.92 ;
      RECT 46.26 1.96 46.9 2.04 ;
      RECT 49.46 0 49.875 0.92 ;
      RECT 50.695 0 51.035 0.92 ;
      RECT 0 0 1.13 114.055 ;
      RECT 1.95 5.72 6.2 59.88 ;
      RECT 6.9 57.62 9.015 59.18 ;
      RECT 6.9 10.145 7.6 57.62 ;
      RECT 6.9 6.54 7.98 10.145 ;
      RECT 7.615 0 7.98 6.54 ;
      RECT 8.3 55.495 47.98 56.92 ;
      RECT 8.315 59.18 9.015 64.715 ;
      RECT 9.205 52.07 47.98 55.495 ;
      RECT 11.355 2.75 40.6 4.5 ;
      RECT 11.355 4.5 41.66 7.505 ;
      RECT 11.355 1.1 14.36 2.75 ;
      RECT 33.935 0.92 40.6 2.75 ;
      RECT 34.755 0 40.6 0.92 ;
      RECT 41.42 0.92 42.48 2.78 ;
      RECT 41.42 2.78 47.32 3.68 ;
      RECT 42.48 3.68 47.32 5.04 ;
      RECT 42.48 5.71 47.98 8.715 ;
      RECT 42.48 5.04 47.58 5.71 ;
      RECT 49.46 0.92 52.465 1.995 ;
      RECT 0 114.055 56 200 ;
      RECT 42.48 0.92 45.88 2.04 ;
      RECT 8.315 64.715 56 68.695 ;
      RECT 8.815 64.715 56 114.055 ;
      RECT 8.815 68.695 56 69.515 ;
      RECT 10.215 63.895 56 64.715 ;
      RECT 1.95 59.88 7.615 114.055 ;
      RECT 1.95 69.515 56 114.055 ;
      RECT 1.95 59.88 7.615 69.515 ;
      RECT 1.95 0 6.795 5.72 ;
      RECT 9.715 56.92 47.98 63.895 ;
      RECT 9.715 56.92 47.98 63.895 ;
      RECT 13.085 0 33.935 0.92 ;
      RECT 13.085 0 33.935 4.5 ;
      RECT 13.085 0 33.935 4.5 ;
      RECT 13.085 0 33.935 4.5 ;
      RECT 9.605 11.365 47.98 52.07 ;
      RECT 11.355 5.755 47.98 11.365 ;
      RECT 42.48 2.04 47.18 2.78 ;
    LAYER li1 ;
      RECT 33.35 63.08 33.52 63.75 ;
      RECT 35.825 59.725 38.665 59.895 ;
      RECT 38.325 63.27 38.495 64.145 ;
      RECT 37.495 63.45 38.025 63.62 ;
      RECT 31.985 60.475 32.89 60.645 ;
      RECT 31.96 61.325 32.13 61.855 ;
      RECT 31.82 62.28 38.235 62.45 ;
      RECT 33.36 60.665 33.53 61.495 ;
      RECT 37.16 60.665 37.33 61.795 ;
      RECT 36.38 60.365 36.55 61.495 ;
      RECT 34.82 60.665 34.99 61.495 ;
      RECT 37.94 60.365 38.11 61.495 ;
      RECT 38.72 60.365 38.89 61.495 ;
      RECT 32.71 61.325 32.88 61.855 ;
      RECT 33.99 60.665 34.16 61.795 ;
      RECT 35.6 60.665 35.77 61.795 ;
      RECT 34.165 68.095 34.335 70.155 ;
      RECT 34.165 64.975 34.335 67.815 ;
      RECT 35.565 64.2 36.095 64.37 ;
      RECT 34.795 68.65 36.095 68.82 ;
      RECT 34.685 67.09 35.645 67.26 ;
      RECT 35.135 69.43 36.015 69.6 ;
      RECT 34.685 65.53 35.645 65.7 ;
      RECT 35.135 64.75 36.035 64.92 ;
      RECT 35.135 66.31 36.035 66.48 ;
      RECT 35.135 67.87 36.015 68.04 ;
      RECT 33.35 64.03 33.52 66.87 ;
      RECT 33.35 67.15 33.52 69.99 ;
      RECT 39.075 68.095 39.245 70.155 ;
      RECT 39.075 64.975 39.245 67.815 ;
      RECT 37.525 65.53 38.715 65.7 ;
      RECT 37.115 66.31 38.315 66.48 ;
      RECT 37.535 67.09 38.715 67.26 ;
      RECT 37.605 68.65 38.315 68.82 ;
      RECT 37.65 70.21 38.315 70.38 ;
      RECT 37.115 67.87 38.315 68.04 ;
      RECT 37.115 69.43 38.315 69.6 ;
      RECT 37.115 64.2 37.645 64.37 ;
      RECT 35.135 70.21 36.095 70.38 ;
      RECT 37.195 64.75 38.605 64.92 ;
      RECT 38.12 71.335 38.29 72.01 ;
      RECT 34.86 75.185 37.18 75.355 ;
      RECT 35.72 75.965 37.82 76.135 ;
      RECT 38.12 72.29 38.29 78.25 ;
      RECT 35.72 71.285 37.82 71.455 ;
      RECT 34.86 72.065 37.18 72.235 ;
      RECT 35.72 72.845 37.82 73.015 ;
      RECT 34.86 73.625 37.18 73.795 ;
      RECT 35.72 74.405 37.82 74.575 ;
      RECT 38.12 90.55 38.29 96.51 ;
      RECT 38.12 96.79 38.29 98.07 ;
      RECT 38.12 89.595 38.29 90.27 ;
      RECT 31.865 96.585 32.035 99.425 ;
      RECT 31.865 93.465 32.035 96.305 ;
      RECT 31.865 92.515 32.035 93.185 ;
      RECT 38.12 87.66 38.29 88.94 ;
      RECT 35.58 79.085 37.68 79.255 ;
      RECT 35.72 77.525 37.82 77.695 ;
      RECT 34.86 79.865 37.82 80.035 ;
      RECT 38.12 81.42 38.29 87.38 ;
      RECT 35.72 80.415 37.82 80.585 ;
      RECT 34.86 81.195 37.18 81.365 ;
      RECT 35.72 81.975 37.82 82.145 ;
      RECT 34.86 82.755 37.18 82.925 ;
      RECT 35.72 83.535 37.82 83.705 ;
      RECT 34.86 84.315 37.18 84.485 ;
      RECT 35.72 85.095 37.82 85.265 ;
      RECT 35.58 88.215 37.68 88.385 ;
      RECT 35.72 86.655 37.82 86.825 ;
      RECT 34.86 88.995 37.82 89.165 ;
      RECT 35.72 89.545 37.82 89.715 ;
      RECT 34.86 90.325 37.18 90.495 ;
      RECT 35.72 91.105 37.82 91.275 ;
      RECT 34.86 91.885 37.18 92.055 ;
      RECT 35.72 92.665 37.82 92.835 ;
      RECT 34.86 93.445 37.18 93.615 ;
      RECT 35.72 94.225 37.82 94.395 ;
      RECT 35.58 97.345 37.82 97.515 ;
      RECT 35.72 95.785 37.82 95.955 ;
      RECT 38.12 78.53 38.29 79.81 ;
      RECT 38.12 80.46 38.29 81.14 ;
      RECT 34.86 87.435 37.18 87.605 ;
      RECT 34.86 78.305 37.18 78.475 ;
      RECT 34.86 96.565 37.18 96.735 ;
      RECT 34.86 95.005 37.18 95.175 ;
      RECT 34.86 85.875 37.18 86.045 ;
      RECT 34.86 76.745 37.18 76.915 ;
      RECT 34.86 98.125 37.82 98.295 ;
      RECT 18.66 121.735 30.96 122.585 ;
      RECT 16.34 136.12 17.11 136.65 ;
      RECT 26.975 136.115 27.72 136.645 ;
      RECT 38.58 71.23 38.75 98.33 ;
      RECT 38.58 12.385 38.75 39.465 ;
      RECT 12.95 137.325 40.01 139.535 ;
      RECT 30.275 112.49 40.01 116.23 ;
      RECT 35.415 134.77 35.925 137.325 ;
      RECT 30.28 116.23 38.84 116.28 ;
      RECT 35.37 116.28 35.96 134.77 ;
      RECT 14.215 8.11 17.53 8.44 ;
      RECT 35.72 12.42 37.82 12.59 ;
      RECT 38.12 13.085 38.29 13.145 ;
      RECT 38.125 12.445 38.295 12.475 ;
      RECT 38.12 12.475 38.295 13.085 ;
      RECT 38.12 13.425 38.29 19.385 ;
      RECT 34.86 13.2 37.18 13.37 ;
      RECT 35.22 11.55 39.63 11.58 ;
      RECT 35.22 0.2 40.01 7.725 ;
      RECT 35.22 9 40.01 11.55 ;
      RECT 35.355 7.725 40.01 9 ;
      RECT 38.12 19.665 38.29 20.945 ;
      RECT 38.12 21.6 38.29 22.275 ;
      RECT 38.12 28.795 38.29 30.075 ;
      RECT 38.12 31.685 38.29 37.645 ;
      RECT 38.12 30.73 38.29 31.405 ;
      RECT 22.765 17.785 25.605 17.955 ;
      RECT 21.815 17.785 22.485 17.955 ;
      RECT 25.885 17.785 28.725 17.955 ;
      RECT 38.12 22.555 38.29 28.515 ;
      RECT 34.86 34.58 37.18 34.75 ;
      RECT 35.72 33.8 37.82 33.97 ;
      RECT 34.86 33.02 37.18 33.19 ;
      RECT 35.72 32.24 37.82 32.41 ;
      RECT 34.86 31.46 37.18 31.63 ;
      RECT 35.72 30.68 37.82 30.85 ;
      RECT 34.86 30.13 37.82 30.3 ;
      RECT 35.72 27.79 37.82 27.96 ;
      RECT 35.72 29.35 37.82 29.52 ;
      RECT 34.86 25.45 37.18 25.62 ;
      RECT 35.72 24.67 37.82 24.84 ;
      RECT 35.72 26.23 37.82 26.4 ;
      RECT 34.86 23.89 37.18 24.06 ;
      RECT 35.72 23.11 37.82 23.28 ;
      RECT 34.86 22.33 37.18 22.5 ;
      RECT 35.72 21.55 37.82 21.72 ;
      RECT 35.72 20.22 37.82 20.39 ;
      RECT 35.72 18.66 37.82 18.83 ;
      RECT 34.86 14.76 37.18 14.93 ;
      RECT 34.86 16.32 37.18 16.49 ;
      RECT 35.72 15.54 37.82 15.71 ;
      RECT 34.86 17.88 37.18 18.05 ;
      RECT 34.86 19.44 37.18 19.61 ;
      RECT 34.86 21 37.82 21.17 ;
      RECT 35.72 13.98 37.54 14.15 ;
      RECT 35.72 17.1 37.82 17.27 ;
      RECT 34.86 28.57 37.18 28.74 ;
      RECT 34.86 27.01 37.18 27.18 ;
      RECT 15.72 55.42 16.39 55.59 ;
      RECT 16.67 55.42 19.51 55.59 ;
      RECT 15.575 53.89 22.96 54.06 ;
      RECT 15.525 48.845 32.195 49.135 ;
      RECT 14.21 39.4 33.72 39.63 ;
      RECT 38.12 37.925 38.29 39.205 ;
      RECT 24.94 53.4 31.27 53.57 ;
      RECT 19.79 55.42 22.63 55.59 ;
      RECT 34.86 39.26 37.82 39.43 ;
      RECT 35.72 36.92 37.82 37.09 ;
      RECT 35.72 38.48 37.82 38.65 ;
      RECT 35.72 35.36 37.82 35.53 ;
      RECT 34.18 54.46 34.71 54.63 ;
      RECT 34.18 50.01 35.37 50.18 ;
      RECT 34.18 51.57 35.37 51.74 ;
      RECT 34.62 49.23 35.78 49.4 ;
      RECT 34.605 50.79 35.78 50.96 ;
      RECT 34.61 52.35 35.37 52.52 ;
      RECT 34.18 53.13 35.37 53.3 ;
      RECT 34.615 53.92 35.78 54.09 ;
      RECT 28.86 55.69 31.7 55.86 ;
      RECT 26.52 55.69 28.58 55.86 ;
      RECT 25.02 55.69 25.69 55.86 ;
      RECT 26.36 54.68 26.53 55.25 ;
      RECT 27.075 54.37 27.245 55.39 ;
      RECT 27.855 54.68 28.025 55.39 ;
      RECT 29.415 54.82 29.585 55.39 ;
      RECT 30.975 54.82 31.145 55.39 ;
      RECT 28.635 53.99 28.805 55.01 ;
      RECT 30.195 53.985 30.365 55.01 ;
      RECT 25.745 54.48 25.915 55.01 ;
      RECT 24.995 54.48 25.165 55.01 ;
      RECT 36.14 51.795 36.31 53.855 ;
      RECT 31.755 54.08 31.925 55.01 ;
      RECT 34.86 37.7 37.18 37.87 ;
      RECT 34.86 36.14 37.18 36.31 ;
      RECT 35.39 41.465 35.56 42.385 ;
      RECT 34.18 43.77 35.37 43.94 ;
      RECT 34.18 41.66 34.71 41.83 ;
      RECT 34.18 48.45 35.37 48.62 ;
      RECT 34.18 46.89 35.37 47.06 ;
      RECT 34.62 44.55 35.78 44.72 ;
      RECT 34.62 42.99 35.78 43.16 ;
      RECT 34.555 42.44 35.085 42.61 ;
      RECT 36.14 45.555 36.31 48.395 ;
      RECT 36.14 43.22 36.31 45.275 ;
      RECT 34.62 47.67 35.78 47.84 ;
      RECT 34.62 46.11 35.78 46.28 ;
      RECT 33.585 42.185 33.755 55.305 ;
      RECT 34.18 45.33 35.37 45.5 ;
      RECT 36.14 48.675 36.31 51.515 ;
      RECT 35.39 54.685 35.56 55.355 ;
      RECT 34.18 55.21 34.71 55.38 ;
      RECT 14.145 66.575 30.57 66.855 ;
      RECT 31.82 62.935 31.99 70.32 ;
      RECT 36.52 63.395 36.69 69.725 ;
      RECT 34.715 63.24 34.885 64.145 ;
      RECT 35.115 63.45 35.645 63.62 ;
      RECT 33.485 59.725 35.545 59.895 ;
    LAYER met3 ;
      RECT 0 3.555 7.615 200 ;
      RECT 7.515 0 7.615 3.555 ;
      RECT 12.215 136.71 12.905 137.3 ;
      RECT 12.215 0 12.905 136.71 ;
      RECT 12.805 137.3 12.905 200 ;
      RECT 28.715 0 28.815 200 ;
      RECT 33.415 34.215 34.7 63.505 ;
      RECT 33.925 33.705 34.7 34.215 ;
      RECT 33.925 0 34.7 33.705 ;
      RECT 39.43 59.52 56 59.93 ;
      RECT 39.43 58.695 56 59.52 ;
      RECT 39.89 58.235 56 58.695 ;
      RECT 39.49 49.11 56 49.51 ;
      RECT 39.49 47.24 56 49.11 ;
      RECT 39.89 46.84 56 47.24 ;
      RECT 39.84 59.93 56 200 ;
      RECT 39.89 49.51 56 58.235 ;
      RECT 39.89 0 56 46.84 ;
      RECT 39.53 58.735 39.94 59.48 ;
      RECT 39.59 47.28 39.99 49.07 ;
      RECT 42.99 3.0 53.0 48.125 ;
      RECT 39.94 58.275 56 200 ;
      RECT 39.99 0 56 200 ;
      RECT 39.99 0 56 200 ;
      RECT 42.94 59.57 53.0 197.0 ;
      RECT 42.99 48.225 53.0 59.52 ;
      RECT 39.99 58.275 56 58.425 ;
      RECT 39.84 58.425 56 58.575 ;
      RECT 39.69 58.575 56 58.725 ;
      RECT 39.54 58.725 56 58.735 ;
      RECT 39.68 59.48 56 59.63 ;
      RECT 39.83 59.63 56 59.78 ;
      RECT 39.94 59.78 56 59.89 ;
      RECT 39.99 46.88 56 47.03 ;
      RECT 39.84 47.03 56 47.18 ;
      RECT 39.69 47.18 56 47.28 ;
      RECT 39.74 49.07 56 49.22 ;
      RECT 39.89 49.22 56 49.37 ;
      RECT 39.99 49.37 56 49.47 ;
      RECT 42.99 59.52 53.0 59.545 ;
      RECT 42.965 59.545 53.0 59.57 ;
      RECT 42.965 48.175 53.0 48.2 ;
      RECT 42.99 48.2 53.0 48.225 ;
      RECT 42.99 48.125 53.0 48.15 ;
      RECT 42.965 48.15 53.0 48.175 ;
      RECT 42.965 48.175 53.0 48.2 ;
      RECT 42.99 48.2 53.0 48.225 ;
      RECT 42.99 48.125 53.0 48.15 ;
      RECT 42.965 48.15 53.0 48.175 ;
      RECT 42.99 59.52 53.0 59.545 ;
      RECT 42.965 59.545 53.0 59.57 ;
      RECT 0 0 1.01 3.555 ;
      RECT 0 3.555 7.515 200 ;
      RECT 12.315 0 12.905 136.67 ;
      RECT 12.465 136.67 12.905 136.82 ;
      RECT 12.615 136.82 12.905 136.97 ;
      RECT 12.765 136.97 12.905 137.12 ;
      RECT 33.515 34.255 34.6 63.465 ;
      RECT 34.025 0 34.6 33.745 ;
      RECT 33.515 63.465 34.45 63.615 ;
      RECT 33.515 63.615 34.3 63.765 ;
      RECT 33.515 63.765 34.15 63.915 ;
      RECT 33.515 63.915 34.0 64.065 ;
      RECT 33.515 64.065 33.85 64.215 ;
      RECT 33.515 64.215 33.7 64.365 ;
      RECT 33.515 64.365 33.55 64.515 ;
      RECT 34.025 33.745 34.6 33.895 ;
      RECT 33.875 33.895 34.6 34.045 ;
      RECT 33.725 34.045 34.6 34.195 ;
      RECT 33.575 34.195 34.6 34.255 ;
  END
END sky130_fd_io__top_pwrdetv2


END LIBRARY
