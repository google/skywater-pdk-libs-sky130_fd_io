# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_io__top_sio_macro
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 480 BY  253.7150 ;
  SYMMETRY R90 ;
  PIN AMUXBUS_A
    ANTENNAPARTIALCUTAREA  0.280000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.905000 0.000000 448.165000 83.360000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 106.840000 480.000000 109.820000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    ANTENNAPARTIALCUTAREA  0.080000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.655000 0.000000 448.915000 83.360000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 102.080000 480.000000 105.060000 ;
    END
  END AMUXBUS_B
  PIN DFT_REFGEN
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.245000 238.950000 449.560000 239.005000 ;
        RECT 449.245000 239.005000 449.505000 239.060000 ;
        RECT 449.245000 239.060000 449.505000 245.815000 ;
        RECT 449.305000 238.890000 449.615000 238.950000 ;
        RECT 449.375000 238.820000 449.675000 238.890000 ;
        RECT 449.445000 238.750000 449.745000 238.820000 ;
        RECT 449.515000 238.680000 449.815000 238.750000 ;
        RECT 449.585000 238.610000 449.885000 238.680000 ;
        RECT 449.655000 238.540000 449.955000 238.610000 ;
        RECT 449.725000 238.470000 450.025000 238.540000 ;
        RECT 449.795000 238.400000 450.095000 238.470000 ;
        RECT 449.865000 238.330000 450.165000 238.400000 ;
        RECT 449.935000 238.260000 450.235000 238.330000 ;
        RECT 450.005000 238.190000 450.305000 238.260000 ;
        RECT 450.075000 238.120000 450.375000 238.190000 ;
        RECT 450.145000 238.050000 450.445000 238.120000 ;
        RECT 450.215000 237.980000 450.515000 238.050000 ;
        RECT 450.285000 237.910000 450.585000 237.980000 ;
        RECT 450.355000 237.840000 450.655000 237.910000 ;
        RECT 450.425000 237.770000 450.725000 237.840000 ;
        RECT 450.495000 237.700000 450.795000 237.770000 ;
        RECT 450.565000 237.630000 450.865000 237.700000 ;
        RECT 450.635000 237.560000 450.935000 237.630000 ;
        RECT 450.705000 237.490000 451.005000 237.560000 ;
        RECT 450.775000 237.420000 451.075000 237.490000 ;
        RECT 450.845000 237.350000 451.145000 237.420000 ;
        RECT 450.915000 237.280000 451.215000 237.350000 ;
        RECT 450.985000 237.210000 451.285000 237.280000 ;
        RECT 451.055000 237.140000 451.355000 237.210000 ;
        RECT 451.125000 237.070000 451.425000 237.140000 ;
        RECT 451.195000 237.000000 451.495000 237.070000 ;
        RECT 451.265000 236.930000 451.565000 237.000000 ;
        RECT 451.335000 236.860000 451.635000 236.930000 ;
        RECT 451.405000 236.790000 451.705000 236.860000 ;
        RECT 451.475000 236.720000 451.775000 236.790000 ;
        RECT 451.545000 236.650000 451.845000 236.720000 ;
        RECT 451.600000 236.595000 451.915000 236.650000 ;
        RECT 451.655000   0.000000 451.915000 236.540000 ;
        RECT 451.655000 236.540000 451.915000 236.595000 ;
    END
  END DFT_REFGEN
  PIN DM0[0]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.380000 0.000000 156.640000 33.095000 ;
    END
  END DM0[0]
  PIN DM0[1]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.980000 0.000000 156.240000 33.835000 ;
    END
  END DM0[1]
  PIN DM0[2]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.810000  0.000000 154.070000 41.985000 ;
        RECT 153.810000 41.985000 154.070000 41.990000 ;
        RECT 153.810000 41.990000 154.075000 41.995000 ;
        RECT 153.810000 41.995000 154.080000 42.095000 ;
        RECT 153.815000 42.095000 154.080000 42.100000 ;
        RECT 153.820000 42.100000 154.080000 42.105000 ;
        RECT 153.820000 42.105000 154.080000 42.910000 ;
    END
  END DM0[2]
  PIN DM1[0]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.365000 0.000000 233.625000 33.095000 ;
    END
  END DM1[0]
  PIN DM1[1]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.765000 0.000000 234.025000 33.835000 ;
    END
  END DM1[1]
  PIN DM1[2]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.925000 41.995000 236.195000 42.095000 ;
        RECT 235.925000 42.095000 236.190000 42.100000 ;
        RECT 235.925000 42.100000 236.185000 42.105000 ;
        RECT 235.925000 42.105000 236.185000 42.910000 ;
        RECT 235.930000 41.990000 236.195000 41.995000 ;
        RECT 235.935000  0.000000 236.195000 41.985000 ;
        RECT 235.935000 41.985000 236.195000 41.990000 ;
    END
  END DM1[2]
  PIN ENABLE_H
    ANTENNAPARTIALCUTAREA  0.240000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.390000 2.235000 153.670000  3.005000 ;
        RECT 153.400000 2.225000 153.670000  2.235000 ;
        RECT 153.400000 3.005000 153.670000  3.015000 ;
        RECT 153.410000 0.000000 153.670000  2.215000 ;
        RECT 153.410000 2.215000 153.670000  2.225000 ;
        RECT 153.410000 3.015000 153.670000  3.025000 ;
        RECT 153.410000 3.025000 153.670000 34.945000 ;
    END
    PORT
      LAYER met2 ;
        RECT 236.335000 0.000000 236.595000  2.190000 ;
        RECT 236.335000 2.190000 236.595000  2.210000 ;
        RECT 236.335000 2.210000 236.615000  2.230000 ;
        RECT 236.335000 2.230000 236.635000  2.235000 ;
        RECT 236.335000 2.235000 236.640000  3.005000 ;
        RECT 236.335000 3.005000 236.620000  3.025000 ;
        RECT 236.335000 3.025000 236.600000  3.045000 ;
        RECT 236.335000 3.045000 236.595000  3.050000 ;
        RECT 236.335000 3.050000 236.595000 34.945000 ;
    END
  END ENABLE_H
  PIN ENABLE_VDDA_H
    ANTENNAGATEAREA  19.20000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.995000 239.270000 450.310000 239.325000 ;
        RECT 449.995000 239.325000 450.255000 239.380000 ;
        RECT 449.995000 239.380000 450.255000 240.715000 ;
        RECT 450.055000 239.210000 450.365000 239.270000 ;
        RECT 450.125000 239.140000 450.425000 239.210000 ;
        RECT 450.195000 239.070000 450.495000 239.140000 ;
        RECT 450.265000 239.000000 450.565000 239.070000 ;
        RECT 450.335000 238.930000 450.635000 239.000000 ;
        RECT 450.405000 238.860000 450.705000 238.930000 ;
        RECT 450.475000 238.790000 450.775000 238.860000 ;
        RECT 450.545000 238.720000 450.845000 238.790000 ;
        RECT 450.615000 238.650000 450.915000 238.720000 ;
        RECT 450.685000 238.580000 450.985000 238.650000 ;
        RECT 450.755000 238.510000 451.055000 238.580000 ;
        RECT 450.825000 238.440000 451.125000 238.510000 ;
        RECT 450.895000 238.370000 451.195000 238.440000 ;
        RECT 450.965000 238.300000 451.265000 238.370000 ;
        RECT 451.035000 238.230000 451.335000 238.300000 ;
        RECT 451.105000 238.160000 451.405000 238.230000 ;
        RECT 451.175000 238.090000 451.475000 238.160000 ;
        RECT 451.245000 238.020000 451.545000 238.090000 ;
        RECT 451.315000 237.950000 451.615000 238.020000 ;
        RECT 451.385000 237.880000 451.685000 237.950000 ;
        RECT 451.455000 237.810000 451.755000 237.880000 ;
        RECT 451.525000 237.740000 451.825000 237.810000 ;
        RECT 451.595000 237.670000 451.895000 237.740000 ;
        RECT 451.665000 237.600000 451.965000 237.670000 ;
        RECT 451.735000 237.530000 452.035000 237.600000 ;
        RECT 451.805000 237.460000 452.105000 237.530000 ;
        RECT 451.875000 237.390000 452.175000 237.460000 ;
        RECT 451.945000 237.320000 452.245000 237.390000 ;
        RECT 452.015000 237.250000 452.315000 237.320000 ;
        RECT 452.085000 237.180000 452.385000 237.250000 ;
        RECT 452.155000 237.110000 452.455000 237.180000 ;
        RECT 452.225000 237.040000 452.525000 237.110000 ;
        RECT 452.295000 236.970000 452.595000 237.040000 ;
        RECT 452.350000 236.915000 452.665000 236.970000 ;
        RECT 452.405000   0.000000 452.665000 236.860000 ;
        RECT 452.405000 236.860000 452.665000 236.915000 ;
    END
  END ENABLE_VDDA_H
  PIN HLD_H_N[0]
    ANTENNAGATEAREA  2.400000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.195000 36.690000 135.835000 36.950000 ;
        RECT 135.455000 36.685000 135.835000 36.690000 ;
        RECT 135.515000 36.625000 135.835000 36.685000 ;
        RECT 135.575000  0.000000 135.835000 36.565000 ;
        RECT 135.575000 36.565000 135.835000 36.625000 ;
    END
  END HLD_H_N[0]
  PIN HLD_H_N[1]
    ANTENNAGATEAREA  2.400000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.170000  0.000000 254.430000 36.565000 ;
        RECT 254.170000 36.565000 254.430000 36.625000 ;
        RECT 254.170000 36.625000 254.490000 36.685000 ;
        RECT 254.170000 36.685000 254.550000 36.690000 ;
        RECT 254.170000 36.690000 254.810000 36.950000 ;
    END
  END HLD_H_N[1]
  PIN HLD_H_N_REFGEN
    ANTENNAGATEAREA  2.400000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.955000 14.810000 405.595000 15.070000 ;
        RECT 404.975000 14.790000 405.360000 14.810000 ;
        RECT 404.995000  0.000000 405.255000 14.685000 ;
        RECT 404.995000 14.685000 405.255000 14.725000 ;
        RECT 404.995000 14.725000 405.295000 14.765000 ;
        RECT 404.995000 14.765000 405.335000 14.770000 ;
        RECT 404.995000 14.770000 405.340000 14.790000 ;
    END
  END HLD_H_N_REFGEN
  PIN HLD_OVR[0]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.995000 2.085000 141.635000 2.345000 ;
        RECT 141.040000 2.040000 141.590000 2.085000 ;
        RECT 141.085000 1.995000 141.545000 2.040000 ;
        RECT 141.090000 1.990000 141.545000 1.995000 ;
        RECT 141.145000 1.935000 141.545000 1.990000 ;
        RECT 141.200000 0.000000 141.545000 1.880000 ;
        RECT 141.200000 1.880000 141.545000 1.935000 ;
    END
  END HLD_OVR[0]
  PIN HLD_OVR[1]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.370000 2.085000 249.010000 2.345000 ;
        RECT 248.415000 2.040000 248.965000 2.085000 ;
        RECT 248.460000 0.000000 248.805000 1.880000 ;
        RECT 248.460000 1.880000 248.805000 1.935000 ;
        RECT 248.460000 1.935000 248.860000 1.990000 ;
        RECT 248.460000 1.990000 248.915000 1.995000 ;
        RECT 248.460000 1.995000 248.920000 2.040000 ;
    END
  END HLD_OVR[1]
  PIN IBUF_SEL[0]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.755000 29.985000 134.820000 30.055000 ;
        RECT 133.755000 30.055000 134.750000 30.125000 ;
        RECT 133.755000 30.125000 134.680000 30.195000 ;
        RECT 133.755000 30.195000 134.630000 30.245000 ;
        RECT 134.070000 30.245000 134.460000 30.305000 ;
        RECT 134.130000 30.305000 134.400000 30.365000 ;
        RECT 134.135000 30.365000 134.395000 30.370000 ;
        RECT 134.135000 30.370000 134.395000 42.740000 ;
        RECT 134.525000 29.980000 134.890000 29.985000 ;
        RECT 134.530000 29.975000 134.895000 29.980000 ;
        RECT 134.535000 29.970000 134.900000 29.975000 ;
        RECT 134.590000 29.915000 134.905000 29.970000 ;
        RECT 134.645000 29.370000 134.960000 29.425000 ;
        RECT 134.645000 29.425000 134.905000 29.480000 ;
        RECT 134.645000 29.480000 134.905000 29.860000 ;
        RECT 134.645000 29.860000 134.905000 29.915000 ;
        RECT 134.715000 29.300000 135.015000 29.370000 ;
        RECT 134.785000 29.230000 135.085000 29.300000 ;
        RECT 134.855000 29.160000 135.155000 29.230000 ;
        RECT 134.925000 29.090000 135.225000 29.160000 ;
        RECT 134.995000 29.020000 135.295000 29.090000 ;
        RECT 135.065000 28.950000 135.365000 29.020000 ;
        RECT 135.120000 28.895000 135.435000 28.950000 ;
        RECT 135.175000  0.000000 135.435000 28.840000 ;
        RECT 135.175000 28.840000 135.435000 28.895000 ;
    END
  END IBUF_SEL[0]
  PIN IBUF_SEL[1]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.570000  0.000000 254.830000 28.840000 ;
        RECT 254.570000 28.840000 254.830000 28.895000 ;
        RECT 254.570000 28.895000 254.885000 28.950000 ;
        RECT 254.640000 28.950000 254.940000 29.020000 ;
        RECT 254.710000 29.020000 255.010000 29.090000 ;
        RECT 254.780000 29.090000 255.080000 29.160000 ;
        RECT 254.850000 29.160000 255.150000 29.230000 ;
        RECT 254.920000 29.230000 255.220000 29.300000 ;
        RECT 254.990000 29.300000 255.290000 29.370000 ;
        RECT 255.045000 29.370000 255.360000 29.425000 ;
        RECT 255.100000 29.425000 255.360000 29.480000 ;
        RECT 255.100000 29.480000 255.360000 29.860000 ;
        RECT 255.100000 29.860000 255.360000 29.915000 ;
        RECT 255.100000 29.915000 255.415000 29.970000 ;
        RECT 255.105000 29.970000 255.470000 29.975000 ;
        RECT 255.110000 29.975000 255.475000 29.980000 ;
        RECT 255.115000 29.980000 255.480000 29.985000 ;
        RECT 255.185000 29.985000 256.250000 30.055000 ;
        RECT 255.255000 30.055000 256.250000 30.125000 ;
        RECT 255.325000 30.125000 256.250000 30.195000 ;
        RECT 255.375000 30.195000 256.250000 30.245000 ;
        RECT 255.545000 30.245000 255.935000 30.305000 ;
        RECT 255.605000 30.305000 255.875000 30.365000 ;
        RECT 255.610000 30.365000 255.870000 30.370000 ;
        RECT 255.610000 30.370000 255.870000 42.740000 ;
    END
  END IBUF_SEL[1]
  PIN IBUF_SEL_REFGEN
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.690000 0.000000 422.950000 23.140000 ;
    END
  END IBUF_SEL_REFGEN
  PIN IN[0]
    ANTENNAPARTIALMETALSIDEAREA  11.31440 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.005000 0.000000 142.265000 7.580000 ;
    END
  END IN[0]
  PIN IN[1]
    ANTENNAPARTIALMETALSIDEAREA  11.31440 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.740000 0.000000 248.000000 7.580000 ;
    END
  END IN[1]
  PIN INP_DIS[0]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.710000 0.000000 106.970000  1.240000 ;
        RECT 106.710000 1.240000 106.970000  1.295000 ;
        RECT 106.710000 1.295000 107.025000  1.350000 ;
        RECT 106.780000 1.350000 107.080000  1.420000 ;
        RECT 106.850000 1.420000 107.150000  1.490000 ;
        RECT 106.920000 1.490000 107.220000  1.560000 ;
        RECT 106.990000 1.560000 107.290000  1.630000 ;
        RECT 107.060000 1.630000 107.360000  1.700000 ;
        RECT 107.130000 1.700000 107.430000  1.770000 ;
        RECT 107.200000 1.770000 107.500000  1.840000 ;
        RECT 107.270000 1.840000 107.570000  1.910000 ;
        RECT 107.315000 1.910000 107.640000  1.955000 ;
        RECT 107.370000 1.955000 107.685000  2.010000 ;
        RECT 107.425000 2.010000 107.685000  2.065000 ;
        RECT 107.425000 2.065000 107.685000 18.155000 ;
    END
  END INP_DIS[0]
  PIN INP_DIS[1]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.320000 1.955000 282.635000  2.010000 ;
        RECT 282.320000 2.010000 282.580000  2.065000 ;
        RECT 282.320000 2.065000 282.580000 18.155000 ;
        RECT 282.365000 1.910000 282.690000  1.955000 ;
        RECT 282.435000 1.840000 282.735000  1.910000 ;
        RECT 282.505000 1.770000 282.805000  1.840000 ;
        RECT 282.575000 1.700000 282.875000  1.770000 ;
        RECT 282.645000 1.630000 282.945000  1.700000 ;
        RECT 282.715000 1.560000 283.015000  1.630000 ;
        RECT 282.785000 1.490000 283.085000  1.560000 ;
        RECT 282.855000 1.420000 283.155000  1.490000 ;
        RECT 282.925000 1.350000 283.225000  1.420000 ;
        RECT 282.980000 1.295000 283.295000  1.350000 ;
        RECT 283.035000 0.000000 283.295000  1.240000 ;
        RECT 283.035000 1.240000 283.295000  1.295000 ;
    END
  END INP_DIS[1]
  PIN IN_H[0]
    ANTENNAPARTIALMETALSIDEAREA  7.199500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.405000 0.000000 142.665000 10.590000 ;
    END
  END IN_H[0]
  PIN IN_H[1]
    ANTENNAPARTIALMETALSIDEAREA  7.199500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.340000 0.000000 247.600000 10.590000 ;
    END
  END IN_H[1]
  PIN OE_N[0]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.255000 49.355000 145.895000 49.615000 ;
        RECT 145.515000 49.350000 145.895000 49.355000 ;
        RECT 145.575000 49.290000 145.895000 49.350000 ;
        RECT 145.635000 28.390000 145.950000 28.445000 ;
        RECT 145.635000 28.445000 145.895000 28.500000 ;
        RECT 145.635000 28.500000 145.895000 49.230000 ;
        RECT 145.635000 49.230000 145.895000 49.290000 ;
        RECT 145.705000 28.320000 146.005000 28.390000 ;
        RECT 145.775000 28.250000 146.075000 28.320000 ;
        RECT 145.845000 28.180000 146.145000 28.250000 ;
        RECT 145.915000 28.110000 146.215000 28.180000 ;
        RECT 145.985000 28.040000 146.285000 28.110000 ;
        RECT 146.055000 27.970000 146.355000 28.040000 ;
        RECT 146.125000 27.900000 146.425000 27.970000 ;
        RECT 146.195000 27.830000 146.495000 27.900000 ;
        RECT 146.265000 27.760000 146.565000 27.830000 ;
        RECT 146.335000 27.690000 146.635000 27.760000 ;
        RECT 146.405000 27.620000 146.705000 27.690000 ;
        RECT 146.475000 27.550000 146.775000 27.620000 ;
        RECT 146.545000 27.480000 146.845000 27.550000 ;
        RECT 146.615000 27.410000 146.915000 27.480000 ;
        RECT 146.685000 27.340000 146.985000 27.410000 ;
        RECT 146.755000 27.270000 147.055000 27.340000 ;
        RECT 146.825000 27.200000 147.125000 27.270000 ;
        RECT 146.895000 27.130000 147.195000 27.200000 ;
        RECT 146.965000 27.060000 147.265000 27.130000 ;
        RECT 147.035000 26.990000 147.335000 27.060000 ;
        RECT 147.105000 26.920000 147.405000 26.990000 ;
        RECT 147.160000 26.865000 147.475000 26.920000 ;
        RECT 147.215000  0.000000 147.475000 26.810000 ;
        RECT 147.215000 26.810000 147.475000 26.865000 ;
    END
  END OE_N[0]
  PIN OE_N[1]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.530000  0.000000 242.790000 26.810000 ;
        RECT 242.530000 26.810000 242.790000 26.865000 ;
        RECT 242.530000 26.865000 242.845000 26.920000 ;
        RECT 242.600000 26.920000 242.900000 26.990000 ;
        RECT 242.670000 26.990000 242.970000 27.060000 ;
        RECT 242.740000 27.060000 243.040000 27.130000 ;
        RECT 242.810000 27.130000 243.110000 27.200000 ;
        RECT 242.880000 27.200000 243.180000 27.270000 ;
        RECT 242.950000 27.270000 243.250000 27.340000 ;
        RECT 243.020000 27.340000 243.320000 27.410000 ;
        RECT 243.090000 27.410000 243.390000 27.480000 ;
        RECT 243.160000 27.480000 243.460000 27.550000 ;
        RECT 243.230000 27.550000 243.530000 27.620000 ;
        RECT 243.300000 27.620000 243.600000 27.690000 ;
        RECT 243.370000 27.690000 243.670000 27.760000 ;
        RECT 243.440000 27.760000 243.740000 27.830000 ;
        RECT 243.510000 27.830000 243.810000 27.900000 ;
        RECT 243.580000 27.900000 243.880000 27.970000 ;
        RECT 243.650000 27.970000 243.950000 28.040000 ;
        RECT 243.720000 28.040000 244.020000 28.110000 ;
        RECT 243.790000 28.110000 244.090000 28.180000 ;
        RECT 243.860000 28.180000 244.160000 28.250000 ;
        RECT 243.930000 28.250000 244.230000 28.320000 ;
        RECT 244.000000 28.320000 244.300000 28.390000 ;
        RECT 244.055000 28.390000 244.370000 28.445000 ;
        RECT 244.110000 28.445000 244.370000 28.500000 ;
        RECT 244.110000 28.500000 244.370000 49.230000 ;
        RECT 244.110000 49.230000 244.370000 49.290000 ;
        RECT 244.110000 49.290000 244.430000 49.350000 ;
        RECT 244.110000 49.350000 244.490000 49.355000 ;
        RECT 244.110000 49.355000 244.750000 49.615000 ;
    END
  END OE_N[1]
  PIN OUT[0]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.455000  0.000000 121.715000 45.840000 ;
        RECT 121.455000 45.840000 121.715000 45.910000 ;
        RECT 121.455000 45.910000 121.785000 45.980000 ;
        RECT 121.455000 45.980000 121.855000 46.020000 ;
        RECT 121.455000 46.020000 124.575000 46.090000 ;
        RECT 121.455000 46.090000 124.645000 46.160000 ;
        RECT 121.455000 46.160000 124.715000 46.230000 ;
        RECT 121.455000 46.230000 124.785000 46.280000 ;
        RECT 124.535000 46.280000 124.835000 46.350000 ;
        RECT 124.605000 46.350000 124.905000 46.420000 ;
        RECT 124.675000 46.420000 124.975000 46.490000 ;
        RECT 124.745000 46.490000 125.045000 46.560000 ;
        RECT 124.815000 46.560000 125.115000 46.630000 ;
        RECT 124.885000 46.630000 125.185000 46.700000 ;
        RECT 124.955000 46.700000 125.255000 46.770000 ;
        RECT 125.025000 46.770000 125.325000 46.840000 ;
        RECT 125.095000 46.840000 125.395000 46.910000 ;
        RECT 125.165000 46.910000 125.465000 46.980000 ;
        RECT 125.235000 46.980000 125.535000 47.050000 ;
        RECT 125.305000 47.050000 125.605000 47.120000 ;
        RECT 125.350000 48.970000 126.055000 51.845000 ;
        RECT 125.375000 47.120000 125.675000 47.190000 ;
        RECT 125.420000 48.900000 125.985000 48.970000 ;
        RECT 125.445000 47.190000 125.745000 47.260000 ;
        RECT 125.490000 48.830000 125.915000 48.900000 ;
        RECT 125.515000 47.260000 125.815000 47.330000 ;
        RECT 125.515000 48.805000 125.915000 48.830000 ;
        RECT 125.545000 47.330000 125.885000 47.360000 ;
        RECT 125.585000 48.735000 125.915000 48.805000 ;
        RECT 125.600000 47.360000 125.915000 47.415000 ;
        RECT 125.655000 47.415000 125.915000 47.470000 ;
        RECT 125.655000 47.470000 125.915000 48.665000 ;
        RECT 125.655000 48.665000 125.915000 48.735000 ;
    END
  END OUT[0]
  PIN OUT[1]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.950000 48.970000 264.655000 51.845000 ;
        RECT 264.020000 48.900000 264.585000 48.970000 ;
        RECT 264.090000 47.360000 264.405000 47.415000 ;
        RECT 264.090000 47.415000 264.350000 47.470000 ;
        RECT 264.090000 47.470000 264.350000 48.665000 ;
        RECT 264.090000 48.665000 264.350000 48.735000 ;
        RECT 264.090000 48.735000 264.420000 48.805000 ;
        RECT 264.090000 48.805000 264.490000 48.830000 ;
        RECT 264.090000 48.830000 264.515000 48.900000 ;
        RECT 264.120000 47.330000 264.460000 47.360000 ;
        RECT 264.190000 47.260000 264.490000 47.330000 ;
        RECT 264.260000 47.190000 264.560000 47.260000 ;
        RECT 264.330000 47.120000 264.630000 47.190000 ;
        RECT 264.400000 47.050000 264.700000 47.120000 ;
        RECT 264.470000 46.980000 264.770000 47.050000 ;
        RECT 264.540000 46.910000 264.840000 46.980000 ;
        RECT 264.610000 46.840000 264.910000 46.910000 ;
        RECT 264.680000 46.770000 264.980000 46.840000 ;
        RECT 264.750000 46.700000 265.050000 46.770000 ;
        RECT 264.820000 46.630000 265.120000 46.700000 ;
        RECT 264.890000 46.560000 265.190000 46.630000 ;
        RECT 264.960000 46.490000 265.260000 46.560000 ;
        RECT 265.030000 46.420000 265.330000 46.490000 ;
        RECT 265.100000 46.350000 265.400000 46.420000 ;
        RECT 265.170000 46.280000 265.470000 46.350000 ;
        RECT 265.220000 46.230000 268.550000 46.280000 ;
        RECT 265.290000 46.160000 268.550000 46.230000 ;
        RECT 265.360000 46.090000 268.550000 46.160000 ;
        RECT 265.430000 46.020000 268.550000 46.090000 ;
        RECT 268.150000 45.980000 268.550000 46.020000 ;
        RECT 268.220000 45.910000 268.550000 45.980000 ;
        RECT 268.290000  0.000000 268.550000 45.840000 ;
        RECT 268.290000 45.840000 268.550000 45.910000 ;
    END
  END OUT[1]
  PIN PAD[0]
    ANTENNAPARTIALMETALSIDEAREA  200.9870 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 105.790000 132.205000 171.190000 194.545000 ;
        RECT 105.920000 132.075000 171.060000 132.205000 ;
        RECT 106.190000 194.545000 170.790000 194.945000 ;
        RECT 106.320000 131.675000 170.660000 132.075000 ;
        RECT 106.590000 194.945000 170.390000 195.345000 ;
        RECT 106.720000 131.275000 170.260000 131.675000 ;
        RECT 106.990000 195.345000 169.990000 195.745000 ;
        RECT 107.120000 130.875000 169.860000 131.275000 ;
        RECT 107.390000 195.745000 169.590000 196.145000 ;
        RECT 107.520000 130.475000 169.460000 130.875000 ;
        RECT 107.790000 196.145000 169.190000 196.545000 ;
        RECT 107.920000 130.075000 169.060000 130.475000 ;
        RECT 108.190000 196.545000 168.790000 196.945000 ;
        RECT 108.320000 129.675000 168.660000 130.075000 ;
        RECT 108.590000 196.945000 168.390000 197.345000 ;
        RECT 108.720000 129.275000 168.260000 129.675000 ;
        RECT 108.990000 197.345000 167.990000 197.745000 ;
        RECT 109.120000 128.875000 167.860000 129.275000 ;
        RECT 109.390000 197.745000 167.590000 198.145000 ;
        RECT 109.520000 128.475000 167.460000 128.875000 ;
        RECT 109.790000 198.145000 167.190000 198.545000 ;
        RECT 109.920000 128.075000 167.060000 128.475000 ;
        RECT 110.190000 198.545000 166.790000 198.945000 ;
        RECT 110.320000 127.675000 166.660000 128.075000 ;
        RECT 110.590000 198.945000 166.390000 199.345000 ;
        RECT 110.720000 127.275000 166.260000 127.675000 ;
        RECT 110.990000 199.345000 165.990000 199.745000 ;
        RECT 111.120000 126.875000 165.860000 127.275000 ;
        RECT 111.390000 199.745000 165.590000 200.145000 ;
        RECT 111.520000 126.475000 165.460000 126.875000 ;
        RECT 111.790000 200.145000 165.190000 200.545000 ;
        RECT 111.920000 126.075000 165.060000 126.475000 ;
        RECT 112.190000 200.545000 164.790000 200.945000 ;
        RECT 112.320000 125.675000 164.660000 126.075000 ;
        RECT 112.320000 200.945000 164.660000 201.075000 ;
    END
  END PAD[0]
  PIN PAD[1]
    ANTENNAPARTIALMETALSIDEAREA  200.9870 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 218.815000 132.205000 284.215000 194.545000 ;
        RECT 218.945000 132.075000 284.085000 132.205000 ;
        RECT 219.215000 194.545000 283.815000 194.945000 ;
        RECT 219.345000 131.675000 283.685000 132.075000 ;
        RECT 219.615000 194.945000 283.415000 195.345000 ;
        RECT 219.745000 131.275000 283.285000 131.675000 ;
        RECT 220.015000 195.345000 283.015000 195.745000 ;
        RECT 220.145000 130.875000 282.885000 131.275000 ;
        RECT 220.415000 195.745000 282.615000 196.145000 ;
        RECT 220.545000 130.475000 282.485000 130.875000 ;
        RECT 220.815000 196.145000 282.215000 196.545000 ;
        RECT 220.945000 130.075000 282.085000 130.475000 ;
        RECT 221.215000 196.545000 281.815000 196.945000 ;
        RECT 221.345000 129.675000 281.685000 130.075000 ;
        RECT 221.615000 196.945000 281.415000 197.345000 ;
        RECT 221.745000 129.275000 281.285000 129.675000 ;
        RECT 222.015000 197.345000 281.015000 197.745000 ;
        RECT 222.145000 128.875000 280.885000 129.275000 ;
        RECT 222.415000 197.745000 280.615000 198.145000 ;
        RECT 222.545000 128.475000 280.485000 128.875000 ;
        RECT 222.815000 198.145000 280.215000 198.545000 ;
        RECT 222.945000 128.075000 280.085000 128.475000 ;
        RECT 223.215000 198.545000 279.815000 198.945000 ;
        RECT 223.345000 127.675000 279.685000 128.075000 ;
        RECT 223.615000 198.945000 279.415000 199.345000 ;
        RECT 223.745000 127.275000 279.285000 127.675000 ;
        RECT 224.015000 199.345000 279.015000 199.745000 ;
        RECT 224.145000 126.875000 278.885000 127.275000 ;
        RECT 224.415000 199.745000 278.615000 200.145000 ;
        RECT 224.545000 126.475000 278.485000 126.875000 ;
        RECT 224.815000 200.145000 278.215000 200.545000 ;
        RECT 224.945000 126.075000 278.085000 126.475000 ;
        RECT 225.215000 200.545000 277.815000 200.945000 ;
        RECT 225.345000 125.675000 277.685000 126.075000 ;
        RECT 225.345000 200.945000 277.685000 201.075000 ;
    END
  END PAD[1]
  PIN PAD_A_ESD_0_H[0]
    ANTENNAPARTIALMETALSIDEAREA  21.16800 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.260000 0.000000 86.105000 30.545000 ;
    END
  END PAD_A_ESD_0_H[0]
  PIN PAD_A_ESD_0_H[1]
    ANTENNAPARTIALMETALSIDEAREA  21.16800 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.900000 0.000000 304.745000 30.545000 ;
    END
  END PAD_A_ESD_0_H[1]
  PIN PAD_A_ESD_1_H[0]
    ANTENNAPARTIALMETALSIDEAREA  16.74750 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.990000 0.000000 178.990000 24.230000 ;
    END
  END PAD_A_ESD_1_H[0]
  PIN PAD_A_ESD_1_H[1]
    ANTENNAPARTIALMETALSIDEAREA  16.74750 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.015000 0.000000 213.015000 24.230000 ;
    END
  END PAD_A_ESD_1_H[1]
  PIN PAD_A_NOESD_H[0]
    ANTENNAPARTIALMETALSIDEAREA  23.05100 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.245000 0.000000 87.095000 33.235000 ;
    END
  END PAD_A_NOESD_H[0]
  PIN PAD_A_NOESD_H[1]
    ANTENNAPARTIALMETALSIDEAREA  23.05450 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.910000 0.000000 303.760000 33.235000 ;
    END
  END PAD_A_NOESD_H[1]
  PIN SLOW[0]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.615000 0.000000 147.875000 46.135000 ;
    END
  END SLOW[0]
  PIN SLOW[1]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.130000 0.000000 242.390000 46.135000 ;
    END
  END SLOW[1]
  PIN TIE_LO_ESD[0]
    ANTENNAGATEAREA  2.400000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  92.305000 102.985000  92.635000 103.025000 ;
        RECT  92.305000 103.025000  92.595000 103.065000 ;
        RECT  92.305000 103.065000  92.595000 111.375000 ;
        RECT  92.305000 111.375000  92.595000 111.435000 ;
        RECT  92.305000 111.435000  92.655000 111.495000 ;
        RECT  92.305000 111.495000  92.715000 111.500000 ;
        RECT  92.305000 111.500000  93.345000 111.600000 ;
        RECT  92.350000 102.940000  92.675000 102.985000 ;
        RECT  92.375000 111.600000  93.345000 111.670000 ;
        RECT  92.420000 102.870000  92.720000 102.940000 ;
        RECT  92.445000 111.670000  93.345000 111.740000 ;
        RECT  92.465000 111.740000  93.345000 111.760000 ;
        RECT  92.490000 102.800000  92.790000 102.870000 ;
        RECT  92.560000 102.730000  92.860000 102.800000 ;
        RECT  92.630000 102.660000  92.930000 102.730000 ;
        RECT  92.700000 102.590000  93.000000 102.660000 ;
        RECT  92.770000 102.520000  93.070000 102.590000 ;
        RECT  92.840000 102.450000  93.140000 102.520000 ;
        RECT  92.910000 102.380000  93.210000 102.450000 ;
        RECT  92.980000 102.310000  93.280000 102.380000 ;
        RECT  93.015000 111.760000  93.345000 111.830000 ;
        RECT  93.050000 102.240000  93.350000 102.310000 ;
        RECT  93.085000 111.830000  93.345000 111.900000 ;
        RECT  93.085000 111.900000  93.345000 112.140000 ;
        RECT  93.120000 102.170000  93.420000 102.240000 ;
        RECT  93.190000 102.100000  93.490000 102.170000 ;
        RECT  93.260000 102.030000  93.560000 102.100000 ;
        RECT  93.330000 101.960000  93.630000 102.030000 ;
        RECT  93.400000 101.890000  93.700000 101.960000 ;
        RECT  93.470000 101.820000  93.770000 101.890000 ;
        RECT  93.540000 101.750000  93.840000 101.820000 ;
        RECT  93.610000 101.680000  93.910000 101.750000 ;
        RECT  93.680000 101.610000  93.980000 101.680000 ;
        RECT  93.750000 101.540000  94.050000 101.610000 ;
        RECT  93.820000 101.470000  94.120000 101.540000 ;
        RECT  93.890000 101.400000  94.190000 101.470000 ;
        RECT  93.960000 101.330000  94.260000 101.400000 ;
        RECT  94.030000 101.260000  94.330000 101.330000 ;
        RECT  94.100000 101.190000  94.400000 101.260000 ;
        RECT  94.170000 101.120000  94.470000 101.190000 ;
        RECT  94.240000 101.050000  94.540000 101.120000 ;
        RECT  94.310000 100.980000  94.610000 101.050000 ;
        RECT  94.380000 100.910000  94.680000 100.980000 ;
        RECT  94.450000 100.840000  94.750000 100.910000 ;
        RECT  94.520000 100.770000  94.820000 100.840000 ;
        RECT  94.590000 100.700000  94.890000 100.770000 ;
        RECT  94.660000 100.630000  94.960000 100.700000 ;
        RECT  94.730000 100.560000  95.030000 100.630000 ;
        RECT  94.800000 100.490000  95.100000 100.560000 ;
        RECT  94.870000 100.420000  95.170000 100.490000 ;
        RECT  94.940000 100.350000  95.240000 100.420000 ;
        RECT  95.010000 100.280000  95.310000 100.350000 ;
        RECT  95.080000 100.210000  95.380000 100.280000 ;
        RECT  95.150000 100.140000  95.450000 100.210000 ;
        RECT  95.220000 100.070000  95.520000 100.140000 ;
        RECT  95.290000 100.000000  95.590000 100.070000 ;
        RECT  95.360000  99.930000  95.660000 100.000000 ;
        RECT  95.430000  99.860000  95.730000  99.930000 ;
        RECT  95.500000  99.790000  95.800000  99.860000 ;
        RECT  95.570000  99.720000  95.870000  99.790000 ;
        RECT  95.640000  99.650000  95.940000  99.720000 ;
        RECT  95.710000  99.580000  96.010000  99.650000 ;
        RECT  95.780000  99.510000  96.080000  99.580000 ;
        RECT  95.850000  99.440000  96.150000  99.510000 ;
        RECT  95.920000  99.370000  96.220000  99.440000 ;
        RECT  95.990000  99.300000  96.290000  99.370000 ;
        RECT  96.060000  99.230000  96.360000  99.300000 ;
        RECT  96.130000  99.160000  96.430000  99.230000 ;
        RECT  96.200000  99.090000  96.500000  99.160000 ;
        RECT  96.270000  99.020000  96.570000  99.090000 ;
        RECT  96.340000  98.950000  96.640000  99.020000 ;
        RECT  96.410000  98.880000  96.710000  98.950000 ;
        RECT  96.480000  98.810000  96.780000  98.880000 ;
        RECT  96.550000  98.740000  96.850000  98.810000 ;
        RECT  96.620000  98.670000  96.920000  98.740000 ;
        RECT  96.690000  98.600000  96.990000  98.670000 ;
        RECT  96.760000  98.530000  97.060000  98.600000 ;
        RECT  96.830000  98.460000  97.130000  98.530000 ;
        RECT  96.900000  98.390000  97.200000  98.460000 ;
        RECT  96.970000  98.320000  97.270000  98.390000 ;
        RECT  97.040000  98.250000  97.340000  98.320000 ;
        RECT  97.110000  98.180000  97.410000  98.250000 ;
        RECT  97.180000  98.110000  97.480000  98.180000 ;
        RECT  97.250000  98.040000  97.550000  98.110000 ;
        RECT  97.320000  97.970000  97.620000  98.040000 ;
        RECT  97.390000  97.900000  97.690000  97.970000 ;
        RECT  97.460000  97.830000  97.760000  97.900000 ;
        RECT  97.530000  97.760000  97.830000  97.830000 ;
        RECT  97.600000  97.690000  97.900000  97.760000 ;
        RECT  97.670000  97.620000  97.970000  97.690000 ;
        RECT  97.740000  97.550000  98.040000  97.620000 ;
        RECT  97.810000  97.480000  98.110000  97.550000 ;
        RECT  97.880000  97.410000  98.180000  97.480000 ;
        RECT  97.950000  97.340000  98.250000  97.410000 ;
        RECT  98.020000  97.270000  98.320000  97.340000 ;
        RECT  98.090000  97.200000  98.390000  97.270000 ;
        RECT  98.160000  97.130000  98.460000  97.200000 ;
        RECT  98.230000  97.060000  98.530000  97.130000 ;
        RECT  98.300000  96.990000  98.600000  97.060000 ;
        RECT  98.370000  96.920000  98.670000  96.990000 ;
        RECT  98.440000  96.850000  98.740000  96.920000 ;
        RECT  98.510000  96.780000  98.810000  96.850000 ;
        RECT  98.580000  96.710000  98.880000  96.780000 ;
        RECT  98.650000  96.640000  98.950000  96.710000 ;
        RECT  98.720000  96.570000  99.020000  96.640000 ;
        RECT  98.790000  96.500000  99.090000  96.570000 ;
        RECT  98.860000  96.430000  99.160000  96.500000 ;
        RECT  98.930000  96.360000  99.230000  96.430000 ;
        RECT  99.000000  96.290000  99.300000  96.360000 ;
        RECT  99.070000  96.220000  99.370000  96.290000 ;
        RECT  99.140000  96.150000  99.440000  96.220000 ;
        RECT  99.210000  96.080000  99.510000  96.150000 ;
        RECT  99.280000  96.010000  99.580000  96.080000 ;
        RECT  99.350000  95.940000  99.650000  96.010000 ;
        RECT  99.420000  95.870000  99.720000  95.940000 ;
        RECT  99.490000  95.800000  99.790000  95.870000 ;
        RECT  99.560000  95.730000  99.860000  95.800000 ;
        RECT  99.630000  95.660000  99.930000  95.730000 ;
        RECT  99.700000  95.590000 100.000000  95.660000 ;
        RECT  99.770000  95.520000 100.070000  95.590000 ;
        RECT  99.840000  95.450000 100.140000  95.520000 ;
        RECT  99.910000  95.380000 100.210000  95.450000 ;
        RECT  99.980000  95.310000 100.280000  95.380000 ;
        RECT 100.050000  95.240000 100.350000  95.310000 ;
        RECT 100.120000  95.170000 100.420000  95.240000 ;
        RECT 100.190000  95.100000 100.490000  95.170000 ;
        RECT 100.260000  95.030000 100.560000  95.100000 ;
        RECT 100.330000  94.960000 100.630000  95.030000 ;
        RECT 100.380000  94.910000 105.385000  94.960000 ;
        RECT 100.450000  94.840000 105.435000  94.910000 ;
        RECT 100.520000  94.770000 105.505000  94.840000 ;
        RECT 100.590000  94.700000 105.575000  94.770000 ;
        RECT 105.305000  94.670000 105.645000  94.700000 ;
        RECT 105.375000  94.600000 105.675000  94.670000 ;
        RECT 105.445000  94.530000 105.745000  94.600000 ;
        RECT 105.515000  94.460000 105.815000  94.530000 ;
        RECT 105.585000  94.390000 105.885000  94.460000 ;
        RECT 105.655000  94.320000 105.955000  94.390000 ;
        RECT 105.725000  94.250000 106.025000  94.320000 ;
        RECT 105.730000  94.245000 106.095000  94.250000 ;
        RECT 105.770000  94.205000 106.095000  94.245000 ;
        RECT 105.810000  89.480000 106.140000  89.520000 ;
        RECT 105.810000  89.520000 106.100000  89.560000 ;
        RECT 105.810000  89.560000 106.095000  89.565000 ;
        RECT 105.810000  89.565000 106.095000  94.165000 ;
        RECT 105.810000  94.165000 106.095000  94.205000 ;
        RECT 105.820000  89.470000 106.180000  89.480000 ;
        RECT 105.890000  89.400000 106.190000  89.470000 ;
        RECT 105.960000  89.330000 106.260000  89.400000 ;
        RECT 106.030000  89.260000 106.330000  89.330000 ;
        RECT 106.100000  89.190000 106.400000  89.260000 ;
        RECT 106.170000  89.120000 106.470000  89.190000 ;
        RECT 106.240000  89.050000 106.540000  89.120000 ;
        RECT 106.310000  88.980000 106.610000  89.050000 ;
        RECT 106.380000  88.910000 106.680000  88.980000 ;
        RECT 106.450000  88.840000 106.750000  88.910000 ;
        RECT 106.520000  88.770000 106.820000  88.840000 ;
        RECT 106.590000  88.700000 106.890000  88.770000 ;
        RECT 106.660000  88.630000 106.960000  88.700000 ;
        RECT 106.730000  88.560000 107.030000  88.630000 ;
        RECT 106.800000  88.490000 107.100000  88.560000 ;
        RECT 106.870000  88.420000 107.170000  88.490000 ;
        RECT 106.940000  88.350000 107.240000  88.420000 ;
        RECT 107.010000  88.280000 107.310000  88.350000 ;
        RECT 107.080000  88.210000 107.380000  88.280000 ;
        RECT 107.150000  88.140000 107.450000  88.210000 ;
        RECT 107.220000  88.070000 107.520000  88.140000 ;
        RECT 107.290000  88.000000 107.590000  88.070000 ;
        RECT 107.360000  87.930000 107.660000  88.000000 ;
        RECT 107.430000  87.860000 107.730000  87.930000 ;
        RECT 107.500000  87.790000 107.800000  87.860000 ;
        RECT 107.570000  87.720000 107.870000  87.790000 ;
        RECT 107.640000  87.650000 107.940000  87.720000 ;
        RECT 107.695000  87.595000 108.010000  87.650000 ;
        RECT 107.750000  76.510000 108.065000  76.565000 ;
        RECT 107.750000  76.565000 108.010000  76.620000 ;
        RECT 107.750000  76.620000 108.010000  87.540000 ;
        RECT 107.750000  87.540000 108.010000  87.595000 ;
        RECT 107.800000  76.460000 108.120000  76.510000 ;
        RECT 107.870000  76.390000 108.170000  76.460000 ;
        RECT 107.940000  76.320000 108.240000  76.390000 ;
        RECT 108.010000  76.250000 108.310000  76.320000 ;
        RECT 108.080000  76.180000 108.380000  76.250000 ;
        RECT 108.150000  76.110000 108.450000  76.180000 ;
        RECT 108.220000  76.040000 108.520000  76.110000 ;
        RECT 108.290000  75.970000 108.590000  76.040000 ;
        RECT 108.360000  75.900000 108.660000  75.970000 ;
        RECT 108.430000  75.830000 108.730000  75.900000 ;
        RECT 108.500000  75.760000 108.800000  75.830000 ;
        RECT 108.570000  47.460000 108.885000  47.515000 ;
        RECT 108.570000  47.515000 108.830000  47.570000 ;
        RECT 108.570000  47.570000 108.830000  56.455000 ;
        RECT 108.570000  56.455000 108.830000  56.510000 ;
        RECT 108.570000  56.510000 108.885000  56.565000 ;
        RECT 108.570000  75.690000 108.870000  75.760000 ;
        RECT 108.585000  47.445000 108.940000  47.460000 ;
        RECT 108.640000  56.565000 108.940000  56.635000 ;
        RECT 108.640000  75.620000 108.940000  75.690000 ;
        RECT 108.655000  47.375000 108.955000  47.445000 ;
        RECT 108.710000  56.635000 109.010000  56.705000 ;
        RECT 108.710000  75.550000 109.010000  75.620000 ;
        RECT 108.725000  47.305000 109.025000  47.375000 ;
        RECT 108.780000  56.705000 109.080000  56.775000 ;
        RECT 108.780000  75.480000 109.080000  75.550000 ;
        RECT 108.795000  47.235000 109.095000  47.305000 ;
        RECT 108.850000  56.775000 109.150000  56.845000 ;
        RECT 108.850000  75.410000 109.150000  75.480000 ;
        RECT 108.865000  47.165000 109.165000  47.235000 ;
        RECT 108.920000  56.845000 109.220000  56.915000 ;
        RECT 108.920000  75.340000 109.220000  75.410000 ;
        RECT 108.935000  47.095000 109.235000  47.165000 ;
        RECT 108.990000  56.915000 109.290000  56.985000 ;
        RECT 108.990000  75.270000 109.290000  75.340000 ;
        RECT 109.005000  47.025000 109.305000  47.095000 ;
        RECT 109.060000  56.985000 109.360000  57.055000 ;
        RECT 109.060000  75.200000 109.360000  75.270000 ;
        RECT 109.075000  46.955000 109.375000  47.025000 ;
        RECT 109.130000  57.055000 109.430000  57.125000 ;
        RECT 109.130000  75.130000 109.430000  75.200000 ;
        RECT 109.145000  46.885000 109.445000  46.955000 ;
        RECT 109.200000  57.125000 109.500000  57.195000 ;
        RECT 109.200000  75.060000 109.500000  75.130000 ;
        RECT 109.215000  46.815000 109.515000  46.885000 ;
        RECT 109.270000  57.195000 109.570000  57.265000 ;
        RECT 109.270000  74.990000 109.570000  75.060000 ;
        RECT 109.285000  46.745000 109.585000  46.815000 ;
        RECT 109.325000  57.265000 109.640000  57.320000 ;
        RECT 109.325000  74.935000 109.640000  74.990000 ;
        RECT 109.355000  46.675000 109.655000  46.745000 ;
        RECT 109.380000  57.320000 109.640000  57.375000 ;
        RECT 109.380000  57.375000 109.640000  74.880000 ;
        RECT 109.380000  74.880000 109.640000  74.935000 ;
        RECT 109.410000  46.620000 109.725000  46.675000 ;
        RECT 109.465000  45.850000 109.780000  45.905000 ;
        RECT 109.465000  45.905000 109.725000  45.960000 ;
        RECT 109.465000  45.960000 109.725000  46.565000 ;
        RECT 109.465000  46.565000 109.725000  46.620000 ;
        RECT 109.515000  45.800000 109.835000  45.850000 ;
        RECT 109.585000  45.730000 109.885000  45.800000 ;
        RECT 109.655000  45.660000 109.955000  45.730000 ;
        RECT 109.725000  45.590000 110.025000  45.660000 ;
        RECT 109.780000  45.535000 110.095000  45.590000 ;
        RECT 109.815000  17.630000 110.130000  17.685000 ;
        RECT 109.815000  17.685000 110.075000  17.740000 ;
        RECT 109.815000  17.740000 110.075000  36.300000 ;
        RECT 109.815000  36.300000 110.075000  36.310000 ;
        RECT 109.815000  36.310000 110.085000  36.320000 ;
        RECT 109.815000  36.320000 110.095000  36.410000 ;
        RECT 109.825000  36.410000 110.095000  36.420000 ;
        RECT 109.835000  36.420000 110.095000  36.430000 ;
        RECT 109.835000  36.430000 110.095000  45.480000 ;
        RECT 109.835000  45.480000 110.095000  45.535000 ;
        RECT 109.840000  17.605000 110.185000  17.630000 ;
        RECT 109.910000  17.535000 110.210000  17.605000 ;
        RECT 109.980000  17.465000 110.280000  17.535000 ;
        RECT 110.035000  17.410000 110.350000  17.465000 ;
        RECT 110.090000   0.000000 110.350000  17.355000 ;
        RECT 110.090000  17.355000 110.350000  17.410000 ;
    END
  END TIE_LO_ESD[0]
  PIN TIE_LO_ESD[1]
    ANTENNAGATEAREA  2.400000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.655000   0.000000 279.915000  17.355000 ;
        RECT 279.655000  17.355000 279.915000  17.410000 ;
        RECT 279.655000  17.410000 279.970000  17.465000 ;
        RECT 279.725000  17.465000 280.025000  17.535000 ;
        RECT 279.795000  17.535000 280.095000  17.605000 ;
        RECT 279.820000  17.605000 280.165000  17.630000 ;
        RECT 279.875000  17.630000 280.190000  17.685000 ;
        RECT 279.910000  36.320000 280.190000  36.410000 ;
        RECT 279.910000  36.410000 280.180000  36.420000 ;
        RECT 279.910000  36.420000 280.170000  36.430000 ;
        RECT 279.910000  36.430000 280.170000  45.480000 ;
        RECT 279.910000  45.480000 280.170000  45.535000 ;
        RECT 279.910000  45.535000 280.225000  45.590000 ;
        RECT 279.920000  36.310000 280.190000  36.320000 ;
        RECT 279.930000  17.685000 280.190000  17.740000 ;
        RECT 279.930000  17.740000 280.190000  36.300000 ;
        RECT 279.930000  36.300000 280.190000  36.310000 ;
        RECT 279.980000  45.590000 280.280000  45.660000 ;
        RECT 280.050000  45.660000 280.350000  45.730000 ;
        RECT 280.120000  45.730000 280.420000  45.800000 ;
        RECT 280.170000  45.800000 280.490000  45.850000 ;
        RECT 280.225000  45.850000 280.540000  45.905000 ;
        RECT 280.280000  45.905000 280.540000  45.960000 ;
        RECT 280.280000  45.960000 280.540000  46.565000 ;
        RECT 280.280000  46.565000 280.540000  46.620000 ;
        RECT 280.280000  46.620000 280.595000  46.675000 ;
        RECT 280.350000  46.675000 280.650000  46.745000 ;
        RECT 280.365000  57.265000 280.680000  57.320000 ;
        RECT 280.365000  57.320000 280.625000  57.375000 ;
        RECT 280.365000  57.375000 280.625000  74.880000 ;
        RECT 280.365000  74.880000 280.625000  74.935000 ;
        RECT 280.365000  74.935000 280.680000  74.990000 ;
        RECT 280.420000  46.745000 280.720000  46.815000 ;
        RECT 280.435000  57.195000 280.735000  57.265000 ;
        RECT 280.435000  74.990000 280.735000  75.060000 ;
        RECT 280.490000  46.815000 280.790000  46.885000 ;
        RECT 280.505000  57.125000 280.805000  57.195000 ;
        RECT 280.505000  75.060000 280.805000  75.130000 ;
        RECT 280.560000  46.885000 280.860000  46.955000 ;
        RECT 280.575000  57.055000 280.875000  57.125000 ;
        RECT 280.575000  75.130000 280.875000  75.200000 ;
        RECT 280.630000  46.955000 280.930000  47.025000 ;
        RECT 280.645000  56.985000 280.945000  57.055000 ;
        RECT 280.645000  75.200000 280.945000  75.270000 ;
        RECT 280.700000  47.025000 281.000000  47.095000 ;
        RECT 280.715000  56.915000 281.015000  56.985000 ;
        RECT 280.715000  75.270000 281.015000  75.340000 ;
        RECT 280.770000  47.095000 281.070000  47.165000 ;
        RECT 280.785000  56.845000 281.085000  56.915000 ;
        RECT 280.785000  75.340000 281.085000  75.410000 ;
        RECT 280.840000  47.165000 281.140000  47.235000 ;
        RECT 280.855000  56.775000 281.155000  56.845000 ;
        RECT 280.855000  75.410000 281.155000  75.480000 ;
        RECT 280.910000  47.235000 281.210000  47.305000 ;
        RECT 280.925000  56.705000 281.225000  56.775000 ;
        RECT 280.925000  75.480000 281.225000  75.550000 ;
        RECT 280.980000  47.305000 281.280000  47.375000 ;
        RECT 280.995000  56.635000 281.295000  56.705000 ;
        RECT 280.995000  75.550000 281.295000  75.620000 ;
        RECT 281.050000  47.375000 281.350000  47.445000 ;
        RECT 281.065000  47.445000 281.420000  47.460000 ;
        RECT 281.065000  56.565000 281.365000  56.635000 ;
        RECT 281.065000  75.620000 281.365000  75.690000 ;
        RECT 281.120000  47.460000 281.435000  47.515000 ;
        RECT 281.120000  56.510000 281.435000  56.565000 ;
        RECT 281.135000  75.690000 281.435000  75.760000 ;
        RECT 281.175000  47.515000 281.435000  47.570000 ;
        RECT 281.175000  47.570000 281.435000  56.455000 ;
        RECT 281.175000  56.455000 281.435000  56.510000 ;
        RECT 281.205000  75.760000 281.505000  75.830000 ;
        RECT 281.275000  75.830000 281.575000  75.900000 ;
        RECT 281.345000  75.900000 281.645000  75.970000 ;
        RECT 281.415000  75.970000 281.715000  76.040000 ;
        RECT 281.485000  76.040000 281.785000  76.110000 ;
        RECT 281.555000  76.110000 281.855000  76.180000 ;
        RECT 281.625000  76.180000 281.925000  76.250000 ;
        RECT 281.695000  76.250000 281.995000  76.320000 ;
        RECT 281.765000  76.320000 282.065000  76.390000 ;
        RECT 281.835000  76.390000 282.135000  76.460000 ;
        RECT 281.885000  76.460000 282.205000  76.510000 ;
        RECT 281.940000  76.510000 282.255000  76.565000 ;
        RECT 281.995000  76.565000 282.255000  76.620000 ;
        RECT 281.995000  76.620000 282.255000  87.540000 ;
        RECT 281.995000  87.540000 282.255000  87.595000 ;
        RECT 281.995000  87.595000 282.310000  87.650000 ;
        RECT 282.065000  87.650000 282.365000  87.720000 ;
        RECT 282.135000  87.720000 282.435000  87.790000 ;
        RECT 282.205000  87.790000 282.505000  87.860000 ;
        RECT 282.275000  87.860000 282.575000  87.930000 ;
        RECT 282.345000  87.930000 282.645000  88.000000 ;
        RECT 282.415000  88.000000 282.715000  88.070000 ;
        RECT 282.485000  88.070000 282.785000  88.140000 ;
        RECT 282.555000  88.140000 282.855000  88.210000 ;
        RECT 282.625000  88.210000 282.925000  88.280000 ;
        RECT 282.695000  88.280000 282.995000  88.350000 ;
        RECT 282.765000  88.350000 283.065000  88.420000 ;
        RECT 282.835000  88.420000 283.135000  88.490000 ;
        RECT 282.905000  88.490000 283.205000  88.560000 ;
        RECT 282.975000  88.560000 283.275000  88.630000 ;
        RECT 283.045000  88.630000 283.345000  88.700000 ;
        RECT 283.115000  88.700000 283.415000  88.770000 ;
        RECT 283.185000  88.770000 283.485000  88.840000 ;
        RECT 283.255000  88.840000 283.555000  88.910000 ;
        RECT 283.325000  88.910000 283.625000  88.980000 ;
        RECT 283.395000  88.980000 283.695000  89.050000 ;
        RECT 283.465000  89.050000 283.765000  89.120000 ;
        RECT 283.535000  89.120000 283.835000  89.190000 ;
        RECT 283.605000  89.190000 283.905000  89.260000 ;
        RECT 283.675000  89.260000 283.975000  89.330000 ;
        RECT 283.745000  89.330000 284.045000  89.400000 ;
        RECT 283.815000  89.400000 284.115000  89.470000 ;
        RECT 283.825000  89.470000 284.185000  89.480000 ;
        RECT 283.865000  89.480000 284.195000  89.520000 ;
        RECT 283.905000  89.520000 284.195000  89.560000 ;
        RECT 283.910000  89.560000 284.195000  89.565000 ;
        RECT 283.910000  89.565000 284.195000  94.165000 ;
        RECT 283.910000  94.165000 284.195000  94.205000 ;
        RECT 283.910000  94.205000 284.235000  94.245000 ;
        RECT 283.910000  94.245000 284.275000  94.250000 ;
        RECT 283.980000  94.250000 284.280000  94.320000 ;
        RECT 284.050000  94.320000 284.350000  94.390000 ;
        RECT 284.120000  94.390000 284.420000  94.460000 ;
        RECT 284.190000  94.460000 284.490000  94.530000 ;
        RECT 284.260000  94.530000 284.560000  94.600000 ;
        RECT 284.330000  94.600000 284.630000  94.670000 ;
        RECT 284.360000  94.670000 284.700000  94.700000 ;
        RECT 284.430000  94.700000 289.415000  94.770000 ;
        RECT 284.500000  94.770000 289.485000  94.840000 ;
        RECT 284.570000  94.840000 289.555000  94.910000 ;
        RECT 284.620000  94.910000 289.625000  94.960000 ;
        RECT 289.375000  94.960000 289.675000  95.030000 ;
        RECT 289.445000  95.030000 289.745000  95.100000 ;
        RECT 289.515000  95.100000 289.815000  95.170000 ;
        RECT 289.585000  95.170000 289.885000  95.240000 ;
        RECT 289.655000  95.240000 289.955000  95.310000 ;
        RECT 289.725000  95.310000 290.025000  95.380000 ;
        RECT 289.795000  95.380000 290.095000  95.450000 ;
        RECT 289.865000  95.450000 290.165000  95.520000 ;
        RECT 289.935000  95.520000 290.235000  95.590000 ;
        RECT 290.005000  95.590000 290.305000  95.660000 ;
        RECT 290.075000  95.660000 290.375000  95.730000 ;
        RECT 290.145000  95.730000 290.445000  95.800000 ;
        RECT 290.215000  95.800000 290.515000  95.870000 ;
        RECT 290.285000  95.870000 290.585000  95.940000 ;
        RECT 290.355000  95.940000 290.655000  96.010000 ;
        RECT 290.425000  96.010000 290.725000  96.080000 ;
        RECT 290.495000  96.080000 290.795000  96.150000 ;
        RECT 290.565000  96.150000 290.865000  96.220000 ;
        RECT 290.635000  96.220000 290.935000  96.290000 ;
        RECT 290.705000  96.290000 291.005000  96.360000 ;
        RECT 290.775000  96.360000 291.075000  96.430000 ;
        RECT 290.845000  96.430000 291.145000  96.500000 ;
        RECT 290.915000  96.500000 291.215000  96.570000 ;
        RECT 290.985000  96.570000 291.285000  96.640000 ;
        RECT 291.055000  96.640000 291.355000  96.710000 ;
        RECT 291.125000  96.710000 291.425000  96.780000 ;
        RECT 291.195000  96.780000 291.495000  96.850000 ;
        RECT 291.265000  96.850000 291.565000  96.920000 ;
        RECT 291.335000  96.920000 291.635000  96.990000 ;
        RECT 291.405000  96.990000 291.705000  97.060000 ;
        RECT 291.475000  97.060000 291.775000  97.130000 ;
        RECT 291.545000  97.130000 291.845000  97.200000 ;
        RECT 291.615000  97.200000 291.915000  97.270000 ;
        RECT 291.685000  97.270000 291.985000  97.340000 ;
        RECT 291.755000  97.340000 292.055000  97.410000 ;
        RECT 291.825000  97.410000 292.125000  97.480000 ;
        RECT 291.895000  97.480000 292.195000  97.550000 ;
        RECT 291.965000  97.550000 292.265000  97.620000 ;
        RECT 292.035000  97.620000 292.335000  97.690000 ;
        RECT 292.105000  97.690000 292.405000  97.760000 ;
        RECT 292.175000  97.760000 292.475000  97.830000 ;
        RECT 292.245000  97.830000 292.545000  97.900000 ;
        RECT 292.315000  97.900000 292.615000  97.970000 ;
        RECT 292.385000  97.970000 292.685000  98.040000 ;
        RECT 292.455000  98.040000 292.755000  98.110000 ;
        RECT 292.525000  98.110000 292.825000  98.180000 ;
        RECT 292.595000  98.180000 292.895000  98.250000 ;
        RECT 292.665000  98.250000 292.965000  98.320000 ;
        RECT 292.735000  98.320000 293.035000  98.390000 ;
        RECT 292.805000  98.390000 293.105000  98.460000 ;
        RECT 292.875000  98.460000 293.175000  98.530000 ;
        RECT 292.945000  98.530000 293.245000  98.600000 ;
        RECT 293.015000  98.600000 293.315000  98.670000 ;
        RECT 293.085000  98.670000 293.385000  98.740000 ;
        RECT 293.155000  98.740000 293.455000  98.810000 ;
        RECT 293.225000  98.810000 293.525000  98.880000 ;
        RECT 293.295000  98.880000 293.595000  98.950000 ;
        RECT 293.365000  98.950000 293.665000  99.020000 ;
        RECT 293.435000  99.020000 293.735000  99.090000 ;
        RECT 293.505000  99.090000 293.805000  99.160000 ;
        RECT 293.575000  99.160000 293.875000  99.230000 ;
        RECT 293.645000  99.230000 293.945000  99.300000 ;
        RECT 293.715000  99.300000 294.015000  99.370000 ;
        RECT 293.785000  99.370000 294.085000  99.440000 ;
        RECT 293.855000  99.440000 294.155000  99.510000 ;
        RECT 293.925000  99.510000 294.225000  99.580000 ;
        RECT 293.995000  99.580000 294.295000  99.650000 ;
        RECT 294.065000  99.650000 294.365000  99.720000 ;
        RECT 294.135000  99.720000 294.435000  99.790000 ;
        RECT 294.205000  99.790000 294.505000  99.860000 ;
        RECT 294.275000  99.860000 294.575000  99.930000 ;
        RECT 294.345000  99.930000 294.645000 100.000000 ;
        RECT 294.415000 100.000000 294.715000 100.070000 ;
        RECT 294.485000 100.070000 294.785000 100.140000 ;
        RECT 294.555000 100.140000 294.855000 100.210000 ;
        RECT 294.625000 100.210000 294.925000 100.280000 ;
        RECT 294.695000 100.280000 294.995000 100.350000 ;
        RECT 294.765000 100.350000 295.065000 100.420000 ;
        RECT 294.835000 100.420000 295.135000 100.490000 ;
        RECT 294.905000 100.490000 295.205000 100.560000 ;
        RECT 294.975000 100.560000 295.275000 100.630000 ;
        RECT 295.045000 100.630000 295.345000 100.700000 ;
        RECT 295.115000 100.700000 295.415000 100.770000 ;
        RECT 295.185000 100.770000 295.485000 100.840000 ;
        RECT 295.255000 100.840000 295.555000 100.910000 ;
        RECT 295.325000 100.910000 295.625000 100.980000 ;
        RECT 295.395000 100.980000 295.695000 101.050000 ;
        RECT 295.465000 101.050000 295.765000 101.120000 ;
        RECT 295.535000 101.120000 295.835000 101.190000 ;
        RECT 295.605000 101.190000 295.905000 101.260000 ;
        RECT 295.675000 101.260000 295.975000 101.330000 ;
        RECT 295.745000 101.330000 296.045000 101.400000 ;
        RECT 295.815000 101.400000 296.115000 101.470000 ;
        RECT 295.885000 101.470000 296.185000 101.540000 ;
        RECT 295.955000 101.540000 296.255000 101.610000 ;
        RECT 296.025000 101.610000 296.325000 101.680000 ;
        RECT 296.095000 101.680000 296.395000 101.750000 ;
        RECT 296.165000 101.750000 296.465000 101.820000 ;
        RECT 296.235000 101.820000 296.535000 101.890000 ;
        RECT 296.305000 101.890000 296.605000 101.960000 ;
        RECT 296.375000 101.960000 296.675000 102.030000 ;
        RECT 296.445000 102.030000 296.745000 102.100000 ;
        RECT 296.515000 102.100000 296.815000 102.170000 ;
        RECT 296.585000 102.170000 296.885000 102.240000 ;
        RECT 296.655000 102.240000 296.955000 102.310000 ;
        RECT 296.660000 111.500000 297.700000 111.600000 ;
        RECT 296.660000 111.600000 297.630000 111.670000 ;
        RECT 296.660000 111.670000 297.560000 111.740000 ;
        RECT 296.660000 111.740000 297.540000 111.760000 ;
        RECT 296.660000 111.760000 296.990000 111.830000 ;
        RECT 296.660000 111.830000 296.920000 111.900000 ;
        RECT 296.660000 111.900000 296.920000 112.140000 ;
        RECT 296.725000 102.310000 297.025000 102.380000 ;
        RECT 296.795000 102.380000 297.095000 102.450000 ;
        RECT 296.865000 102.450000 297.165000 102.520000 ;
        RECT 296.935000 102.520000 297.235000 102.590000 ;
        RECT 297.005000 102.590000 297.305000 102.660000 ;
        RECT 297.075000 102.660000 297.375000 102.730000 ;
        RECT 297.145000 102.730000 297.445000 102.800000 ;
        RECT 297.215000 102.800000 297.515000 102.870000 ;
        RECT 297.285000 102.870000 297.585000 102.940000 ;
        RECT 297.290000 111.495000 297.700000 111.500000 ;
        RECT 297.330000 102.940000 297.655000 102.985000 ;
        RECT 297.350000 111.435000 297.700000 111.495000 ;
        RECT 297.370000 102.985000 297.700000 103.025000 ;
        RECT 297.410000 103.025000 297.700000 103.065000 ;
        RECT 297.410000 103.065000 297.700000 111.375000 ;
        RECT 297.410000 111.375000 297.700000 111.435000 ;
    END
  END TIE_LO_ESD[1]
  PIN VINREF_DFT
    ANTENNAPARTIALMETALSIDEAREA  42.13650 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.030000 0.000000 466.670000 60.295000 ;
    END
  END VINREF_DFT
  PIN VOHREF
    ANTENNAPARTIALMETALSIDEAREA  58.06500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.445000 0.000000 419.705000 5.035000 ;
    END
  END VOHREF
  PIN VOH_SEL[0]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.920000 244.355000 447.560000 244.615000 ;
        RECT 446.945000 244.330000 447.505000 244.355000 ;
        RECT 447.015000 244.260000 447.435000 244.330000 ;
        RECT 447.085000  85.835000 447.400000  85.890000 ;
        RECT 447.085000  85.890000 447.345000  85.945000 ;
        RECT 447.085000  85.945000 447.345000 244.170000 ;
        RECT 447.085000 244.170000 447.345000 244.180000 ;
        RECT 447.085000 244.180000 447.355000 244.190000 ;
        RECT 447.085000 244.190000 447.365000 244.260000 ;
        RECT 447.125000  85.795000 447.455000  85.835000 ;
        RECT 447.195000  85.725000 447.495000  85.795000 ;
        RECT 447.265000  85.655000 447.565000  85.725000 ;
        RECT 447.335000  85.585000 447.635000  85.655000 ;
        RECT 447.405000  85.515000 447.705000  85.585000 ;
        RECT 447.475000  85.445000 447.775000  85.515000 ;
        RECT 447.545000  85.375000 447.845000  85.445000 ;
        RECT 447.615000  85.305000 447.915000  85.375000 ;
        RECT 447.685000  85.235000 447.985000  85.305000 ;
        RECT 447.755000  85.165000 448.055000  85.235000 ;
        RECT 447.825000  85.095000 448.125000  85.165000 ;
        RECT 447.895000  85.025000 448.195000  85.095000 ;
        RECT 447.965000  84.955000 448.265000  85.025000 ;
        RECT 448.035000  84.885000 448.335000  84.955000 ;
        RECT 448.105000  84.815000 448.405000  84.885000 ;
        RECT 448.175000  84.745000 448.475000  84.815000 ;
        RECT 448.245000  84.675000 448.545000  84.745000 ;
        RECT 448.315000  84.605000 448.615000  84.675000 ;
        RECT 448.385000  84.535000 448.685000  84.605000 ;
        RECT 448.455000  84.465000 448.755000  84.535000 ;
        RECT 448.525000  84.395000 448.825000  84.465000 ;
        RECT 448.595000  84.325000 448.895000  84.395000 ;
        RECT 448.665000  84.255000 448.965000  84.325000 ;
        RECT 448.735000  84.185000 449.035000  84.255000 ;
        RECT 448.805000  84.115000 449.105000  84.185000 ;
        RECT 448.875000  84.045000 449.175000  84.115000 ;
        RECT 448.945000  83.975000 449.245000  84.045000 ;
        RECT 449.015000  83.905000 449.315000  83.975000 ;
        RECT 449.085000  83.835000 449.385000  83.905000 ;
        RECT 449.155000  83.765000 449.455000  83.835000 ;
        RECT 449.225000  83.695000 449.525000  83.765000 ;
        RECT 449.295000  83.625000 449.595000  83.695000 ;
        RECT 449.350000  83.570000 449.665000  83.625000 ;
        RECT 449.405000   0.000000 449.665000  83.515000 ;
        RECT 449.405000  83.515000 449.665000  83.570000 ;
    END
  END VOH_SEL[0]
  PIN VOH_SEL[1]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.745000 238.310000 448.060000 238.365000 ;
        RECT 447.745000 238.365000 448.005000 238.420000 ;
        RECT 447.745000 238.420000 448.005000 245.015000 ;
        RECT 447.805000 238.250000 448.115000 238.310000 ;
        RECT 447.875000 238.180000 448.175000 238.250000 ;
        RECT 447.945000 238.110000 448.245000 238.180000 ;
        RECT 448.015000 238.040000 448.315000 238.110000 ;
        RECT 448.085000 237.970000 448.385000 238.040000 ;
        RECT 448.155000 237.900000 448.455000 237.970000 ;
        RECT 448.225000 237.830000 448.525000 237.900000 ;
        RECT 448.295000 237.760000 448.595000 237.830000 ;
        RECT 448.365000 237.690000 448.665000 237.760000 ;
        RECT 448.435000 237.620000 448.735000 237.690000 ;
        RECT 448.505000 237.550000 448.805000 237.620000 ;
        RECT 448.575000 237.480000 448.875000 237.550000 ;
        RECT 448.645000 237.410000 448.945000 237.480000 ;
        RECT 448.715000 237.340000 449.015000 237.410000 ;
        RECT 448.785000 237.270000 449.085000 237.340000 ;
        RECT 448.855000 237.200000 449.155000 237.270000 ;
        RECT 448.925000 237.130000 449.225000 237.200000 ;
        RECT 448.995000 237.060000 449.295000 237.130000 ;
        RECT 449.065000 236.990000 449.365000 237.060000 ;
        RECT 449.135000 236.920000 449.435000 236.990000 ;
        RECT 449.205000 236.850000 449.505000 236.920000 ;
        RECT 449.275000 236.780000 449.575000 236.850000 ;
        RECT 449.345000 236.710000 449.645000 236.780000 ;
        RECT 449.415000 236.640000 449.715000 236.710000 ;
        RECT 449.485000 236.570000 449.785000 236.640000 ;
        RECT 449.555000 236.500000 449.855000 236.570000 ;
        RECT 449.625000 236.430000 449.925000 236.500000 ;
        RECT 449.695000 236.360000 449.995000 236.430000 ;
        RECT 449.765000 236.290000 450.065000 236.360000 ;
        RECT 449.835000 236.220000 450.135000 236.290000 ;
        RECT 449.905000 236.150000 450.205000 236.220000 ;
        RECT 449.975000 236.080000 450.275000 236.150000 ;
        RECT 450.045000 236.010000 450.345000 236.080000 ;
        RECT 450.100000 235.955000 450.415000 236.010000 ;
        RECT 450.155000   0.000000 450.415000 235.900000 ;
        RECT 450.155000 235.900000 450.415000 235.955000 ;
    END
  END VOH_SEL[1]
  PIN VOH_SEL[2]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.495000 238.630000 448.810000 238.685000 ;
        RECT 448.495000 238.685000 448.755000 238.740000 ;
        RECT 448.495000 238.740000 448.755000 245.415000 ;
        RECT 448.555000 238.570000 448.865000 238.630000 ;
        RECT 448.625000 238.500000 448.925000 238.570000 ;
        RECT 448.695000 238.430000 448.995000 238.500000 ;
        RECT 448.765000 238.360000 449.065000 238.430000 ;
        RECT 448.835000 238.290000 449.135000 238.360000 ;
        RECT 448.905000 238.220000 449.205000 238.290000 ;
        RECT 448.975000 238.150000 449.275000 238.220000 ;
        RECT 449.045000 238.080000 449.345000 238.150000 ;
        RECT 449.115000 238.010000 449.415000 238.080000 ;
        RECT 449.185000 237.940000 449.485000 238.010000 ;
        RECT 449.255000 237.870000 449.555000 237.940000 ;
        RECT 449.325000 237.800000 449.625000 237.870000 ;
        RECT 449.395000 237.730000 449.695000 237.800000 ;
        RECT 449.465000 237.660000 449.765000 237.730000 ;
        RECT 449.535000 237.590000 449.835000 237.660000 ;
        RECT 449.605000 237.520000 449.905000 237.590000 ;
        RECT 449.675000 237.450000 449.975000 237.520000 ;
        RECT 449.745000 237.380000 450.045000 237.450000 ;
        RECT 449.815000 237.310000 450.115000 237.380000 ;
        RECT 449.885000 237.240000 450.185000 237.310000 ;
        RECT 449.955000 237.170000 450.255000 237.240000 ;
        RECT 450.025000 237.100000 450.325000 237.170000 ;
        RECT 450.095000 237.030000 450.395000 237.100000 ;
        RECT 450.165000 236.960000 450.465000 237.030000 ;
        RECT 450.235000 236.890000 450.535000 236.960000 ;
        RECT 450.305000 236.820000 450.605000 236.890000 ;
        RECT 450.375000 236.750000 450.675000 236.820000 ;
        RECT 450.445000 236.680000 450.745000 236.750000 ;
        RECT 450.515000 236.610000 450.815000 236.680000 ;
        RECT 450.585000 236.540000 450.885000 236.610000 ;
        RECT 450.655000 236.470000 450.955000 236.540000 ;
        RECT 450.725000 236.400000 451.025000 236.470000 ;
        RECT 450.795000 236.330000 451.095000 236.400000 ;
        RECT 450.850000 236.275000 451.165000 236.330000 ;
        RECT 450.905000   0.000000 451.165000 236.220000 ;
        RECT 450.905000 236.220000 451.165000 236.275000 ;
    END
  END VOH_SEL[2]
  PIN VOUTREF_DFT
    ANTENNAPARTIALMETALSIDEAREA  42.13650 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.530000 0.000000 465.170000 60.295000 ;
    END
  END VOUTREF_DFT
  PIN VREF_SEL[0]
    ANTENNAGATEAREA  0.999000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.745000 239.590000 451.060000 239.645000 ;
        RECT 450.745000 239.645000 451.005000 239.700000 ;
        RECT 450.745000 239.700000 451.005000 241.785000 ;
        RECT 450.805000 239.530000 451.115000 239.590000 ;
        RECT 450.875000 239.460000 451.175000 239.530000 ;
        RECT 450.945000 239.390000 451.245000 239.460000 ;
        RECT 451.015000 239.320000 451.315000 239.390000 ;
        RECT 451.085000 239.250000 451.385000 239.320000 ;
        RECT 451.155000 239.180000 451.455000 239.250000 ;
        RECT 451.225000 239.110000 451.525000 239.180000 ;
        RECT 451.295000 239.040000 451.595000 239.110000 ;
        RECT 451.365000 238.970000 451.665000 239.040000 ;
        RECT 451.435000 238.900000 451.735000 238.970000 ;
        RECT 451.505000 238.830000 451.805000 238.900000 ;
        RECT 451.575000 238.760000 451.875000 238.830000 ;
        RECT 451.645000 238.690000 451.945000 238.760000 ;
        RECT 451.715000 238.620000 452.015000 238.690000 ;
        RECT 451.785000 238.550000 452.085000 238.620000 ;
        RECT 451.855000 238.480000 452.155000 238.550000 ;
        RECT 451.925000 238.410000 452.225000 238.480000 ;
        RECT 451.995000 238.340000 452.295000 238.410000 ;
        RECT 452.065000 238.270000 452.365000 238.340000 ;
        RECT 452.135000 238.200000 452.435000 238.270000 ;
        RECT 452.205000 238.130000 452.505000 238.200000 ;
        RECT 452.275000 238.060000 452.575000 238.130000 ;
        RECT 452.345000 237.990000 452.645000 238.060000 ;
        RECT 452.415000 237.920000 452.715000 237.990000 ;
        RECT 452.485000 237.850000 452.785000 237.920000 ;
        RECT 452.555000 237.780000 452.855000 237.850000 ;
        RECT 452.625000 237.710000 452.925000 237.780000 ;
        RECT 452.695000 237.640000 452.995000 237.710000 ;
        RECT 452.765000 237.570000 453.065000 237.640000 ;
        RECT 452.835000 237.500000 453.135000 237.570000 ;
        RECT 452.905000 237.430000 453.205000 237.500000 ;
        RECT 452.975000 237.360000 453.275000 237.430000 ;
        RECT 453.045000 237.290000 453.345000 237.360000 ;
        RECT 453.100000 237.235000 453.415000 237.290000 ;
        RECT 453.155000   0.000000 453.415000 237.180000 ;
        RECT 453.155000 237.180000 453.415000 237.235000 ;
    END
  END VREF_SEL[0]
  PIN VREF_SEL[1]
    ANTENNAGATEAREA  0.999000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.115000 241.965000 451.755000 242.225000 ;
        RECT 451.355000 241.900000 451.755000 241.965000 ;
        RECT 451.425000 241.830000 451.755000 241.900000 ;
        RECT 451.495000 239.910000 451.810000 239.965000 ;
        RECT 451.495000 239.965000 451.755000 240.020000 ;
        RECT 451.495000 240.020000 451.755000 241.760000 ;
        RECT 451.495000 241.760000 451.755000 241.830000 ;
        RECT 451.555000 239.850000 451.865000 239.910000 ;
        RECT 451.625000 239.780000 451.925000 239.850000 ;
        RECT 451.695000 239.710000 451.995000 239.780000 ;
        RECT 451.765000 239.640000 452.065000 239.710000 ;
        RECT 451.835000 239.570000 452.135000 239.640000 ;
        RECT 451.905000 239.500000 452.205000 239.570000 ;
        RECT 451.975000 239.430000 452.275000 239.500000 ;
        RECT 452.045000 239.360000 452.345000 239.430000 ;
        RECT 452.115000 239.290000 452.415000 239.360000 ;
        RECT 452.185000 239.220000 452.485000 239.290000 ;
        RECT 452.255000 239.150000 452.555000 239.220000 ;
        RECT 452.325000 239.080000 452.625000 239.150000 ;
        RECT 452.395000 239.010000 452.695000 239.080000 ;
        RECT 452.465000 238.940000 452.765000 239.010000 ;
        RECT 452.535000 238.870000 452.835000 238.940000 ;
        RECT 452.605000 238.800000 452.905000 238.870000 ;
        RECT 452.675000 238.730000 452.975000 238.800000 ;
        RECT 452.745000 238.660000 453.045000 238.730000 ;
        RECT 452.815000 238.590000 453.115000 238.660000 ;
        RECT 452.885000 238.520000 453.185000 238.590000 ;
        RECT 452.955000 238.450000 453.255000 238.520000 ;
        RECT 453.025000 238.380000 453.325000 238.450000 ;
        RECT 453.095000 238.310000 453.395000 238.380000 ;
        RECT 453.165000 238.240000 453.465000 238.310000 ;
        RECT 453.235000 238.170000 453.535000 238.240000 ;
        RECT 453.305000 238.100000 453.605000 238.170000 ;
        RECT 453.375000 238.030000 453.675000 238.100000 ;
        RECT 453.445000 237.960000 453.745000 238.030000 ;
        RECT 453.515000 237.890000 453.815000 237.960000 ;
        RECT 453.585000 237.820000 453.885000 237.890000 ;
        RECT 453.655000 237.750000 453.955000 237.820000 ;
        RECT 453.725000 237.680000 454.025000 237.750000 ;
        RECT 453.795000 237.610000 454.095000 237.680000 ;
        RECT 453.850000 237.555000 454.165000 237.610000 ;
        RECT 453.905000   0.000000 454.165000 237.500000 ;
        RECT 453.905000 237.500000 454.165000 237.555000 ;
    END
  END VREF_SEL[1]
  PIN VREG_EN[0]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.805000  0.000000 150.065000 27.875000 ;
        RECT 149.805000 27.875000 150.065000 27.945000 ;
        RECT 149.805000 27.945000 150.135000 28.015000 ;
        RECT 149.805000 28.015000 150.205000 28.085000 ;
        RECT 149.805000 28.085000 150.275000 28.155000 ;
        RECT 149.805000 28.155000 150.345000 28.225000 ;
        RECT 149.805000 28.225000 150.415000 28.250000 ;
        RECT 149.805000 31.265000 150.370000 31.335000 ;
        RECT 149.805000 31.335000 150.300000 31.405000 ;
        RECT 149.805000 31.405000 150.230000 31.475000 ;
        RECT 149.805000 31.475000 150.160000 31.545000 ;
        RECT 149.805000 31.545000 150.090000 31.615000 ;
        RECT 149.805000 31.615000 150.065000 31.640000 ;
        RECT 149.805000 31.640000 150.065000 58.140000 ;
        RECT 149.805000 58.140000 150.065000 58.200000 ;
        RECT 149.805000 58.200000 150.125000 58.260000 ;
        RECT 149.805000 58.260000 150.185000 58.265000 ;
        RECT 149.805000 58.265000 150.445000 58.525000 ;
        RECT 149.830000 31.240000 150.440000 31.265000 ;
        RECT 149.875000 28.250000 150.440000 28.320000 ;
        RECT 149.900000 31.170000 150.465000 31.240000 ;
        RECT 149.945000 28.320000 150.510000 28.390000 ;
        RECT 149.970000 28.390000 150.580000 28.415000 ;
        RECT 149.970000 31.100000 150.535000 31.170000 ;
        RECT 149.995000 31.075000 150.605000 31.100000 ;
        RECT 150.040000 28.415000 150.605000 28.485000 ;
        RECT 150.065000 31.005000 150.605000 31.075000 ;
        RECT 150.110000 28.485000 150.605000 28.555000 ;
        RECT 150.135000 30.935000 150.605000 31.005000 ;
        RECT 150.180000 28.555000 150.605000 28.625000 ;
        RECT 150.205000 30.865000 150.605000 30.935000 ;
        RECT 150.250000 28.625000 150.605000 28.695000 ;
        RECT 150.275000 30.795000 150.605000 30.865000 ;
        RECT 150.320000 28.695000 150.605000 28.765000 ;
        RECT 150.345000 28.765000 150.605000 28.790000 ;
        RECT 150.345000 28.790000 150.605000 30.725000 ;
        RECT 150.345000 30.725000 150.605000 30.795000 ;
    END
  END VREG_EN[0]
  PIN VREG_EN[1]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.400000 28.415000 239.965000 28.485000 ;
        RECT 239.400000 28.485000 239.895000 28.555000 ;
        RECT 239.400000 28.555000 239.825000 28.625000 ;
        RECT 239.400000 28.625000 239.755000 28.695000 ;
        RECT 239.400000 28.695000 239.685000 28.765000 ;
        RECT 239.400000 28.765000 239.660000 28.790000 ;
        RECT 239.400000 28.790000 239.660000 30.725000 ;
        RECT 239.400000 30.725000 239.660000 30.795000 ;
        RECT 239.400000 30.795000 239.730000 30.865000 ;
        RECT 239.400000 30.865000 239.800000 30.935000 ;
        RECT 239.400000 30.935000 239.870000 31.005000 ;
        RECT 239.400000 31.005000 239.940000 31.075000 ;
        RECT 239.400000 31.075000 240.010000 31.100000 ;
        RECT 239.425000 28.390000 240.035000 28.415000 ;
        RECT 239.470000 31.100000 240.035000 31.170000 ;
        RECT 239.495000 28.320000 240.060000 28.390000 ;
        RECT 239.540000 31.170000 240.105000 31.240000 ;
        RECT 239.560000 58.265000 240.200000 58.525000 ;
        RECT 239.565000 28.250000 240.130000 28.320000 ;
        RECT 239.565000 31.240000 240.175000 31.265000 ;
        RECT 239.590000 28.225000 240.200000 28.250000 ;
        RECT 239.635000 31.265000 240.200000 31.335000 ;
        RECT 239.660000 28.155000 240.200000 28.225000 ;
        RECT 239.705000 31.335000 240.200000 31.405000 ;
        RECT 239.730000 28.085000 240.200000 28.155000 ;
        RECT 239.775000 31.405000 240.200000 31.475000 ;
        RECT 239.800000 28.015000 240.200000 28.085000 ;
        RECT 239.820000 58.260000 240.200000 58.265000 ;
        RECT 239.845000 31.475000 240.200000 31.545000 ;
        RECT 239.870000 27.945000 240.200000 28.015000 ;
        RECT 239.880000 58.200000 240.200000 58.260000 ;
        RECT 239.915000 31.545000 240.200000 31.615000 ;
        RECT 239.940000  0.000000 240.200000 27.875000 ;
        RECT 239.940000 27.875000 240.200000 27.945000 ;
        RECT 239.940000 31.615000 240.200000 31.640000 ;
        RECT 239.940000 31.640000 240.200000 58.140000 ;
        RECT 239.940000 58.140000 240.200000 58.200000 ;
    END
  END VREG_EN[1]
  PIN VREG_EN_REFGEN
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.840000  0.000000 445.100000 22.305000 ;
        RECT 444.840000 22.305000 445.100000 22.340000 ;
        RECT 444.840000 22.340000 445.135000 22.375000 ;
        RECT 444.840000 22.375000 445.170000 23.015000 ;
    END
  END VREG_EN_REFGEN
  PIN VTRIP_SEL[0]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.260000 10.930000 127.575000 10.985000 ;
        RECT 127.260000 10.985000 127.520000 11.040000 ;
        RECT 127.260000 11.040000 127.520000 23.665000 ;
        RECT 127.260000 23.665000 127.520000 23.720000 ;
        RECT 127.260000 23.720000 127.575000 23.775000 ;
        RECT 127.315000 10.875000 127.630000 10.930000 ;
        RECT 127.330000 23.775000 127.630000 23.845000 ;
        RECT 127.385000 10.805000 127.685000 10.875000 ;
        RECT 127.400000 23.845000 127.700000 23.915000 ;
        RECT 127.455000 10.735000 127.755000 10.805000 ;
        RECT 127.470000 23.915000 127.770000 23.985000 ;
        RECT 127.525000 10.665000 127.825000 10.735000 ;
        RECT 127.540000 23.985000 127.840000 24.055000 ;
        RECT 127.595000 10.595000 127.895000 10.665000 ;
        RECT 127.610000 24.055000 127.910000 24.125000 ;
        RECT 127.665000 10.525000 127.965000 10.595000 ;
        RECT 127.680000 24.125000 127.980000 24.195000 ;
        RECT 127.735000 10.455000 128.035000 10.525000 ;
        RECT 127.750000 24.195000 128.050000 24.265000 ;
        RECT 127.805000 10.385000 128.105000 10.455000 ;
        RECT 127.805000 24.265000 128.120000 24.320000 ;
        RECT 127.860000 24.320000 128.120000 24.375000 ;
        RECT 127.860000 24.375000 128.120000 42.525000 ;
        RECT 127.860000 42.525000 128.120000 42.585000 ;
        RECT 127.860000 42.585000 128.180000 42.645000 ;
        RECT 127.860000 42.645000 128.240000 42.650000 ;
        RECT 127.860000 42.650000 128.880000 42.910000 ;
        RECT 127.875000 10.315000 128.175000 10.385000 ;
        RECT 127.945000 10.245000 128.245000 10.315000 ;
        RECT 128.015000 10.175000 128.315000 10.245000 ;
        RECT 128.070000 10.120000 128.385000 10.175000 ;
        RECT 128.125000  0.000000 128.385000 10.065000 ;
        RECT 128.125000 10.065000 128.385000 10.120000 ;
    END
  END VTRIP_SEL[0]
  PIN VTRIP_SEL[1]
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.125000 42.650000 262.145000 42.910000 ;
        RECT 261.620000  0.000000 261.880000 10.065000 ;
        RECT 261.620000 10.065000 261.880000 10.120000 ;
        RECT 261.620000 10.120000 261.935000 10.175000 ;
        RECT 261.690000 10.175000 261.990000 10.245000 ;
        RECT 261.760000 10.245000 262.060000 10.315000 ;
        RECT 261.765000 42.645000 262.145000 42.650000 ;
        RECT 261.825000 42.585000 262.145000 42.645000 ;
        RECT 261.830000 10.315000 262.130000 10.385000 ;
        RECT 261.885000 24.265000 262.200000 24.320000 ;
        RECT 261.885000 24.320000 262.145000 24.375000 ;
        RECT 261.885000 24.375000 262.145000 42.525000 ;
        RECT 261.885000 42.525000 262.145000 42.585000 ;
        RECT 261.900000 10.385000 262.200000 10.455000 ;
        RECT 261.955000 24.195000 262.255000 24.265000 ;
        RECT 261.970000 10.455000 262.270000 10.525000 ;
        RECT 262.025000 24.125000 262.325000 24.195000 ;
        RECT 262.040000 10.525000 262.340000 10.595000 ;
        RECT 262.095000 24.055000 262.395000 24.125000 ;
        RECT 262.110000 10.595000 262.410000 10.665000 ;
        RECT 262.165000 23.985000 262.465000 24.055000 ;
        RECT 262.180000 10.665000 262.480000 10.735000 ;
        RECT 262.235000 23.915000 262.535000 23.985000 ;
        RECT 262.250000 10.735000 262.550000 10.805000 ;
        RECT 262.305000 23.845000 262.605000 23.915000 ;
        RECT 262.320000 10.805000 262.620000 10.875000 ;
        RECT 262.375000 10.875000 262.690000 10.930000 ;
        RECT 262.375000 23.775000 262.675000 23.845000 ;
        RECT 262.430000 10.930000 262.745000 10.985000 ;
        RECT 262.430000 23.720000 262.745000 23.775000 ;
        RECT 262.485000 10.985000 262.745000 11.040000 ;
        RECT 262.485000 11.040000 262.745000 23.665000 ;
        RECT 262.485000 23.665000 262.745000 23.720000 ;
    END
  END VTRIP_SEL[1]
  PIN VTRIP_SEL_REFGEN
    ANTENNAGATEAREA  0.720000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.840000 0.000000 403.100000 23.140000 ;
    END
  END VTRIP_SEL_REFGEN
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 62.600000 480.000000 67.250000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 62.700000 480.000000 67.150000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 55.750000 480.000000 61.200000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 55.850000 480.000000 61.100000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 68.650000 480.000000 72.100000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 68.750000 480.000000 72.000000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT   0.000000 123.750000  28.815000 123.800000 ;
        RECT   0.000000 123.800000  28.865000 123.850000 ;
        RECT   0.000000 123.850000  28.930000 123.865000 ;
        RECT   0.000000 123.865000  28.930000 124.015000 ;
        RECT   0.000000 124.015000  29.080000 124.165000 ;
        RECT   0.000000 124.165000  29.230000 124.315000 ;
        RECT   0.000000 124.315000  29.380000 124.465000 ;
        RECT   0.000000 124.465000  29.530000 124.615000 ;
        RECT   0.000000 124.615000  29.680000 124.765000 ;
        RECT   0.000000 124.765000  29.830000 124.915000 ;
        RECT   0.000000 124.915000  29.980000 125.065000 ;
        RECT   0.000000 125.065000  30.130000 125.215000 ;
        RECT   0.000000 125.215000  30.280000 125.365000 ;
        RECT   0.000000 125.365000  30.430000 125.515000 ;
        RECT   0.000000 125.515000  30.580000 125.665000 ;
        RECT   0.000000 125.665000  30.730000 125.815000 ;
        RECT   0.000000 125.815000  30.880000 125.965000 ;
        RECT   0.000000 125.965000  31.030000 126.115000 ;
        RECT   0.000000 126.115000  31.180000 126.265000 ;
        RECT   0.000000 126.265000  31.330000 126.415000 ;
        RECT   0.000000 126.415000  31.480000 126.565000 ;
        RECT   0.000000 126.565000  31.630000 126.715000 ;
        RECT   0.000000 126.715000  31.780000 126.865000 ;
        RECT   0.000000 126.865000  31.930000 127.015000 ;
        RECT   0.000000 127.015000  32.080000 127.165000 ;
        RECT   0.000000 127.165000  32.230000 127.315000 ;
        RECT   0.000000 127.315000  32.380000 127.465000 ;
        RECT   0.000000 127.465000  32.530000 127.615000 ;
        RECT   0.000000 127.615000  32.680000 127.765000 ;
        RECT   0.000000 127.765000  32.830000 127.915000 ;
        RECT   0.000000 127.915000  32.980000 128.065000 ;
        RECT   0.000000 128.065000  33.130000 128.215000 ;
        RECT   0.000000 128.215000  33.280000 128.365000 ;
        RECT   0.000000 128.365000  33.430000 128.515000 ;
        RECT   0.000000 128.515000  33.580000 128.665000 ;
        RECT   0.000000 128.665000  33.730000 128.815000 ;
        RECT   0.000000 128.815000  33.880000 128.965000 ;
        RECT   0.000000 128.965000  34.030000 129.115000 ;
        RECT   0.000000 129.115000  34.180000 129.265000 ;
        RECT   0.000000 129.265000  34.330000 129.415000 ;
        RECT   0.000000 129.415000  34.480000 129.565000 ;
        RECT   0.000000 129.565000  34.630000 129.715000 ;
        RECT   0.000000 129.715000  34.780000 129.865000 ;
        RECT   0.000000 129.865000  34.930000 130.015000 ;
        RECT   0.000000 130.015000  35.080000 130.165000 ;
        RECT   0.000000 130.165000  35.230000 130.315000 ;
        RECT   0.000000 130.315000  35.380000 130.465000 ;
        RECT   0.000000 130.465000  35.530000 130.615000 ;
        RECT   0.000000 130.615000  35.680000 130.765000 ;
        RECT   0.000000 130.765000  35.830000 130.915000 ;
        RECT   0.000000 130.915000  35.980000 131.065000 ;
        RECT   0.000000 131.065000  36.130000 131.215000 ;
        RECT   0.000000 131.215000  36.280000 131.365000 ;
        RECT   0.000000 131.365000  36.430000 131.515000 ;
        RECT   0.000000 131.515000  36.580000 131.665000 ;
        RECT   0.000000 131.665000  36.730000 131.815000 ;
        RECT   0.000000 131.815000  36.880000 131.965000 ;
        RECT   0.000000 131.965000  37.030000 132.115000 ;
        RECT   0.000000 132.115000  37.180000 132.265000 ;
        RECT   0.000000 132.265000  37.330000 132.415000 ;
        RECT   0.000000 132.415000  37.480000 132.565000 ;
        RECT   0.000000 132.565000  37.630000 132.715000 ;
        RECT   0.000000 132.715000  37.780000 132.865000 ;
        RECT   0.000000 132.865000  37.930000 133.015000 ;
        RECT   0.000000 133.015000  38.080000 133.165000 ;
        RECT   0.000000 133.165000  38.230000 133.315000 ;
        RECT   0.000000 133.315000  38.380000 133.465000 ;
        RECT   0.000000 133.465000  38.530000 133.615000 ;
        RECT   0.000000 133.615000  38.680000 133.765000 ;
        RECT   0.000000 133.765000  38.830000 133.915000 ;
        RECT   0.000000 133.915000  38.980000 134.065000 ;
        RECT   0.000000 134.065000  39.130000 134.215000 ;
        RECT   0.000000 134.215000  39.280000 134.365000 ;
        RECT   0.000000 134.365000  39.430000 134.515000 ;
        RECT   0.000000 134.515000  39.580000 134.665000 ;
        RECT   0.000000 134.665000  39.730000 134.815000 ;
        RECT   0.000000 134.815000  39.880000 134.965000 ;
        RECT   0.000000 134.965000  40.030000 135.115000 ;
        RECT   0.000000 135.115000  40.180000 135.265000 ;
        RECT   0.000000 135.265000  40.330000 135.415000 ;
        RECT   0.000000 135.415000  40.480000 135.565000 ;
        RECT   0.000000 135.565000  40.630000 135.715000 ;
        RECT   0.000000 135.715000  40.780000 135.865000 ;
        RECT   0.000000 135.865000  40.930000 136.015000 ;
        RECT   0.000000 136.015000  41.080000 136.165000 ;
        RECT   0.000000 136.165000  41.230000 136.315000 ;
        RECT   0.000000 136.315000  41.380000 136.465000 ;
        RECT   0.000000 136.465000  41.530000 136.615000 ;
        RECT   0.000000 136.615000  41.680000 136.765000 ;
        RECT   0.000000 136.765000  41.830000 136.915000 ;
        RECT   0.000000 136.915000  41.980000 137.065000 ;
        RECT   0.000000 137.065000  42.130000 137.215000 ;
        RECT   0.000000 137.215000  42.280000 137.365000 ;
        RECT   0.000000 137.365000  42.430000 137.515000 ;
        RECT   0.000000 137.515000  42.580000 137.665000 ;
        RECT   0.000000 137.665000  42.730000 137.815000 ;
        RECT   0.000000 137.815000  42.880000 137.965000 ;
        RECT   0.000000 137.965000  43.030000 138.115000 ;
        RECT   0.000000 138.115000  43.180000 138.265000 ;
        RECT   0.000000 138.265000  43.330000 138.415000 ;
        RECT   0.000000 138.415000  43.480000 138.565000 ;
        RECT   0.000000 138.565000  43.630000 138.715000 ;
        RECT   0.000000 138.715000  43.780000 138.865000 ;
        RECT   0.000000 138.865000  43.930000 139.015000 ;
        RECT   0.000000 139.015000  44.080000 139.165000 ;
        RECT   0.000000 139.165000  44.230000 139.315000 ;
        RECT   0.000000 139.315000  44.380000 139.465000 ;
        RECT   0.000000 139.465000  44.530000 139.615000 ;
        RECT   0.000000 139.615000  44.680000 139.765000 ;
        RECT   0.000000 139.765000  44.830000 139.915000 ;
        RECT   0.000000 139.915000  44.980000 140.065000 ;
        RECT   0.000000 140.065000  45.130000 140.215000 ;
        RECT   0.000000 140.215000  45.280000 140.365000 ;
        RECT   0.000000 140.365000  45.430000 140.515000 ;
        RECT   0.000000 140.515000  45.580000 140.665000 ;
        RECT   0.000000 140.665000  45.730000 140.815000 ;
        RECT   0.000000 140.815000  45.880000 140.965000 ;
        RECT   0.000000 140.965000  46.030000 141.115000 ;
        RECT   0.000000 141.115000  46.180000 141.265000 ;
        RECT   0.000000 141.265000  46.330000 141.415000 ;
        RECT   0.000000 141.415000  46.480000 141.565000 ;
        RECT   0.000000 141.565000  46.630000 141.715000 ;
        RECT   0.000000 141.715000  46.780000 141.865000 ;
        RECT   0.000000 141.865000  46.930000 142.015000 ;
        RECT   0.000000 142.015000  47.080000 142.165000 ;
        RECT   0.000000 142.165000  47.230000 142.315000 ;
        RECT   0.000000 142.315000  47.380000 142.465000 ;
        RECT   0.000000 142.465000  47.530000 142.615000 ;
        RECT   0.000000 142.615000  47.680000 142.765000 ;
        RECT   0.000000 142.765000  47.830000 142.915000 ;
        RECT   0.000000 142.915000  47.980000 143.065000 ;
        RECT   0.000000 143.065000  48.130000 143.215000 ;
        RECT   0.000000 143.215000  48.280000 143.365000 ;
        RECT   0.000000 143.365000  48.430000 143.515000 ;
        RECT   0.000000 143.515000  48.580000 143.665000 ;
        RECT   0.000000 143.665000  48.730000 143.815000 ;
        RECT   0.000000 143.815000  48.880000 143.965000 ;
        RECT   0.000000 143.965000  49.030000 144.115000 ;
        RECT   0.000000 144.115000  49.180000 144.265000 ;
        RECT   0.000000 144.265000  49.330000 144.415000 ;
        RECT   0.000000 144.415000  49.480000 144.565000 ;
        RECT   0.000000 144.565000  49.630000 144.715000 ;
        RECT   0.000000 144.715000  49.780000 144.865000 ;
        RECT   0.000000 144.865000  49.930000 145.015000 ;
        RECT   0.000000 145.015000  50.080000 145.165000 ;
        RECT   0.000000 145.165000  50.230000 145.315000 ;
        RECT   0.000000 145.315000  50.380000 145.465000 ;
        RECT   0.000000 145.465000  50.530000 145.615000 ;
        RECT   0.000000 145.615000  50.680000 145.765000 ;
        RECT   0.000000 145.765000  50.830000 145.915000 ;
        RECT   0.000000 145.915000  50.980000 146.065000 ;
        RECT   0.000000 146.065000  51.130000 146.215000 ;
        RECT   0.000000 146.215000  51.280000 146.365000 ;
        RECT   0.000000 146.365000  51.430000 146.515000 ;
        RECT   0.000000 146.515000  51.580000 146.665000 ;
        RECT   0.000000 146.665000  51.730000 146.815000 ;
        RECT   0.000000 146.815000  51.880000 146.965000 ;
        RECT   0.000000 146.965000  52.030000 147.115000 ;
        RECT   0.000000 147.115000  52.180000 147.265000 ;
        RECT   0.000000 147.265000  52.330000 147.415000 ;
        RECT   0.000000 147.415000  52.480000 147.565000 ;
        RECT   0.000000 147.565000  52.630000 147.715000 ;
        RECT   0.000000 147.715000  52.780000 147.865000 ;
        RECT   0.000000 147.865000  52.930000 148.015000 ;
        RECT   0.000000 148.015000  53.080000 148.165000 ;
        RECT   0.000000 148.165000  53.230000 148.315000 ;
        RECT   0.000000 148.315000  53.380000 148.465000 ;
        RECT   0.000000 148.465000  53.530000 148.615000 ;
        RECT   0.000000 148.615000  53.680000 148.715000 ;
        RECT  18.740000 148.715000  53.780000 148.865000 ;
        RECT  18.890000 148.865000  53.930000 149.015000 ;
        RECT  18.955000 149.015000  54.080000 149.080000 ;
        RECT  19.105000 149.080000  54.145000 149.230000 ;
        RECT  19.255000 149.230000  54.145000 149.380000 ;
        RECT  19.405000 149.380000  54.145000 149.530000 ;
        RECT  19.555000 149.530000  54.145000 149.680000 ;
        RECT  19.705000 149.680000  54.145000 149.830000 ;
        RECT  19.855000 149.830000  54.145000 149.980000 ;
        RECT  20.005000 149.980000  54.145000 150.130000 ;
        RECT  20.155000 150.130000  54.145000 150.280000 ;
        RECT  20.305000 150.280000  54.145000 150.430000 ;
        RECT  20.455000 150.430000  54.145000 150.580000 ;
        RECT  20.605000 150.580000  54.145000 150.730000 ;
        RECT  20.755000 150.730000  54.145000 150.880000 ;
        RECT  20.905000 150.880000  54.145000 151.030000 ;
        RECT  21.055000 151.030000  54.145000 151.180000 ;
        RECT  21.205000 151.180000  54.145000 151.330000 ;
        RECT  21.355000 151.330000  54.145000 151.480000 ;
        RECT  21.505000 151.480000  54.145000 151.630000 ;
        RECT  21.655000 151.630000  54.145000 151.780000 ;
        RECT  21.805000 151.780000  54.145000 151.930000 ;
        RECT  21.955000 151.930000  54.145000 152.080000 ;
        RECT  22.105000 152.080000  54.145000 152.230000 ;
        RECT  22.255000 152.230000  54.145000 152.380000 ;
        RECT  22.405000 152.380000  54.145000 152.530000 ;
        RECT  22.555000 152.530000  54.145000 152.680000 ;
        RECT  22.705000 152.680000  54.145000 152.830000 ;
        RECT  22.855000 152.830000  54.145000 152.980000 ;
        RECT  23.005000 152.980000  54.145000 153.130000 ;
        RECT  23.155000 153.130000  54.145000 153.280000 ;
        RECT  23.305000 153.280000  54.145000 153.430000 ;
        RECT  23.455000 153.430000  54.145000 153.580000 ;
        RECT  23.605000 153.580000  54.145000 153.730000 ;
        RECT  23.755000 153.730000  54.145000 153.880000 ;
        RECT  23.905000 153.880000  54.145000 154.030000 ;
        RECT  24.055000 154.030000  54.145000 154.180000 ;
        RECT  24.205000 154.180000  54.145000 154.330000 ;
        RECT  24.355000 154.330000  54.145000 154.480000 ;
        RECT  24.505000 154.480000  54.145000 154.630000 ;
        RECT  24.655000 154.630000  54.145000 154.780000 ;
        RECT  24.805000 154.780000  54.145000 154.930000 ;
        RECT  24.955000 154.930000  54.145000 155.080000 ;
        RECT  25.105000 155.080000  54.145000 155.230000 ;
        RECT  25.255000 155.230000  54.145000 155.380000 ;
        RECT  25.405000 155.380000  54.145000 155.530000 ;
        RECT  25.555000 155.530000  54.145000 155.680000 ;
        RECT  25.705000 155.680000  54.145000 155.830000 ;
        RECT  25.855000 155.830000  54.145000 155.980000 ;
        RECT  26.005000 155.980000  54.145000 156.130000 ;
        RECT  26.155000 156.130000  54.145000 156.280000 ;
        RECT  26.305000 156.280000  54.145000 156.430000 ;
        RECT  26.455000 156.430000  54.145000 156.580000 ;
        RECT  26.605000 156.580000  54.145000 156.730000 ;
        RECT  26.755000 156.730000  54.145000 156.880000 ;
        RECT  26.905000 156.880000  54.145000 157.030000 ;
        RECT  27.055000 157.030000  54.145000 157.180000 ;
        RECT  27.205000 157.180000  54.145000 157.330000 ;
        RECT  27.355000 157.330000  54.145000 157.480000 ;
        RECT  27.505000 157.480000  54.145000 157.630000 ;
        RECT  27.655000 157.630000  54.145000 157.780000 ;
        RECT  27.805000 157.780000  54.145000 157.930000 ;
        RECT  27.955000 157.930000  54.145000 158.080000 ;
        RECT  28.105000 158.080000  54.145000 158.230000 ;
        RECT  28.255000 158.230000  54.145000 158.380000 ;
        RECT  28.405000 158.380000  54.145000 158.530000 ;
        RECT  28.555000 158.530000  54.145000 158.680000 ;
        RECT  28.705000 158.680000  54.145000 158.830000 ;
        RECT  28.855000 158.830000  54.145000 158.980000 ;
        RECT  29.005000 158.980000  54.145000 159.130000 ;
        RECT  29.155000 159.130000  54.145000 159.280000 ;
        RECT  29.260000 159.280000  54.145000 159.385000 ;
        RECT  29.260000 159.385000  54.145000 197.600000 ;
        RECT  29.260000 197.600000  54.145000 197.750000 ;
        RECT  29.260000 197.750000  54.295000 197.900000 ;
        RECT  29.260000 197.900000  54.445000 198.050000 ;
        RECT  29.260000 198.050000  54.595000 198.200000 ;
        RECT  29.260000 198.200000  54.745000 198.350000 ;
        RECT  29.260000 198.350000  54.895000 198.500000 ;
        RECT  29.260000 198.500000  55.045000 198.650000 ;
        RECT  29.260000 198.650000  55.195000 198.800000 ;
        RECT  29.260000 198.800000  55.345000 198.950000 ;
        RECT  29.260000 198.950000  55.495000 199.100000 ;
        RECT  29.260000 199.100000  55.645000 199.250000 ;
        RECT  29.260000 199.250000  55.795000 199.400000 ;
        RECT  29.260000 199.400000  55.945000 199.550000 ;
        RECT  29.260000 199.550000  56.095000 199.700000 ;
        RECT  29.260000 199.700000  56.245000 199.850000 ;
        RECT  29.260000 199.850000  56.395000 200.000000 ;
        RECT  29.260000 200.000000  56.545000 200.150000 ;
        RECT  29.260000 200.150000  56.695000 200.300000 ;
        RECT  29.260000 200.300000  56.845000 200.450000 ;
        RECT  29.260000 200.450000  56.995000 200.600000 ;
        RECT  29.260000 200.600000  57.145000 200.750000 ;
        RECT  29.260000 200.750000  57.295000 200.900000 ;
        RECT  29.260000 200.900000  57.445000 201.050000 ;
        RECT  29.260000 201.050000  57.595000 201.200000 ;
        RECT  29.260000 201.200000  57.745000 201.350000 ;
        RECT  29.260000 201.350000  57.895000 201.500000 ;
        RECT  29.260000 201.500000  58.045000 201.650000 ;
        RECT  29.260000 201.650000  58.195000 201.800000 ;
        RECT  29.260000 201.800000  58.345000 201.950000 ;
        RECT  29.260000 201.950000  58.495000 202.100000 ;
        RECT  29.260000 202.100000  58.645000 202.250000 ;
        RECT  29.260000 202.250000  58.795000 202.400000 ;
        RECT  29.260000 202.400000  58.945000 202.550000 ;
        RECT  29.260000 202.550000  59.095000 202.700000 ;
        RECT  29.260000 202.700000  59.245000 202.850000 ;
        RECT  29.260000 202.850000  59.395000 203.000000 ;
        RECT  29.260000 203.000000  59.545000 203.150000 ;
        RECT  29.260000 203.150000  59.695000 203.300000 ;
        RECT  29.260000 203.300000  59.845000 203.450000 ;
        RECT  29.260000 203.450000  59.995000 203.600000 ;
        RECT  29.260000 203.600000  60.145000 203.750000 ;
        RECT  29.260000 203.750000  60.295000 203.900000 ;
        RECT  29.260000 203.900000  60.445000 204.050000 ;
        RECT  29.260000 204.050000  60.595000 204.200000 ;
        RECT  29.260000 204.200000  60.745000 204.350000 ;
        RECT  29.260000 204.350000  60.895000 204.500000 ;
        RECT  29.260000 204.500000  61.045000 204.505000 ;
        RECT  29.260000 204.505000 422.530000 204.655000 ;
        RECT  29.260000 204.655000 422.380000 204.805000 ;
        RECT  29.260000 204.805000 422.230000 204.955000 ;
        RECT  29.260000 204.955000 422.080000 205.105000 ;
        RECT  29.260000 205.105000 421.930000 205.255000 ;
        RECT  29.260000 205.255000 421.780000 205.405000 ;
        RECT  29.260000 205.405000 421.630000 205.555000 ;
        RECT  29.260000 205.555000 421.480000 205.705000 ;
        RECT  29.260000 205.705000 421.330000 205.855000 ;
        RECT  29.260000 205.855000 421.180000 206.005000 ;
        RECT  29.260000 206.005000 421.030000 206.155000 ;
        RECT  29.260000 206.155000 420.880000 206.305000 ;
        RECT  29.260000 206.305000 420.730000 206.455000 ;
        RECT  29.260000 206.455000 420.580000 206.605000 ;
        RECT  29.260000 206.605000 420.430000 206.755000 ;
        RECT  29.260000 206.755000 420.280000 206.905000 ;
        RECT  29.260000 206.905000 420.130000 207.055000 ;
        RECT  29.260000 207.055000 419.980000 207.205000 ;
        RECT  29.260000 207.205000 419.860000 207.325000 ;
        RECT  29.410000 207.325000 419.710000 207.475000 ;
        RECT  29.560000 207.475000 419.560000 207.625000 ;
        RECT  29.710000 207.625000 419.410000 207.775000 ;
        RECT  29.860000 207.775000 419.260000 207.925000 ;
        RECT  30.010000 207.925000 419.110000 208.075000 ;
        RECT  30.160000 208.075000 418.960000 208.225000 ;
        RECT  30.310000 208.225000 418.810000 208.375000 ;
        RECT  30.460000 208.375000 418.660000 208.525000 ;
        RECT  30.610000 208.525000 418.510000 208.675000 ;
        RECT  30.760000 208.675000 418.360000 208.825000 ;
        RECT  30.910000 208.825000 418.210000 208.975000 ;
        RECT  31.060000 208.975000 418.060000 209.125000 ;
        RECT  31.210000 209.125000 417.910000 209.275000 ;
        RECT  31.360000 209.275000 417.760000 209.425000 ;
        RECT  31.510000 209.425000 417.610000 209.575000 ;
        RECT  31.660000 209.575000 417.460000 209.725000 ;
        RECT  31.810000 209.725000 417.310000 209.875000 ;
        RECT  31.960000 209.875000 417.160000 210.025000 ;
        RECT  32.110000 210.025000 417.010000 210.175000 ;
        RECT  32.260000 210.175000 416.860000 210.325000 ;
        RECT  32.410000 210.325000 416.710000 210.475000 ;
        RECT  32.560000 210.475000 416.560000 210.625000 ;
        RECT  32.710000 210.625000 416.410000 210.775000 ;
        RECT  32.860000 210.775000 416.260000 210.925000 ;
        RECT  33.010000 210.925000 416.110000 211.075000 ;
        RECT  33.160000 211.075000 415.960000 211.225000 ;
        RECT  33.310000 211.225000 415.810000 211.375000 ;
        RECT  33.460000 211.375000 415.660000 211.525000 ;
        RECT  33.610000 211.525000 415.510000 211.675000 ;
        RECT  33.760000 211.675000 415.360000 211.825000 ;
        RECT  33.910000 211.825000 415.210000 211.975000 ;
        RECT  34.060000 211.975000 415.060000 212.125000 ;
        RECT  34.210000 212.125000 414.910000 212.275000 ;
        RECT  34.360000 212.275000 414.760000 212.425000 ;
        RECT  34.510000 212.425000 414.610000 212.575000 ;
        RECT  34.660000 212.575000 414.460000 212.725000 ;
        RECT  34.810000 212.725000 414.310000 212.875000 ;
        RECT  34.960000 212.875000 414.160000 213.025000 ;
        RECT  35.110000 213.025000 414.010000 213.175000 ;
        RECT  35.260000 213.175000 413.860000 213.325000 ;
        RECT  35.410000 213.325000 413.710000 213.475000 ;
        RECT  35.560000 213.475000 413.560000 213.625000 ;
        RECT  35.710000 213.625000 413.410000 213.775000 ;
        RECT  35.860000 213.775000 413.260000 213.925000 ;
        RECT  36.010000 213.925000 413.110000 214.075000 ;
        RECT  36.160000 214.075000 412.960000 214.225000 ;
        RECT  36.310000 214.225000 412.810000 214.375000 ;
        RECT  36.460000 214.375000 412.660000 214.525000 ;
        RECT  36.610000 214.525000 412.510000 214.675000 ;
        RECT  36.760000 214.675000 412.360000 214.825000 ;
        RECT  36.910000 214.825000 412.210000 214.975000 ;
        RECT  37.060000 214.975000 412.060000 215.125000 ;
        RECT  37.210000 215.125000 411.910000 215.275000 ;
        RECT  37.360000 215.275000 411.760000 215.425000 ;
        RECT  37.510000 215.425000 411.610000 215.575000 ;
        RECT  37.660000 215.575000 411.460000 215.725000 ;
        RECT  37.810000 215.725000 411.310000 215.875000 ;
        RECT  37.960000 215.875000 411.160000 216.025000 ;
        RECT  38.110000 216.025000 411.010000 216.175000 ;
        RECT  38.260000 216.175000 410.860000 216.325000 ;
        RECT  38.410000 216.325000 410.710000 216.475000 ;
        RECT  38.560000 216.475000 410.560000 216.625000 ;
        RECT  38.710000 216.625000 410.410000 216.775000 ;
        RECT  38.860000 216.775000 410.260000 216.925000 ;
        RECT  39.010000 216.925000 410.110000 217.075000 ;
        RECT  39.160000 217.075000 409.960000 217.225000 ;
        RECT  39.310000 217.225000 409.810000 217.375000 ;
        RECT  39.460000 217.375000 409.660000 217.525000 ;
        RECT  39.610000 217.525000 409.510000 217.675000 ;
        RECT  39.760000 217.675000 409.360000 217.825000 ;
        RECT  39.910000 217.825000 409.210000 217.975000 ;
        RECT  40.060000 217.975000 409.060000 218.125000 ;
        RECT  40.210000 218.125000 408.910000 218.275000 ;
        RECT  40.360000 218.275000 408.760000 218.425000 ;
        RECT  40.510000 218.425000 408.610000 218.575000 ;
        RECT  40.660000 218.575000 408.460000 218.725000 ;
        RECT  40.810000 218.725000 408.310000 218.875000 ;
        RECT  40.960000 218.875000 408.160000 219.025000 ;
        RECT  41.110000 219.025000 408.010000 219.175000 ;
        RECT  41.260000 219.175000 407.860000 219.325000 ;
        RECT  41.410000 219.325000 407.710000 219.475000 ;
        RECT  41.560000 219.475000 407.560000 219.625000 ;
        RECT  41.710000 219.625000 407.410000 219.775000 ;
        RECT  41.860000 219.775000 407.260000 219.925000 ;
        RECT  42.010000 219.925000 407.110000 220.075000 ;
        RECT  42.160000 220.075000 406.960000 220.225000 ;
        RECT  42.310000 220.225000 406.810000 220.375000 ;
        RECT  42.460000 220.375000 406.660000 220.525000 ;
        RECT  42.610000 220.525000 406.510000 220.675000 ;
        RECT  42.760000 220.675000 406.360000 220.825000 ;
        RECT  42.910000 220.825000 406.210000 220.975000 ;
        RECT  43.060000 220.975000 406.060000 221.125000 ;
        RECT  43.210000 221.125000 405.910000 221.275000 ;
        RECT  43.360000 221.275000 405.760000 221.425000 ;
        RECT  43.510000 221.425000 405.610000 221.575000 ;
        RECT  43.660000 221.575000 405.460000 221.725000 ;
        RECT  43.810000 221.725000 405.310000 221.875000 ;
        RECT  43.960000 221.875000 405.160000 222.025000 ;
        RECT  44.110000 222.025000 405.010000 222.175000 ;
        RECT  44.260000 222.175000 404.860000 222.325000 ;
        RECT  44.410000 222.325000 404.710000 222.475000 ;
        RECT  44.560000 222.475000 404.560000 222.625000 ;
        RECT  44.710000 222.625000 404.410000 222.775000 ;
        RECT  44.860000 222.775000 404.260000 222.925000 ;
        RECT  45.010000 222.925000 404.110000 223.075000 ;
        RECT  45.160000 223.075000 403.960000 223.225000 ;
        RECT  45.310000 223.225000 403.810000 223.375000 ;
        RECT  45.460000 223.375000 403.660000 223.525000 ;
        RECT  45.610000 223.525000 403.510000 223.675000 ;
        RECT  45.760000 223.675000 403.360000 223.825000 ;
        RECT  45.910000 223.825000 403.210000 223.975000 ;
        RECT  46.060000 223.975000 403.060000 224.125000 ;
        RECT  46.210000 224.125000 402.910000 224.275000 ;
        RECT  46.360000 224.275000 402.760000 224.425000 ;
        RECT  46.510000 224.425000 402.610000 224.575000 ;
        RECT  46.660000 224.575000 402.460000 224.725000 ;
        RECT  46.810000 224.725000 402.310000 224.875000 ;
        RECT  46.960000 224.875000 402.160000 225.025000 ;
        RECT  47.110000 225.025000 402.010000 225.175000 ;
        RECT  47.260000 225.175000 401.860000 225.325000 ;
        RECT  47.410000 225.325000 401.710000 225.475000 ;
        RECT  47.560000 225.475000 401.560000 225.625000 ;
        RECT  47.710000 225.625000 401.410000 225.775000 ;
        RECT  47.860000 225.775000 401.260000 225.925000 ;
        RECT  48.010000 225.925000 401.110000 226.075000 ;
        RECT  48.160000 226.075000 400.960000 226.225000 ;
        RECT  48.310000 226.225000 400.810000 226.375000 ;
        RECT  48.460000 226.375000 400.660000 226.525000 ;
        RECT  48.610000 226.525000 400.510000 226.675000 ;
        RECT  48.760000 226.675000 400.360000 226.825000 ;
        RECT  48.910000 226.825000 400.210000 226.975000 ;
        RECT  49.060000 226.975000 400.060000 227.125000 ;
        RECT  49.210000 227.125000 399.910000 227.275000 ;
        RECT  49.360000 227.275000 399.760000 227.425000 ;
        RECT  49.510000 227.425000 399.610000 227.575000 ;
        RECT  49.660000 227.575000 399.460000 227.725000 ;
        RECT  49.810000 227.725000 399.310000 227.875000 ;
        RECT  49.835000 227.875000 399.285000 227.900000 ;
        RECT 388.110000 204.365000 422.680000 204.505000 ;
        RECT 388.260000 204.215000 422.820000 204.365000 ;
        RECT 388.410000 204.065000 422.970000 204.215000 ;
        RECT 388.560000 203.915000 423.120000 204.065000 ;
        RECT 388.710000 203.765000 423.270000 203.915000 ;
        RECT 388.860000 203.615000 423.420000 203.765000 ;
        RECT 389.010000 203.465000 423.570000 203.615000 ;
        RECT 389.160000 203.315000 423.720000 203.465000 ;
        RECT 389.310000 203.165000 423.870000 203.315000 ;
        RECT 389.460000 203.015000 424.020000 203.165000 ;
        RECT 389.610000 202.865000 424.170000 203.015000 ;
        RECT 389.760000 202.715000 424.320000 202.865000 ;
        RECT 389.910000 202.565000 424.470000 202.715000 ;
        RECT 390.060000 202.415000 424.620000 202.565000 ;
        RECT 390.210000 202.265000 424.770000 202.415000 ;
        RECT 390.360000 202.115000 424.920000 202.265000 ;
        RECT 390.510000 201.965000 425.070000 202.115000 ;
        RECT 390.660000 201.815000 425.220000 201.965000 ;
        RECT 390.810000 201.665000 425.370000 201.815000 ;
        RECT 390.960000 201.515000 425.520000 201.665000 ;
        RECT 391.110000 201.365000 425.670000 201.515000 ;
        RECT 391.260000 201.215000 425.820000 201.365000 ;
        RECT 391.410000 201.065000 425.970000 201.215000 ;
        RECT 391.560000 200.915000 426.120000 201.065000 ;
        RECT 391.710000 200.765000 426.270000 200.915000 ;
        RECT 391.860000 200.615000 426.420000 200.765000 ;
        RECT 392.010000 200.465000 426.570000 200.615000 ;
        RECT 392.160000 200.315000 426.720000 200.465000 ;
        RECT 392.310000 200.165000 426.870000 200.315000 ;
        RECT 392.460000 200.015000 427.020000 200.165000 ;
        RECT 392.610000 199.865000 427.170000 200.015000 ;
        RECT 392.760000 199.715000 427.320000 199.865000 ;
        RECT 392.910000 199.565000 427.470000 199.715000 ;
        RECT 393.060000 199.415000 427.620000 199.565000 ;
        RECT 393.210000 199.265000 427.770000 199.415000 ;
        RECT 393.360000 199.115000 427.920000 199.265000 ;
        RECT 393.510000 198.965000 428.070000 199.115000 ;
        RECT 393.660000 198.815000 428.220000 198.965000 ;
        RECT 393.810000 198.665000 428.370000 198.815000 ;
        RECT 393.960000 198.515000 428.520000 198.665000 ;
        RECT 394.110000 198.365000 428.670000 198.515000 ;
        RECT 394.260000 198.215000 428.820000 198.365000 ;
        RECT 394.410000 198.065000 428.970000 198.215000 ;
        RECT 394.560000 197.915000 429.120000 198.065000 ;
        RECT 394.710000 197.765000 429.270000 197.915000 ;
        RECT 394.860000 197.615000 429.420000 197.765000 ;
        RECT 395.010000 197.465000 429.570000 197.615000 ;
        RECT 395.160000 197.315000 429.720000 197.465000 ;
        RECT 395.310000 197.165000 429.870000 197.315000 ;
        RECT 395.460000 197.015000 430.020000 197.165000 ;
        RECT 395.610000 196.865000 430.170000 197.015000 ;
        RECT 395.760000 196.715000 430.320000 196.865000 ;
        RECT 395.910000 196.565000 430.470000 196.715000 ;
        RECT 396.060000 196.415000 430.620000 196.565000 ;
        RECT 396.210000 196.265000 430.770000 196.415000 ;
        RECT 396.360000 196.115000 430.920000 196.265000 ;
        RECT 396.510000 195.965000 431.070000 196.115000 ;
        RECT 396.660000 195.815000 431.220000 195.965000 ;
        RECT 396.810000 195.665000 431.370000 195.815000 ;
        RECT 396.960000 195.515000 431.520000 195.665000 ;
        RECT 397.110000 195.365000 431.670000 195.515000 ;
        RECT 397.260000 195.215000 431.820000 195.365000 ;
        RECT 397.410000 195.065000 431.970000 195.215000 ;
        RECT 397.560000 194.915000 432.120000 195.065000 ;
        RECT 397.710000 194.765000 432.270000 194.915000 ;
        RECT 397.860000 194.615000 432.420000 194.765000 ;
        RECT 398.010000 194.465000 432.570000 194.615000 ;
        RECT 398.160000 194.315000 432.720000 194.465000 ;
        RECT 398.310000 194.165000 432.870000 194.315000 ;
        RECT 398.460000 194.015000 433.020000 194.165000 ;
        RECT 398.610000 193.865000 433.170000 194.015000 ;
        RECT 398.760000 193.715000 433.320000 193.865000 ;
        RECT 398.910000 193.565000 433.470000 193.715000 ;
        RECT 399.060000 193.415000 433.620000 193.565000 ;
        RECT 399.210000 193.265000 433.770000 193.415000 ;
        RECT 399.360000 193.115000 433.920000 193.265000 ;
        RECT 399.510000 192.965000 434.070000 193.115000 ;
        RECT 399.660000 192.815000 434.220000 192.965000 ;
        RECT 399.810000 192.665000 434.370000 192.815000 ;
        RECT 399.960000 192.515000 434.520000 192.665000 ;
        RECT 400.110000 192.365000 434.670000 192.515000 ;
        RECT 400.260000 192.215000 434.820000 192.365000 ;
        RECT 400.410000 192.065000 434.970000 192.215000 ;
        RECT 400.560000 191.915000 435.120000 192.065000 ;
        RECT 400.710000 191.765000 435.270000 191.915000 ;
        RECT 400.860000 191.615000 435.420000 191.765000 ;
        RECT 401.010000 191.465000 435.570000 191.615000 ;
        RECT 401.160000 191.315000 435.720000 191.465000 ;
        RECT 401.310000 191.165000 435.870000 191.315000 ;
        RECT 401.460000 191.015000 436.020000 191.165000 ;
        RECT 401.610000 190.865000 436.170000 191.015000 ;
        RECT 401.760000 190.715000 436.320000 190.865000 ;
        RECT 401.910000 190.565000 436.470000 190.715000 ;
        RECT 402.060000 190.415000 436.620000 190.565000 ;
        RECT 402.210000 190.265000 436.770000 190.415000 ;
        RECT 402.360000 190.115000 436.920000 190.265000 ;
        RECT 402.510000 189.965000 437.070000 190.115000 ;
        RECT 402.660000 189.815000 437.220000 189.965000 ;
        RECT 402.810000 189.665000 437.370000 189.815000 ;
        RECT 402.960000 189.515000 437.520000 189.665000 ;
        RECT 403.110000 189.365000 437.670000 189.515000 ;
        RECT 403.260000 189.215000 437.820000 189.365000 ;
        RECT 403.410000 189.065000 437.970000 189.215000 ;
        RECT 403.560000 188.915000 438.120000 189.065000 ;
        RECT 403.710000 188.765000 438.270000 188.915000 ;
        RECT 403.860000 188.615000 438.420000 188.765000 ;
        RECT 404.010000 188.465000 438.570000 188.615000 ;
        RECT 404.160000 188.315000 438.720000 188.465000 ;
        RECT 404.310000 188.165000 438.870000 188.315000 ;
        RECT 404.460000 188.015000 439.020000 188.165000 ;
        RECT 404.610000 187.865000 439.170000 188.015000 ;
        RECT 404.760000 187.715000 439.320000 187.865000 ;
        RECT 404.910000 187.565000 439.470000 187.715000 ;
        RECT 405.060000 187.415000 439.620000 187.565000 ;
        RECT 405.210000 187.265000 439.770000 187.415000 ;
        RECT 405.360000 187.115000 439.920000 187.265000 ;
        RECT 405.510000 186.965000 440.070000 187.115000 ;
        RECT 405.660000 186.815000 440.220000 186.965000 ;
        RECT 405.810000 186.665000 440.370000 186.815000 ;
        RECT 405.960000 186.515000 440.520000 186.665000 ;
        RECT 406.110000 186.365000 440.670000 186.515000 ;
        RECT 406.260000 186.215000 440.820000 186.365000 ;
        RECT 406.410000 186.065000 440.970000 186.215000 ;
        RECT 406.560000 185.915000 441.120000 186.065000 ;
        RECT 406.710000 185.765000 441.270000 185.915000 ;
        RECT 406.860000 185.615000 441.420000 185.765000 ;
        RECT 407.010000 185.465000 441.570000 185.615000 ;
        RECT 407.160000 185.315000 441.720000 185.465000 ;
        RECT 407.310000 185.165000 441.870000 185.315000 ;
        RECT 407.460000 185.015000 442.020000 185.165000 ;
        RECT 407.610000 184.865000 442.170000 185.015000 ;
        RECT 407.760000 184.715000 442.320000 184.865000 ;
        RECT 407.910000 184.565000 442.470000 184.715000 ;
        RECT 408.060000 184.415000 442.620000 184.565000 ;
        RECT 408.210000 184.265000 442.770000 184.415000 ;
        RECT 408.360000 184.115000 442.920000 184.265000 ;
        RECT 408.510000 183.965000 443.070000 184.115000 ;
        RECT 408.660000 183.815000 443.220000 183.965000 ;
        RECT 408.810000 183.665000 443.370000 183.815000 ;
        RECT 408.960000 183.515000 443.520000 183.665000 ;
        RECT 409.110000 183.365000 443.670000 183.515000 ;
        RECT 409.260000 183.215000 443.820000 183.365000 ;
        RECT 409.410000 183.065000 443.970000 183.215000 ;
        RECT 409.560000 182.915000 444.120000 183.065000 ;
        RECT 409.710000 182.765000 444.270000 182.915000 ;
        RECT 409.860000 182.615000 444.420000 182.765000 ;
        RECT 410.010000 182.465000 444.570000 182.615000 ;
        RECT 410.160000 182.315000 444.720000 182.465000 ;
        RECT 410.310000 182.165000 444.870000 182.315000 ;
        RECT 410.460000 182.015000 445.020000 182.165000 ;
        RECT 410.610000 181.865000 445.170000 182.015000 ;
        RECT 410.760000 181.715000 445.320000 181.865000 ;
        RECT 410.910000 181.565000 445.470000 181.715000 ;
        RECT 411.060000 181.415000 445.620000 181.565000 ;
        RECT 411.210000 181.265000 445.770000 181.415000 ;
        RECT 411.360000 181.115000 445.920000 181.265000 ;
        RECT 411.510000 180.965000 446.070000 181.115000 ;
        RECT 411.660000 180.815000 446.220000 180.965000 ;
        RECT 411.810000 180.665000 446.370000 180.815000 ;
        RECT 411.960000 180.515000 446.520000 180.665000 ;
        RECT 412.110000 180.365000 446.670000 180.515000 ;
        RECT 412.260000 180.215000 446.820000 180.365000 ;
        RECT 412.410000 180.065000 446.970000 180.215000 ;
        RECT 412.560000 179.915000 447.120000 180.065000 ;
        RECT 412.710000 179.765000 447.270000 179.915000 ;
        RECT 412.860000 179.615000 447.420000 179.765000 ;
        RECT 413.010000 179.465000 447.570000 179.615000 ;
        RECT 413.160000 179.315000 447.720000 179.465000 ;
        RECT 413.310000 179.165000 447.870000 179.315000 ;
        RECT 413.460000 179.015000 448.020000 179.165000 ;
        RECT 413.610000 178.865000 448.170000 179.015000 ;
        RECT 413.760000 178.715000 448.320000 178.865000 ;
        RECT 413.910000 178.565000 448.470000 178.715000 ;
        RECT 414.060000 178.415000 448.620000 178.565000 ;
        RECT 414.210000 178.265000 448.770000 178.415000 ;
        RECT 414.360000 178.115000 448.920000 178.265000 ;
        RECT 414.510000 177.965000 449.070000 178.115000 ;
        RECT 414.660000 177.815000 449.220000 177.965000 ;
        RECT 414.810000 177.665000 449.370000 177.815000 ;
        RECT 414.960000 177.515000 449.520000 177.665000 ;
        RECT 415.110000 177.365000 449.670000 177.515000 ;
        RECT 415.260000 177.215000 449.820000 177.365000 ;
        RECT 415.410000 177.065000 449.970000 177.215000 ;
        RECT 415.560000 176.915000 450.120000 177.065000 ;
        RECT 415.710000 176.765000 450.270000 176.915000 ;
        RECT 415.860000 176.615000 450.420000 176.765000 ;
        RECT 416.010000 176.465000 450.570000 176.615000 ;
        RECT 416.160000 176.315000 450.720000 176.465000 ;
        RECT 416.310000 176.165000 450.870000 176.315000 ;
        RECT 416.460000 176.015000 451.020000 176.165000 ;
        RECT 416.610000 175.865000 451.170000 176.015000 ;
        RECT 416.760000 175.715000 451.320000 175.865000 ;
        RECT 416.910000 175.565000 451.470000 175.715000 ;
        RECT 417.060000 175.415000 451.620000 175.565000 ;
        RECT 417.210000 175.265000 451.770000 175.415000 ;
        RECT 417.360000 175.115000 451.920000 175.265000 ;
        RECT 417.510000 174.965000 452.070000 175.115000 ;
        RECT 417.660000 174.815000 452.220000 174.965000 ;
        RECT 417.810000 174.665000 452.370000 174.815000 ;
        RECT 417.960000 174.515000 452.520000 174.665000 ;
        RECT 418.110000 174.365000 452.670000 174.515000 ;
        RECT 418.260000 174.215000 452.820000 174.365000 ;
        RECT 418.410000 174.065000 452.970000 174.215000 ;
        RECT 418.560000 173.915000 453.120000 174.065000 ;
        RECT 418.710000 173.765000 453.270000 173.915000 ;
        RECT 418.860000 173.615000 453.420000 173.765000 ;
        RECT 419.010000 173.465000 453.570000 173.615000 ;
        RECT 419.160000 173.315000 453.720000 173.465000 ;
        RECT 419.310000 173.165000 453.870000 173.315000 ;
        RECT 419.460000 173.015000 454.020000 173.165000 ;
        RECT 419.610000 172.865000 454.170000 173.015000 ;
        RECT 419.760000 172.715000 454.320000 172.865000 ;
        RECT 419.910000 172.565000 454.470000 172.715000 ;
        RECT 420.060000 172.415000 454.620000 172.565000 ;
        RECT 420.210000 172.265000 454.770000 172.415000 ;
        RECT 420.360000 172.115000 454.920000 172.265000 ;
        RECT 420.510000 171.965000 455.070000 172.115000 ;
        RECT 420.660000 171.815000 455.220000 171.965000 ;
        RECT 420.810000 171.665000 455.370000 171.815000 ;
        RECT 420.960000 171.515000 455.520000 171.665000 ;
        RECT 421.110000 171.365000 455.670000 171.515000 ;
        RECT 421.260000 171.215000 455.820000 171.365000 ;
        RECT 421.410000 171.065000 455.970000 171.215000 ;
        RECT 421.560000 170.915000 456.120000 171.065000 ;
        RECT 421.710000 170.765000 456.270000 170.915000 ;
        RECT 421.860000 170.615000 456.420000 170.765000 ;
        RECT 422.010000 170.465000 456.570000 170.615000 ;
        RECT 422.160000 170.315000 456.720000 170.465000 ;
        RECT 422.310000 170.165000 456.870000 170.315000 ;
        RECT 422.460000 170.015000 457.020000 170.165000 ;
        RECT 422.610000 169.865000 457.170000 170.015000 ;
        RECT 422.760000 169.715000 457.320000 169.865000 ;
        RECT 422.910000 169.565000 457.470000 169.715000 ;
        RECT 423.060000 169.415000 457.620000 169.565000 ;
        RECT 423.210000 169.265000 457.770000 169.415000 ;
        RECT 423.360000 169.115000 457.920000 169.265000 ;
        RECT 423.510000 168.965000 458.070000 169.115000 ;
        RECT 423.660000 168.815000 458.220000 168.965000 ;
        RECT 423.810000 168.665000 458.370000 168.815000 ;
        RECT 423.960000 168.515000 458.520000 168.665000 ;
        RECT 424.110000 168.365000 458.670000 168.515000 ;
        RECT 424.260000 168.215000 458.820000 168.365000 ;
        RECT 424.410000 168.065000 458.970000 168.215000 ;
        RECT 424.560000 167.915000 459.120000 168.065000 ;
        RECT 424.710000 167.765000 459.270000 167.915000 ;
        RECT 424.860000 167.615000 459.420000 167.765000 ;
        RECT 425.010000 167.465000 459.570000 167.615000 ;
        RECT 425.160000 167.315000 459.720000 167.465000 ;
        RECT 425.310000 167.165000 459.870000 167.315000 ;
        RECT 425.460000 167.015000 460.020000 167.165000 ;
        RECT 425.610000 166.865000 460.170000 167.015000 ;
        RECT 425.760000 166.715000 460.320000 166.865000 ;
        RECT 425.910000 166.565000 460.470000 166.715000 ;
        RECT 426.060000 166.415000 460.620000 166.565000 ;
        RECT 426.210000 166.265000 460.770000 166.415000 ;
        RECT 426.360000 166.115000 460.920000 166.265000 ;
        RECT 426.510000 165.965000 461.070000 166.115000 ;
        RECT 426.660000 165.815000 461.220000 165.965000 ;
        RECT 426.810000 165.665000 461.370000 165.815000 ;
        RECT 426.960000 165.515000 461.520000 165.665000 ;
        RECT 427.110000 165.365000 461.670000 165.515000 ;
        RECT 427.260000 165.215000 461.820000 165.365000 ;
        RECT 427.410000 165.065000 461.970000 165.215000 ;
        RECT 427.560000 164.915000 462.120000 165.065000 ;
        RECT 427.710000 164.765000 462.270000 164.915000 ;
        RECT 427.860000 164.615000 462.420000 164.765000 ;
        RECT 428.010000 164.465000 462.570000 164.615000 ;
        RECT 428.160000 164.315000 462.720000 164.465000 ;
        RECT 428.310000 164.165000 462.870000 164.315000 ;
        RECT 428.460000 164.015000 463.020000 164.165000 ;
        RECT 428.610000 163.865000 463.170000 164.015000 ;
        RECT 428.760000 163.715000 463.320000 163.865000 ;
        RECT 428.910000 163.565000 463.470000 163.715000 ;
        RECT 429.060000 163.415000 463.620000 163.565000 ;
        RECT 429.210000 163.265000 463.770000 163.415000 ;
        RECT 429.360000 163.115000 463.920000 163.265000 ;
        RECT 429.510000 162.965000 464.070000 163.115000 ;
        RECT 429.660000 162.815000 464.220000 162.965000 ;
        RECT 429.810000 162.665000 464.370000 162.815000 ;
        RECT 429.960000 162.515000 464.520000 162.665000 ;
        RECT 430.110000 162.365000 464.670000 162.515000 ;
        RECT 430.260000 162.215000 464.820000 162.365000 ;
        RECT 430.410000 162.065000 464.970000 162.215000 ;
        RECT 430.560000 161.915000 465.120000 162.065000 ;
        RECT 430.710000 161.765000 465.270000 161.915000 ;
        RECT 430.860000 161.615000 465.420000 161.765000 ;
        RECT 431.010000 161.465000 465.570000 161.615000 ;
        RECT 431.160000 161.315000 465.720000 161.465000 ;
        RECT 431.310000 161.165000 465.870000 161.315000 ;
        RECT 431.460000 161.015000 466.020000 161.165000 ;
        RECT 431.610000 160.865000 466.170000 161.015000 ;
        RECT 431.760000 160.715000 466.320000 160.865000 ;
        RECT 431.910000 160.565000 466.470000 160.715000 ;
        RECT 432.060000 160.415000 466.620000 160.565000 ;
        RECT 432.210000 160.265000 466.770000 160.415000 ;
        RECT 432.360000 160.115000 466.920000 160.265000 ;
        RECT 432.510000 159.965000 467.070000 160.115000 ;
        RECT 432.660000 159.815000 467.220000 159.965000 ;
        RECT 432.810000 159.665000 467.370000 159.815000 ;
        RECT 432.960000 159.515000 467.520000 159.665000 ;
        RECT 433.110000 159.365000 467.670000 159.515000 ;
        RECT 433.260000 159.215000 467.820000 159.365000 ;
        RECT 433.410000 159.065000 467.970000 159.215000 ;
        RECT 433.560000 158.915000 468.120000 159.065000 ;
        RECT 433.710000 158.765000 468.270000 158.915000 ;
        RECT 433.860000 158.615000 468.420000 158.765000 ;
        RECT 434.010000 158.465000 468.570000 158.615000 ;
        RECT 434.160000 158.315000 468.720000 158.465000 ;
        RECT 434.310000 158.165000 468.870000 158.315000 ;
        RECT 434.460000 158.015000 469.020000 158.165000 ;
        RECT 434.610000 157.865000 469.170000 158.015000 ;
        RECT 434.760000 157.715000 469.320000 157.865000 ;
        RECT 434.910000 157.565000 469.470000 157.715000 ;
        RECT 435.060000 157.415000 469.620000 157.565000 ;
        RECT 435.210000 157.265000 469.770000 157.415000 ;
        RECT 435.360000 157.115000 469.920000 157.265000 ;
        RECT 435.510000 156.965000 470.070000 157.115000 ;
        RECT 435.660000 156.815000 470.220000 156.965000 ;
        RECT 435.810000 156.665000 470.370000 156.815000 ;
        RECT 435.960000 156.515000 470.520000 156.665000 ;
        RECT 436.110000 156.365000 470.670000 156.515000 ;
        RECT 436.260000 156.215000 470.820000 156.365000 ;
        RECT 436.410000 156.065000 470.970000 156.215000 ;
        RECT 436.560000 155.915000 471.120000 156.065000 ;
        RECT 436.710000 155.765000 471.270000 155.915000 ;
        RECT 436.860000 155.615000 471.420000 155.765000 ;
        RECT 437.010000 155.465000 471.570000 155.615000 ;
        RECT 437.160000 155.315000 471.720000 155.465000 ;
        RECT 437.310000 155.165000 471.870000 155.315000 ;
        RECT 437.460000 155.015000 472.020000 155.165000 ;
        RECT 437.610000 154.865000 472.170000 155.015000 ;
        RECT 437.760000 154.715000 472.320000 154.865000 ;
        RECT 437.910000 154.565000 472.470000 154.715000 ;
        RECT 438.060000 154.415000 472.620000 154.565000 ;
        RECT 438.210000 154.265000 472.770000 154.415000 ;
        RECT 438.360000 154.115000 472.920000 154.265000 ;
        RECT 438.510000 153.965000 473.070000 154.115000 ;
        RECT 438.660000 153.815000 473.220000 153.965000 ;
        RECT 438.810000 153.665000 473.370000 153.815000 ;
        RECT 438.960000 153.515000 473.520000 153.665000 ;
        RECT 439.110000 153.365000 473.670000 153.515000 ;
        RECT 439.260000 153.215000 473.820000 153.365000 ;
        RECT 439.410000 153.065000 473.970000 153.215000 ;
        RECT 439.560000 152.915000 474.120000 153.065000 ;
        RECT 439.710000 152.765000 474.270000 152.915000 ;
        RECT 439.860000 152.615000 474.420000 152.765000 ;
        RECT 440.010000 152.465000 474.570000 152.615000 ;
        RECT 440.160000 152.315000 474.720000 152.465000 ;
        RECT 440.310000 152.165000 474.870000 152.315000 ;
        RECT 440.460000 152.015000 475.020000 152.165000 ;
        RECT 440.610000 151.865000 475.170000 152.015000 ;
        RECT 440.760000 151.715000 475.320000 151.865000 ;
        RECT 440.910000 151.565000 475.470000 151.715000 ;
        RECT 441.060000 151.415000 475.620000 151.565000 ;
        RECT 441.210000 151.265000 475.770000 151.415000 ;
        RECT 441.360000 151.115000 475.920000 151.265000 ;
        RECT 441.510000 150.965000 476.070000 151.115000 ;
        RECT 441.660000 150.815000 476.220000 150.965000 ;
        RECT 441.810000 150.665000 476.370000 150.815000 ;
        RECT 441.960000 150.515000 476.520000 150.665000 ;
        RECT 442.110000 150.365000 476.670000 150.515000 ;
        RECT 442.260000 150.215000 476.820000 150.365000 ;
        RECT 442.410000 150.065000 476.970000 150.215000 ;
        RECT 442.560000 149.915000 477.120000 150.065000 ;
        RECT 442.710000 149.765000 477.270000 149.915000 ;
        RECT 442.860000 149.615000 477.420000 149.765000 ;
        RECT 443.010000 149.465000 477.570000 149.615000 ;
        RECT 443.160000 149.315000 477.720000 149.465000 ;
        RECT 443.310000 149.165000 477.870000 149.315000 ;
        RECT 443.460000 149.015000 478.020000 149.165000 ;
        RECT 443.610000 148.865000 478.170000 149.015000 ;
        RECT 443.760000 148.715000 478.320000 148.865000 ;
        RECT 443.825000 148.650000 480.000000 148.715000 ;
        RECT 443.975000 148.500000 480.000000 148.650000 ;
        RECT 444.125000 148.350000 480.000000 148.500000 ;
        RECT 444.275000 148.200000 480.000000 148.350000 ;
        RECT 444.425000 148.050000 480.000000 148.200000 ;
        RECT 444.575000 147.900000 480.000000 148.050000 ;
        RECT 444.725000 147.750000 480.000000 147.900000 ;
        RECT 444.875000 147.600000 480.000000 147.750000 ;
        RECT 445.025000 147.450000 480.000000 147.600000 ;
        RECT 445.175000 147.300000 480.000000 147.450000 ;
        RECT 445.325000 147.150000 480.000000 147.300000 ;
        RECT 445.475000 147.000000 480.000000 147.150000 ;
        RECT 445.625000 146.850000 480.000000 147.000000 ;
        RECT 445.775000 146.700000 480.000000 146.850000 ;
        RECT 445.925000 146.550000 480.000000 146.700000 ;
        RECT 446.075000 146.400000 480.000000 146.550000 ;
        RECT 446.225000 146.250000 480.000000 146.400000 ;
        RECT 446.375000 146.100000 480.000000 146.250000 ;
        RECT 446.525000 145.950000 480.000000 146.100000 ;
        RECT 446.675000 145.800000 480.000000 145.950000 ;
        RECT 446.825000 145.650000 480.000000 145.800000 ;
        RECT 446.975000 145.500000 480.000000 145.650000 ;
        RECT 447.125000 145.350000 480.000000 145.500000 ;
        RECT 447.275000 145.200000 480.000000 145.350000 ;
        RECT 447.425000 145.050000 480.000000 145.200000 ;
        RECT 447.575000 144.900000 480.000000 145.050000 ;
        RECT 447.725000 144.750000 480.000000 144.900000 ;
        RECT 447.875000 144.600000 480.000000 144.750000 ;
        RECT 448.025000 144.450000 480.000000 144.600000 ;
        RECT 448.175000 144.300000 480.000000 144.450000 ;
        RECT 448.325000 144.150000 480.000000 144.300000 ;
        RECT 448.475000 144.000000 480.000000 144.150000 ;
        RECT 448.625000 143.850000 480.000000 144.000000 ;
        RECT 448.775000 143.700000 480.000000 143.850000 ;
        RECT 448.925000 143.550000 480.000000 143.700000 ;
        RECT 449.075000 143.400000 480.000000 143.550000 ;
        RECT 449.225000 143.250000 480.000000 143.400000 ;
        RECT 449.375000 143.100000 480.000000 143.250000 ;
        RECT 449.525000 142.950000 480.000000 143.100000 ;
        RECT 449.675000 142.800000 480.000000 142.950000 ;
        RECT 449.825000 142.650000 480.000000 142.800000 ;
        RECT 449.975000 142.500000 480.000000 142.650000 ;
        RECT 450.125000 142.350000 480.000000 142.500000 ;
        RECT 450.275000 142.200000 480.000000 142.350000 ;
        RECT 450.425000 142.050000 480.000000 142.200000 ;
        RECT 450.575000 141.900000 480.000000 142.050000 ;
        RECT 450.725000 141.750000 480.000000 141.900000 ;
        RECT 450.875000 141.600000 480.000000 141.750000 ;
        RECT 451.025000 141.450000 480.000000 141.600000 ;
        RECT 451.175000 141.300000 480.000000 141.450000 ;
        RECT 451.325000 141.150000 480.000000 141.300000 ;
        RECT 451.475000 141.000000 480.000000 141.150000 ;
        RECT 451.625000 140.850000 480.000000 141.000000 ;
        RECT 451.775000 140.700000 480.000000 140.850000 ;
        RECT 451.925000 140.550000 480.000000 140.700000 ;
        RECT 452.075000 140.400000 480.000000 140.550000 ;
        RECT 452.225000 140.250000 480.000000 140.400000 ;
        RECT 452.375000 140.100000 480.000000 140.250000 ;
        RECT 452.525000 139.950000 480.000000 140.100000 ;
        RECT 452.675000 139.800000 480.000000 139.950000 ;
        RECT 452.825000 139.650000 480.000000 139.800000 ;
        RECT 452.975000 139.500000 480.000000 139.650000 ;
        RECT 453.125000 139.350000 480.000000 139.500000 ;
        RECT 453.275000 139.200000 480.000000 139.350000 ;
        RECT 453.425000 139.050000 480.000000 139.200000 ;
        RECT 453.575000 138.900000 480.000000 139.050000 ;
        RECT 453.725000 138.750000 480.000000 138.900000 ;
        RECT 453.875000 138.600000 480.000000 138.750000 ;
        RECT 454.025000 138.450000 480.000000 138.600000 ;
        RECT 454.175000 138.300000 480.000000 138.450000 ;
        RECT 454.325000 138.150000 480.000000 138.300000 ;
        RECT 454.475000 138.000000 480.000000 138.150000 ;
        RECT 454.625000 137.850000 480.000000 138.000000 ;
        RECT 454.775000 137.700000 480.000000 137.850000 ;
        RECT 454.925000 137.550000 480.000000 137.700000 ;
        RECT 455.075000 137.400000 480.000000 137.550000 ;
        RECT 455.225000 137.250000 480.000000 137.400000 ;
        RECT 455.375000 137.100000 480.000000 137.250000 ;
        RECT 455.525000 136.950000 480.000000 137.100000 ;
        RECT 455.675000 136.800000 480.000000 136.950000 ;
        RECT 455.825000 136.650000 480.000000 136.800000 ;
        RECT 455.975000 136.500000 480.000000 136.650000 ;
        RECT 456.125000 136.350000 480.000000 136.500000 ;
        RECT 456.275000 136.200000 480.000000 136.350000 ;
        RECT 456.425000 136.050000 480.000000 136.200000 ;
        RECT 456.575000 135.900000 480.000000 136.050000 ;
        RECT 456.725000 135.750000 480.000000 135.900000 ;
        RECT 456.875000 135.600000 480.000000 135.750000 ;
        RECT 457.025000 135.450000 480.000000 135.600000 ;
        RECT 457.175000 135.300000 480.000000 135.450000 ;
        RECT 457.325000 135.150000 480.000000 135.300000 ;
        RECT 457.475000 135.000000 480.000000 135.150000 ;
        RECT 457.625000 134.850000 480.000000 135.000000 ;
        RECT 457.775000 134.700000 480.000000 134.850000 ;
        RECT 457.925000 134.550000 480.000000 134.700000 ;
        RECT 458.075000 134.400000 480.000000 134.550000 ;
        RECT 458.225000 134.250000 480.000000 134.400000 ;
        RECT 458.375000 134.100000 480.000000 134.250000 ;
        RECT 458.525000 133.950000 480.000000 134.100000 ;
        RECT 458.675000 133.800000 480.000000 133.950000 ;
        RECT 458.825000 133.650000 480.000000 133.800000 ;
        RECT 458.975000 133.500000 480.000000 133.650000 ;
        RECT 459.125000 133.350000 480.000000 133.500000 ;
        RECT 459.275000 133.200000 480.000000 133.350000 ;
        RECT 459.425000 133.050000 480.000000 133.200000 ;
        RECT 459.575000 132.900000 480.000000 133.050000 ;
        RECT 459.725000 132.750000 480.000000 132.900000 ;
        RECT 459.875000 132.600000 480.000000 132.750000 ;
        RECT 460.025000 132.450000 480.000000 132.600000 ;
        RECT 460.175000 132.300000 480.000000 132.450000 ;
        RECT 460.325000 132.150000 480.000000 132.300000 ;
        RECT 460.475000 132.000000 480.000000 132.150000 ;
        RECT 460.625000 131.850000 480.000000 132.000000 ;
        RECT 460.775000 131.700000 480.000000 131.850000 ;
        RECT 460.925000 131.550000 480.000000 131.700000 ;
        RECT 461.075000 131.400000 480.000000 131.550000 ;
        RECT 461.225000 131.250000 480.000000 131.400000 ;
        RECT 461.375000 131.100000 480.000000 131.250000 ;
        RECT 461.525000 130.950000 480.000000 131.100000 ;
        RECT 461.675000 130.800000 480.000000 130.950000 ;
        RECT 461.825000 130.650000 480.000000 130.800000 ;
        RECT 461.975000 130.500000 480.000000 130.650000 ;
        RECT 462.125000 130.350000 480.000000 130.500000 ;
        RECT 462.275000 130.200000 480.000000 130.350000 ;
        RECT 462.425000 130.050000 480.000000 130.200000 ;
        RECT 462.575000 129.900000 480.000000 130.050000 ;
        RECT 462.725000 129.750000 480.000000 129.900000 ;
        RECT 462.875000 129.600000 480.000000 129.750000 ;
        RECT 463.025000 129.450000 480.000000 129.600000 ;
        RECT 463.175000 129.300000 480.000000 129.450000 ;
        RECT 463.325000 129.150000 480.000000 129.300000 ;
        RECT 463.475000 129.000000 480.000000 129.150000 ;
        RECT 463.625000 128.850000 480.000000 129.000000 ;
        RECT 463.775000 128.700000 480.000000 128.850000 ;
        RECT 463.925000 128.550000 480.000000 128.700000 ;
        RECT 464.075000 128.400000 480.000000 128.550000 ;
        RECT 464.225000 128.250000 480.000000 128.400000 ;
        RECT 464.375000 128.100000 480.000000 128.250000 ;
        RECT 464.525000 127.950000 480.000000 128.100000 ;
        RECT 464.675000 127.800000 480.000000 127.950000 ;
        RECT 464.825000 127.650000 480.000000 127.800000 ;
        RECT 464.975000 127.500000 480.000000 127.650000 ;
        RECT 465.125000 127.350000 480.000000 127.500000 ;
        RECT 465.275000 127.200000 480.000000 127.350000 ;
        RECT 465.425000 127.050000 480.000000 127.200000 ;
        RECT 465.575000 126.900000 480.000000 127.050000 ;
        RECT 465.725000 126.750000 480.000000 126.900000 ;
        RECT 465.875000 126.600000 480.000000 126.750000 ;
        RECT 466.025000 126.450000 480.000000 126.600000 ;
        RECT 466.175000 126.300000 480.000000 126.450000 ;
        RECT 466.325000 126.150000 480.000000 126.300000 ;
        RECT 466.475000 126.000000 480.000000 126.150000 ;
        RECT 466.625000 125.850000 480.000000 126.000000 ;
        RECT 466.775000 125.700000 480.000000 125.850000 ;
        RECT 466.925000 125.550000 480.000000 125.700000 ;
        RECT 467.075000 125.400000 480.000000 125.550000 ;
        RECT 467.225000 125.250000 480.000000 125.400000 ;
        RECT 467.375000 125.100000 480.000000 125.250000 ;
        RECT 467.525000 124.950000 480.000000 125.100000 ;
        RECT 467.675000 124.800000 480.000000 124.950000 ;
        RECT 467.825000 124.650000 480.000000 124.800000 ;
        RECT 467.975000 124.500000 480.000000 124.650000 ;
        RECT 468.125000 124.350000 480.000000 124.500000 ;
        RECT 468.275000 124.200000 480.000000 124.350000 ;
        RECT 468.425000 124.050000 480.000000 124.200000 ;
        RECT 468.575000 123.900000 480.000000 124.050000 ;
        RECT 468.725000 123.750000 480.000000 123.900000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 73.500000 480.000000 78.150000 ;
        RECT 9.585000 73.495000 458.005000 73.500000 ;
        RECT 9.625000 73.455000 457.965000 73.495000 ;
        RECT 9.665000 73.415000 457.925000 73.455000 ;
    END
    PORT
      LAYER met5 ;
        RECT   0.000000 123.750000  28.815000 124.150000 ;
        RECT   0.000000 124.150000  29.215000 124.550000 ;
        RECT   0.000000 124.550000  29.615000 124.950000 ;
        RECT   0.000000 124.950000  30.015000 125.350000 ;
        RECT   0.000000 125.350000  30.415000 125.750000 ;
        RECT   0.000000 125.750000  30.815000 126.150000 ;
        RECT   0.000000 126.150000  31.215000 126.550000 ;
        RECT   0.000000 126.550000  31.615000 126.950000 ;
        RECT   0.000000 126.950000  32.015000 127.350000 ;
        RECT   0.000000 127.350000  32.415000 127.750000 ;
        RECT   0.000000 127.750000  32.815000 128.150000 ;
        RECT   0.000000 128.150000  33.215000 128.550000 ;
        RECT   0.000000 128.550000  33.615000 128.950000 ;
        RECT   0.000000 128.950000  34.015000 129.350000 ;
        RECT   0.000000 129.350000  34.415000 129.750000 ;
        RECT   0.000000 129.750000  34.815000 130.150000 ;
        RECT   0.000000 130.150000  35.215000 130.550000 ;
        RECT   0.000000 130.550000  35.615000 130.950000 ;
        RECT   0.000000 130.950000  36.015000 131.350000 ;
        RECT   0.000000 131.350000  36.415000 131.750000 ;
        RECT   0.000000 131.750000  36.815000 132.150000 ;
        RECT   0.000000 132.150000  37.215000 132.550000 ;
        RECT   0.000000 132.550000  37.615000 132.950000 ;
        RECT   0.000000 132.950000  38.015000 133.350000 ;
        RECT   0.000000 133.350000  38.480000 133.415000 ;
        RECT   0.000000 133.415000  38.480000 133.815000 ;
        RECT   0.000000 133.815000  38.880000 134.215000 ;
        RECT   0.000000 134.215000  39.280000 134.615000 ;
        RECT   0.000000 134.615000  39.680000 135.015000 ;
        RECT   0.000000 135.015000  40.080000 135.415000 ;
        RECT   0.000000 135.415000  40.480000 135.815000 ;
        RECT   0.000000 135.815000  40.880000 136.215000 ;
        RECT   0.000000 136.215000  41.280000 136.615000 ;
        RECT   0.000000 136.615000  41.680000 137.015000 ;
        RECT   0.000000 137.015000  42.080000 137.415000 ;
        RECT   0.000000 137.415000  42.480000 137.815000 ;
        RECT   0.000000 137.815000  42.880000 138.215000 ;
        RECT   0.000000 138.215000  43.280000 138.615000 ;
        RECT   0.000000 138.615000  43.680000 139.015000 ;
        RECT   0.000000 139.015000  44.080000 139.415000 ;
        RECT   0.000000 139.415000  44.480000 139.815000 ;
        RECT   0.000000 139.815000  44.880000 140.215000 ;
        RECT   0.000000 140.215000  45.280000 140.615000 ;
        RECT   0.000000 140.615000  45.680000 141.015000 ;
        RECT   0.000000 141.015000  46.080000 141.415000 ;
        RECT   0.000000 141.415000  46.480000 141.815000 ;
        RECT   0.000000 141.815000  46.880000 142.215000 ;
        RECT   0.000000 142.215000  47.280000 142.615000 ;
        RECT   0.000000 142.615000  47.680000 143.015000 ;
        RECT   0.000000 143.015000  48.080000 143.415000 ;
        RECT   0.000000 143.415000  48.480000 143.815000 ;
        RECT   0.000000 143.815000  48.880000 144.215000 ;
        RECT   0.000000 144.215000  49.280000 144.615000 ;
        RECT   0.000000 144.615000  49.680000 145.015000 ;
        RECT   0.000000 145.015000  50.080000 145.415000 ;
        RECT   0.000000 145.415000  50.480000 145.815000 ;
        RECT   0.000000 145.815000  50.880000 145.905000 ;
        RECT   0.000000 145.905000  50.990000 145.925000 ;
        RECT   0.000000 145.925000  50.990000 146.325000 ;
        RECT   0.000000 146.325000  51.390000 146.725000 ;
        RECT   0.000000 146.725000  51.790000 147.125000 ;
        RECT   0.000000 147.125000  52.190000 147.525000 ;
        RECT   0.000000 147.525000  52.590000 147.925000 ;
        RECT   0.000000 147.925000  52.990000 148.325000 ;
        RECT   0.000000 148.325000  53.390000 148.715000 ;
        RECT  18.770000 148.715000  53.780000 148.895000 ;
        RECT  18.950000 148.895000  53.960000 149.075000 ;
        RECT  18.955000 149.075000  54.140000 149.080000 ;
        RECT  19.355000 149.080000  54.145000 149.480000 ;
        RECT  19.755000 149.480000  54.145000 149.880000 ;
        RECT  20.155000 149.880000  54.145000 150.280000 ;
        RECT  20.555000 150.280000  54.145000 150.680000 ;
        RECT  20.955000 150.680000  54.145000 151.080000 ;
        RECT  21.355000 151.080000  54.145000 151.480000 ;
        RECT  21.755000 151.480000  54.145000 151.880000 ;
        RECT  22.155000 151.880000  54.145000 152.280000 ;
        RECT  22.555000 152.280000  54.145000 152.680000 ;
        RECT  22.955000 152.680000  54.145000 153.080000 ;
        RECT  23.355000 153.080000  54.145000 153.480000 ;
        RECT  23.755000 153.480000  54.145000 153.880000 ;
        RECT  24.155000 153.880000  54.145000 154.280000 ;
        RECT  24.555000 154.280000  54.145000 154.680000 ;
        RECT  24.955000 154.680000  54.145000 155.080000 ;
        RECT  25.355000 155.080000  54.145000 155.480000 ;
        RECT  25.755000 155.480000  54.145000 155.880000 ;
        RECT  26.155000 155.880000  54.145000 156.280000 ;
        RECT  26.555000 156.280000  54.145000 156.680000 ;
        RECT  26.955000 156.680000  54.145000 157.080000 ;
        RECT  27.355000 157.080000  54.145000 157.480000 ;
        RECT  27.755000 157.480000  54.145000 157.880000 ;
        RECT  28.155000 157.880000  54.145000 158.280000 ;
        RECT  28.555000 158.280000  54.145000 158.680000 ;
        RECT  28.955000 158.680000  54.145000 159.080000 ;
        RECT  29.260000 159.080000  54.145000 159.385000 ;
        RECT  29.260000 159.385000  54.145000 197.600000 ;
        RECT  29.260000 197.600000  54.145000 198.000000 ;
        RECT  29.260000 198.000000  54.545000 198.400000 ;
        RECT  29.260000 198.400000  54.945000 198.800000 ;
        RECT  29.260000 198.800000  55.345000 199.200000 ;
        RECT  29.260000 199.200000  55.745000 199.600000 ;
        RECT  29.260000 199.600000  56.145000 200.000000 ;
        RECT  29.260000 200.000000  56.545000 200.400000 ;
        RECT  29.260000 200.400000  56.945000 200.800000 ;
        RECT  29.260000 200.800000  57.345000 201.200000 ;
        RECT  29.260000 201.200000  57.745000 201.600000 ;
        RECT  29.260000 201.600000  58.145000 202.000000 ;
        RECT  29.260000 202.000000  58.545000 202.400000 ;
        RECT  29.260000 202.400000  58.945000 202.800000 ;
        RECT  29.260000 202.800000  59.345000 203.200000 ;
        RECT  29.260000 203.200000  59.745000 203.600000 ;
        RECT  29.260000 203.600000  60.145000 204.000000 ;
        RECT  29.260000 204.000000  60.545000 204.400000 ;
        RECT  29.260000 204.400000  60.945000 204.490000 ;
        RECT  29.260000 204.490000 422.295000 204.890000 ;
        RECT  29.260000 204.890000 421.895000 205.290000 ;
        RECT  29.260000 205.290000 421.495000 205.690000 ;
        RECT  29.260000 205.690000 421.095000 206.090000 ;
        RECT  29.260000 206.090000 420.695000 206.490000 ;
        RECT  29.260000 206.490000 420.295000 206.890000 ;
        RECT  29.260000 206.890000 419.895000 207.290000 ;
        RECT  29.260000 207.290000 419.860000 207.325000 ;
        RECT  29.660000 207.325000 419.460000 207.725000 ;
        RECT  30.060000 207.725000 419.060000 208.125000 ;
        RECT  30.460000 208.125000 418.660000 208.525000 ;
        RECT  30.860000 208.525000 418.260000 208.925000 ;
        RECT  31.260000 208.925000 417.860000 209.325000 ;
        RECT  31.660000 209.325000 417.460000 209.725000 ;
        RECT  32.060000 209.725000 417.060000 210.125000 ;
        RECT  32.460000 210.125000 416.660000 210.525000 ;
        RECT  32.860000 210.525000 416.260000 210.925000 ;
        RECT  33.260000 210.925000 415.860000 211.325000 ;
        RECT  33.660000 211.325000 415.460000 211.725000 ;
        RECT  34.060000 211.725000 415.060000 212.125000 ;
        RECT  34.460000 212.125000 414.660000 212.525000 ;
        RECT  34.860000 212.525000 414.260000 212.925000 ;
        RECT  35.260000 212.925000 413.860000 213.325000 ;
        RECT  35.660000 213.325000 413.460000 213.725000 ;
        RECT  36.060000 213.725000 413.060000 214.125000 ;
        RECT  36.460000 214.125000 412.660000 214.525000 ;
        RECT  36.860000 214.525000 412.260000 214.925000 ;
        RECT  37.260000 214.925000 411.860000 215.325000 ;
        RECT  37.660000 215.325000 411.460000 215.725000 ;
        RECT  38.060000 215.725000 411.060000 216.125000 ;
        RECT  38.460000 216.125000 410.660000 216.525000 ;
        RECT  38.860000 216.525000 410.260000 216.925000 ;
        RECT  39.260000 216.925000 409.860000 217.325000 ;
        RECT  39.660000 217.325000 409.460000 217.725000 ;
        RECT  40.060000 217.725000 409.060000 218.125000 ;
        RECT  40.460000 218.125000 408.660000 218.525000 ;
        RECT  40.860000 218.525000 408.260000 218.925000 ;
        RECT  41.260000 218.925000 407.860000 219.325000 ;
        RECT  41.660000 219.325000 407.460000 219.725000 ;
        RECT  42.060000 219.725000 407.060000 220.125000 ;
        RECT  42.460000 220.125000 406.660000 220.525000 ;
        RECT  42.860000 220.525000 406.260000 220.925000 ;
        RECT  43.260000 220.925000 405.860000 221.325000 ;
        RECT  43.660000 221.325000 405.460000 221.725000 ;
        RECT  44.060000 221.725000 405.060000 222.125000 ;
        RECT  44.460000 222.125000 404.660000 222.525000 ;
        RECT  44.860000 222.525000 404.260000 222.925000 ;
        RECT  45.260000 222.925000 403.860000 223.325000 ;
        RECT  45.660000 223.325000 403.460000 223.725000 ;
        RECT  46.060000 223.725000 403.060000 224.125000 ;
        RECT  46.460000 224.125000 402.660000 224.525000 ;
        RECT  46.860000 224.525000 402.260000 224.925000 ;
        RECT  47.260000 224.925000 401.860000 225.325000 ;
        RECT  47.660000 225.325000 401.460000 225.725000 ;
        RECT  48.060000 225.725000 401.060000 226.125000 ;
        RECT  48.460000 226.125000 400.660000 226.525000 ;
        RECT  48.860000 226.525000 400.260000 226.925000 ;
        RECT  49.260000 226.925000 399.860000 227.325000 ;
        RECT  49.660000 227.325000 399.460000 227.725000 ;
        RECT  49.835000 227.725000 399.285000 227.900000 ;
        RECT 388.290000 204.170000 422.695000 204.490000 ;
        RECT 388.690000 203.770000 423.015000 204.170000 ;
        RECT 389.090000 203.370000 423.415000 203.770000 ;
        RECT 389.490000 202.970000 423.815000 203.370000 ;
        RECT 389.890000 202.570000 424.215000 202.970000 ;
        RECT 390.290000 202.170000 424.615000 202.570000 ;
        RECT 390.690000 201.770000 425.015000 202.170000 ;
        RECT 391.090000 201.370000 425.415000 201.770000 ;
        RECT 391.490000 200.970000 425.815000 201.370000 ;
        RECT 391.890000 200.570000 426.215000 200.970000 ;
        RECT 392.290000 200.170000 426.615000 200.570000 ;
        RECT 392.690000 199.770000 427.015000 200.170000 ;
        RECT 393.090000 199.370000 427.415000 199.770000 ;
        RECT 393.490000 198.970000 427.815000 199.370000 ;
        RECT 393.890000 198.570000 428.215000 198.970000 ;
        RECT 394.290000 198.170000 428.615000 198.570000 ;
        RECT 394.690000 197.770000 429.015000 198.170000 ;
        RECT 395.090000 197.370000 429.415000 197.770000 ;
        RECT 395.490000 196.970000 429.815000 197.370000 ;
        RECT 395.890000 196.570000 430.215000 196.970000 ;
        RECT 396.290000 196.170000 430.615000 196.570000 ;
        RECT 396.690000 195.770000 431.015000 196.170000 ;
        RECT 397.090000 195.370000 431.415000 195.770000 ;
        RECT 397.490000 194.970000 431.815000 195.370000 ;
        RECT 397.890000 194.570000 432.215000 194.970000 ;
        RECT 398.290000 194.170000 432.615000 194.570000 ;
        RECT 398.690000 193.770000 433.015000 194.170000 ;
        RECT 399.090000 193.370000 433.415000 193.770000 ;
        RECT 399.490000 192.970000 433.815000 193.370000 ;
        RECT 399.890000 192.570000 434.215000 192.970000 ;
        RECT 400.290000 192.170000 434.615000 192.570000 ;
        RECT 400.690000 191.770000 435.015000 192.170000 ;
        RECT 401.090000 191.370000 435.415000 191.770000 ;
        RECT 401.490000 190.970000 435.815000 191.370000 ;
        RECT 401.890000 190.570000 436.215000 190.970000 ;
        RECT 402.290000 190.170000 436.615000 190.570000 ;
        RECT 402.690000 189.770000 437.015000 190.170000 ;
        RECT 403.090000 189.370000 437.415000 189.770000 ;
        RECT 403.490000 188.970000 437.815000 189.370000 ;
        RECT 403.890000 188.570000 438.215000 188.970000 ;
        RECT 404.290000 188.170000 438.615000 188.570000 ;
        RECT 404.690000 187.770000 439.015000 188.170000 ;
        RECT 405.090000 187.370000 439.415000 187.770000 ;
        RECT 405.490000 186.970000 439.815000 187.370000 ;
        RECT 405.890000 186.570000 440.215000 186.970000 ;
        RECT 406.290000 186.170000 440.615000 186.570000 ;
        RECT 406.690000 185.770000 441.015000 186.170000 ;
        RECT 407.090000 185.370000 441.415000 185.770000 ;
        RECT 407.490000 184.970000 441.815000 185.370000 ;
        RECT 407.890000 184.570000 442.215000 184.970000 ;
        RECT 408.290000 184.170000 442.615000 184.570000 ;
        RECT 408.690000 183.770000 443.015000 184.170000 ;
        RECT 409.090000 183.370000 443.415000 183.770000 ;
        RECT 409.490000 182.970000 443.815000 183.370000 ;
        RECT 409.890000 182.570000 444.215000 182.970000 ;
        RECT 410.290000 182.170000 444.615000 182.570000 ;
        RECT 410.690000 181.770000 445.015000 182.170000 ;
        RECT 411.090000 181.370000 445.415000 181.770000 ;
        RECT 411.490000 180.970000 445.815000 181.370000 ;
        RECT 411.890000 180.570000 446.215000 180.970000 ;
        RECT 412.290000 180.170000 446.615000 180.570000 ;
        RECT 412.690000 179.770000 447.015000 180.170000 ;
        RECT 413.090000 179.370000 447.415000 179.770000 ;
        RECT 413.490000 178.970000 447.815000 179.370000 ;
        RECT 413.890000 178.570000 448.215000 178.970000 ;
        RECT 414.290000 178.170000 448.615000 178.570000 ;
        RECT 414.690000 177.770000 449.015000 178.170000 ;
        RECT 415.090000 177.370000 449.415000 177.770000 ;
        RECT 415.490000 176.970000 449.815000 177.370000 ;
        RECT 415.890000 176.570000 450.215000 176.970000 ;
        RECT 416.290000 176.170000 450.615000 176.570000 ;
        RECT 416.690000 175.770000 451.015000 176.170000 ;
        RECT 417.090000 175.370000 451.415000 175.770000 ;
        RECT 417.490000 174.970000 451.815000 175.370000 ;
        RECT 417.890000 174.570000 452.215000 174.970000 ;
        RECT 418.290000 174.170000 452.615000 174.570000 ;
        RECT 418.690000 173.770000 453.015000 174.170000 ;
        RECT 419.090000 173.370000 453.415000 173.770000 ;
        RECT 419.490000 172.970000 453.815000 173.370000 ;
        RECT 419.890000 172.570000 454.215000 172.970000 ;
        RECT 420.290000 172.170000 454.615000 172.570000 ;
        RECT 420.690000 171.770000 455.015000 172.170000 ;
        RECT 421.090000 171.370000 455.415000 171.770000 ;
        RECT 421.490000 170.970000 455.815000 171.370000 ;
        RECT 421.890000 170.570000 456.215000 170.970000 ;
        RECT 422.290000 170.170000 456.615000 170.570000 ;
        RECT 422.690000 169.770000 457.015000 170.170000 ;
        RECT 423.090000 169.370000 457.415000 169.770000 ;
        RECT 423.490000 168.970000 457.815000 169.370000 ;
        RECT 423.890000 168.570000 458.215000 168.970000 ;
        RECT 424.290000 168.170000 458.615000 168.570000 ;
        RECT 424.690000 167.770000 459.015000 168.170000 ;
        RECT 425.090000 167.370000 459.415000 167.770000 ;
        RECT 425.490000 166.970000 459.815000 167.370000 ;
        RECT 425.890000 166.570000 460.215000 166.970000 ;
        RECT 426.290000 166.170000 460.615000 166.570000 ;
        RECT 426.690000 165.770000 461.015000 166.170000 ;
        RECT 427.090000 165.370000 461.415000 165.770000 ;
        RECT 427.490000 164.970000 461.815000 165.370000 ;
        RECT 427.890000 164.570000 462.215000 164.970000 ;
        RECT 428.290000 164.170000 462.615000 164.570000 ;
        RECT 428.690000 163.770000 463.015000 164.170000 ;
        RECT 429.090000 163.370000 463.415000 163.770000 ;
        RECT 429.490000 162.970000 463.815000 163.370000 ;
        RECT 429.890000 162.570000 464.215000 162.970000 ;
        RECT 430.290000 162.170000 464.615000 162.570000 ;
        RECT 430.690000 161.770000 465.015000 162.170000 ;
        RECT 431.090000 161.370000 465.415000 161.770000 ;
        RECT 431.490000 160.970000 465.815000 161.370000 ;
        RECT 431.890000 160.570000 466.215000 160.970000 ;
        RECT 432.290000 160.170000 466.615000 160.570000 ;
        RECT 432.690000 159.770000 467.015000 160.170000 ;
        RECT 433.090000 159.370000 467.415000 159.770000 ;
        RECT 433.490000 158.970000 467.815000 159.370000 ;
        RECT 433.890000 158.570000 468.215000 158.970000 ;
        RECT 434.290000 158.170000 468.615000 158.570000 ;
        RECT 434.690000 157.770000 469.015000 158.170000 ;
        RECT 435.090000 157.370000 469.415000 157.770000 ;
        RECT 435.490000 156.970000 469.815000 157.370000 ;
        RECT 435.890000 156.570000 470.215000 156.970000 ;
        RECT 436.290000 156.170000 470.615000 156.570000 ;
        RECT 436.690000 155.770000 471.015000 156.170000 ;
        RECT 437.090000 155.370000 471.415000 155.770000 ;
        RECT 437.490000 154.970000 471.815000 155.370000 ;
        RECT 437.890000 154.570000 472.215000 154.970000 ;
        RECT 438.290000 154.170000 472.615000 154.570000 ;
        RECT 438.690000 153.770000 473.015000 154.170000 ;
        RECT 439.090000 153.370000 473.415000 153.770000 ;
        RECT 439.490000 152.970000 473.815000 153.370000 ;
        RECT 439.890000 152.570000 474.215000 152.970000 ;
        RECT 440.290000 152.170000 474.615000 152.570000 ;
        RECT 440.690000 151.750000 475.425000 151.760000 ;
        RECT 440.690000 151.760000 475.415000 151.770000 ;
        RECT 440.690000 151.770000 475.015000 152.170000 ;
        RECT 440.960000 151.500000 475.435000 151.750000 ;
        RECT 441.360000 151.100000 475.685000 151.500000 ;
        RECT 441.760000 150.700000 476.085000 151.100000 ;
        RECT 442.160000 150.300000 476.485000 150.700000 ;
        RECT 442.560000 149.900000 476.885000 150.300000 ;
        RECT 442.960000 149.500000 477.285000 149.900000 ;
        RECT 443.360000 149.100000 477.685000 149.500000 ;
        RECT 443.760000 148.700000 478.085000 149.100000 ;
        RECT 444.090000 148.370000 480.000000 148.700000 ;
        RECT 444.490000 147.970000 480.000000 148.370000 ;
        RECT 444.890000 147.570000 480.000000 147.970000 ;
        RECT 445.290000 147.170000 480.000000 147.570000 ;
        RECT 445.690000 146.770000 480.000000 147.170000 ;
        RECT 446.090000 146.370000 480.000000 146.770000 ;
        RECT 446.490000 145.970000 480.000000 146.370000 ;
        RECT 446.890000 145.510000 480.000000 145.570000 ;
        RECT 446.890000 145.570000 480.000000 145.970000 ;
        RECT 447.110000 145.350000 480.000000 145.510000 ;
        RECT 447.510000 144.950000 480.000000 145.350000 ;
        RECT 447.910000 144.550000 480.000000 144.950000 ;
        RECT 448.310000 144.150000 480.000000 144.550000 ;
        RECT 448.710000 143.750000 480.000000 144.150000 ;
        RECT 449.110000 143.350000 480.000000 143.750000 ;
        RECT 449.510000 142.950000 480.000000 143.350000 ;
        RECT 449.910000 142.550000 480.000000 142.950000 ;
        RECT 450.310000 142.150000 480.000000 142.550000 ;
        RECT 450.710000 141.750000 480.000000 142.150000 ;
        RECT 451.110000 141.350000 480.000000 141.750000 ;
        RECT 451.510000 140.950000 480.000000 141.350000 ;
        RECT 451.910000 140.550000 480.000000 140.950000 ;
        RECT 452.310000 140.150000 480.000000 140.550000 ;
        RECT 452.710000 139.750000 480.000000 140.150000 ;
        RECT 453.110000 139.350000 480.000000 139.750000 ;
        RECT 453.510000 138.950000 480.000000 139.350000 ;
        RECT 453.910000 138.550000 480.000000 138.950000 ;
        RECT 454.310000 138.150000 480.000000 138.550000 ;
        RECT 454.710000 137.750000 480.000000 138.150000 ;
        RECT 455.110000 137.350000 480.000000 137.750000 ;
        RECT 455.510000 136.950000 480.000000 137.350000 ;
        RECT 455.910000 136.550000 480.000000 136.950000 ;
        RECT 456.310000 136.150000 480.000000 136.550000 ;
        RECT 456.710000 135.750000 480.000000 136.150000 ;
        RECT 457.110000 135.350000 480.000000 135.750000 ;
        RECT 457.510000 134.950000 480.000000 135.350000 ;
        RECT 457.910000 134.550000 480.000000 134.950000 ;
        RECT 458.310000 134.150000 480.000000 134.550000 ;
        RECT 458.710000 133.750000 480.000000 134.150000 ;
        RECT 459.110000 133.350000 480.000000 133.750000 ;
        RECT 459.510000 132.950000 480.000000 133.350000 ;
        RECT 459.910000 132.550000 480.000000 132.950000 ;
        RECT 460.310000 132.150000 480.000000 132.550000 ;
        RECT 460.710000 131.750000 480.000000 132.150000 ;
        RECT 461.110000 131.350000 480.000000 131.750000 ;
        RECT 461.510000 130.950000 480.000000 131.350000 ;
        RECT 461.910000 130.550000 480.000000 130.950000 ;
        RECT 462.310000 130.150000 480.000000 130.550000 ;
        RECT 462.710000 129.750000 480.000000 130.150000 ;
        RECT 463.110000 129.350000 480.000000 129.750000 ;
        RECT 463.510000 128.950000 480.000000 129.350000 ;
        RECT 463.910000 128.550000 480.000000 128.950000 ;
        RECT 464.310000 128.150000 480.000000 128.550000 ;
        RECT 464.710000 127.750000 480.000000 128.150000 ;
        RECT 465.110000 127.350000 480.000000 127.750000 ;
        RECT 465.510000 126.950000 480.000000 127.350000 ;
        RECT 465.910000 126.550000 480.000000 126.950000 ;
        RECT 466.310000 126.150000 480.000000 126.550000 ;
        RECT 466.710000 125.750000 480.000000 126.150000 ;
        RECT 467.110000 125.350000 480.000000 125.750000 ;
        RECT 467.510000 124.950000 480.000000 125.350000 ;
        RECT 467.910000 124.550000 480.000000 124.950000 ;
        RECT 468.310000 124.150000 480.000000 124.550000 ;
        RECT 468.710000 123.750000 480.000000 124.150000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 73.600000 480.000000 78.050000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 117.800000 480.000000 122.250000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 117.900000 480.000000 122.150000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 101.450000 480.000000 101.780000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 105.360000 480.000000 106.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 110.120000 480.000000 110.450000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 90.450000 480.000000 93.900000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 101.450000 480.000000 110.450000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 90.550000 480.000000 93.800000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 95.300000 480.000000 99.950000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 95.400000 480.000000 99.850000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 229.500000 480.000000 253.715000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 79.550000 480.000000 84.200000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 229.500000 480.000000 253.715000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 79.650000 480.000000 84.100000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 111.950000 480.000000 116.400000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 112.050000 480.000000 116.300000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 85.600000 480.000000 89.050000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 85.700000 480.000000 88.950000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT   1.120000   0.335000   9.380000  17.505000 ;
      RECT   1.130000  17.505000  10.440000  40.640000 ;
      RECT   1.130000  40.640000   7.130000 187.555000 ;
      RECT   1.175000 187.555000  19.475000 195.580000 ;
      RECT   1.175000 195.580000  40.820000 202.710000 ;
      RECT   1.175000 202.710000  16.405000 227.215000 ;
      RECT   1.175000 227.215000  24.380000 250.140000 ;
      RECT   1.175000 250.140000  40.820000 253.385000 ;
      RECT   7.780000  41.695000  11.680000  41.725000 ;
      RECT   7.780000  41.725000  14.480000  41.895000 ;
      RECT   7.780000  41.895000  11.680000  41.925000 ;
      RECT   7.780000  41.925000   8.010000 184.540000 ;
      RECT   7.780000 184.540000  17.240000 184.770000 ;
      RECT   8.455000  65.275000   8.870000  65.865000 ;
      RECT   9.350000  65.275000   9.680000  65.865000 ;
      RECT  10.160000 136.140000  10.490000 136.730000 ;
      RECT  10.160000 182.950000  10.490000 183.540000 ;
      RECT  10.900000   2.965000  29.245000   3.135000 ;
      RECT  10.900000   3.135000  11.070000  16.245000 ;
      RECT  10.900000  16.245000  29.245000  16.415000 ;
      RECT  10.970000 182.950000  11.300000 183.550000 ;
      RECT  11.780000 182.950000  12.110000 183.550000 ;
      RECT  11.830000   3.905000  14.340000   4.075000 ;
      RECT  11.830000   4.075000  12.000000  15.315000 ;
      RECT  11.830000  15.315000  14.340000  15.485000 ;
      RECT  12.410000   4.675000  12.580000  14.565000 ;
      RECT  12.590000 182.950000  12.920000 183.550000 ;
      RECT  12.635000   4.315000  13.535000   4.485000 ;
      RECT  12.635000  14.905000  13.945000  15.075000 ;
      RECT  12.700000  17.350000  14.720000  18.100000 ;
      RECT  12.700000  27.930000  14.720000  28.680000 ;
      RECT  12.750000   4.485000  13.420000  14.905000 ;
      RECT  13.400000 182.950000  13.730000 183.550000 ;
      RECT  13.590000   4.675000  13.760000  14.525000 ;
      RECT  14.170000   4.075000  14.340000  15.315000 ;
      RECT  14.210000  43.425000  14.540000  44.015000 ;
      RECT  14.210000 182.950000  14.540000 183.555000 ;
      RECT  14.310000  41.895000  14.480000  42.790000 ;
      RECT  14.310000  42.790000  15.270000  42.960000 ;
      RECT  14.665000  29.675000  24.335000  29.845000 ;
      RECT  14.665000  29.845000  21.100000  29.880000 ;
      RECT  14.665000  29.880000  14.835000  35.050000 ;
      RECT  14.665000  35.050000  21.100000  36.400000 ;
      RECT  14.665000  36.400000  14.835000  41.570000 ;
      RECT  14.665000  41.570000  21.100000  41.605000 ;
      RECT  14.665000  41.605000  24.335000  41.775000 ;
      RECT  15.100000   3.135000  29.245000   3.665000 ;
      RECT  15.100000   3.665000  16.055000  13.725000 ;
      RECT  15.100000  13.725000  29.245000  14.425000 ;
      RECT  15.100000  14.425000  15.270000  16.045000 ;
      RECT  15.100000  16.045000  29.245000  16.245000 ;
      RECT  15.100000  42.960000  15.270000  53.700000 ;
      RECT  15.100000  53.700000  17.210000  53.870000 ;
      RECT  15.140000  54.165000  15.790000  56.710000 ;
      RECT  15.140000  56.710000  15.670000  58.050000 ;
      RECT  15.355000  16.415000  29.245000  16.745000 ;
      RECT  15.355000  16.745000  16.055000  26.805000 ;
      RECT  15.355000  26.805000  29.245000  27.505000 ;
      RECT  15.600000  30.645000  19.570000  30.815000 ;
      RECT  15.600000  30.815000  15.770000  34.085000 ;
      RECT  15.600000  37.365000  15.770000  40.635000 ;
      RECT  15.600000  40.635000  19.515000  40.805000 ;
      RECT  15.685000  41.775000  16.020000  42.710000 ;
      RECT  15.850000  42.710000  16.020000  53.095000 ;
      RECT  15.850000  53.095000  24.335000  53.265000 ;
      RECT  16.045000  34.345000  18.730000  34.515000 ;
      RECT  16.045000  36.935000  18.730000  37.105000 ;
      RECT  16.080000  31.065000  16.250000  33.775000 ;
      RECT  16.080000  37.675000  16.250000  40.385000 ;
      RECT  16.150000  56.710000  16.480000  58.300000 ;
      RECT  16.430000  42.415000  16.600000  52.305000 ;
      RECT  16.470000  34.325000  17.140000  34.345000 ;
      RECT  16.470000  37.105000  17.140000  37.125000 ;
      RECT  16.655000  42.025000  17.780000  42.195000 ;
      RECT  16.655000  52.675000  17.780000  52.845000 ;
      RECT  16.815000   4.425000  21.190000   5.135000 ;
      RECT  16.815000   5.135000  17.515000  12.265000 ;
      RECT  16.815000  12.265000  21.190000  12.965000 ;
      RECT  16.815000  17.505000  21.190000  18.205000 ;
      RECT  16.815000  18.205000  17.515000  25.335000 ;
      RECT  16.815000  25.335000  21.190000  26.045000 ;
      RECT  17.010000  82.505000  17.240000 184.540000 ;
      RECT  17.040000  53.870000  17.210000  82.505000 ;
      RECT  17.360000  31.065000  17.530000  33.775000 ;
      RECT  17.360000  37.675000  17.530000  40.385000 ;
      RECT  17.610000  42.195000  17.780000  52.675000 ;
      RECT  17.645000 134.865000  30.945000 141.545000 ;
      RECT  17.645000 141.545000  19.675000 161.195000 ;
      RECT  17.645000 161.195000  60.940000 162.215000 ;
      RECT  17.645000 162.215000  18.775000 164.565000 ;
      RECT  17.650000  56.665000  25.215000  56.835000 ;
      RECT  17.650000  56.835000  17.820000  70.255000 ;
      RECT  17.650000  70.255000  25.215000  70.425000 ;
      RECT  17.720000  34.325000  18.730000  34.345000 ;
      RECT  17.720000  37.105000  18.730000  37.125000 ;
      RECT  17.820000  71.830000  84.585000  72.420000 ;
      RECT  17.820000  72.420000  27.645000  72.730000 ;
      RECT  17.885000  71.560000  84.585000  71.830000 ;
      RECT  17.990000   6.000000  18.530000  11.395000 ;
      RECT  17.990000  19.075000  18.530000  24.470000 ;
      RECT  18.060000 172.935000  18.680000 173.750000 ;
      RECT  18.060000 173.750000  18.965000 174.835000 ;
      RECT  18.060000 174.835000  48.865000 176.430000 ;
      RECT  18.060000 176.430000  21.780000 177.695000 ;
      RECT  18.060000 177.695000  22.280000 178.695000 ;
      RECT  18.060000 178.695000  21.780000 181.365000 ;
      RECT  18.060000 181.365000  22.490000 185.455000 ;
      RECT  18.060000 185.455000  22.205000 186.105000 ;
      RECT  18.060000 186.105000  40.820000 186.695000 ;
      RECT  18.060000 186.695000  19.475000 187.555000 ;
      RECT  18.070000 165.335000  18.580000 165.425000 ;
      RECT  18.070000 165.425000  19.065000 171.430000 ;
      RECT  18.070000 171.430000  22.745000 171.990000 ;
      RECT  18.070000 171.990000  19.065000 172.100000 ;
      RECT  18.140000  31.065000  18.310000  33.775000 ;
      RECT  18.140000  37.675000  18.310000  40.385000 ;
      RECT  18.330000  41.775000  19.340000  53.095000 ;
      RECT  18.335000   5.420000  19.660000   5.830000 ;
      RECT  18.335000  24.640000  19.660000  25.050000 ;
      RECT  18.465000  57.685000  18.635000  62.535000 ;
      RECT  18.465000  64.050000  18.635000  68.900000 ;
      RECT  18.850000  84.375000  28.260000  84.545000 ;
      RECT  18.850000  84.545000  24.180000  86.190000 ;
      RECT  18.850000  86.190000  19.020000 104.255000 ;
      RECT  18.850000 104.255000  20.190000 107.995000 ;
      RECT  18.850000 107.995000  19.020000 125.215000 ;
      RECT  18.850000 125.215000  26.295000 125.365000 ;
      RECT  18.850000 125.365000  28.290000 125.415000 ;
      RECT  18.850000 125.415000  20.160000 127.705000 ;
      RECT  18.850000 127.705000  28.290000 127.755000 ;
      RECT  18.850000 127.755000  26.295000 127.905000 ;
      RECT  18.850000 127.905000  19.020000 133.775000 ;
      RECT  18.850000 133.775000  28.260000 133.945000 ;
      RECT  18.865000 203.475000  45.520000 204.335000 ;
      RECT  18.865000 204.335000  19.725000 225.590000 ;
      RECT  18.865000 225.590000  42.430000 226.440000 ;
      RECT  18.865000 226.440000  26.000000 226.450000 ;
      RECT  18.875000  63.270000  19.545000  63.440000 ;
      RECT  18.880000 173.020000  19.050000 173.040000 ;
      RECT  18.880000 173.040000  19.565000 173.110000 ;
      RECT  18.880000 173.110000  26.240000 173.480000 ;
      RECT  18.880000 173.480000  19.565000 173.550000 ;
      RECT  18.920000  31.065000  19.090000  33.775000 ;
      RECT  18.920000  37.675000  19.090000  40.385000 ;
      RECT  19.235000 163.330000  19.565000 163.400000 ;
      RECT  19.235000 163.400000  25.975000 163.770000 ;
      RECT  19.235000 163.770000  19.565000 163.840000 ;
      RECT  19.235000 164.210000  19.565000 164.280000 ;
      RECT  19.235000 164.280000  25.975000 164.650000 ;
      RECT  19.235000 164.650000  19.565000 164.720000 ;
      RECT  19.235000 165.640000  19.565000 165.710000 ;
      RECT  19.235000 165.710000  25.975000 166.080000 ;
      RECT  19.235000 166.080000  19.565000 166.150000 ;
      RECT  19.235000 166.520000  19.565000 166.590000 ;
      RECT  19.235000 166.590000  25.975000 166.960000 ;
      RECT  19.235000 166.960000  19.565000 167.030000 ;
      RECT  19.235000 168.020000  19.565000 168.090000 ;
      RECT  19.235000 168.090000  26.485000 168.190000 ;
      RECT  19.235000 168.190000  25.975000 168.460000 ;
      RECT  19.235000 168.460000  19.565000 168.530000 ;
      RECT  19.235000 168.900000  19.565000 168.970000 ;
      RECT  19.235000 168.970000  25.975000 169.340000 ;
      RECT  19.235000 169.340000  19.565000 169.410000 ;
      RECT  19.235000 169.850000  19.565000 169.920000 ;
      RECT  19.235000 169.920000  26.315000 170.290000 ;
      RECT  19.235000 170.290000  19.565000 170.360000 ;
      RECT  19.235000 170.730000  19.565000 170.800000 ;
      RECT  19.235000 170.800000  25.975000 171.170000 ;
      RECT  19.235000 171.170000  19.565000 171.260000 ;
      RECT  19.235000 172.160000  19.565000 172.230000 ;
      RECT  19.235000 172.230000  25.975000 172.600000 ;
      RECT  19.235000 172.600000  19.565000 172.690000 ;
      RECT  19.330000  87.565000  19.500000  88.310000 ;
      RECT  19.330000  88.310000  19.530000  93.725000 ;
      RECT  19.330000  93.725000  19.500000  94.355000 ;
      RECT  19.330000 117.835000  19.500000 118.465000 ;
      RECT  19.330000 118.465000  19.530000 123.880000 ;
      RECT  19.330000 123.880000  19.500000 124.625000 ;
      RECT  19.400000  30.815000  19.570000  34.085000 ;
      RECT  19.465000   6.000000  20.005000  11.395000 ;
      RECT  19.465000  19.075000  20.005000  24.470000 ;
      RECT  19.555000  87.175000  27.555000  87.345000 ;
      RECT  19.555000  94.825000  27.555000  94.995000 ;
      RECT  19.555000 117.195000  27.555000 117.365000 ;
      RECT  19.555000 124.845000  27.555000 125.015000 ;
      RECT  19.650000  99.615000  20.600000  99.785000 ;
      RECT  19.650000  99.785000  19.820000 103.265000 ;
      RECT  19.650000 103.265000  20.600000 103.435000 ;
      RECT  19.650000 109.205000  19.820000 111.915000 ;
      RECT  19.690000 128.155000  19.860000 132.905000 ;
      RECT  19.700000  87.345000  27.440000  94.825000 ;
      RECT  19.700000 117.365000  27.440000 124.845000 ;
      RECT  19.705000 108.815000  20.375000 108.985000 ;
      RECT  19.730000 163.060000  25.475000 163.230000 ;
      RECT  19.730000 164.820000  25.475000 164.890000 ;
      RECT  19.730000 164.890000  26.485000 165.060000 ;
      RECT  19.730000 165.370000  25.475000 165.540000 ;
      RECT  19.730000 167.130000  25.475000 167.300000 ;
      RECT  19.730000 167.680000  22.745000 167.850000 ;
      RECT  19.730000 170.460000  25.350000 170.630000 ;
      RECT  19.730000 172.770000  25.350000 172.940000 ;
      RECT  19.745000  57.685000  19.915000  62.535000 ;
      RECT  19.745000  64.050000  19.915000  68.900000 ;
      RECT  19.755000 174.020000  38.150000 174.220000 ;
      RECT  19.890000  42.025000  21.015000  42.195000 ;
      RECT  19.890000  42.195000  20.060000  52.675000 ;
      RECT  19.890000  52.675000  21.015000  52.845000 ;
      RECT  19.915000 133.405000  26.615000 133.415000 ;
      RECT  19.915000 133.415000  26.675000 133.585000 ;
      RECT  19.930000 125.185000  26.295000 125.215000 ;
      RECT  19.930000 127.905000  26.295000 127.935000 ;
      RECT  19.960000 187.220000  21.200000 187.550000 ;
      RECT  20.005000 190.495000  20.255000 193.230000 ;
      RECT  20.020000 108.535000  20.190000 108.815000 ;
      RECT  20.020000 108.985000  20.190000 113.005000 ;
      RECT  20.020000 113.005000  20.845000 113.175000 ;
      RECT  20.035000 163.940000  22.745000 164.110000 ;
      RECT  20.035000 166.250000  22.745000 166.420000 ;
      RECT  20.035000 169.580000  22.745000 169.750000 ;
      RECT  20.035000 171.340000  22.745000 171.430000 ;
      RECT  20.035000 171.990000  22.745000 172.060000 ;
      RECT  20.035000 173.650000  22.745000 173.820000 ;
      RECT  20.060000 193.230000  20.230000 195.580000 ;
      RECT  20.120000  95.425000  21.070000  95.595000 ;
      RECT  20.120000  95.595000  20.290000  99.075000 ;
      RECT  20.120000  99.075000  21.070000  99.245000 ;
      RECT  20.120000 113.725000  20.290000 116.435000 ;
      RECT  20.130000  73.910000  22.520000  74.080000 ;
      RECT  20.130000  74.080000  20.300000  80.160000 ;
      RECT  20.130000  80.160000  22.520000  80.330000 ;
      RECT  20.135000  57.265000  20.805000  57.435000 ;
      RECT  20.135000  69.340000  20.805000  69.510000 ;
      RECT  20.155000  63.270000  22.105000  63.440000 ;
      RECT  20.175000 116.655000  20.845000 116.825000 ;
      RECT  20.335000  29.880000  21.100000  32.905000 ;
      RECT  20.335000  32.905000  20.505000  34.025000 ;
      RECT  20.335000  34.025000  21.100000  35.050000 ;
      RECT  20.335000  36.400000  21.100000  36.775000 ;
      RECT  20.335000  36.775000  20.505000  38.545000 ;
      RECT  20.335000  38.545000  21.100000  41.570000 ;
      RECT  20.375000 187.770000  24.525000 187.940000 ;
      RECT  20.415000 104.730000  20.585000 104.850000 ;
      RECT  20.415000 104.850000  26.235000 105.120000 ;
      RECT  20.415000 105.120000  20.585000 105.630000 ;
      RECT  20.415000 105.630000  26.235000 105.900000 ;
      RECT  20.415000 105.900000  20.585000 106.410000 ;
      RECT  20.415000 106.410000  26.235000 106.680000 ;
      RECT  20.415000 106.680000  20.585000 107.190000 ;
      RECT  20.415000 107.190000  26.235000 107.460000 ;
      RECT  20.415000 107.460000  20.585000 107.570000 ;
      RECT  20.415000 125.920000  20.585000 127.200000 ;
      RECT  20.430000  99.785000  20.600000 103.265000 ;
      RECT  20.430000 109.205000  20.600000 111.915000 ;
      RECT  20.460000 113.175000  20.630000 116.655000 ;
      RECT  20.485000 205.120000  40.820000 206.330000 ;
      RECT  20.485000 206.330000  21.690000 223.340000 ;
      RECT  20.490000   5.135000  21.190000  12.265000 ;
      RECT  20.490000  18.205000  21.190000  25.335000 ;
      RECT  20.490000 147.690000  35.590000 147.710000 ;
      RECT  20.490000 147.710000  35.650000 147.880000 ;
      RECT  20.490000 147.880000  20.660000 159.775000 ;
      RECT  20.490000 159.775000  35.650000 159.945000 ;
      RECT  20.490000 205.100000  40.820000 205.120000 ;
      RECT  20.490000 223.340000  21.690000 223.550000 ;
      RECT  20.490000 223.550000  40.820000 224.820000 ;
      RECT  20.545000 162.445000  38.050000 162.645000 ;
      RECT  20.545000 162.645000  21.135000 162.860000 ;
      RECT  20.570000 128.135000  20.740000 132.905000 ;
      RECT  20.625000 194.005000  21.635000 194.175000 ;
      RECT  20.625000 194.885000  21.635000 195.055000 ;
      RECT  20.640000 190.360000  20.810000 191.370000 ;
      RECT  20.640000 192.220000  20.810000 193.230000 ;
      RECT  20.680000 194.175000  21.525000 194.180000 ;
      RECT  20.710000  74.510000  20.880000  79.470000 ;
      RECT  20.770000  99.615000  21.880000  99.785000 ;
      RECT  20.770000 103.265000  21.880000 103.435000 ;
      RECT  20.770000 108.815000  21.880000 108.985000 ;
      RECT  20.770000 112.465000  21.880000 112.635000 ;
      RECT  20.805000 125.695000  25.555000 125.865000 ;
      RECT  20.805000 126.475000  25.555000 126.645000 ;
      RECT  20.805000 127.255000  25.555000 127.425000 ;
      RECT  20.850000  99.785000  21.460000  99.815000 ;
      RECT  20.850000 108.985000  21.460000 109.015000 ;
      RECT  20.865000 191.620000  28.865000 191.790000 ;
      RECT  20.865000 193.480000  28.865000 193.650000 ;
      RECT  20.875000 104.510000  25.845000 104.680000 ;
      RECT  20.875000 106.070000  25.845000 106.240000 ;
      RECT  20.875000 107.630000  25.845000 107.800000 ;
      RECT  20.885000 105.290000  25.845000 105.460000 ;
      RECT  20.885000 106.850000  25.845000 107.020000 ;
      RECT  20.885000 126.645000  25.475000 126.650000 ;
      RECT  20.900000  95.595000  21.070000  99.075000 ;
      RECT  20.900000 113.725000  21.070000 116.435000 ;
      RECT  20.955000  79.690000  22.180000  79.860000 ;
      RECT  21.005000 168.630000  25.475000 168.800000 ;
      RECT  21.025000  57.685000  21.195000  62.535000 ;
      RECT  21.025000  64.050000  21.195000  68.900000 ;
      RECT  21.045000 174.405000  38.520000 174.605000 ;
      RECT  21.070000  42.415000  21.240000  52.305000 ;
      RECT  21.070000 152.010000  21.240000 154.720000 ;
      RECT  21.140000 142.760000  25.440000 142.930000 ;
      RECT  21.140000 142.930000  21.310000 144.580000 ;
      RECT  21.140000 144.580000  25.440000 144.750000 ;
      RECT  21.145000 155.270000  24.535000 155.440000 ;
      RECT  21.155000  33.455000  22.635000  33.625000 ;
      RECT  21.155000  37.285000  22.155000  37.455000 ;
      RECT  21.155000  37.825000  22.635000  37.995000 ;
      RECT  21.240000  74.720000  21.410000  79.470000 ;
      RECT  21.240000  95.425000  22.010000  95.595000 ;
      RECT  21.240000  99.075000  25.850000  99.245000 ;
      RECT  21.240000 113.005000  25.850000 113.175000 ;
      RECT  21.240000 116.655000  22.010000 116.825000 ;
      RECT  21.295000  42.025000  22.420000  42.195000 ;
      RECT  21.295000  52.675000  22.420000  52.845000 ;
      RECT  21.320000  99.045000  21.930000  99.075000 ;
      RECT  21.320000 113.175000  21.930000 113.205000 ;
      RECT  21.415000  57.265000  22.085000  57.435000 ;
      RECT  21.415000  69.340000  22.085000  69.510000 ;
      RECT  21.450000 128.155000  21.620000 132.905000 ;
      RECT  21.540000  95.595000  21.710000  99.045000 ;
      RECT  21.540000 113.205000  21.710000 116.655000 ;
      RECT  21.550000 143.240000  24.300000 143.410000 ;
      RECT  21.550000 144.100000  24.300000 144.270000 ;
      RECT  21.590000 143.670000  24.300000 143.840000 ;
      RECT  21.710000  99.785000  21.880000 103.265000 ;
      RECT  21.710000 108.985000  21.880000 112.465000 ;
      RECT  21.715000  38.385000  21.980000  41.255000 ;
      RECT  21.745000  30.195000  21.980000  33.065000 ;
      RECT  21.755000  28.980000  25.065000  29.150000 ;
      RECT  21.755000  29.150000  22.285000  29.490000 ;
      RECT  21.770000  74.510000  21.940000  79.470000 ;
      RECT  21.795000 189.160000  22.325000 189.330000 ;
      RECT  21.845000 156.170000  22.015000 158.880000 ;
      RECT  21.855000 194.230000  22.025000 194.900000 ;
      RECT  21.945000 152.890000  22.120000 154.890000 ;
      RECT  21.945000 154.890000  23.880000 155.015000 ;
      RECT  21.950000   3.665000  22.650000  13.725000 ;
      RECT  21.950000  16.745000  22.650000  26.805000 ;
      RECT  21.950000 152.010000  22.120000 152.890000 ;
      RECT  21.950000 155.015000  23.880000 155.060000 ;
      RECT  21.990000 189.080000  22.160000 189.160000 ;
      RECT  21.990000 189.330000  22.160000 189.410000 ;
      RECT  22.050000  99.615000  23.160000  99.785000 ;
      RECT  22.050000 103.265000  23.160000 103.435000 ;
      RECT  22.050000 108.815000  23.160000 108.985000 ;
      RECT  22.050000 112.465000  23.160000 112.635000 ;
      RECT  22.070000 159.100000  22.740000 159.270000 ;
      RECT  22.110000 159.270000  22.640000 159.285000 ;
      RECT  22.120000 179.455000  22.290000 179.895000 ;
      RECT  22.120000 179.895000  23.310000 180.360000 ;
      RECT  22.120000 180.360000  22.870000 180.975000 ;
      RECT  22.175000 186.950000  22.705000 187.120000 ;
      RECT  22.180000  95.485000  22.350000  98.855000 ;
      RECT  22.180000 113.725000  22.350000 116.765000 ;
      RECT  22.185000 187.120000  22.465000 187.555000 ;
      RECT  22.210000  34.025000  22.380000  36.735000 ;
      RECT  22.215000 189.630000  24.215000 189.800000 ;
      RECT  22.250000  42.195000  22.420000  52.675000 ;
      RECT  22.285000 189.800000  24.155000 189.810000 ;
      RECT  22.305000  57.685000  22.475000  62.535000 ;
      RECT  22.305000  64.050000  22.475000  68.900000 ;
      RECT  22.330000 128.135000  22.500000 132.905000 ;
      RECT  22.350000  74.080000  22.520000  80.160000 ;
      RECT  22.420000 148.630000  22.590000 151.500000 ;
      RECT  22.435000  37.285000  23.435000  37.455000 ;
      RECT  22.450000 208.335000  36.680000 209.185000 ;
      RECT  22.450000 209.185000  25.000000 213.440000 ;
      RECT  22.450000 213.440000  36.680000 213.950000 ;
      RECT  22.450000 213.950000  24.145000 218.200000 ;
      RECT  22.450000 218.200000  36.680000 219.330000 ;
      RECT  22.480000 177.675000  22.780000 178.685000 ;
      RECT  22.480000 178.685000  22.740000 179.395000 ;
      RECT  22.480000 179.395000  22.990000 179.725000 ;
      RECT  22.480000 219.330000  36.680000 219.390000 ;
      RECT  22.480000 219.390000  32.945000 219.455000 ;
      RECT  22.520000  95.425000  23.290000  95.595000 ;
      RECT  22.520000 116.655000  23.290000 116.825000 ;
      RECT  22.545000  29.320000  24.705000  29.490000 ;
      RECT  22.590000  42.025000  23.375000  42.195000 ;
      RECT  22.590000  52.675000  23.375000  52.845000 ;
      RECT  22.595000  99.045000  23.205000  99.075000 ;
      RECT  22.595000 113.175000  23.205000 113.205000 ;
      RECT  22.620000 148.070000  34.850000 148.240000 ;
      RECT  22.640000 207.860000  36.680000 208.335000 ;
      RECT  22.650000  42.195000  23.200000  42.495000 ;
      RECT  22.685000  39.040000  22.860000  41.130000 ;
      RECT  22.690000  30.195000  22.860000  32.905000 ;
      RECT  22.690000  38.545000  22.860000  39.040000 ;
      RECT  22.690000  41.130000  22.860000  41.605000 ;
      RECT  22.715000  63.270000  23.385000  63.440000 ;
      RECT  22.815000  95.595000  22.985000  99.045000 ;
      RECT  22.815000 113.205000  22.985000 116.655000 ;
      RECT  22.830000 152.010000  23.000000 154.720000 ;
      RECT  22.910000 178.855000  23.420000 179.185000 ;
      RECT  22.915000  33.455000  23.585000  33.625000 ;
      RECT  22.915000  37.825000  23.585000  37.995000 ;
      RECT  22.915000 163.940000  23.245000 164.110000 ;
      RECT  22.915000 166.250000  23.445000 166.420000 ;
      RECT  22.915000 167.680000  23.445000 167.850000 ;
      RECT  22.915000 169.580000  23.445000 169.750000 ;
      RECT  22.915000 173.650000  23.445000 173.820000 ;
      RECT  22.990000  99.785000  23.160000 103.265000 ;
      RECT  22.990000 108.985000  23.160000 112.465000 ;
      RECT  23.000000 182.465000  23.425000 182.795000 ;
      RECT  23.070000 181.885000  24.830000 182.265000 ;
      RECT  23.115000 179.845000  23.340000 179.865000 ;
      RECT  23.115000 179.865000  23.330000 179.885000 ;
      RECT  23.115000 179.885000  23.310000 179.895000 ;
      RECT  23.120000 179.835000  23.355000 179.845000 ;
      RECT  23.125000 155.440000  23.295000 158.740000 ;
      RECT  23.125000 158.740000  23.655000 159.270000 ;
      RECT  23.130000  73.910000  33.380000  74.080000 ;
      RECT  23.130000  74.080000  23.300000  75.580000 ;
      RECT  23.130000  76.640000  23.300000  78.760000 ;
      RECT  23.130000  78.760000  35.330000  78.930000 ;
      RECT  23.130000  79.190000  35.330000  79.595000 ;
      RECT  23.130000  79.595000  34.900000  82.420000 ;
      RECT  23.135000 179.815000  23.355000 179.835000 ;
      RECT  23.140000 183.275000  23.425000 183.945000 ;
      RECT  23.145000 179.795000  23.355000 179.815000 ;
      RECT  23.160000 179.185000  23.355000 179.795000 ;
      RECT  23.190000  78.930000  35.330000  79.190000 ;
      RECT  23.200000 148.630000  23.370000 151.500000 ;
      RECT  23.210000 128.155000  23.380000 132.905000 ;
      RECT  23.255000 182.795000  23.425000 183.275000 ;
      RECT  23.255000 183.945000  23.425000 184.645000 ;
      RECT  23.255000 184.645000  23.610000 185.655000 ;
      RECT  23.295000 171.340000  25.475000 171.410000 ;
      RECT  23.295000 171.410000  26.315000 171.580000 ;
      RECT  23.295000 171.820000  33.225000 171.990000 ;
      RECT  23.295000 171.990000  25.475000 172.060000 ;
      RECT  23.330000  99.615000  24.440000  99.785000 ;
      RECT  23.330000 103.265000  24.100000 103.435000 ;
      RECT  23.330000 108.815000  24.440000 108.985000 ;
      RECT  23.330000 112.465000  24.445000 112.635000 ;
      RECT  23.390000 177.675000  23.560000 177.785000 ;
      RECT  23.390000 177.785000  24.570000 177.955000 ;
      RECT  23.390000 177.955000  23.560000 178.685000 ;
      RECT  23.410000   4.425000  27.785000   5.135000 ;
      RECT  23.410000   5.135000  24.110000  12.265000 ;
      RECT  23.410000  12.265000  27.785000  12.965000 ;
      RECT  23.410000  17.505000  27.785000  18.205000 ;
      RECT  23.410000  18.205000  24.110000  25.335000 ;
      RECT  23.410000  25.335000  27.785000  26.045000 ;
      RECT  23.430000  42.415000  23.600000  52.305000 ;
      RECT  23.460000  96.145000  23.630000  98.855000 ;
      RECT  23.460000 113.725000  23.630000 116.435000 ;
      RECT  23.480000 179.965000  23.830000 180.975000 ;
      RECT  23.490000  34.025000  23.660000  36.775000 ;
      RECT  23.570000  30.195000  23.740000  32.905000 ;
      RECT  23.570000  38.545000  23.740000  41.255000 ;
      RECT  23.585000  57.685000  23.755000  62.535000 ;
      RECT  23.585000  64.050000  23.755000  68.900000 ;
      RECT  23.590000 178.855000  23.900000 179.130000 ;
      RECT  23.590000 179.130000  23.830000 179.965000 ;
      RECT  23.665000 183.385000  25.710000 183.555000 ;
      RECT  23.710000  74.590000  23.880000  75.600000 ;
      RECT  23.710000  76.650000  23.880000  77.660000 ;
      RECT  23.710000 152.010000  23.880000 154.890000 ;
      RECT  23.730000 178.125000  24.215000 178.455000 ;
      RECT  23.730000 178.455000  23.900000 178.855000 ;
      RECT  23.780000 182.265000  24.830000 182.895000 ;
      RECT  23.800000  95.425000  24.570000  95.595000 ;
      RECT  23.800000 116.655000  24.570000 116.825000 ;
      RECT  23.820000 183.785000  24.350000 183.955000 ;
      RECT  23.820000 183.955000  23.990000 185.625000 ;
      RECT  23.865000 163.940000  25.475000 164.110000 ;
      RECT  23.865000 166.250000  25.475000 166.420000 ;
      RECT  23.865000 167.680000  25.475000 167.850000 ;
      RECT  23.865000 169.580000  25.475000 169.750000 ;
      RECT  23.865000 173.650000  25.475000 173.820000 ;
      RECT  23.880000  99.045000  24.490000  99.075000 ;
      RECT  23.880000 113.175000  24.490000 113.205000 ;
      RECT  23.980000 148.790000  24.150000 151.500000 ;
      RECT  24.000000 179.300000  24.240000 180.975000 ;
      RECT  24.040000  30.350000  24.335000  37.025000 ;
      RECT  24.040000  39.135000  24.335000  41.605000 ;
      RECT  24.040000  41.775000  24.335000  51.935000 ;
      RECT  24.040000  52.565000  24.335000  53.095000 ;
      RECT  24.070000 178.625000  24.570000 178.795000 ;
      RECT  24.070000 178.795000  24.240000 179.300000 ;
      RECT  24.090000 128.135000  24.260000 132.905000 ;
      RECT  24.100000  95.595000  24.270000  99.045000 ;
      RECT  24.100000 113.205000  24.270000 116.655000 ;
      RECT  24.120000 187.325000  24.690000 187.495000 ;
      RECT  24.165000  29.845000  24.335000  30.350000 ;
      RECT  24.165000  37.025000  24.335000  39.135000 ;
      RECT  24.165000  51.935000  24.335000  52.565000 ;
      RECT  24.270000  99.785000  24.440000 102.485000 ;
      RECT  24.270000 102.485000  24.445000 102.715000 ;
      RECT  24.270000 108.985000  24.440000 111.685000 ;
      RECT  24.270000 111.685000  24.445000 111.915000 ;
      RECT  24.270000 188.455000  24.440000 189.410000 ;
      RECT  24.275000 102.715000  24.445000 103.375000 ;
      RECT  24.275000 111.915000  24.445000 112.465000 ;
      RECT  24.300000 184.645000  24.830000 185.655000 ;
      RECT  24.370000 184.125000  25.340000 184.375000 ;
      RECT  24.385000 177.955000  24.570000 178.625000 ;
      RECT  24.405000 156.170000  24.575000 158.880000 ;
      RECT  24.410000 178.965000  25.935000 179.455000 ;
      RECT  24.425000 163.770000  25.975000 163.840000 ;
      RECT  24.425000 163.840000  25.475000 163.940000 ;
      RECT  24.490000 143.270000  25.020000 143.440000 ;
      RECT  24.490000 184.635000  24.660000 184.645000 ;
      RECT  24.520000 187.220000  24.690000 187.325000 ;
      RECT  24.520000 187.495000  24.690000 187.550000 ;
      RECT  24.535000  29.490000  24.705000  30.665000 ;
      RECT  24.535000  30.665000  26.150000  30.835000 ;
      RECT  24.590000 152.010000  24.760000 154.720000 ;
      RECT  24.595000   6.000000  25.135000  11.395000 ;
      RECT  24.595000  19.075000  25.135000  24.470000 ;
      RECT  24.610000  99.615000  25.720000  99.785000 ;
      RECT  24.610000 108.815000  25.720000 108.985000 ;
      RECT  24.615000 103.265000  25.720000 103.435000 ;
      RECT  24.615000 112.465000  25.720000 112.635000 ;
      RECT  24.630000 159.100000  25.300000 159.270000 ;
      RECT  24.670000 214.380000  24.840000 217.340000 ;
      RECT  24.740000  95.485000  24.910000  98.855000 ;
      RECT  24.740000 113.725000  24.910000 116.765000 ;
      RECT  24.760000 148.630000  24.930000 151.500000 ;
      RECT  24.800000  85.175000  27.510000  85.345000 ;
      RECT  24.800000  86.455000  27.510000  86.625000 ;
      RECT  24.850000 143.440000  25.020000 144.135000 ;
      RECT  24.895000  29.150000  25.065000  30.295000 ;
      RECT  24.895000  30.295000  26.150000  30.465000 ;
      RECT  24.895000 217.560000  27.175000 217.730000 ;
      RECT  24.905000 177.785000  26.715000 177.955000 ;
      RECT  24.905000 177.955000  25.075000 178.455000 ;
      RECT  24.940000   5.420000  26.265000   5.830000 ;
      RECT  24.940000  24.640000  26.265000  25.050000 ;
      RECT  24.970000 128.155000  25.140000 132.905000 ;
      RECT  24.985000 179.625000  25.155000 181.145000 ;
      RECT  24.985000 181.145000  26.715000 181.315000 ;
      RECT  24.990000  74.590000  25.160000  77.660000 ;
      RECT  25.030000 184.375000  25.340000 185.455000 ;
      RECT  25.030000 185.455000  26.080000 185.625000 ;
      RECT  25.045000  56.835000  25.215000  70.255000 ;
      RECT  25.080000  95.425000  25.850000  95.595000 ;
      RECT  25.080000 116.655000  25.850000 116.825000 ;
      RECT  25.090000 183.555000  25.710000 183.725000 ;
      RECT  25.100000  45.925000  27.010000  46.095000 ;
      RECT  25.100000  46.095000  25.270000  53.095000 ;
      RECT  25.100000  53.095000  30.145000  53.175000 ;
      RECT  25.100000  53.175000  33.120000  53.265000 ;
      RECT  25.130000  53.265000  33.120000  53.345000 ;
      RECT  25.150000 226.450000  26.000000 248.525000 ;
      RECT  25.150000 248.525000  42.430000 249.375000 ;
      RECT  25.160000  99.045000  25.770000  99.075000 ;
      RECT  25.160000 113.175000  25.770000 113.205000 ;
      RECT  25.270000 142.930000  25.440000 144.580000 ;
      RECT  25.285000 155.105000  26.295000 155.440000 ;
      RECT  25.285000 155.440000  25.455000 158.880000 ;
      RECT  25.330000  75.820000  27.360000  75.990000 ;
      RECT  25.380000  95.595000  25.550000  99.045000 ;
      RECT  25.380000 113.205000  25.550000 116.655000 ;
      RECT  25.470000 152.010000  25.640000 154.865000 ;
      RECT  25.540000 148.790000  25.710000 151.500000 ;
      RECT  25.540000 181.885000  25.710000 183.385000 ;
      RECT  25.540000 183.725000  25.710000 184.585000 ;
      RECT  25.540000 184.585000  26.110000 184.915000 ;
      RECT  25.550000  99.785000  25.720000 103.265000 ;
      RECT  25.550000 108.985000  25.720000 112.465000 ;
      RECT  25.580000  46.445000  25.750000  47.795000 ;
      RECT  25.580000  48.245000  25.750000  49.595000 ;
      RECT  25.580000  50.575000  25.750000  51.925000 ;
      RECT  25.600000 209.800000  25.770000 212.510000 ;
      RECT  25.610000  76.620000  25.780000  77.970000 ;
      RECT  25.635000  50.005000  26.305000  50.175000 ;
      RECT  25.645000 163.330000  25.975000 163.400000 ;
      RECT  25.645000 164.190000  25.815000 164.210000 ;
      RECT  25.645000 164.210000  25.975000 164.280000 ;
      RECT  25.645000 164.650000  25.975000 164.720000 ;
      RECT  25.645000 165.060000  25.975000 165.710000 ;
      RECT  25.645000 166.080000  25.975000 166.150000 ;
      RECT  25.645000 166.520000  25.975000 166.590000 ;
      RECT  25.645000 166.960000  25.975000 167.030000 ;
      RECT  25.645000 168.020000  26.485000 168.090000 ;
      RECT  25.645000 168.460000  25.975000 168.530000 ;
      RECT  25.645000 168.900000  25.975000 168.970000 ;
      RECT  25.645000 169.340000  25.975000 169.410000 ;
      RECT  25.645000 169.850000  26.315000 169.920000 ;
      RECT  25.645000 170.290000  26.315000 170.360000 ;
      RECT  25.645000 170.730000  25.975000 170.800000 ;
      RECT  25.645000 171.170000  25.975000 171.240000 ;
      RECT  25.645000 172.160000  25.975000 172.230000 ;
      RECT  25.645000 172.600000  25.975000 172.670000 ;
      RECT  25.645000 173.025000  26.240000 173.110000 ;
      RECT  25.645000 173.480000  26.240000 173.555000 ;
      RECT  25.755000 212.730000  26.425000 212.900000 ;
      RECT  25.765000 178.125000  25.935000 178.965000 ;
      RECT  25.765000 179.455000  25.935000 180.975000 ;
      RECT  25.775000 217.730000  26.770000 217.735000 ;
      RECT  25.850000 128.135000  26.020000 132.905000 ;
      RECT  25.890000  52.335000  26.220000  52.845000 ;
      RECT  25.890000  99.615000  26.660000  99.785000 ;
      RECT  25.890000 103.265000  26.660000 103.435000 ;
      RECT  25.890000 108.815000  26.660000 108.985000 ;
      RECT  25.890000 112.465000  26.660000 112.635000 ;
      RECT  25.920000 183.275000  26.450000 183.945000 ;
      RECT  25.925000  50.175000  26.190000  52.335000 ;
      RECT  25.940000 184.915000  26.110000 184.975000 ;
      RECT  25.945000  39.575000  53.345000  39.745000 ;
      RECT  25.945000  39.745000  26.260000  43.980000 ;
      RECT  25.945000  43.980000  34.955000  44.145000 ;
      RECT  25.950000 214.630000  26.120000 217.340000 ;
      RECT  25.960000  78.350000  27.990000  78.520000 ;
      RECT  25.970000  99.785000  26.580000  99.815000 ;
      RECT  25.970000 108.985000  26.580000 109.015000 ;
      RECT  26.005000 188.125000  28.965000 188.295000 ;
      RECT  26.020000  95.425000  26.970000  95.595000 ;
      RECT  26.020000  95.595000  26.190000  99.075000 ;
      RECT  26.020000  99.075000  26.970000  99.245000 ;
      RECT  26.020000 113.005000  26.970000 113.175000 ;
      RECT  26.020000 113.175000  26.190000 116.655000 ;
      RECT  26.020000 116.655000  26.970000 116.825000 ;
      RECT  26.040000 187.245000  28.965000 187.415000 ;
      RECT  26.065000 104.675000  26.235000 104.850000 ;
      RECT  26.065000 105.120000  26.235000 105.630000 ;
      RECT  26.065000 105.900000  26.235000 106.410000 ;
      RECT  26.065000 106.680000  26.235000 107.190000 ;
      RECT  26.065000 107.460000  26.235000 107.575000 ;
      RECT  26.065000 125.415000  28.290000 126.035000 ;
      RECT  26.065000 127.040000  28.290000 127.705000 ;
      RECT  26.070000   6.000000  26.610000  11.395000 ;
      RECT  26.070000  19.075000  26.610000  24.470000 ;
      RECT  26.080000 155.700000  26.710000 155.870000 ;
      RECT  26.080000 155.870000  26.250000 156.845000 ;
      RECT  26.090000  44.145000  34.955000  44.150000 ;
      RECT  26.090000 182.465000  26.450000 182.795000 ;
      RECT  26.095000 126.035000  28.290000 127.040000 ;
      RECT  26.105000 179.035000  27.270000 179.205000 ;
      RECT  26.120000 181.885000  27.540000 182.265000 ;
      RECT  26.145000 169.500000  32.730000 169.670000 ;
      RECT  26.145000 169.670000  26.315000 169.850000 ;
      RECT  26.145000 170.730000  26.815000 170.800000 ;
      RECT  26.145000 170.800000  33.225000 171.170000 ;
      RECT  26.145000 171.170000  26.815000 171.240000 ;
      RECT  26.145000 171.240000  26.315000 171.410000 ;
      RECT  26.255000 189.005000  28.965000 189.175000 ;
      RECT  26.270000  74.590000  26.440000  75.600000 ;
      RECT  26.280000 182.795000  26.450000 183.275000 ;
      RECT  26.280000 183.945000  26.450000 184.675000 ;
      RECT  26.280000 184.675000  26.660000 185.685000 ;
      RECT  26.315000 163.705000  29.495000 163.875000 ;
      RECT  26.315000 163.875000  26.485000 164.890000 ;
      RECT  26.315000 166.820000  28.855000 166.990000 ;
      RECT  26.315000 166.990000  26.485000 168.020000 ;
      RECT  26.320000 148.630000  26.490000 151.500000 ;
      RECT  26.350000 152.010000  26.520000 154.720000 ;
      RECT  26.360000  46.445000  26.530000  47.795000 ;
      RECT  26.360000  48.245000  26.530000  49.595000 ;
      RECT  26.360000  50.575000  26.530000  51.925000 ;
      RECT  26.440000  28.185000  30.125000  28.365000 ;
      RECT  26.440000  28.365000  26.620000  37.515000 ;
      RECT  26.440000  37.515000  51.980000  37.695000 ;
      RECT  26.480000 209.800000  26.650000 212.510000 ;
      RECT  26.485000 169.840000  26.815000 169.920000 ;
      RECT  26.485000 169.920000  33.225000 170.290000 ;
      RECT  26.485000 170.290000  26.815000 170.370000 ;
      RECT  26.485000 171.610000  26.815000 171.680000 ;
      RECT  26.485000 171.680000  33.225000 171.820000 ;
      RECT  26.485000 171.990000  33.225000 172.050000 ;
      RECT  26.485000 172.050000  26.815000 172.120000 ;
      RECT  26.485000 173.040000  26.815000 173.110000 ;
      RECT  26.485000 173.110000  33.225000 173.260000 ;
      RECT  26.485000 173.260000  37.760000 173.460000 ;
      RECT  26.485000 173.460000  33.225000 173.480000 ;
      RECT  26.485000 173.480000  26.815000 173.550000 ;
      RECT  26.510000 156.170000  26.680000 158.880000 ;
      RECT  26.540000 155.270000  27.210000 155.440000 ;
      RECT  26.540000 155.440000  26.710000 155.700000 ;
      RECT  26.545000 177.955000  26.715000 178.455000 ;
      RECT  26.545000 179.625000  26.715000 181.145000 ;
      RECT  26.560000 104.365000  28.285000 105.115000 ;
      RECT  26.560000 107.090000  28.285000 107.840000 ;
      RECT  26.585000  50.005000  28.430000  50.175000 ;
      RECT  26.635000  40.130000  53.130000  40.460000 ;
      RECT  26.635000  40.760000  27.305000  41.720000 ;
      RECT  26.635000  42.020000  27.305000  42.980000 ;
      RECT  26.635000  43.280000  36.095000  43.610000 ;
      RECT  26.665000  50.000000  28.370000  50.005000 ;
      RECT  26.670000  52.195000  27.000000  52.845000 ;
      RECT  26.705000 182.265000  27.540000 182.795000 ;
      RECT  26.705000 212.730000  28.185000 212.900000 ;
      RECT  26.720000 105.675000  27.390000 105.850000 ;
      RECT  26.720000 106.460000  27.390000 106.630000 ;
      RECT  26.730000 128.155000  26.900000 132.905000 ;
      RECT  26.750000 183.145000  27.280000 183.725000 ;
      RECT  26.770000  74.590000  27.720000  74.760000 ;
      RECT  26.800000  95.595000  26.970000  99.075000 ;
      RECT  26.800000 113.175000  26.970000 116.655000 ;
      RECT  26.830000 100.005000  27.000000 100.795000 ;
      RECT  26.830000 100.795000  27.440000 100.965000 ;
      RECT  26.830000 100.965000  27.000000 102.715000 ;
      RECT  26.830000 109.205000  27.000000 109.995000 ;
      RECT  26.830000 109.995000  27.440000 110.165000 ;
      RECT  26.830000 110.165000  27.000000 111.915000 ;
      RECT  26.840000  46.095000  27.010000  46.800000 ;
      RECT  26.840000  46.800000  33.120000  46.970000 ;
      RECT  26.885000 133.415000  27.555000 133.585000 ;
      RECT  26.885000 176.655000  27.835000 176.985000 ;
      RECT  26.885000 176.985000  27.155000 179.035000 ;
      RECT  26.890000  76.620000  27.720000  76.790000 ;
      RECT  26.890000  76.790000  27.060000  77.970000 ;
      RECT  26.935000 183.725000  27.105000 185.625000 ;
      RECT  26.945000 133.405000  27.515000 133.415000 ;
      RECT  26.955000  66.305000  44.940000  68.100000 ;
      RECT  26.955000  68.100000  64.075000  68.330000 ;
      RECT  26.955000  68.330000  64.045000  70.420000 ;
      RECT  26.955000  70.420000  97.970000  71.040000 ;
      RECT  26.955000  71.040000  84.585000  71.560000 ;
      RECT  26.955000 163.270000  28.005000 163.440000 ;
      RECT  26.955000 164.150000  27.965000 164.360000 ;
      RECT  26.955000 164.360000  30.175000 164.530000 ;
      RECT  26.970000  56.030000  32.665000  56.200000 ;
      RECT  26.970000  56.200000  27.140000  64.455000 ;
      RECT  26.970000  64.455000  32.665000  64.625000 ;
      RECT  26.985000 165.980000  27.995000 166.150000 ;
      RECT  26.985000 166.150000  28.005000 166.320000 ;
      RECT  26.985000 166.320000  27.995000 166.510000 ;
      RECT  26.985000 167.200000  27.995000 167.385000 ;
      RECT  26.985000 167.385000  30.175000 167.555000 ;
      RECT  26.985000 169.670000  32.730000 169.750000 ;
      RECT  26.985000 170.460000  28.050000 170.630000 ;
      RECT  26.985000 172.220000  28.805000 172.390000 ;
      RECT  26.985000 172.770000  32.730000 172.940000 ;
      RECT  26.985000 173.650000  28.035000 173.820000 ;
      RECT  27.015000 164.730000  27.185000 165.470000 ;
      RECT  27.015000 165.470000  28.515000 165.780000 ;
      RECT  27.015000 167.780000  27.185000 168.320000 ;
      RECT  27.015000 168.320000  28.885000 168.490000 ;
      RECT  27.055000  99.615000  27.780000  99.785000 ;
      RECT  27.055000 103.265000  27.780000 103.435000 ;
      RECT  27.055000 112.465000  27.780000 112.635000 ;
      RECT  27.085000   5.135000  27.785000  12.265000 ;
      RECT  27.085000  18.205000  27.785000  25.335000 ;
      RECT  27.100000 148.790000  27.270000 151.500000 ;
      RECT  27.110000 171.340000  32.730000 171.510000 ;
      RECT  27.115000 169.030000  28.005000 169.200000 ;
      RECT  27.120000  51.140000  27.310000  51.925000 ;
      RECT  27.120000  51.925000  27.290000  52.025000 ;
      RECT  27.140000  48.245000  27.310000  49.595000 ;
      RECT  27.140000  50.575000  27.310000  51.140000 ;
      RECT  27.150000 227.595000  40.485000 228.345000 ;
      RECT  27.150000 228.345000  27.900000 246.620000 ;
      RECT  27.150000 246.620000  40.485000 247.375000 ;
      RECT  27.230000 152.010000  27.400000 154.720000 ;
      RECT  27.230000 214.380000  27.400000 217.340000 ;
      RECT  27.295000 179.575000  27.465000 179.625000 ;
      RECT  27.295000 179.625000  27.495000 180.825000 ;
      RECT  27.325000 177.155000  27.495000 178.595000 ;
      RECT  27.325000 180.825000  27.495000 180.975000 ;
      RECT  27.360000 209.800000  27.530000 212.510000 ;
      RECT  27.370000 184.635000  27.540000 185.685000 ;
      RECT  27.390000 155.945000  27.560000 158.880000 ;
      RECT  27.450000  52.195000  27.780000  52.230000 ;
      RECT  27.450000  52.230000  28.060000  52.400000 ;
      RECT  27.450000  52.400000  27.780000  52.845000 ;
      RECT  27.455000 155.270000  28.125000 155.440000 ;
      RECT  27.455000 217.560000  29.735000 217.730000 ;
      RECT  27.475000  30.255000  51.470000  30.425000 ;
      RECT  27.475000  30.425000  27.645000  36.580000 ;
      RECT  27.475000  36.580000  50.100000  36.590000 ;
      RECT  27.475000  36.590000  51.470000  36.750000 ;
      RECT  27.520000  77.070000  27.690000  78.350000 ;
      RECT  27.550000  74.560000  27.720000  74.590000 ;
      RECT  27.550000  74.760000  27.720000  75.120000 ;
      RECT  27.550000  75.120000  28.020000  75.650000 ;
      RECT  27.550000  75.650000  27.720000  76.620000 ;
      RECT  27.610000  87.565000  27.780000  94.355000 ;
      RECT  27.610000  99.785000  27.780000 103.265000 ;
      RECT  27.610000 108.815000  27.780000 112.465000 ;
      RECT  27.610000 117.835000  27.780000 124.625000 ;
      RECT  27.610000 128.155000  27.780000 132.905000 ;
      RECT  27.665000 164.700000  28.055000 164.870000 ;
      RECT  27.665000 167.750000  27.995000 167.980000 ;
      RECT  27.665000 167.980000  30.755000 168.150000 ;
      RECT  27.665000 179.320000  28.090000 179.850000 ;
      RECT  27.705000  48.245000  27.875000  49.595000 ;
      RECT  27.715000 159.100000  28.245000 159.270000 ;
      RECT  27.725000 164.870000  28.055000 165.100000 ;
      RECT  27.725000 165.100000  30.755000 165.270000 ;
      RECT  27.730000  85.420000  27.900000  86.400000 ;
      RECT  27.730000 105.820000  27.900000 106.490000 ;
      RECT  27.880000 148.630000  28.050000 151.500000 ;
      RECT  27.890000  75.820000  28.960000  75.990000 ;
      RECT  27.890000 155.440000  28.100000 159.100000 ;
      RECT  27.890000 159.270000  28.100000 159.440000 ;
      RECT  27.895000  56.945000  31.725000  57.175000 ;
      RECT  27.895000  57.175000  28.125000  63.485000 ;
      RECT  27.895000  63.485000  28.715000  63.515000 ;
      RECT  27.895000  63.515000  31.755000  63.685000 ;
      RECT  27.895000  63.685000  28.715000  63.715000 ;
      RECT  27.920000  50.575000  28.090000  51.925000 ;
      RECT  27.920000 177.155000  28.090000 179.320000 ;
      RECT  27.920000 179.850000  28.090000 182.900000 ;
      RECT  27.950000 184.215000  40.820000 186.105000 ;
      RECT  28.090000  84.545000  28.260000 103.825000 ;
      RECT  28.090000 103.825000  28.285000 104.365000 ;
      RECT  28.090000 105.115000  28.285000 107.090000 ;
      RECT  28.090000 107.840000  28.285000 108.450000 ;
      RECT  28.090000 108.450000  28.260000 117.400000 ;
      RECT  28.090000 117.400000  28.290000 125.365000 ;
      RECT  28.090000 127.755000  28.290000 133.100000 ;
      RECT  28.090000 133.100000  28.260000 133.775000 ;
      RECT  28.100000  31.485000  28.270000  32.155000 ;
      RECT  28.100000  32.665000  28.270000  33.335000 ;
      RECT  28.100000  33.845000  28.270000  34.515000 ;
      RECT  28.100000  35.025000  28.270000  35.695000 ;
      RECT  28.110000 152.010000  28.280000 154.720000 ;
      RECT  28.170000  76.620000  28.340000  77.970000 ;
      RECT  28.190000  74.080000  28.360000  75.580000 ;
      RECT  28.190000 176.655000  28.700000 176.690000 ;
      RECT  28.190000 176.690000  28.720000 176.860000 ;
      RECT  28.190000 176.860000  28.700000 176.985000 ;
      RECT  28.190000 183.065000  28.700000 183.395000 ;
      RECT  28.220000 170.460000  28.795000 170.630000 ;
      RECT  28.230000  52.195000  28.560000  52.845000 ;
      RECT  28.240000 209.800000  28.410000 212.510000 ;
      RECT  28.260000 176.985000  28.630000 183.065000 ;
      RECT  28.265000 165.780000  28.515000 166.440000 ;
      RECT  28.265000 173.650000  28.795000 173.820000 ;
      RECT  28.270000 156.170000  28.440000 158.880000 ;
      RECT  28.415000 159.100000  31.805000 159.270000 ;
      RECT  28.485000  48.100000  28.655000  49.595000 ;
      RECT  28.510000 214.630000  28.680000 217.340000 ;
      RECT  28.515000  57.980000  28.685000  62.830000 ;
      RECT  28.520000  31.155000  38.410000  31.325000 ;
      RECT  28.520000  32.335000  38.410000  32.505000 ;
      RECT  28.520000  33.515000  38.410000  33.685000 ;
      RECT  28.520000  34.695000  38.410000  34.865000 ;
      RECT  28.520000  35.875000  38.410000  36.045000 ;
      RECT  28.520000  78.350000  30.550000  78.520000 ;
      RECT  28.540000  47.675000  29.210000  47.845000 ;
      RECT  28.545000   3.665000  29.245000  13.725000 ;
      RECT  28.545000  16.745000  29.245000  26.805000 ;
      RECT  28.625000 229.105000  38.920000 229.275000 ;
      RECT  28.625000 229.275000  28.835000 245.690000 ;
      RECT  28.625000 245.690000  38.920000 245.865000 ;
      RECT  28.660000 148.790000  28.830000 151.500000 ;
      RECT  28.660000 152.010000  28.830000 154.735000 ;
      RECT  28.680000  51.135000  28.870000  51.925000 ;
      RECT  28.680000  51.925000  28.850000  52.025000 ;
      RECT  28.680000 217.730000  29.675000 217.735000 ;
      RECT  28.685000 166.305000  28.855000 166.820000 ;
      RECT  28.695000 164.530000  29.365000 164.890000 ;
      RECT  28.695000 167.555000  29.365000 167.670000 ;
      RECT  28.700000  50.575000  28.870000  51.135000 ;
      RECT  28.790000  74.590000  29.740000  74.760000 ;
      RECT  28.790000  74.760000  28.960000  75.820000 ;
      RECT  28.790000  75.990000  28.960000  76.620000 ;
      RECT  28.790000  76.620000  29.620000  76.790000 ;
      RECT  28.800000 177.155000  28.970000 178.205000 ;
      RECT  28.800000 178.435000  28.970000 178.765000 ;
      RECT  28.800000 179.385000  28.970000 179.715000 ;
      RECT  28.800000 179.885000  28.970000 182.595000 ;
      RECT  28.820000  77.070000  28.990000  78.350000 ;
      RECT  28.875000  47.845000  29.045000  48.780000 ;
      RECT  28.885000 155.270000  34.995000 155.440000 ;
      RECT  28.905000  57.400000  29.575000  57.570000 ;
      RECT  28.915000 163.530000  29.495000 163.705000 ;
      RECT  28.915000 163.875000  29.495000 164.060000 ;
      RECT  28.915000 165.270000  29.255000 165.720000 ;
      RECT  28.920000 190.360000  29.090000 191.370000 ;
      RECT  28.920000 192.220000  29.090000 193.230000 ;
      RECT  28.975000  57.390000  29.505000  57.400000 ;
      RECT  29.010000  52.195000  29.340000  52.230000 ;
      RECT  29.010000  52.230000  29.620000  52.400000 ;
      RECT  29.010000  52.400000  29.340000  52.845000 ;
      RECT  29.070000 176.655000  29.580000 176.985000 ;
      RECT  29.070000 183.065000  29.580000 183.395000 ;
      RECT  29.085000 165.720000  29.255000 167.145000 ;
      RECT  29.130000  75.120000  29.300000  75.820000 ;
      RECT  29.130000  75.820000  31.180000  75.990000 ;
      RECT  29.140000 176.985000  29.510000 183.065000 ;
      RECT  29.145000  86.645000  30.035000  88.205000 ;
      RECT  29.145000  89.825000  30.035000  94.985000 ;
      RECT  29.145000  97.085000  30.035000  99.415000 ;
      RECT  29.145000 103.775000  30.035000 108.215000 ;
      RECT  29.145000 112.835000  30.035000 115.480000 ;
      RECT  29.145000 117.405000  30.035000 122.700000 ;
      RECT  29.145000 125.500000  30.035000 127.655000 ;
      RECT  29.145000 128.425000  30.035000 129.725000 ;
      RECT  29.145000 130.805000  30.035000 134.385000 ;
      RECT  29.145000 191.620000  33.145000 191.790000 ;
      RECT  29.145000 193.480000  33.145000 193.650000 ;
      RECT  29.145000 230.095000  29.315000 245.125000 ;
      RECT  29.150000 155.945000  29.320000 158.880000 ;
      RECT  29.165000  84.410000  30.015000  86.645000 ;
      RECT  29.165000  88.205000  30.015000  89.825000 ;
      RECT  29.165000  94.985000  30.015000  97.085000 ;
      RECT  29.165000  99.415000  30.015000 103.775000 ;
      RECT  29.165000 108.215000  30.015000 112.835000 ;
      RECT  29.165000 115.480000  30.015000 117.405000 ;
      RECT  29.165000 122.700000  30.015000 125.500000 ;
      RECT  29.165000 127.655000  30.015000 128.425000 ;
      RECT  29.165000 129.725000  30.015000 130.805000 ;
      RECT  29.165000 134.385000  30.015000 134.865000 ;
      RECT  29.185000 187.400000  29.355000 188.070000 ;
      RECT  29.185000 188.350000  29.355000 189.020000 ;
      RECT  29.215000 170.460000  29.545000 170.630000 ;
      RECT  29.215000 173.650000  29.545000 173.820000 ;
      RECT  29.265000  48.245000  29.435000  49.595000 ;
      RECT  29.285000 229.695000  30.735000 229.865000 ;
      RECT  29.415000 168.150000  30.755000 168.320000 ;
      RECT  29.415000 168.320000  29.585000 168.540000 ;
      RECT  29.440000 148.630000  29.610000 151.500000 ;
      RECT  29.440000 151.670000  34.290000 151.840000 ;
      RECT  29.440000 151.840000  29.610000 154.735000 ;
      RECT  29.450000  76.790000  29.620000  77.970000 ;
      RECT  29.480000  50.575000  29.650000  51.925000 ;
      RECT  29.490000  47.675000  32.270000  47.845000 ;
      RECT  29.680000 177.155000  29.850000 182.900000 ;
      RECT  29.715000 170.460000  32.425000 170.630000 ;
      RECT  29.715000 172.220000  32.425000 172.390000 ;
      RECT  29.715000 173.650000  32.425000 173.820000 ;
      RECT  29.745000 165.980000  30.755000 166.070000 ;
      RECT  29.745000 166.070000  32.895000 166.240000 ;
      RECT  29.745000 166.240000  37.440000 166.410000 ;
      RECT  29.745000 166.410000  32.895000 166.580000 ;
      RECT  29.745000 166.580000  30.755000 167.030000 ;
      RECT  29.745000 169.030000  30.755000 169.200000 ;
      RECT  29.755000 168.670000  30.755000 169.030000 ;
      RECT  29.785000 209.185000  30.295000 213.440000 ;
      RECT  29.790000 214.380000  29.960000 217.340000 ;
      RECT  29.795000  58.080000  29.965000  62.830000 ;
      RECT  29.845000 163.270000  30.755000 164.105000 ;
      RECT  29.845000 164.530000  30.175000 164.720000 ;
      RECT  29.845000 167.555000  30.175000 167.810000 ;
      RECT  29.925000 230.175000  30.095000 245.125000 ;
      RECT  29.945000   0.750000  71.625000   0.930000 ;
      RECT  29.945000   0.930000  30.125000  28.185000 ;
      RECT  29.975000  50.370000  33.120000  50.540000 ;
      RECT  29.975000  50.540000  30.960000  50.820000 ;
      RECT  29.975000  50.820000  30.145000  51.305000 ;
      RECT  29.975000  51.305000  30.300000  52.535000 ;
      RECT  29.975000  52.535000  30.145000  53.095000 ;
      RECT  30.015000 217.560000  32.295000 217.730000 ;
      RECT  30.030000 156.170000  30.200000 158.880000 ;
      RECT  30.045000  48.245000  30.215000  49.740000 ;
      RECT  30.070000  74.590000  30.240000  75.600000 ;
      RECT  30.185000  57.400000  30.855000  57.570000 ;
      RECT  30.220000 148.790000  30.390000 151.500000 ;
      RECT  30.220000 152.010000  30.390000 154.720000 ;
      RECT  30.230000 177.155000  30.400000 178.205000 ;
      RECT  30.230000 178.435000  30.400000 178.765000 ;
      RECT  30.230000 179.385000  30.400000 179.715000 ;
      RECT  30.230000 179.885000  30.400000 182.595000 ;
      RECT  30.255000  57.390000  30.785000  57.400000 ;
      RECT  30.375000 164.105000  30.755000 164.690000 ;
      RECT  30.375000 167.030000  30.755000 167.740000 ;
      RECT  30.500000 176.655000  31.010000 176.985000 ;
      RECT  30.500000 183.065000  31.010000 183.395000 ;
      RECT  30.565000  63.485000  31.755000  63.515000 ;
      RECT  30.565000  63.685000  31.755000  63.715000 ;
      RECT  30.570000 176.985000  30.940000 183.065000 ;
      RECT  30.580000 156.170000  30.750000 156.455000 ;
      RECT  30.580000 156.455000  31.110000 156.985000 ;
      RECT  30.580000 156.985000  30.750000 158.880000 ;
      RECT  30.705000 230.095000  30.875000 245.125000 ;
      RECT  30.730000  76.620000  30.900000  77.970000 ;
      RECT  30.865000  29.320000  71.625000  29.490000 ;
      RECT  30.920000 209.680000  31.090000 210.690000 ;
      RECT  30.920000 212.245000  31.090000 213.115000 ;
      RECT  31.000000 148.630000  31.170000 151.500000 ;
      RECT  31.000000 151.840000  31.170000 154.735000 ;
      RECT  31.070000 214.630000  31.240000 217.340000 ;
      RECT  31.075000  57.980000  31.245000  62.830000 ;
      RECT  31.075000 211.785000  31.745000 211.955000 ;
      RECT  31.110000 177.155000  31.280000 182.900000 ;
      RECT  31.145000 210.910000  32.625000 211.080000 ;
      RECT  31.160000 158.675000  31.690000 159.100000 ;
      RECT  31.185000 229.275000  31.355000 245.690000 ;
      RECT  31.190000 217.730000  31.955000 217.735000 ;
      RECT  31.300000   5.235000  47.515000   5.415000 ;
      RECT  31.300000   5.415000  31.480000  15.485000 ;
      RECT  31.300000  15.485000  31.500000  16.910000 ;
      RECT  31.300000  16.910000  31.480000  28.375000 ;
      RECT  31.300000  28.375000  70.680000  28.555000 ;
      RECT  31.315000 163.450000  31.645000 165.560000 ;
      RECT  31.315000 165.560000  33.760000 165.830000 ;
      RECT  31.315000 166.820000  33.760000 167.090000 ;
      RECT  31.315000 167.090000  31.645000 169.200000 ;
      RECT  31.350000  74.590000  31.520000  77.660000 ;
      RECT  31.380000 176.655000  32.770000 176.985000 ;
      RECT  31.380000 183.065000  32.770000 183.395000 ;
      RECT  31.405000  83.975000  89.205000  84.825000 ;
      RECT  31.405000  84.825000  31.575000  96.855000 ;
      RECT  31.405000  96.855000  79.175000  97.145000 ;
      RECT  31.405000  97.145000  31.575000 106.160000 ;
      RECT  31.405000 106.160000  71.755000 106.360000 ;
      RECT  31.405000 106.360000  31.575000 115.375000 ;
      RECT  31.405000 115.375000  79.175000 115.675000 ;
      RECT  31.405000 115.675000  31.575000 127.885000 ;
      RECT  31.405000 127.885000  90.225000 128.205000 ;
      RECT  31.450000 176.985000  31.820000 183.065000 ;
      RECT  31.470000   2.235000  31.980000   2.905000 ;
      RECT  31.490000   3.925000  32.000000   4.595000 ;
      RECT  31.525000  57.920000  31.755000  63.485000 ;
      RECT  31.555000  57.175000  31.725000  57.920000 ;
      RECT  31.665000 230.095000  31.835000 245.125000 ;
      RECT  31.710000 128.205000  32.560000 143.885000 ;
      RECT  31.710000 143.885000  39.450000 145.100000 ;
      RECT  31.720000  21.575000  31.900000  22.110000 ;
      RECT  31.730000   6.305000  32.000000   6.500000 ;
      RECT  31.730000   6.500000  32.025000   9.840000 ;
      RECT  31.730000   9.840000  32.000000   9.915000 ;
      RECT  31.730000   9.915000  31.900000  10.035000 ;
      RECT  31.730000  10.605000  31.900000  12.565000 ;
      RECT  31.730000  13.165000  31.900000  20.525000 ;
      RECT  31.730000  21.155000  31.900000  21.575000 ;
      RECT  31.730000  22.110000  31.900000  22.505000 ;
      RECT  31.730000  23.385000  31.900000  23.580000 ;
      RECT  31.730000  23.580000  32.025000  26.920000 ;
      RECT  31.730000  26.920000  31.900000  27.115000 ;
      RECT  31.780000 148.790000  31.950000 151.500000 ;
      RECT  31.780000 152.010000  31.950000 154.720000 ;
      RECT  31.800000 209.680000  31.970000 210.690000 ;
      RECT  31.800000 212.245000  31.970000 213.115000 ;
      RECT  31.805000 229.695000  33.255000 229.865000 ;
      RECT  31.860000 155.830000  33.790000 156.000000 ;
      RECT  31.860000 156.000000  32.030000 158.880000 ;
      RECT  31.865000 164.015000  32.035000 165.025000 ;
      RECT  31.990000 177.155000  32.160000 178.205000 ;
      RECT  31.990000 178.435000  32.160000 178.765000 ;
      RECT  31.990000 179.385000  32.160000 179.715000 ;
      RECT  31.990000 179.885000  32.160000 182.595000 ;
      RECT  32.025000 211.785000  32.695000 211.955000 ;
      RECT  32.120000   5.945000  34.830000   6.115000 ;
      RECT  32.120000  10.225000  34.830000  10.395000 ;
      RECT  32.120000  11.505000  34.830000  11.675000 ;
      RECT  32.120000  12.785000  34.830000  12.955000 ;
      RECT  32.120000  14.065000  34.830000  14.235000 ;
      RECT  32.120000  15.345000  34.830000  15.515000 ;
      RECT  32.120000  16.625000  34.830000  16.795000 ;
      RECT  32.120000  17.905000  34.830000  18.075000 ;
      RECT  32.120000  19.185000  34.830000  19.355000 ;
      RECT  32.120000  20.465000  34.830000  20.635000 ;
      RECT  32.120000  21.745000  34.830000  21.915000 ;
      RECT  32.120000  23.025000  34.830000  23.195000 ;
      RECT  32.120000  27.305000  34.830000  27.475000 ;
      RECT  32.325000  48.245000  32.495000  49.740000 ;
      RECT  32.330000 176.985000  32.700000 183.065000 ;
      RECT  32.350000 214.380000  32.520000 217.340000 ;
      RECT  32.380000 159.045000  32.910000 159.575000 ;
      RECT  32.425000 172.560000  33.680000 172.745000 ;
      RECT  32.425000 172.745000  32.730000 172.770000 ;
      RECT  32.445000 230.175000  32.615000 245.125000 ;
      RECT  32.495000  56.200000  32.665000  64.455000 ;
      RECT  32.560000 148.630000  32.730000 151.500000 ;
      RECT  32.560000 151.840000  32.730000 154.735000 ;
      RECT  32.565000 163.450000  32.895000 163.460000 ;
      RECT  32.565000 163.460000  35.725000 163.730000 ;
      RECT  32.565000 163.730000  32.895000 163.960000 ;
      RECT  32.565000 168.690000  32.895000 168.920000 ;
      RECT  32.565000 168.920000  35.725000 169.190000 ;
      RECT  32.565000 169.190000  32.895000 169.200000 ;
      RECT  32.575000 217.560000  34.855000 217.730000 ;
      RECT  32.595000 172.415000  33.680000 172.560000 ;
      RECT  32.630000  74.590000  32.800000  75.600000 ;
      RECT  32.630000  76.650000  32.800000  77.660000 ;
      RECT  32.635000 217.730000  33.630000 217.735000 ;
      RECT  32.680000 209.680000  32.850000 210.690000 ;
      RECT  32.680000 212.185000  32.850000 212.915000 ;
      RECT  32.740000 156.170000  32.910000 159.045000 ;
      RECT  32.870000 177.155000  33.040000 182.900000 ;
      RECT  32.875000  89.620000  33.765000  94.495000 ;
      RECT  32.875000 118.025000  33.765000 122.900000 ;
      RECT  32.895000 169.850000  33.225000 169.920000 ;
      RECT  32.895000 170.290000  33.225000 170.360000 ;
      RECT  32.895000 170.730000  33.225000 170.800000 ;
      RECT  32.895000 171.170000  33.225000 171.240000 ;
      RECT  32.895000 171.610000  33.225000 171.680000 ;
      RECT  32.895000 172.050000  33.225000 172.120000 ;
      RECT  32.895000 173.040000  33.225000 173.110000 ;
      RECT  32.895000 173.480000  33.225000 173.550000 ;
      RECT  32.915000  85.710000  33.765000  89.620000 ;
      RECT  32.915000  94.495000  33.765000  95.620000 ;
      RECT  32.915000  95.620000  33.085000  95.730000 ;
      RECT  32.915000 116.790000  33.085000 116.900000 ;
      RECT  32.915000 116.900000  33.765000 118.025000 ;
      RECT  32.915000 122.900000  33.765000 126.810000 ;
      RECT  32.950000  46.970000  33.120000  50.370000 ;
      RECT  32.950000  50.540000  33.120000  53.175000 ;
      RECT  33.035000 164.425000  33.365000 165.090000 ;
      RECT  33.035000 165.090000  37.280000 165.260000 ;
      RECT  33.035000 167.390000  37.280000 167.560000 ;
      RECT  33.035000 167.560000  33.365000 168.225000 ;
      RECT  33.140000 176.655000  33.650000 176.985000 ;
      RECT  33.140000 183.065000  33.650000 183.395000 ;
      RECT  33.155000 159.100000  34.845000 159.270000 ;
      RECT  33.200000 190.360000  33.370000 190.940000 ;
      RECT  33.200000 190.940000  33.785000 191.110000 ;
      RECT  33.200000 191.110000  33.370000 191.370000 ;
      RECT  33.200000 192.220000  33.370000 193.230000 ;
      RECT  33.210000  74.080000  33.380000  75.580000 ;
      RECT  33.210000  76.640000  35.330000  78.760000 ;
      RECT  33.210000  98.390000  70.340000  98.560000 ;
      RECT  33.210000  98.560000  33.380000 104.760000 ;
      RECT  33.210000 104.760000  70.340000 104.930000 ;
      RECT  33.210000 107.590000  70.340000 107.760000 ;
      RECT  33.210000 107.760000  33.380000 113.960000 ;
      RECT  33.210000 113.960000  70.340000 114.130000 ;
      RECT  33.210000 176.985000  33.580000 183.065000 ;
      RECT  33.225000 230.095000  33.395000 245.125000 ;
      RECT  33.325000 129.450000  48.575000 129.620000 ;
      RECT  33.325000 129.620000  33.495000 131.490000 ;
      RECT  33.325000 131.490000  48.575000 131.660000 ;
      RECT  33.325000 131.660000  33.495000 142.950000 ;
      RECT  33.325000 142.950000  40.385000 143.120000 ;
      RECT  33.340000 148.790000  33.510000 151.500000 ;
      RECT  33.340000 152.010000  33.510000 154.720000 ;
      RECT  33.430000 165.830000  41.700000 166.070000 ;
      RECT  33.430000 166.580000  41.700000 166.785000 ;
      RECT  33.430000 166.785000  39.270000 166.795000 ;
      RECT  33.430000 166.795000  33.760000 166.820000 ;
      RECT  33.530000   3.925000  36.835000   4.595000 ;
      RECT  33.620000 156.000000  33.790000 158.880000 ;
      RECT  33.630000 214.630000  33.800000 217.340000 ;
      RECT  33.705000 229.275000  33.875000 245.690000 ;
      RECT  33.750000 130.240000  33.920000 130.400000 ;
      RECT  33.750000 130.400000  34.380000 130.570000 ;
      RECT  33.750000 130.570000  33.920000 130.910000 ;
      RECT  33.750000 177.155000  33.920000 178.205000 ;
      RECT  33.750000 178.435000  33.920000 178.765000 ;
      RECT  33.750000 179.385000  33.920000 179.715000 ;
      RECT  33.750000 179.885000  33.920000 182.595000 ;
      RECT  33.780000 101.080000  33.960000 101.970000 ;
      RECT  33.780000 110.280000  33.960000 111.170000 ;
      RECT  33.790000  98.800000  34.420000  98.970000 ;
      RECT  33.790000  98.970000  33.960000 101.080000 ;
      RECT  33.790000 101.970000  33.960000 104.350000 ;
      RECT  33.790000 104.350000  34.420000 104.520000 ;
      RECT  33.790000 108.000000  34.420000 108.170000 ;
      RECT  33.790000 108.170000  33.960000 110.280000 ;
      RECT  33.790000 111.170000  33.960000 113.550000 ;
      RECT  33.790000 113.550000  34.420000 113.720000 ;
      RECT  33.820000  85.370000  37.820000  85.540000 ;
      RECT  33.820000  95.920000  37.820000  96.090000 ;
      RECT  33.820000 116.430000  37.820000 116.600000 ;
      RECT  33.820000 126.980000  37.820000 127.150000 ;
      RECT  33.935000  85.540000  37.705000  95.920000 ;
      RECT  33.935000 116.600000  37.705000 126.980000 ;
      RECT  33.960000 173.630000  36.670000 173.800000 ;
      RECT  33.980000 163.120000  36.940000 163.290000 ;
      RECT  33.980000 164.680000  36.940000 164.850000 ;
      RECT  33.980000 167.800000  36.940000 167.970000 ;
      RECT  33.980000 169.360000  36.940000 169.530000 ;
      RECT  33.980000 170.920000  36.940000 171.090000 ;
      RECT  33.980000 172.480000  36.940000 172.650000 ;
      RECT  34.025000 132.010000  34.195000 141.970000 ;
      RECT  34.045000 192.515000  40.820000 195.580000 ;
      RECT  34.050000  73.725000  35.330000  76.640000 ;
      RECT  34.120000 148.630000  34.290000 151.500000 ;
      RECT  34.120000 151.840000  34.290000 154.735000 ;
      RECT  34.170000  98.970000  34.340000 104.350000 ;
      RECT  34.170000 108.170000  34.340000 113.550000 ;
      RECT  34.185000 230.095000  34.355000 245.125000 ;
      RECT  34.230000 163.900000  36.940000 164.070000 ;
      RECT  34.230000 165.460000  36.940000 165.630000 ;
      RECT  34.230000 167.020000  36.940000 167.190000 ;
      RECT  34.230000 168.580000  36.940000 168.750000 ;
      RECT  34.230000 170.140000  41.700000 170.310000 ;
      RECT  34.230000 171.700000  36.940000 171.870000 ;
      RECT  34.250000 142.270000  47.840000 142.440000 ;
      RECT  34.325000 229.695000  35.775000 229.865000 ;
      RECT  34.420000 130.030000  37.135000 130.200000 ;
      RECT  34.420000 130.910000  37.135000 131.080000 ;
      RECT  34.495000  44.150000  34.955000  45.835000 ;
      RECT  34.495000  45.835000  36.205000  46.165000 ;
      RECT  34.495000  46.165000  34.955000  46.705000 ;
      RECT  34.495000  46.705000  63.260000  46.875000 ;
      RECT  34.535000  63.565000  44.940000  66.305000 ;
      RECT  34.540000 156.345000  35.070000 156.875000 ;
      RECT  34.550000  58.790000  64.075000  58.960000 ;
      RECT  34.550000  58.960000  44.940000  59.000000 ;
      RECT  34.550000  59.000000  34.760000  60.035000 ;
      RECT  34.550000  60.035000  44.940000  62.505000 ;
      RECT  34.550000  62.505000  34.760000  63.355000 ;
      RECT  34.550000  63.355000  44.940000  63.565000 ;
      RECT  34.570000  99.140000  34.740000 103.890000 ;
      RECT  34.570000 108.340000  34.740000 113.090000 ;
      RECT  34.680000 178.435000  35.210000 178.605000 ;
      RECT  34.795000  98.800000  38.795000  98.970000 ;
      RECT  34.795000 104.350000  38.795000 104.520000 ;
      RECT  34.795000 108.000000  38.795000 108.170000 ;
      RECT  34.795000 113.550000  38.795000 113.720000 ;
      RECT  34.800000 176.430000  34.970000 178.435000 ;
      RECT  34.800000 178.605000  34.970000 183.390000 ;
      RECT  34.900000 148.790000  35.070000 151.500000 ;
      RECT  34.900000 152.010000  35.070000 154.720000 ;
      RECT  34.900000 155.975000  35.070000 156.345000 ;
      RECT  34.900000 156.875000  35.070000 158.880000 ;
      RECT  34.910000 214.380000  35.080000 217.340000 ;
      RECT  34.965000 230.175000  35.135000 245.125000 ;
      RECT  35.135000 172.890000  38.520000 172.935000 ;
      RECT  35.135000 172.935000  39.625000 173.060000 ;
      RECT  35.300000 218.195000  36.680000 218.200000 ;
      RECT  35.320000  59.795000  35.490000  60.035000 ;
      RECT  35.380000   6.305000  35.550000  10.035000 ;
      RECT  35.380000  13.175000  35.550000  14.955000 ;
      RECT  35.380000  14.955000  35.970000  15.125000 ;
      RECT  35.380000  15.125000  35.550000  15.735000 ;
      RECT  35.380000  15.735000  35.970000  15.905000 ;
      RECT  35.380000  15.905000  35.550000  17.515000 ;
      RECT  35.380000  17.515000  35.970000  17.685000 ;
      RECT  35.380000  17.685000  35.550000  18.295000 ;
      RECT  35.380000  18.295000  35.970000  18.465000 ;
      RECT  35.380000  18.465000  35.550000  27.115000 ;
      RECT  35.380000 177.270000  35.550000 179.980000 ;
      RECT  35.380000 180.740000  35.550000 183.450000 ;
      RECT  35.415000  43.610000  36.095000  44.275000 ;
      RECT  35.415000  44.575000  36.085000  45.535000 ;
      RECT  35.415000 171.285000  38.520000 171.455000 ;
      RECT  35.480000 147.880000  35.650000 159.775000 ;
      RECT  35.490000 209.185000  36.680000 213.440000 ;
      RECT  35.490000 213.950000  36.680000 218.195000 ;
      RECT  35.545000  59.435000  43.825000  59.605000 ;
      RECT  35.605000  59.390000  43.690000  59.435000 ;
      RECT  35.605000 176.600000  42.115000 176.770000 ;
      RECT  35.605000 183.620000  42.115000 183.790000 ;
      RECT  35.700000  47.905000  41.215000  47.935000 ;
      RECT  35.700000  47.935000  41.925000  48.105000 ;
      RECT  35.700000  48.105000  35.875000  49.955000 ;
      RECT  35.700000  49.955000  41.925000  50.125000 ;
      RECT  35.700000  50.125000  41.810000  50.135000 ;
      RECT  35.745000 230.095000  35.915000 245.125000 ;
      RECT  35.770000   5.945000  38.480000   6.115000 ;
      RECT  35.770000  10.225000  38.480000  10.395000 ;
      RECT  35.770000  11.505000  38.480000  11.675000 ;
      RECT  35.770000  12.785000  38.480000  12.955000 ;
      RECT  35.770000  14.065000  38.480000  14.235000 ;
      RECT  35.770000  15.345000  38.480000  15.515000 ;
      RECT  35.770000  16.625000  38.480000  16.795000 ;
      RECT  35.770000  17.905000  38.480000  18.075000 ;
      RECT  35.770000  19.185000  38.480000  19.355000 ;
      RECT  35.770000  20.465000  38.480000  20.635000 ;
      RECT  35.770000  21.745000  38.480000  21.915000 ;
      RECT  35.770000  23.025000  38.480000  23.195000 ;
      RECT  35.770000  27.305000  38.480000  27.475000 ;
      RECT  35.895000  73.985000  38.305000  74.155000 ;
      RECT  35.895000  74.155000  36.065000  80.160000 ;
      RECT  35.895000  80.160000  38.305000  80.360000 ;
      RECT  36.035000   5.930000  38.480000   5.945000 ;
      RECT  36.035000   6.115000  38.480000  10.225000 ;
      RECT  36.035000  10.395000  38.480000  11.505000 ;
      RECT  36.035000  11.675000  38.480000  12.785000 ;
      RECT  36.075000  48.640000  36.245000  49.420000 ;
      RECT  36.080000 186.695000  40.820000 192.515000 ;
      RECT  36.095000  21.915000  38.480000  23.025000 ;
      RECT  36.095000  23.195000  38.480000  27.305000 ;
      RECT  36.145000  51.195000  44.705000  54.460000 ;
      RECT  36.145000  54.460000  63.260000  54.670000 ;
      RECT  36.145000  54.670000  36.355000  58.790000 ;
      RECT  36.145000  98.970000  37.440000 104.350000 ;
      RECT  36.145000 108.170000  37.440000 113.550000 ;
      RECT  36.160000 177.270000  36.330000 183.450000 ;
      RECT  36.210000 163.885000  36.740000 163.900000 ;
      RECT  36.225000 229.275000  36.395000 245.690000 ;
      RECT  36.305000 132.010000  36.475000 141.860000 ;
      RECT  36.375000  74.405000  36.545000  79.155000 ;
      RECT  36.465000  48.415000  41.215000  48.585000 ;
      RECT  36.465000  48.945000  41.215000  49.115000 ;
      RECT  36.465000  49.475000  41.215000  49.645000 ;
      RECT  36.510000  49.465000  41.215000  49.475000 ;
      RECT  36.705000 230.095000  36.875000 245.125000 ;
      RECT  36.720000  79.665000  37.530000  79.835000 ;
      RECT  36.785000  55.340000  62.640000  58.050000 ;
      RECT  36.845000 229.695000  38.295000 229.865000 ;
      RECT  36.940000 177.270000  37.110000 179.980000 ;
      RECT  36.940000 180.740000  37.110000 183.450000 ;
      RECT  37.010000  54.980000  62.410000  55.150000 ;
      RECT  37.075000 176.770000  42.115000 176.800000 ;
      RECT  37.110000 163.175000  37.440000 163.730000 ;
      RECT  37.110000 164.815000  39.565000 164.985000 ;
      RECT  37.110000 164.985000  37.280000 165.090000 ;
      RECT  37.110000 167.560000  37.280000 167.665000 ;
      RECT  37.110000 167.665000  39.265000 167.835000 ;
      RECT  37.130000 205.070000  40.565000 205.100000 ;
      RECT  37.130000 206.330000  40.820000 217.345000 ;
      RECT  37.140000 168.020000  37.470000 168.575000 ;
      RECT  37.460000 164.305000  41.700000 164.575000 ;
      RECT  37.485000 230.175000  37.655000 245.125000 ;
      RECT  37.490000 177.270000  37.660000 179.980000 ;
      RECT  37.490000 180.740000  37.660000 183.450000 ;
      RECT  37.530000 217.345000  40.820000 223.550000 ;
      RECT  37.590000 166.965000  37.760000 166.990000 ;
      RECT  37.590000 166.990000  38.520000 167.160000 ;
      RECT  37.590000 167.160000  37.760000 167.495000 ;
      RECT  37.590000 168.930000  37.760000 169.160000 ;
      RECT  37.590000 169.160000  38.520000 169.330000 ;
      RECT  37.590000 169.330000  37.760000 169.595000 ;
      RECT  37.590000 170.540000  42.270000 170.740000 ;
      RECT  37.590000 170.740000  37.760000 171.115000 ;
      RECT  37.590000 173.460000  37.760000 173.790000 ;
      RECT  37.655000  74.405000  37.825000  79.155000 ;
      RECT  37.850000 162.645000  38.050000 163.965000 ;
      RECT  37.850000 163.965000  38.520000 164.135000 ;
      RECT  37.850000 168.515000  38.520000 168.685000 ;
      RECT  37.870000 168.155000  38.040000 168.515000 ;
      RECT  37.875000  85.710000  39.195000  95.620000 ;
      RECT  37.875000 116.900000  39.195000 126.810000 ;
      RECT  38.060000 169.635000  38.440000 169.970000 ;
      RECT  38.135000  74.155000  38.305000  80.160000 ;
      RECT  38.180000   3.925000  38.875000   4.595000 ;
      RECT  38.190000 170.915000  38.520000 171.285000 ;
      RECT  38.190000 171.455000  38.520000 171.555000 ;
      RECT  38.190000 171.555000  39.355000 171.885000 ;
      RECT  38.190000 173.060000  39.625000 173.265000 ;
      RECT  38.190000 173.265000  38.520000 173.850000 ;
      RECT  38.265000 230.095000  38.435000 245.125000 ;
      RECT  38.270000 177.270000  38.440000 180.150000 ;
      RECT  38.270000 180.150000  41.560000 180.570000 ;
      RECT  38.270000 180.570000  38.440000 183.450000 ;
      RECT  38.320000 174.080000  42.270000 174.280000 ;
      RECT  38.320000 174.280000  38.520000 174.405000 ;
      RECT  38.550000 162.215000  60.940000 162.385000 ;
      RECT  38.580000 147.070000  39.470000 147.600000 ;
      RECT  38.580000 148.365000  39.470000 149.940000 ;
      RECT  38.580000 150.570000  39.470000 151.610000 ;
      RECT  38.580000 152.350000  39.470000 154.015000 ;
      RECT  38.585000 132.010000  38.755000 141.970000 ;
      RECT  38.600000 145.100000  39.450000 147.070000 ;
      RECT  38.600000 147.600000  39.450000 148.365000 ;
      RECT  38.600000 149.940000  39.450000 150.570000 ;
      RECT  38.600000 151.610000  39.450000 152.350000 ;
      RECT  38.600000 154.015000  39.450000 159.150000 ;
      RECT  38.600000 159.150000  90.225000 160.000000 ;
      RECT  38.600000 160.000000  88.140000 160.220000 ;
      RECT  38.680000 169.635000  41.700000 169.970000 ;
      RECT  38.705000 172.575000  41.065000 172.745000 ;
      RECT  38.745000 229.275000  38.920000 245.690000 ;
      RECT  38.810000  31.485000  38.980000  32.155000 ;
      RECT  38.810000  32.665000  38.980000  33.335000 ;
      RECT  38.810000  33.845000  38.980000  34.515000 ;
      RECT  38.810000  35.025000  38.980000  35.695000 ;
      RECT  38.850000  99.140000  39.020000 103.890000 ;
      RECT  38.850000 108.340000  39.020000 113.090000 ;
      RECT  38.945000 172.075000  39.615000 172.405000 ;
      RECT  38.990000 162.845000  41.700000 163.015000 ;
      RECT  38.990000 163.625000  41.700000 163.795000 ;
      RECT  38.990000 165.185000  41.700000 165.355000 ;
      RECT  38.990000 166.070000  41.700000 166.135000 ;
      RECT  38.990000 166.515000  41.700000 166.580000 ;
      RECT  38.990000 167.295000  41.700000 167.465000 ;
      RECT  38.990000 168.075000  42.580000 168.245000 ;
      RECT  38.990000 168.855000  41.700000 169.025000 ;
      RECT  38.990000 170.310000  41.700000 170.355000 ;
      RECT  38.990000 171.065000  41.700000 171.235000 ;
      RECT  38.990000 173.585000  41.700000 173.755000 ;
      RECT  38.990000 174.465000  42.610000 174.635000 ;
      RECT  39.030000   6.305000  39.200000  14.955000 ;
      RECT  39.030000  14.955000  39.620000  15.125000 ;
      RECT  39.030000  15.125000  39.200000  15.735000 ;
      RECT  39.030000  15.735000  39.620000  15.905000 ;
      RECT  39.030000  15.905000  39.200000  17.515000 ;
      RECT  39.030000  17.515000  39.620000  17.685000 ;
      RECT  39.030000  17.685000  39.200000  18.295000 ;
      RECT  39.030000  18.295000  39.620000  18.465000 ;
      RECT  39.030000  18.465000  39.200000  27.115000 ;
      RECT  39.050000 177.270000  39.220000 179.980000 ;
      RECT  39.050000 180.740000  39.220000 183.450000 ;
      RECT  39.075000  98.800000  43.075000  98.970000 ;
      RECT  39.075000 104.350000  43.075000 104.520000 ;
      RECT  39.075000 108.000000  43.075000 108.170000 ;
      RECT  39.075000 113.550000  43.075000 113.720000 ;
      RECT  39.250000  85.370000  43.250000  85.540000 ;
      RECT  39.250000  95.920000  43.250000  96.090000 ;
      RECT  39.250000 116.430000  43.250000 116.600000 ;
      RECT  39.250000 126.980000  43.250000 127.150000 ;
      RECT  39.365000  85.540000  43.135000  95.920000 ;
      RECT  39.365000 116.600000  43.005000 126.980000 ;
      RECT  39.420000   5.945000  42.130000   6.115000 ;
      RECT  39.420000  10.225000  42.130000  10.395000 ;
      RECT  39.420000  11.505000  42.130000  11.675000 ;
      RECT  39.420000  12.785000  42.130000  12.955000 ;
      RECT  39.420000  14.065000  42.130000  14.235000 ;
      RECT  39.420000  15.345000  42.130000  15.515000 ;
      RECT  39.420000  16.625000  42.130000  16.795000 ;
      RECT  39.420000  17.905000  42.130000  18.075000 ;
      RECT  39.420000  19.185000  42.130000  19.355000 ;
      RECT  39.420000  20.465000  42.130000  20.635000 ;
      RECT  39.420000  21.745000  42.130000  21.915000 ;
      RECT  39.420000  23.025000  42.130000  23.195000 ;
      RECT  39.420000  27.305000  42.130000  27.475000 ;
      RECT  39.600000  59.795000  39.770000  60.035000 ;
      RECT  39.660000 166.955000  46.915000 167.125000 ;
      RECT  39.690000  31.485000  39.860000  32.155000 ;
      RECT  39.690000  32.665000  39.860000  33.335000 ;
      RECT  39.690000  33.845000  39.860000  34.515000 ;
      RECT  39.690000  35.025000  39.860000  35.695000 ;
      RECT  39.735000 228.345000  40.485000 246.620000 ;
      RECT  39.830000 177.270000  40.000000 180.150000 ;
      RECT  39.830000 180.570000  40.000000 183.450000 ;
      RECT  39.845000 173.165000  40.015000 173.585000 ;
      RECT  39.855000   3.925000  40.630000   4.595000 ;
      RECT  39.940000 164.815000  46.915000 164.985000 ;
      RECT  40.110000  31.155000  50.000000  31.325000 ;
      RECT  40.110000  32.335000  50.000000  32.505000 ;
      RECT  40.110000  33.515000  50.000000  33.685000 ;
      RECT  40.110000  34.695000  50.000000  34.865000 ;
      RECT  40.110000  35.875000  50.000000  36.045000 ;
      RECT  40.215000 143.120000  40.385000 148.365000 ;
      RECT  40.215000 148.365000  43.865000 148.535000 ;
      RECT  40.215000 148.535000  40.385000 152.335000 ;
      RECT  40.215000 152.335000  43.865000 152.505000 ;
      RECT  40.215000 152.505000  40.385000 154.645000 ;
      RECT  40.215000 154.645000  43.865000 154.815000 ;
      RECT  40.215000 154.815000  40.385000 158.215000 ;
      RECT  40.215000 158.215000  48.575000 158.590000 ;
      RECT  40.330000 171.235000  40.500000 171.655000 ;
      RECT  40.375000   2.335000  40.905000   2.505000 ;
      RECT  40.385000   2.235000  40.895000   2.335000 ;
      RECT  40.385000   2.505000  40.895000   2.905000 ;
      RECT  40.395000 172.415000  41.065000 172.575000 ;
      RECT  40.425000  98.970000  41.720000 104.350000 ;
      RECT  40.425000 108.170000  41.720000 113.550000 ;
      RECT  40.610000 177.270000  40.780000 179.980000 ;
      RECT  40.610000 180.740000  40.780000 183.450000 ;
      RECT  40.825000 156.075000  43.820000 156.245000 ;
      RECT  40.825000 156.855000  43.535000 157.025000 ;
      RECT  40.825000 157.635000  43.535000 157.805000 ;
      RECT  40.855000 155.525000  43.865000 155.695000 ;
      RECT  40.865000 132.010000  41.035000 141.860000 ;
      RECT  40.865000 153.215000  43.865000 153.385000 ;
      RECT  41.000000 171.555000  41.405000 171.885000 ;
      RECT  41.000000 172.935000  41.405000 173.265000 ;
      RECT  41.030000 145.725000  43.865000 145.895000 ;
      RECT  41.085000 153.765000  43.865000 153.935000 ;
      RECT  41.115000 143.300000  45.865000 143.795000 ;
      RECT  41.115000 144.405000  46.255000 144.575000 ;
      RECT  41.155000 146.605000  43.865000 146.775000 ;
      RECT  41.155000 147.485000  43.865000 147.655000 ;
      RECT  41.155000 149.245000  43.865000 149.415000 ;
      RECT  41.155000 149.795000  43.865000 149.965000 ;
      RECT  41.155000 150.575000  44.255000 150.745000 ;
      RECT  41.155000 151.455000  43.865000 151.625000 ;
      RECT  41.235000 171.885000  41.405000 172.935000 ;
      RECT  41.255000  74.465000  87.720000  75.120000 ;
      RECT  41.255000  75.120000  42.110000  82.955000 ;
      RECT  41.255000  82.955000  87.720000  83.975000 ;
      RECT  41.390000 177.270000  41.560000 180.150000 ;
      RECT  41.390000 180.570000  41.560000 183.450000 ;
      RECT  41.580000 184.190000  44.535000 200.645000 ;
      RECT  41.580000 200.645000  45.520000 203.475000 ;
      RECT  41.580000 204.335000  45.520000 215.530000 ;
      RECT  41.580000 215.530000  45.375000 215.970000 ;
      RECT  41.580000 215.970000  42.430000 225.590000 ;
      RECT  41.580000 226.440000  42.430000 248.525000 ;
      RECT  41.580000 249.375000  42.430000 252.535000 ;
      RECT  41.580000 252.535000 175.920000 253.385000 ;
      RECT  41.755000  48.105000  41.925000  48.825000 ;
      RECT  41.755000  49.185000  41.925000  49.955000 ;
      RECT  41.780000  44.015000  42.310000  44.185000 ;
      RECT  41.780000  44.640000  42.310000  44.810000 ;
      RECT  41.780000  45.270000  42.310000  45.440000 ;
      RECT  41.790000  43.945000  42.300000  44.015000 ;
      RECT  41.790000  44.185000  42.300000  44.275000 ;
      RECT  41.790000  44.575000  42.300000  44.640000 ;
      RECT  41.790000  44.810000  42.300000  44.905000 ;
      RECT  41.790000  45.205000  42.300000  45.270000 ;
      RECT  41.790000  45.440000  42.300000  45.535000 ;
      RECT  41.920000 162.900000  42.190000 163.570000 ;
      RECT  41.920000 165.410000  42.190000 166.080000 ;
      RECT  41.945000  45.835000  62.940000  46.165000 ;
      RECT  41.985000   3.925000  42.670000   4.595000 ;
      RECT  42.020000 163.570000  42.190000 164.100000 ;
      RECT  42.100000 168.580000  42.270000 170.540000 ;
      RECT  42.100000 170.740000  42.270000 171.290000 ;
      RECT  42.100000 171.570000  42.270000 174.080000 ;
      RECT  42.170000 177.270000  42.340000 179.980000 ;
      RECT  42.170000 180.740000  42.340000 183.450000 ;
      RECT  42.440000 168.825000  42.610000 169.005000 ;
      RECT  42.440000 169.005000  45.530000 169.175000 ;
      RECT  42.440000 169.175000  42.610000 169.355000 ;
      RECT  42.440000 170.385000  42.610000 170.565000 ;
      RECT  42.440000 170.565000  45.530000 170.735000 ;
      RECT  42.440000 170.735000  42.610000 170.915000 ;
      RECT  42.440000 171.945000  42.610000 172.125000 ;
      RECT  42.440000 172.125000  45.530000 172.295000 ;
      RECT  42.440000 172.295000  42.610000 172.475000 ;
      RECT  42.440000 173.505000  42.610000 173.685000 ;
      RECT  42.440000 173.685000  45.530000 173.855000 ;
      RECT  42.440000 173.855000  42.610000 174.465000 ;
      RECT  42.460000 163.295000  46.915000 163.625000 ;
      RECT  42.460000 163.625000  43.040000 164.015000 ;
      RECT  42.460000 164.015000  46.915000 164.345000 ;
      RECT  42.460000 164.735000  46.915000 164.815000 ;
      RECT  42.460000 164.985000  46.915000 165.065000 ;
      RECT  42.460000 165.455000  46.915000 165.785000 ;
      RECT  42.460000 165.785000  43.040000 166.175000 ;
      RECT  42.460000 166.175000  46.915000 166.505000 ;
      RECT  42.460000 166.895000  46.915000 166.955000 ;
      RECT  42.460000 167.125000  46.915000 167.225000 ;
      RECT  42.510000 178.435000  43.040000 178.605000 ;
      RECT  42.565000   6.500000  42.850000   9.840000 ;
      RECT  42.565000  23.580000  42.850000  26.920000 ;
      RECT  42.680000   6.305000  42.850000   6.500000 ;
      RECT  42.680000   9.840000  42.850000  23.580000 ;
      RECT  42.680000  26.920000  42.850000  27.115000 ;
      RECT  42.750000 176.430000  42.920000 178.435000 ;
      RECT  42.750000 178.605000  42.920000 183.390000 ;
      RECT  42.820000 168.225000  48.865000 168.395000 ;
      RECT  42.820000 169.785000  48.865000 169.955000 ;
      RECT  42.820000 171.345000  48.865000 171.515000 ;
      RECT  42.820000 172.905000  48.865000 173.485000 ;
      RECT  42.820000 174.055000  48.865000 174.835000 ;
      RECT  42.855000  77.110000  43.055000  80.650000 ;
      RECT  42.870000  75.880000  85.820000  76.050000 ;
      RECT  42.870000  76.050000  43.040000  77.110000 ;
      RECT  42.870000  80.650000  43.040000  82.020000 ;
      RECT  42.870000  82.020000  85.820000  82.190000 ;
      RECT  43.130000  99.140000  43.300000 103.890000 ;
      RECT  43.130000 108.340000  43.300000 113.090000 ;
      RECT  43.145000 132.010000  43.315000 141.970000 ;
      RECT  43.185000 162.755000  59.495000 163.075000 ;
      RECT  43.200000   5.415000  43.370000  28.375000 ;
      RECT  43.210000  46.875000  44.705000  51.195000 ;
      RECT  43.305000  85.710000  43.475000  95.560000 ;
      RECT  43.305000 116.960000  43.475000 126.810000 ;
      RECT  43.355000  98.800000  47.355000  98.970000 ;
      RECT  43.355000 104.350000  47.355000 104.520000 ;
      RECT  43.355000 108.000000  47.355000 108.170000 ;
      RECT  43.355000 113.550000  47.355000 113.720000 ;
      RECT  43.435000  77.110000  43.635000  80.650000 ;
      RECT  43.450000  76.400000  43.620000  77.110000 ;
      RECT  43.450000  80.650000  43.620000  81.150000 ;
      RECT  43.465000  81.610000  44.175000  81.780000 ;
      RECT  43.485000 216.295000  51.300000 219.215000 ;
      RECT  43.485000 219.215000 172.950000 220.065000 ;
      RECT  43.485000 220.065000 140.900000 220.085000 ;
      RECT  43.485000 220.085000  47.855000 247.105000 ;
      RECT  43.485000 247.105000 165.290000 251.735000 ;
      RECT  43.485000 251.735000 164.155000 251.760000 ;
      RECT  43.530000  85.370000  47.530000  85.540000 ;
      RECT  43.530000  95.920000  47.530000  96.090000 ;
      RECT  43.530000 116.430000  47.530000 116.600000 ;
      RECT  43.530000 126.980000  47.530000 127.150000 ;
      RECT  43.645000  85.540000  47.415000  95.920000 ;
      RECT  43.645000 116.600000  47.285000 126.980000 ;
      RECT  43.665000 145.285000  44.255000 145.455000 ;
      RECT  43.685000 176.600000  90.225000 177.450000 ;
      RECT  43.685000 177.450000  44.535000 184.190000 ;
      RECT  43.725000 157.250000  44.255000 157.420000 ;
      RECT  43.850000  80.880000  44.020000  81.610000 ;
      RECT  43.870000   3.925000  44.525000   4.595000 ;
      RECT  43.880000  59.795000  44.050000  60.035000 ;
      RECT  44.035000 145.455000  44.255000 146.960000 ;
      RECT  44.035000 151.455000  44.565000 151.625000 ;
      RECT  44.085000 147.840000  44.255000 149.335000 ;
      RECT  44.085000 149.335000  44.795000 149.505000 ;
      RECT  44.085000 149.850000  44.255000 150.575000 ;
      RECT  44.085000 151.200000  44.255000 151.455000 ;
      RECT  44.085000 151.625000  44.255000 154.590000 ;
      RECT  44.085000 154.870000  44.795000 155.540000 ;
      RECT  44.085000 156.300000  44.255000 157.250000 ;
      RECT  44.085000 157.420000  44.255000 157.650000 ;
      RECT  44.205000   6.340000  44.375000  16.190000 ;
      RECT  44.205000  17.340000  44.375000  27.190000 ;
      RECT  44.230000  76.400000  44.400000  77.050000 ;
      RECT  44.230000  77.050000  44.435000  80.250000 ;
      RECT  44.230000  80.250000  44.400000  81.150000 ;
      RECT  44.265000 147.335000  44.795000 147.505000 ;
      RECT  44.455000  81.555000  49.295000  81.835000 ;
      RECT  44.455000 144.575000  46.255000 145.440000 ;
      RECT  44.540000   5.820000  45.210000   5.990000 ;
      RECT  44.540000  27.400000  45.210000  27.900000 ;
      RECT  44.600000 149.780000  44.795000 150.310000 ;
      RECT  44.610000 153.765000  45.140000 153.935000 ;
      RECT  44.625000 146.610000  44.795000 147.335000 ;
      RECT  44.625000 147.675000  44.795000 148.350000 ;
      RECT  44.625000 148.350000  45.155000 148.520000 ;
      RECT  44.625000 148.520000  44.795000 149.025000 ;
      RECT  44.625000 149.505000  44.795000 149.780000 ;
      RECT  44.625000 150.310000  44.795000 150.870000 ;
      RECT  44.625000 151.960000  44.795000 152.320000 ;
      RECT  44.625000 152.320000  45.215000 152.490000 ;
      RECT  44.625000 152.490000  44.795000 152.630000 ;
      RECT  44.625000 153.240000  44.795000 153.765000 ;
      RECT  44.625000 155.540000  44.795000 157.580000 ;
      RECT  44.705000  98.970000  46.000000 104.350000 ;
      RECT  44.705000 108.170000  46.000000 113.550000 ;
      RECT  44.770000  59.000000  44.940000  59.635000 ;
      RECT  44.770000  59.635000  46.120000  59.885000 ;
      RECT  44.770000  59.885000  44.940000  60.035000 ;
      RECT  44.770000  62.505000  44.940000  63.355000 ;
      RECT  45.015000 154.515000  48.065000 154.685000 ;
      RECT  45.015000 155.295000  47.725000 155.465000 ;
      RECT  45.015000 156.075000  48.065000 156.245000 ;
      RECT  45.015000 156.855000  47.725000 157.025000 ;
      RECT  45.015000 157.635000  48.065000 157.805000 ;
      RECT  45.070000 147.335000  48.575000 147.505000 ;
      RECT  45.220000 146.455000  48.055000 146.625000 ;
      RECT  45.220000 149.095000  48.055000 149.265000 ;
      RECT  45.220000 149.645000  48.055000 149.815000 ;
      RECT  45.300000 178.210000 160.800000 178.905000 ;
      RECT  45.300000 178.905000  95.640000 182.950000 ;
      RECT  45.300000 182.950000  46.440000 196.425000 ;
      RECT  45.300000 196.425000 172.950000 197.275000 ;
      RECT  45.300000 197.275000  51.300000 199.885000 ;
      RECT  45.305000  47.305000  62.640000  50.015000 ;
      RECT  45.305000  50.955000  62.640000  53.665000 ;
      RECT  45.345000 148.215000  48.055000 148.385000 ;
      RECT  45.345000 150.925000  48.575000 151.095000 ;
      RECT  45.345000 151.805000  48.055000 151.975000 ;
      RECT  45.345000 152.685000  48.575000 152.855000 ;
      RECT  45.345000 153.965000  48.055000 154.135000 ;
      RECT  45.370000  65.035000  46.080000  65.285000 ;
      RECT  45.385000   6.340000  45.555000  16.190000 ;
      RECT  45.385000  17.340000  45.555000  27.190000 ;
      RECT  45.425000 132.010000  45.595000 141.860000 ;
      RECT  45.495000  77.110000  45.695000  80.920000 ;
      RECT  45.510000  76.400000  45.680000  77.110000 ;
      RECT  45.510000  80.920000  45.680000  81.555000 ;
      RECT  45.590000  50.560000  62.410000  50.730000 ;
      RECT  45.630000  50.530000  62.355000  50.560000 ;
      RECT  45.720000   5.815000  46.390000   5.985000 ;
      RECT  45.720000  27.400000  46.390000  27.900000 ;
      RECT  45.730000 173.485000  48.865000 174.055000 ;
      RECT  45.830000  59.595000  46.040000  59.635000 ;
      RECT  45.830000  59.885000  46.040000  59.925000 ;
      RECT  45.830000  64.995000  46.000000  65.035000 ;
      RECT  45.830000  65.285000  46.000000  65.325000 ;
      RECT  45.990000 167.705000  60.940000 167.875000 ;
      RECT  46.055000   3.925000  46.600000   4.595000 ;
      RECT  46.085000 144.010000  46.255000 144.405000 ;
      RECT  46.280000 199.885000  51.300000 216.295000 ;
      RECT  46.535000 167.875000  48.865000 168.225000 ;
      RECT  46.535000 168.395000  48.865000 169.785000 ;
      RECT  46.535000 169.955000  48.865000 171.345000 ;
      RECT  46.535000 171.515000  48.865000 172.905000 ;
      RECT  46.565000   6.340000  46.735000  16.190000 ;
      RECT  46.565000  17.340000  46.735000  27.190000 ;
      RECT  46.625000 142.930000  47.155000 143.100000 ;
      RECT  46.625000 143.100000  46.795000 145.850000 ;
      RECT  46.775000  77.050000  46.975000  80.860000 ;
      RECT  46.790000  76.400000  46.960000  77.050000 ;
      RECT  46.790000  80.860000  46.960000  81.150000 ;
      RECT  46.920000  67.005000  47.630000  67.255000 ;
      RECT  47.045000 143.300000  48.055000 143.795000 ;
      RECT  47.045000 145.905000  48.055000 146.075000 ;
      RECT  47.165000 163.295000  55.535000 163.625000 ;
      RECT  47.165000 164.015000  55.535000 164.345000 ;
      RECT  47.165000 164.735000  55.535000 165.065000 ;
      RECT  47.165000 165.455000  55.535000 165.785000 ;
      RECT  47.165000 166.175000  55.535000 166.505000 ;
      RECT  47.165000 166.895000  55.535000 167.225000 ;
      RECT  47.200000 183.710000 121.065000 185.670000 ;
      RECT  47.200000 185.670000  48.050000 187.450000 ;
      RECT  47.200000 187.450000 101.370000 187.620000 ;
      RECT  47.200000 187.620000  48.050000 189.190000 ;
      RECT  47.200000 189.190000 101.370000 189.360000 ;
      RECT  47.200000 189.360000  48.050000 190.930000 ;
      RECT  47.200000 190.930000 101.370000 191.100000 ;
      RECT  47.200000 191.100000  48.050000 192.815000 ;
      RECT  47.200000 192.815000  80.130000 192.985000 ;
      RECT  47.200000 192.985000  67.620000 194.500000 ;
      RECT  47.200000 194.500000 101.370000 194.595000 ;
      RECT  47.200000 194.595000 158.850000 195.440000 ;
      RECT  47.200000 195.440000 114.160000 195.445000 ;
      RECT  47.335000   4.010000  70.680000   4.190000 ;
      RECT  47.335000   4.190000  47.515000   5.235000 ;
      RECT  47.335000   5.415000  47.515000  10.480000 ;
      RECT  47.335000  10.480000  70.680000  10.990000 ;
      RECT  47.335000  10.990000  47.515000  11.865000 ;
      RECT  47.335000  11.865000  48.280000  12.535000 ;
      RECT  47.335000  12.535000  47.515000  19.635000 ;
      RECT  47.335000  19.635000  48.280000  20.305000 ;
      RECT  47.335000  20.305000  47.515000  21.175000 ;
      RECT  47.335000  21.175000  70.680000  21.685000 ;
      RECT  47.335000  21.685000  47.515000  28.375000 ;
      RECT  47.380000  66.965000  47.550000  67.005000 ;
      RECT  47.380000  67.255000  47.550000  67.295000 ;
      RECT  47.410000  99.140000  47.580000 103.890000 ;
      RECT  47.410000 108.340000  47.580000 113.090000 ;
      RECT  47.585000  85.710000  48.905000  95.620000 ;
      RECT  47.585000 116.900000  48.905000 126.810000 ;
      RECT  47.615000  28.555000  70.645000  28.565000 ;
      RECT  47.635000  98.800000  51.635000  98.970000 ;
      RECT  47.635000 104.350000  51.635000 104.520000 ;
      RECT  47.635000 108.000000  51.635000 108.170000 ;
      RECT  47.635000 113.550000  51.635000 113.720000 ;
      RECT  47.705000 132.010000  47.875000 141.970000 ;
      RECT  47.805000  21.165000  69.605000  21.175000 ;
      RECT  47.805000  21.685000  69.605000  21.695000 ;
      RECT  47.895000 154.685000  48.065000 156.075000 ;
      RECT  47.895000 156.245000  48.065000 157.635000 ;
      RECT  48.055000  77.110000  48.255000  80.920000 ;
      RECT  48.070000  76.400000  48.240000  77.110000 ;
      RECT  48.070000  80.920000  48.240000  81.555000 ;
      RECT  48.075000  44.025000  48.605000  44.195000 ;
      RECT  48.075000  44.640000  48.605000  44.810000 ;
      RECT  48.075000  45.270000  48.605000  45.440000 ;
      RECT  48.085000  43.945000  48.595000  44.025000 ;
      RECT  48.085000  44.195000  48.595000  44.275000 ;
      RECT  48.085000  44.575000  48.595000  44.640000 ;
      RECT  48.085000  44.810000  48.595000  44.905000 ;
      RECT  48.085000  45.205000  48.595000  45.270000 ;
      RECT  48.085000  45.440000  48.595000  45.535000 ;
      RECT  48.110000  13.665000  48.280000  13.705000 ;
      RECT  48.110000  13.705000  48.700000  13.875000 ;
      RECT  48.110000  13.875000  48.280000  14.335000 ;
      RECT  48.110000  14.845000  48.280000  15.095000 ;
      RECT  48.110000  15.095000  48.810000  15.265000 ;
      RECT  48.110000  15.265000  48.280000  15.515000 ;
      RECT  48.110000  16.655000  48.585000  16.720000 ;
      RECT  48.110000  16.720000  49.115000  16.890000 ;
      RECT  48.110000  16.890000  48.585000  17.325000 ;
      RECT  48.110000  17.835000  48.280000  18.120000 ;
      RECT  48.110000  18.120000  48.810000  18.290000 ;
      RECT  48.110000  18.290000  48.280000  18.505000 ;
      RECT  48.160000   4.620000  48.810000   4.950000 ;
      RECT  48.160000   5.250000  48.810000   5.580000 ;
      RECT  48.160000   5.880000  48.810000   6.210000 ;
      RECT  48.160000   6.510000  48.810000   6.840000 ;
      RECT  48.160000   7.140000  48.810000   7.470000 ;
      RECT  48.160000   7.770000  48.810000   8.100000 ;
      RECT  48.160000   8.400000  48.810000   8.730000 ;
      RECT  48.160000   9.030000  48.810000   9.360000 ;
      RECT  48.160000   9.660000  48.810000   9.990000 ;
      RECT  48.160000  22.635000  48.810000  22.965000 ;
      RECT  48.160000  23.265000  48.810000  23.595000 ;
      RECT  48.160000  23.895000  48.810000  24.225000 ;
      RECT  48.160000  24.525000  48.810000  24.855000 ;
      RECT  48.160000  25.155000  48.810000  25.485000 ;
      RECT  48.160000  25.785000  48.810000  26.115000 ;
      RECT  48.160000  26.415000  48.810000  26.745000 ;
      RECT  48.160000  27.045000  48.810000  27.375000 ;
      RECT  48.160000  27.675000  48.810000  28.005000 ;
      RECT  48.240000 186.330000  48.410000 186.475000 ;
      RECT  48.240000 186.475000  48.425000 187.000000 ;
      RECT  48.240000 188.070000  48.410000 188.140000 ;
      RECT  48.240000 188.140000  48.425000 188.670000 ;
      RECT  48.240000 188.670000  48.410000 188.740000 ;
      RECT  48.240000 189.810000  48.410000 189.880000 ;
      RECT  48.240000 189.880000  48.425000 190.410000 ;
      RECT  48.240000 190.410000  48.410000 190.480000 ;
      RECT  48.240000 191.550000  48.410000 191.620000 ;
      RECT  48.240000 191.620000  48.425000 192.150000 ;
      RECT  48.240000 192.150000  48.410000 192.220000 ;
      RECT  48.255000 187.000000  48.425000 187.005000 ;
      RECT  48.405000 129.620000  48.575000 131.490000 ;
      RECT  48.405000 131.660000  48.575000 147.335000 ;
      RECT  48.405000 147.505000  48.575000 150.925000 ;
      RECT  48.405000 151.095000  48.575000 152.685000 ;
      RECT  48.405000 152.855000  48.575000 158.215000 ;
      RECT  48.500000  11.525000  58.390000  11.695000 ;
      RECT  48.500000  12.705000  58.390000  12.875000 ;
      RECT  48.500000  13.325000  58.390000  13.495000 ;
      RECT  48.500000  14.505000  58.390000  14.675000 ;
      RECT  48.500000  15.685000  58.390000  15.855000 ;
      RECT  48.500000  16.315000  58.390000  16.485000 ;
      RECT  48.500000  17.495000  58.390000  17.665000 ;
      RECT  48.500000  18.675000  58.390000  18.845000 ;
      RECT  48.500000  19.295000  58.390000  19.465000 ;
      RECT  48.500000  20.475000  58.390000  20.645000 ;
      RECT  48.630000 186.190000  63.580000 186.360000 ;
      RECT  48.630000 186.970000  63.580000 187.140000 ;
      RECT  48.630000 187.930000  63.580000 188.100000 ;
      RECT  48.630000 188.710000  63.580000 188.880000 ;
      RECT  48.630000 189.670000  63.580000 189.840000 ;
      RECT  48.630000 190.450000  63.580000 190.620000 ;
      RECT  48.630000 191.410000  63.580000 191.580000 ;
      RECT  48.630000 192.190000  63.580000 192.360000 ;
      RECT  48.760000  85.370000  52.960000  85.540000 ;
      RECT  48.760000  95.920000  52.960000  96.090000 ;
      RECT  48.855000 221.230000 139.285000 222.080000 ;
      RECT  48.855000 222.080000  49.705000 245.255000 ;
      RECT  48.855000 245.255000 139.285000 246.105000 ;
      RECT  48.960000 116.430000  52.960000 116.600000 ;
      RECT  48.960000 126.980000  52.960000 127.150000 ;
      RECT  48.985000  98.970000  50.280000 104.350000 ;
      RECT  48.985000 108.170000  50.280000 113.550000 ;
      RECT  49.075000  85.540000  52.845000  95.920000 ;
      RECT  49.075000 116.600000  52.845000 126.980000 ;
      RECT  49.305000 146.790000  50.195000 147.135000 ;
      RECT  49.305000 148.365000  50.195000 151.055000 ;
      RECT  49.305000 152.475000  50.195000 157.925000 ;
      RECT  49.335000  77.050000  49.535000  80.860000 ;
      RECT  49.340000 128.205000  49.990000 143.735000 ;
      RECT  49.340000 143.735000  90.225000 143.905000 ;
      RECT  49.340000 143.905000  50.190000 146.790000 ;
      RECT  49.340000 147.135000  50.190000 148.365000 ;
      RECT  49.340000 151.055000  50.190000 152.475000 ;
      RECT  49.340000 157.925000  50.190000 159.150000 ;
      RECT  49.350000  76.400000  49.520000  77.050000 ;
      RECT  49.350000  80.860000  49.520000  81.150000 ;
      RECT  49.575000  81.610000  50.300000  81.780000 ;
      RECT  49.625000 168.645000  61.085000 169.345000 ;
      RECT  49.625000 169.345000  50.325000 175.240000 ;
      RECT  49.625000 175.240000  61.085000 175.940000 ;
      RECT  49.990000  36.750000  51.470000  36.760000 ;
      RECT  50.115000  77.050000  50.315000  80.860000 ;
      RECT  50.130000  76.400000  50.300000  77.050000 ;
      RECT  50.130000  80.860000  50.300000  81.610000 ;
      RECT  50.400000  31.485000  50.570000  32.155000 ;
      RECT  50.400000  32.665000  50.570000  33.335000 ;
      RECT  50.400000  33.845000  50.570000  34.515000 ;
      RECT  50.400000  35.025000  50.570000  35.695000 ;
      RECT  50.470000 222.845000 137.670000 223.695000 ;
      RECT  50.470000 223.695000  51.320000 243.640000 ;
      RECT  50.470000 243.640000 137.670000 244.490000 ;
      RECT  50.680000  76.400000  50.850000  81.150000 ;
      RECT  50.905000  81.315000  51.290000  81.320000 ;
      RECT  50.905000  81.320000  53.745000  81.780000 ;
      RECT  50.905000  82.390000  51.435000  82.560000 ;
      RECT  50.955000 145.155000  86.525000 145.325000 ;
      RECT  50.955000 145.325000  51.125000 158.215000 ;
      RECT  50.955000 158.215000  86.525000 158.385000 ;
      RECT  51.020000  80.750000  51.290000  81.315000 ;
      RECT  51.085000 170.105000  59.625000 170.805000 ;
      RECT  51.085000 170.805000  51.785000 173.780000 ;
      RECT  51.085000 173.780000  59.625000 174.480000 ;
      RECT  51.300000  30.425000  51.470000  36.590000 ;
      RECT  51.460000  76.400000  51.630000  81.150000 ;
      RECT  51.495000 129.450000  87.790000 129.620000 ;
      RECT  51.495000 129.620000  51.665000 142.385000 ;
      RECT  51.525000 129.415000  87.730000 129.450000 ;
      RECT  51.535000 147.505000  51.705000 157.355000 ;
      RECT  51.690000  99.140000  51.860000 103.890000 ;
      RECT  51.690000 108.340000  51.860000 113.090000 ;
      RECT  51.800000  34.290000  71.625000  34.470000 ;
      RECT  51.800000  34.470000  51.980000  37.515000 ;
      RECT  51.800000  80.750000  52.070000  81.320000 ;
      RECT  51.890000 146.815000  54.260000 146.985000 ;
      RECT  51.915000  98.800000  55.915000  98.970000 ;
      RECT  51.915000 104.350000  55.915000 104.520000 ;
      RECT  51.915000 108.000000  55.915000 108.170000 ;
      RECT  51.915000 113.550000  55.915000 113.720000 ;
      RECT  52.070000 130.030000  52.400000 130.540000 ;
      RECT  52.070000 135.540000  53.030000 136.050000 ;
      RECT  52.070000 136.430000  52.400000 136.940000 ;
      RECT  52.070000 141.940000  53.030000 142.450000 ;
      RECT  52.090000 224.125000  62.090000 226.445000 ;
      RECT  52.090000 228.735000  62.090000 230.645000 ;
      RECT  52.090000 232.935000  62.090000 235.255000 ;
      RECT  52.090000 236.415000  62.090000 238.735000 ;
      RECT  52.090000 241.700000  62.090000 242.935000 ;
      RECT  52.150000 130.540000  52.320000 130.600000 ;
      RECT  52.150000 136.940000  52.320000 137.000000 ;
      RECT  52.240000  76.400000  52.410000  81.150000 ;
      RECT  52.460000  40.760000  54.485000  41.090000 ;
      RECT  52.460000  41.390000  54.485000  41.720000 ;
      RECT  52.460000  42.020000  54.485000  42.350000 ;
      RECT  52.460000  42.650000  53.130000  43.610000 ;
      RECT  52.480000 198.455000  79.190000 199.305000 ;
      RECT  52.480000 199.305000  53.790000 199.985000 ;
      RECT  52.480000 199.985000  54.010000 214.935000 ;
      RECT  52.480000 214.935000  53.790000 215.605000 ;
      RECT  52.480000 215.605000  79.190000 218.285000 ;
      RECT  52.580000  29.490000  52.750000  34.290000 ;
      RECT  52.580000  80.750000  52.850000  81.320000 ;
      RECT  52.585000  45.270000  53.115000  45.440000 ;
      RECT  52.595000  45.205000  53.105000  45.270000 ;
      RECT  52.595000  45.440000  53.105000  45.535000 ;
      RECT  52.655000 171.280000  58.050000 171.820000 ;
      RECT  52.655000 172.755000  58.050000 173.295000 ;
      RECT  52.700000 130.030000  53.660000 130.540000 ;
      RECT  52.700000 136.430000  53.660000 136.940000 ;
      RECT  52.715000 147.505000  52.885000 157.355000 ;
      RECT  52.785000   2.755000  53.315000   2.925000 ;
      RECT  52.805000   2.235000  53.315000   2.755000 ;
      RECT  53.015000  85.710000  53.865000  89.620000 ;
      RECT  53.015000  89.620000  53.905000  94.495000 ;
      RECT  53.015000  94.495000  53.865000  95.620000 ;
      RECT  53.015000 116.900000  53.865000 118.025000 ;
      RECT  53.015000 118.025000  53.905000 122.900000 ;
      RECT  53.015000 122.900000  53.865000 126.810000 ;
      RECT  53.020000  76.400000  53.190000  81.150000 ;
      RECT  53.060000  36.440000  80.710000  36.610000 ;
      RECT  53.060000  36.610000  53.345000  39.575000 ;
      RECT  53.265000  98.970000  54.560000 104.350000 ;
      RECT  53.265000 108.170000  54.560000 113.550000 ;
      RECT  53.265000 147.505000  53.435000 157.355000 ;
      RECT  53.330000  58.760000  64.075000  58.790000 ;
      RECT  53.330000  58.960000  64.075000  58.990000 ;
      RECT  53.330000 135.540000  54.290000 136.050000 ;
      RECT  53.330000 141.940000  54.290000 142.450000 ;
      RECT  53.360000  80.750000  53.630000  81.320000 ;
      RECT  53.625000  30.880000  56.195000  31.050000 ;
      RECT  53.625000  31.050000  53.795000  33.355000 ;
      RECT  53.625000  33.355000  56.195000  33.525000 ;
      RECT  53.695000  36.980000  54.505000  37.310000 ;
      RECT  53.695000  37.610000  54.485000  37.940000 ;
      RECT  53.695000  38.240000  54.485000  39.200000 ;
      RECT  53.695000  39.500000  54.485000  40.460000 ;
      RECT  53.695000  42.650000  54.490000  42.980000 ;
      RECT  53.695000  95.620000  53.865000  95.730000 ;
      RECT  53.695000 116.790000  53.865000 116.900000 ;
      RECT  53.800000  76.400000  53.970000  77.050000 ;
      RECT  53.800000  77.050000  53.980000  80.460000 ;
      RECT  53.800000  80.460000  53.970000  81.150000 ;
      RECT  53.960000 130.030000  54.920000 130.540000 ;
      RECT  53.960000 136.430000  54.920000 136.940000 ;
      RECT  54.065000 199.505000  56.905000 199.675000 ;
      RECT  54.065000 215.155000  56.905000 215.385000 ;
      RECT  54.130000  31.890000  54.300000  32.560000 ;
      RECT  54.350000  76.400000  54.520000  81.610000 ;
      RECT  54.350000  81.610000  55.455000  81.780000 ;
      RECT  54.370000  44.020000  54.900000  44.190000 ;
      RECT  54.370000  44.640000  54.900000  44.810000 ;
      RECT  54.380000  43.945000  54.890000  44.020000 ;
      RECT  54.380000  44.190000  54.890000  44.275000 ;
      RECT  54.380000  44.575000  54.890000  44.640000 ;
      RECT  54.380000  44.810000  54.890000  44.905000 ;
      RECT  54.445000 147.505000  54.615000 157.355000 ;
      RECT  54.550000  31.575000  55.560000  31.745000 ;
      RECT  54.550000  32.755000  55.560000  32.925000 ;
      RECT  54.590000 135.540000  55.550000 136.050000 ;
      RECT  54.590000 141.940000  55.550000 142.450000 ;
      RECT  54.620000 199.965000  54.790000 214.935000 ;
      RECT  55.165000 145.325000  55.335000 158.215000 ;
      RECT  55.205000  84.825000  55.375000  96.855000 ;
      RECT  55.205000 115.675000  55.375000 127.885000 ;
      RECT  55.220000 130.030000  56.180000 130.540000 ;
      RECT  55.220000 136.430000  56.180000 136.940000 ;
      RECT  55.400000 199.985000  55.570000 214.985000 ;
      RECT  55.530000   8.400000  56.180000   8.730000 ;
      RECT  55.530000  23.895000  56.180000  24.225000 ;
      RECT  55.565000 146.390000  56.095000 146.560000 ;
      RECT  55.630000  76.400000  55.800000  81.150000 ;
      RECT  55.765000 146.560000  56.095000 147.065000 ;
      RECT  55.765000 151.465000  56.095000 152.865000 ;
      RECT  55.765000 157.265000  56.725000 157.775000 ;
      RECT  55.785000 163.295000  60.940000 163.625000 ;
      RECT  55.785000 164.015000  60.240000 164.345000 ;
      RECT  55.785000 164.735000  60.240000 165.065000 ;
      RECT  55.785000 165.455000  60.940000 165.785000 ;
      RECT  55.785000 166.175000  60.240000 166.505000 ;
      RECT  55.785000 166.895000  60.240000 167.225000 ;
      RECT  55.850000 135.540000  56.810000 136.050000 ;
      RECT  55.850000 141.940000  56.810000 142.450000 ;
      RECT  55.925000  81.610000  56.735000  81.780000 ;
      RECT  55.970000  99.140000  56.140000 103.890000 ;
      RECT  55.970000 108.340000  56.140000 113.090000 ;
      RECT  56.025000  31.050000  56.195000  33.355000 ;
      RECT  56.085000  81.180000  56.615000  81.610000 ;
      RECT  56.180000 199.965000  56.350000 214.935000 ;
      RECT  56.195000  98.800000  60.195000  98.970000 ;
      RECT  56.195000 104.350000  60.195000 104.520000 ;
      RECT  56.195000 108.000000  60.195000 108.170000 ;
      RECT  56.195000 113.550000  60.195000 113.720000 ;
      RECT  56.395000 146.555000  57.355000 147.065000 ;
      RECT  56.395000 151.465000  56.725000 152.865000 ;
      RECT  56.480000 130.030000  57.440000 130.540000 ;
      RECT  56.480000 136.430000  57.440000 136.940000 ;
      RECT  56.530000   7.770000  57.180000   8.100000 ;
      RECT  56.530000  24.525000  57.180000  24.855000 ;
      RECT  56.595000  43.945000  61.910000  44.275000 ;
      RECT  56.595000  44.575000  61.910000  44.905000 ;
      RECT  56.675000  88.500000  57.565000  93.375000 ;
      RECT  56.675000 119.145000  57.565000 124.020000 ;
      RECT  56.685000 163.075000  58.295000 163.125000 ;
      RECT  56.715000  85.710000  57.565000  88.500000 ;
      RECT  56.715000  93.375000  57.565000  95.620000 ;
      RECT  56.715000  95.620000  56.885000  95.730000 ;
      RECT  56.715000 116.790000  56.885000 116.900000 ;
      RECT  56.715000 116.900000  57.565000 119.145000 ;
      RECT  56.715000 124.020000  57.565000 126.810000 ;
      RECT  56.910000  76.400000  57.080000  81.150000 ;
      RECT  56.930000   9.030000  57.580000   9.360000 ;
      RECT  56.930000  23.265000  57.580000  23.595000 ;
      RECT  56.960000   8.400000  57.610000   8.730000 ;
      RECT  56.960000  23.895000  57.610000  24.225000 ;
      RECT  56.960000 199.985000  58.150000 214.935000 ;
      RECT  57.025000 151.465000  57.355000 152.865000 ;
      RECT  57.025000 157.265000  57.985000 157.775000 ;
      RECT  57.075000 199.305000  58.035000 199.985000 ;
      RECT  57.075000 214.935000  58.035000 215.605000 ;
      RECT  57.095000  45.270000  57.625000  45.440000 ;
      RECT  57.105000  45.205000  57.615000  45.270000 ;
      RECT  57.105000  45.440000  57.615000  45.535000 ;
      RECT  57.110000 135.540000  58.070000 136.050000 ;
      RECT  57.110000 141.940000  58.070000 142.450000 ;
      RECT  57.205000  81.610000  58.015000  81.780000 ;
      RECT  57.365000  81.180000  57.895000  81.610000 ;
      RECT  57.545000  98.970000  58.840000 104.350000 ;
      RECT  57.545000 108.170000  58.840000 113.550000 ;
      RECT  57.595000  29.490000  57.765000  34.290000 ;
      RECT  57.620000  85.370000  61.620000  85.540000 ;
      RECT  57.620000  95.920000  61.620000  96.090000 ;
      RECT  57.620000 116.430000  61.750000 116.600000 ;
      RECT  57.620000 126.980000  61.750000 127.150000 ;
      RECT  57.655000 146.555000  58.745000 146.560000 ;
      RECT  57.655000 146.560000  58.615000 147.065000 ;
      RECT  57.655000 151.465000  57.985000 152.865000 ;
      RECT  57.735000  85.540000  61.505000  95.920000 ;
      RECT  57.735000 116.600000  61.505000 126.980000 ;
      RECT  57.740000 130.030000  58.700000 130.540000 ;
      RECT  57.740000 136.430000  58.700000 136.940000 ;
      RECT  58.075000  37.610000  80.190000  37.940000 ;
      RECT  58.075000  38.240000  80.190000  38.570000 ;
      RECT  58.075000  38.870000  80.190000  39.200000 ;
      RECT  58.075000  39.500000  80.190000  39.830000 ;
      RECT  58.075000  40.130000  80.190000  40.460000 ;
      RECT  58.075000  40.760000  80.190000  41.090000 ;
      RECT  58.075000  41.390000  80.190000  41.720000 ;
      RECT  58.075000  42.020000  80.190000  42.350000 ;
      RECT  58.190000  76.400000  58.360000  81.150000 ;
      RECT  58.205000 199.505000  61.045000 199.675000 ;
      RECT  58.205000 215.155000  61.050000 215.385000 ;
      RECT  58.215000 146.390000  58.745000 146.555000 ;
      RECT  58.220000 171.625000  58.630000 172.950000 ;
      RECT  58.230000  13.705000  58.930000  13.875000 ;
      RECT  58.230000  15.285000  58.930000  15.455000 ;
      RECT  58.230000  16.720000  58.930000  16.890000 ;
      RECT  58.230000  18.120000  58.930000  18.290000 ;
      RECT  58.285000 151.465000  58.615000 152.865000 ;
      RECT  58.285000 157.265000  59.245000 157.775000 ;
      RECT  58.370000 135.540000  59.330000 136.050000 ;
      RECT  58.370000 141.940000  59.330000 142.450000 ;
      RECT  58.485000  81.610000  59.295000  81.780000 ;
      RECT  58.645000  81.180000  59.175000  81.610000 ;
      RECT  58.760000  13.665000  58.930000  13.705000 ;
      RECT  58.760000  13.875000  58.930000  15.285000 ;
      RECT  58.760000  15.455000  58.930000  15.515000 ;
      RECT  58.760000  16.655000  58.930000  16.720000 ;
      RECT  58.760000  16.890000  58.930000  18.120000 ;
      RECT  58.760000  18.290000  58.930000  18.505000 ;
      RECT  58.760000 199.965000  58.930000 214.935000 ;
      RECT  58.780000  37.055000  59.310000  37.225000 ;
      RECT  58.780000  42.755000  59.310000  42.925000 ;
      RECT  58.865000 244.490000 137.510000 244.520000 ;
      RECT  58.915000 146.555000  59.875000 147.065000 ;
      RECT  58.915000 151.465000  59.245000 152.865000 ;
      RECT  58.915000 170.805000  59.625000 173.780000 ;
      RECT  58.930000   7.140000  59.580000   7.470000 ;
      RECT  58.930000  25.155000  59.580000  25.485000 ;
      RECT  59.000000 130.030000  59.960000 130.540000 ;
      RECT  59.000000 136.430000  59.960000 136.940000 ;
      RECT  59.225000  30.880000  61.845000  31.050000 ;
      RECT  59.275000  31.050000  59.445000  33.355000 ;
      RECT  59.275000  33.355000  61.845000  33.525000 ;
      RECT  59.300000  13.665000  59.470000  13.725000 ;
      RECT  59.300000  13.725000  60.000000  13.895000 ;
      RECT  59.300000  13.895000  59.470000  14.915000 ;
      RECT  59.300000  14.915000  60.000000  15.085000 ;
      RECT  59.300000  15.085000  59.470000  15.515000 ;
      RECT  59.300000  16.655000  59.470000  16.710000 ;
      RECT  59.300000  16.710000  60.000000  16.880000 ;
      RECT  59.300000  16.880000  59.470000  18.275000 ;
      RECT  59.300000  18.275000  60.000000  18.445000 ;
      RECT  59.300000  18.445000  59.470000  18.505000 ;
      RECT  59.470000  76.400000  59.640000  81.150000 ;
      RECT  59.540000 199.985000  59.710000 214.985000 ;
      RECT  59.545000 151.465000  59.875000 152.865000 ;
      RECT  59.545000 157.265000  60.505000 157.775000 ;
      RECT  59.630000 135.540000  60.590000 136.050000 ;
      RECT  59.630000 141.940000  60.590000 142.450000 ;
      RECT  59.660000 164.345000  60.240000 164.735000 ;
      RECT  59.660000 166.505000  60.240000 166.895000 ;
      RECT  59.765000  81.610000  60.575000  81.780000 ;
      RECT  59.810000  31.890000  59.980000  32.560000 ;
      RECT  59.840000  11.525000  69.730000  11.695000 ;
      RECT  59.840000  12.705000  69.730000  12.875000 ;
      RECT  59.840000  13.325000  69.730000  13.495000 ;
      RECT  59.840000  14.505000  69.730000  14.675000 ;
      RECT  59.840000  15.685000  69.730000  15.855000 ;
      RECT  59.840000  16.315000  69.730000  16.485000 ;
      RECT  59.840000  17.495000  69.730000  17.665000 ;
      RECT  59.840000  18.675000  69.730000  18.845000 ;
      RECT  59.840000  19.295000  69.730000  19.465000 ;
      RECT  59.840000  20.475000  69.730000  20.645000 ;
      RECT  59.925000  81.180000  60.455000  81.610000 ;
      RECT  60.175000 146.555000  61.265000 146.560000 ;
      RECT  60.175000 146.560000  61.135000 147.065000 ;
      RECT  60.175000 151.465000  60.505000 152.865000 ;
      RECT  60.220000   7.770000  60.870000   7.850000 ;
      RECT  60.220000   7.850000  60.950000   8.020000 ;
      RECT  60.220000   8.020000  60.870000   8.100000 ;
      RECT  60.220000  24.525000  60.870000  24.605000 ;
      RECT  60.220000  24.605000  60.950000  24.775000 ;
      RECT  60.220000  24.775000  60.870000  24.855000 ;
      RECT  60.230000  31.575000  61.240000  31.745000 ;
      RECT  60.230000  32.755000  61.240000  32.925000 ;
      RECT  60.250000  99.140000  60.420000 103.890000 ;
      RECT  60.250000 108.340000  60.420000 113.090000 ;
      RECT  60.260000 130.030000  61.220000 130.540000 ;
      RECT  60.260000 136.430000  61.220000 136.940000 ;
      RECT  60.320000 199.965000  60.490000 214.935000 ;
      RECT  60.385000 169.345000  61.085000 175.240000 ;
      RECT  60.390000   8.480000  60.980000   8.650000 ;
      RECT  60.390000  23.975000  60.980000  24.145000 ;
      RECT  60.470000   8.400000  60.980000   8.480000 ;
      RECT  60.470000   8.650000  60.980000   8.730000 ;
      RECT  60.470000  23.895000  60.980000  23.975000 ;
      RECT  60.470000  24.145000  60.980000  24.225000 ;
      RECT  60.475000  98.800000  64.475000  98.970000 ;
      RECT  60.475000 104.350000  64.475000 104.520000 ;
      RECT  60.475000 108.000000  64.475000 108.170000 ;
      RECT  60.475000 113.550000  64.475000 113.720000 ;
      RECT  60.640000 130.540000  60.810000 130.600000 ;
      RECT  60.640000 136.940000  60.810000 137.000000 ;
      RECT  60.735000 146.390000  61.265000 146.555000 ;
      RECT  60.750000  76.400000  60.920000  81.150000 ;
      RECT  60.770000 162.385000  60.940000 163.295000 ;
      RECT  60.770000 163.625000  60.940000 165.455000 ;
      RECT  60.770000 165.785000  60.940000 167.705000 ;
      RECT  60.805000 151.465000  61.135000 152.865000 ;
      RECT  60.805000 157.265000  61.765000 157.775000 ;
      RECT  60.890000 135.540000  61.850000 136.050000 ;
      RECT  60.890000 141.940000  61.850000 142.450000 ;
      RECT  60.930000   6.510000  61.580000   6.840000 ;
      RECT  60.930000  25.785000  61.580000  26.115000 ;
      RECT  61.045000  81.610000  61.855000  81.780000 ;
      RECT  61.100000 199.985000  62.290000 214.935000 ;
      RECT  61.120000  45.205000  61.510000  45.245000 ;
      RECT  61.120000  45.245000  61.910000  45.495000 ;
      RECT  61.120000  45.495000  61.510000  45.535000 ;
      RECT  61.205000  81.180000  61.735000  81.610000 ;
      RECT  61.215000 199.305000  62.175000 199.985000 ;
      RECT  61.220000 214.935000  62.175000 215.605000 ;
      RECT  61.240000  44.275000  61.910000  44.575000 ;
      RECT  61.360000   8.400000  61.530000   8.480000 ;
      RECT  61.360000   8.480000  61.950000   8.650000 ;
      RECT  61.360000   8.650000  61.530000   8.730000 ;
      RECT  61.360000   9.030000  62.010000   9.360000 ;
      RECT  61.360000  23.265000  62.010000  23.595000 ;
      RECT  61.360000  23.895000  61.530000  23.975000 ;
      RECT  61.360000  23.975000  61.950000  24.145000 ;
      RECT  61.360000  24.145000  61.530000  24.225000 ;
      RECT  61.435000 146.555000  62.395000 147.065000 ;
      RECT  61.435000 151.465000  61.765000 152.865000 ;
      RECT  61.520000 130.030000  62.480000 130.540000 ;
      RECT  61.520000 136.430000  62.480000 136.940000 ;
      RECT  61.675000  31.050000  61.845000  33.355000 ;
      RECT  61.675000  85.710000  62.995000  95.620000 ;
      RECT  61.675000 116.900000  62.995000 126.810000 ;
      RECT  61.685000  65.805000  62.395000  66.055000 ;
      RECT  61.700000   8.400000  61.870000   8.480000 ;
      RECT  61.700000   8.650000  61.870000   8.730000 ;
      RECT  61.700000  23.895000  61.870000  23.975000 ;
      RECT  61.700000  24.145000  61.870000  24.225000 ;
      RECT  61.715000   1.885000  62.525000   2.985000 ;
      RECT  61.745000 160.220000  62.595000 176.600000 ;
      RECT  61.765000  65.765000  61.940000  65.805000 ;
      RECT  61.765000  66.055000  61.940000  66.095000 ;
      RECT  61.825000  98.970000  63.120000 104.350000 ;
      RECT  61.825000 108.170000  63.120000 113.550000 ;
      RECT  61.960000   6.510000  62.610000   6.840000 ;
      RECT  61.960000  25.785000  62.610000  26.115000 ;
      RECT  62.030000  76.400000  62.200000  81.150000 ;
      RECT  62.065000 151.465000  62.395000 152.865000 ;
      RECT  62.065000 157.265000  63.025000 157.775000 ;
      RECT  62.150000 135.540000  63.110000 136.050000 ;
      RECT  62.150000 141.940000  63.110000 142.450000 ;
      RECT  62.180000  42.650000  80.190000  42.980000 ;
      RECT  62.245000  36.980000  80.190000  37.310000 ;
      RECT  62.325000  81.610000  63.135000  81.780000 ;
      RECT  62.345000 199.505000  65.185000 199.675000 ;
      RECT  62.345000 215.155000  65.185000 215.385000 ;
      RECT  62.440000 223.865000  63.235000 224.035000 ;
      RECT  62.440000 224.035000  62.805000 233.745000 ;
      RECT  62.485000  81.180000  63.015000  81.610000 ;
      RECT  62.540000 237.925000  63.505000 239.225000 ;
      RECT  62.635000  43.350000  80.710000  43.520000 ;
      RECT  62.635000  43.520000  62.940000  45.835000 ;
      RECT  62.635000  46.165000  62.940000  46.610000 ;
      RECT  62.635000  46.610000  63.260000  46.705000 ;
      RECT  62.645000  29.490000  62.815000  34.290000 ;
      RECT  62.695000 146.390000  63.225000 146.560000 ;
      RECT  62.695000 146.560000  63.025000 147.065000 ;
      RECT  62.695000 151.465000  63.025000 152.865000 ;
      RECT  62.730000 239.805000  64.600000 242.540000 ;
      RECT  62.730000 242.540000  89.595000 243.460000 ;
      RECT  62.760000 243.460000  89.595000 243.640000 ;
      RECT  62.780000 130.030000  63.740000 130.540000 ;
      RECT  62.780000 136.430000  63.740000 136.940000 ;
      RECT  62.900000 199.965000  63.070000 214.935000 ;
      RECT  62.975000 224.205000  63.965000 224.735000 ;
      RECT  62.975000 224.735000  63.505000 237.925000 ;
      RECT  63.050000  46.875000  63.260000  54.460000 ;
      RECT  63.050000  54.670000  63.260000  58.760000 ;
      RECT  63.050000  85.370000  67.050000  85.540000 ;
      RECT  63.050000  95.920000  67.050000  96.090000 ;
      RECT  63.050000 116.430000  67.050000 116.600000 ;
      RECT  63.050000 126.980000  67.050000 127.150000 ;
      RECT  63.165000  85.540000  66.935000  95.920000 ;
      RECT  63.165000 116.600000  66.935000 126.980000 ;
      RECT  63.310000  76.400000  63.480000  81.150000 ;
      RECT  63.355000 161.460000  88.445000 162.310000 ;
      RECT  63.355000 162.310000  64.205000 174.990000 ;
      RECT  63.355000 174.990000  88.445000 175.840000 ;
      RECT  63.395000 145.325000  63.985000 158.215000 ;
      RECT  63.405000 223.865000  63.965000 224.205000 ;
      RECT  63.410000 135.540000  64.370000 136.050000 ;
      RECT  63.410000 141.940000  64.370000 142.450000 ;
      RECT  63.585000  30.880000  66.155000  31.050000 ;
      RECT  63.585000  31.050000  63.755000  33.355000 ;
      RECT  63.585000  33.355000  66.155000  33.525000 ;
      RECT  63.605000  81.610000  64.415000  81.780000 ;
      RECT  63.680000 199.985000  63.850000 214.985000 ;
      RECT  63.750000 224.905000  63.920000 230.570000 ;
      RECT  63.750000 230.570000  64.600000 239.805000 ;
      RECT  63.765000  81.180000  64.295000  81.610000 ;
      RECT  63.845000  58.990000  64.075000  68.100000 ;
      RECT  64.040000 130.030000  65.000000 130.540000 ;
      RECT  64.040000 136.430000  65.000000 136.940000 ;
      RECT  64.100000  31.890000  64.270000  32.560000 ;
      RECT  64.160000  51.410000  66.730000  54.780000 ;
      RECT  64.160000  54.780000 110.720000  55.295000 ;
      RECT  64.160000  55.295000  92.285000  55.645000 ;
      RECT  64.160000  55.645000  77.280000  56.075000 ;
      RECT  64.160000  56.075000  65.660000  58.085000 ;
      RECT  64.160000 223.865000  64.695000 224.035000 ;
      RECT  64.160000 224.035000  64.585000 224.760000 ;
      RECT  64.160000 224.760000  64.690000 230.315000 ;
      RECT  64.345000 186.190000  79.375000 186.360000 ;
      RECT  64.345000 186.970000  79.375000 187.140000 ;
      RECT  64.345000 187.930000  79.295000 188.100000 ;
      RECT  64.345000 188.710000  79.375000 188.880000 ;
      RECT  64.345000 189.670000  79.295000 189.840000 ;
      RECT  64.345000 190.450000  79.375000 190.620000 ;
      RECT  64.345000 191.410000  79.295000 191.580000 ;
      RECT  64.345000 192.190000  79.375000 192.360000 ;
      RECT  64.375000 146.750000  64.545000 156.600000 ;
      RECT  64.445000 166.450000  64.615000 170.850000 ;
      RECT  64.460000 199.965000  64.630000 214.935000 ;
      RECT  64.520000  31.575000  65.530000  31.745000 ;
      RECT  64.520000  32.755000  65.530000  32.925000 ;
      RECT  64.530000  99.140000  64.700000 103.890000 ;
      RECT  64.530000 108.340000  64.700000 113.090000 ;
      RECT  64.560000  44.300000  94.960000  44.470000 ;
      RECT  64.560000  44.470000  64.730000  50.440000 ;
      RECT  64.560000  50.440000  67.085000  50.610000 ;
      RECT  64.590000  76.400000  64.760000  81.150000 ;
      RECT  64.600000 157.010000  72.880000 157.180000 ;
      RECT  64.670000 135.540000  65.630000 136.050000 ;
      RECT  64.670000 141.940000  65.630000 142.450000 ;
      RECT  64.715000 146.360000  68.485000 146.530000 ;
      RECT  64.730000   7.770000  65.380000   8.100000 ;
      RECT  64.730000   8.400000  65.380000   8.730000 ;
      RECT  64.730000   9.030000  65.380000   9.360000 ;
      RECT  64.730000  23.265000  65.380000  23.595000 ;
      RECT  64.730000  23.895000  65.380000  24.225000 ;
      RECT  64.730000  24.525000  65.380000  24.855000 ;
      RECT  64.755000  98.800000  68.755000  98.970000 ;
      RECT  64.755000 104.350000  68.755000 104.520000 ;
      RECT  64.755000 108.000000  68.755000 108.170000 ;
      RECT  64.755000 113.550000  68.755000 113.720000 ;
      RECT  64.755000 224.260000  65.285000 224.590000 ;
      RECT  64.800000 199.675000  65.070000 215.155000 ;
      RECT  64.860000 224.590000  65.190000 240.725000 ;
      RECT  64.885000  81.610000  65.695000  81.780000 ;
      RECT  65.045000  81.180000  65.575000  81.610000 ;
      RECT  65.080000 162.480000  75.080000 165.195000 ;
      RECT  65.080000 172.105000  75.080000 174.820000 ;
      RECT  65.140000  44.820000  65.310000  48.355000 ;
      RECT  65.140000  48.355000  65.670000  48.525000 ;
      RECT  65.140000  48.525000  65.310000  49.570000 ;
      RECT  65.240000 199.985000  66.430000 214.935000 ;
      RECT  65.300000 130.030000  66.260000 130.540000 ;
      RECT  65.300000 136.430000  66.260000 136.940000 ;
      RECT  65.355000 199.305000  66.315000 199.985000 ;
      RECT  65.355000 214.935000  66.315000 215.605000 ;
      RECT  65.360000 226.750000  65.990000 228.050000 ;
      RECT  65.360000 234.660000  65.990000 235.960000 ;
      RECT  65.360000 237.100000  65.695000 238.400000 ;
      RECT  65.415000  50.080000  68.125000  50.250000 ;
      RECT  65.460000 228.830000  76.630000 229.680000 ;
      RECT  65.460000 229.680000  65.990000 232.355000 ;
      RECT  65.460000 232.355000  76.630000 232.985000 ;
      RECT  65.460000 233.170000  65.990000 234.660000 ;
      RECT  65.475000  50.610000  67.085000  50.665000 ;
      RECT  65.490000  58.085000  65.660000  69.665000 ;
      RECT  65.490000  69.665000  78.330000  69.835000 ;
      RECT  65.525000 224.340000  66.055000 224.510000 ;
      RECT  65.525000 224.510000  65.990000 226.750000 ;
      RECT  65.525000 238.400000  65.695000 239.795000 ;
      RECT  65.525000 239.795000  66.055000 239.965000 ;
      RECT  65.525000 240.135000  77.310000 240.705000 ;
      RECT  65.730000  47.970000  66.260000  48.140000 ;
      RECT  65.760000   7.770000  66.410000   8.100000 ;
      RECT  65.760000   8.400000  66.410000   8.730000 ;
      RECT  65.760000   9.030000  66.410000   9.360000 ;
      RECT  65.760000  23.265000  66.410000  23.595000 ;
      RECT  65.760000  23.895000  66.410000  24.225000 ;
      RECT  65.760000  24.525000  66.410000  24.855000 ;
      RECT  65.870000  76.400000  66.040000  81.150000 ;
      RECT  65.920000  44.820000  66.090000  47.970000 ;
      RECT  65.920000  48.140000  66.090000  49.570000 ;
      RECT  65.930000 135.540000  66.890000 136.050000 ;
      RECT  65.930000 141.940000  66.890000 142.450000 ;
      RECT  65.985000  31.050000  66.155000  33.355000 ;
      RECT  66.105000  98.970000  67.400000 104.350000 ;
      RECT  66.105000 108.170000  67.400000 113.550000 ;
      RECT  66.160000 225.160000  76.160000 227.480000 ;
      RECT  66.160000 230.445000  76.160000 232.185000 ;
      RECT  66.160000 235.150000  76.160000 237.910000 ;
      RECT  66.160000 240.875000  76.160000 242.110000 ;
      RECT  66.165000  81.610000  66.975000  81.780000 ;
      RECT  66.225000 239.845000  77.310000 240.135000 ;
      RECT  66.255000 224.260000  75.985000 224.590000 ;
      RECT  66.315000 232.985000  76.630000 233.560000 ;
      RECT  66.315000 233.560000 136.095000 234.410000 ;
      RECT  66.320000  61.640000  66.490000  64.350000 ;
      RECT  66.325000  81.180000  66.855000  81.610000 ;
      RECT  66.485000  57.285000  66.655000  59.995000 ;
      RECT  66.485000 199.505000  69.325000 199.675000 ;
      RECT  66.485000 215.155000  69.325000 215.385000 ;
      RECT  66.525000  48.355000  67.055000  48.525000 ;
      RECT  66.560000 130.030000  67.520000 130.540000 ;
      RECT  66.560000 136.430000  67.520000 136.940000 ;
      RECT  66.600000 199.675000  66.870000 215.155000 ;
      RECT  66.700000  44.820000  66.870000  48.355000 ;
      RECT  66.700000  48.525000  66.870000  49.570000 ;
      RECT  66.710000  61.250000  67.380000  61.420000 ;
      RECT  66.780000  61.235000  67.310000  61.250000 ;
      RECT  66.905000  56.500000  67.575000  56.670000 ;
      RECT  66.945000  29.490000  67.115000  34.290000 ;
      RECT  67.040000 199.965000  67.210000 214.935000 ;
      RECT  67.105000  85.710000  67.275000  95.560000 ;
      RECT  67.105000 116.960000  67.275000 126.810000 ;
      RECT  67.140000  51.720000  67.310000  54.780000 ;
      RECT  67.150000  76.400000  67.320000  81.150000 ;
      RECT  67.190000 135.540000  68.150000 136.050000 ;
      RECT  67.190000 141.940000  68.150000 142.450000 ;
      RECT  67.275000  50.250000  68.125000  51.000000 ;
      RECT  67.275000  51.000000  68.790000  51.170000 ;
      RECT  67.290000  47.970000  67.820000  48.140000 ;
      RECT  67.330000  85.370000  71.330000  85.540000 ;
      RECT  67.330000  95.920000  71.330000  96.090000 ;
      RECT  67.330000 116.430000  71.330000 116.600000 ;
      RECT  67.330000 126.980000  71.330000 127.150000 ;
      RECT  67.445000  81.610000  68.255000  81.780000 ;
      RECT  67.445000  85.540000  71.215000  95.920000 ;
      RECT  67.445000 116.600000  71.215000 126.980000 ;
      RECT  67.480000  44.820000  67.650000  47.970000 ;
      RECT  67.480000  48.140000  67.650000  49.570000 ;
      RECT  67.600000  61.640000  67.770000  64.350000 ;
      RECT  67.605000  81.180000  68.135000  81.610000 ;
      RECT  67.765000  57.285000  67.935000  59.995000 ;
      RECT  67.820000 130.030000  68.780000 130.540000 ;
      RECT  67.820000 136.430000  68.780000 136.940000 ;
      RECT  67.820000 199.985000  67.990000 214.985000 ;
      RECT  67.830000  52.180000  68.360000  52.350000 ;
      RECT  67.985000  30.880000  70.555000  31.050000 ;
      RECT  67.985000  31.050000  68.155000  33.355000 ;
      RECT  67.985000  33.355000  70.555000  33.525000 ;
      RECT  67.990000  61.250000  68.660000  61.420000 ;
      RECT  68.020000  51.720000  68.190000  52.180000 ;
      RECT  68.020000  52.350000  68.190000  54.430000 ;
      RECT  68.060000  61.235000  68.590000  61.250000 ;
      RECT  68.090000  48.355000  68.620000  48.525000 ;
      RECT  68.130000 193.685000  68.690000 193.855000 ;
      RECT  68.180000 193.605000  68.690000 193.685000 ;
      RECT  68.180000 193.855000  68.690000 193.935000 ;
      RECT  68.185000  56.500000  68.855000  56.670000 ;
      RECT  68.260000  44.820000  68.430000  48.355000 ;
      RECT  68.260000  48.525000  68.430000  49.570000 ;
      RECT  68.430000  76.400000  68.600000  81.150000 ;
      RECT  68.450000 135.540000  69.410000 136.050000 ;
      RECT  68.450000 141.940000  69.410000 142.450000 ;
      RECT  68.515000  31.890000  68.685000  32.560000 ;
      RECT  68.530000   9.660000  69.180000   9.990000 ;
      RECT  68.530000  22.635000  69.180000  22.965000 ;
      RECT  68.555000  50.095000  71.305000  50.250000 ;
      RECT  68.555000  50.250000  71.245000  50.265000 ;
      RECT  68.595000  50.080000  71.305000  50.095000 ;
      RECT  68.600000 199.965000  68.770000 214.935000 ;
      RECT  68.655000 146.750000  68.825000 156.600000 ;
      RECT  68.725000  81.610000  69.535000  81.780000 ;
      RECT  68.810000  99.140000  68.980000 103.890000 ;
      RECT  68.810000 108.340000  68.980000 113.090000 ;
      RECT  68.870000  47.555000  69.400000  47.725000 ;
      RECT  68.880000  61.640000  69.050000  64.350000 ;
      RECT  68.885000  81.180000  69.415000  81.610000 ;
      RECT  68.900000  51.720000  69.070000  54.780000 ;
      RECT  68.935000  31.575000  69.945000  31.745000 ;
      RECT  68.935000  32.755000  69.945000  32.925000 ;
      RECT  68.985000  13.665000  70.120000  14.335000 ;
      RECT  68.995000 146.360000  72.765000 146.530000 ;
      RECT  69.040000  44.820000  69.210000  47.555000 ;
      RECT  69.040000  47.725000  69.210000  49.570000 ;
      RECT  69.045000  57.285000  69.215000  59.995000 ;
      RECT  69.080000 130.030000  69.410000 130.540000 ;
      RECT  69.080000 136.430000  69.410000 136.940000 ;
      RECT  69.110000  98.800000  69.760000  98.970000 ;
      RECT  69.110000 104.350000  69.760000 104.520000 ;
      RECT  69.110000 108.000000  69.760000 108.170000 ;
      RECT  69.110000 113.550000  69.760000 113.720000 ;
      RECT  69.130000   7.770000  69.780000   8.100000 ;
      RECT  69.130000   9.030000  69.780000   9.360000 ;
      RECT  69.130000  23.265000  69.780000  23.595000 ;
      RECT  69.130000  24.525000  69.780000  24.855000 ;
      RECT  69.160000 130.540000  69.330000 130.600000 ;
      RECT  69.160000 136.940000  69.330000 137.000000 ;
      RECT  69.190000   8.480000  69.920000   8.650000 ;
      RECT  69.190000  23.975000  69.920000  24.145000 ;
      RECT  69.190000  98.970000  69.360000 104.350000 ;
      RECT  69.190000 108.170000  69.360000 113.550000 ;
      RECT  69.200000  50.265000  70.550000  51.170000 ;
      RECT  69.270000   8.400000  69.920000   8.480000 ;
      RECT  69.270000   8.650000  69.920000   8.730000 ;
      RECT  69.270000  23.895000  69.920000  23.975000 ;
      RECT  69.270000  24.145000  69.920000  24.225000 ;
      RECT  69.300000   4.620000  69.980000   4.950000 ;
      RECT  69.300000  27.675000  69.980000  28.005000 ;
      RECT  69.330000   5.250000  69.980000   5.580000 ;
      RECT  69.330000   5.880000  69.980000   6.210000 ;
      RECT  69.330000   6.510000  69.980000   6.840000 ;
      RECT  69.330000  25.785000  69.980000  26.115000 ;
      RECT  69.330000  26.415000  69.980000  26.745000 ;
      RECT  69.330000  27.045000  69.980000  27.375000 ;
      RECT  69.380000 199.985000  70.570000 214.935000 ;
      RECT  69.495000 199.305000  70.455000 199.985000 ;
      RECT  69.495000 214.935000  70.455000 215.605000 ;
      RECT  69.530000  15.020000  70.120000  15.190000 ;
      RECT  69.530000  16.710000  70.120000  16.880000 ;
      RECT  69.530000  18.085000  70.120000  18.255000 ;
      RECT  69.590000  52.180000  70.120000  52.350000 ;
      RECT  69.590000  98.970000  69.760000 101.080000 ;
      RECT  69.590000 101.080000  69.770000 101.970000 ;
      RECT  69.590000 101.970000  69.760000 104.350000 ;
      RECT  69.590000 108.170000  69.760000 110.280000 ;
      RECT  69.590000 110.280000  69.770000 111.170000 ;
      RECT  69.590000 111.170000  69.760000 113.550000 ;
      RECT  69.650000  48.355000  70.180000  48.525000 ;
      RECT  69.710000  76.400000  69.880000  81.150000 ;
      RECT  69.780000  51.720000  69.950000  52.180000 ;
      RECT  69.780000  52.350000  69.950000  54.430000 ;
      RECT  69.820000  44.820000  69.990000  48.355000 ;
      RECT  69.820000  48.525000  69.990000  49.570000 ;
      RECT  69.840000 130.030000  70.170000 130.540000 ;
      RECT  69.840000 135.540000  70.800000 136.050000 ;
      RECT  69.840000 136.430000  70.170000 136.940000 ;
      RECT  69.840000 141.940000  70.800000 142.450000 ;
      RECT  69.920000 130.540000  70.090000 130.600000 ;
      RECT  69.920000 136.940000  70.090000 137.000000 ;
      RECT  69.950000  11.865000  70.680000  12.535000 ;
      RECT  69.950000  14.845000  70.120000  15.020000 ;
      RECT  69.950000  15.190000  70.120000  15.515000 ;
      RECT  69.950000  16.680000  70.120000  16.710000 ;
      RECT  69.950000  16.880000  70.120000  17.350000 ;
      RECT  69.950000  17.860000  70.120000  18.085000 ;
      RECT  69.950000  18.255000  70.120000  18.530000 ;
      RECT  69.950000  19.635000  70.680000  20.305000 ;
      RECT  70.005000  81.610000  70.815000  81.780000 ;
      RECT  70.105000  58.795000  70.275000  68.685000 ;
      RECT  70.165000  81.180000  70.695000  81.610000 ;
      RECT  70.170000  98.560000  70.340000 104.760000 ;
      RECT  70.170000 107.760000  70.340000 113.960000 ;
      RECT  70.385000  31.050000  70.555000  33.355000 ;
      RECT  70.430000  47.555000  70.960000  47.725000 ;
      RECT  70.455000  58.375000  71.125000  58.545000 ;
      RECT  70.455000  69.085000  71.125000  69.255000 ;
      RECT  70.470000 130.030000  71.430000 130.540000 ;
      RECT  70.470000 136.430000  71.430000 136.940000 ;
      RECT  70.500000   4.190000  70.680000  10.480000 ;
      RECT  70.500000  10.990000  70.680000  11.865000 ;
      RECT  70.500000  12.535000  70.680000  19.635000 ;
      RECT  70.500000  20.305000  70.680000  21.175000 ;
      RECT  70.500000  21.685000  70.680000  28.375000 ;
      RECT  70.600000  44.820000  70.770000  47.555000 ;
      RECT  70.600000  47.725000  70.770000  49.570000 ;
      RECT  70.625000 199.505000  73.465000 199.675000 ;
      RECT  70.625000 215.155000  73.465000 215.385000 ;
      RECT  70.660000  51.720000  70.830000  54.780000 ;
      RECT  70.960000  50.660000  72.310000  51.170000 ;
      RECT  70.990000  76.400000  71.160000  81.150000 ;
      RECT  71.020000  48.355000  71.550000  48.525000 ;
      RECT  71.100000 135.540000  72.060000 136.050000 ;
      RECT  71.100000 141.940000  72.060000 142.450000 ;
      RECT  71.180000 199.965000  71.350000 214.935000 ;
      RECT  71.285000  58.795000  71.455000  68.685000 ;
      RECT  71.285000  81.610000  72.095000  81.780000 ;
      RECT  71.350000  52.180000  71.880000  52.350000 ;
      RECT  71.380000  44.820000  71.550000  48.355000 ;
      RECT  71.380000  48.525000  71.550000  49.570000 ;
      RECT  71.385000  85.710000  72.705000  95.620000 ;
      RECT  71.385000 116.900000  72.705000 126.810000 ;
      RECT  71.445000   0.930000  71.625000  25.605000 ;
      RECT  71.445000  25.605000  72.025000  26.000000 ;
      RECT  71.445000  26.000000  71.625000  29.320000 ;
      RECT  71.445000  29.490000  71.625000  34.290000 ;
      RECT  71.445000  81.180000  71.975000  81.610000 ;
      RECT  71.540000  51.720000  71.710000  52.180000 ;
      RECT  71.540000  52.350000  71.710000  54.430000 ;
      RECT  71.585000  97.145000  71.755000 106.160000 ;
      RECT  71.585000 106.360000  71.755000 115.375000 ;
      RECT  71.605000  50.250000  78.650000  50.265000 ;
      RECT  71.605000  50.265000  72.310000  50.660000 ;
      RECT  71.635000  58.375000  72.305000  58.545000 ;
      RECT  71.635000  69.085000  72.305000  69.255000 ;
      RECT  71.640000  50.095000  78.805000  50.250000 ;
      RECT  71.675000  50.080000  78.805000  50.095000 ;
      RECT  71.730000 130.030000  72.690000 130.540000 ;
      RECT  71.730000 136.430000  72.690000 136.940000 ;
      RECT  71.930000  44.470000  72.100000  49.570000 ;
      RECT  71.960000 199.985000  72.130000 214.985000 ;
      RECT  72.270000  76.400000  72.440000  81.150000 ;
      RECT  72.360000 135.540000  73.320000 136.050000 ;
      RECT  72.360000 141.940000  73.320000 142.450000 ;
      RECT  72.420000  51.720000  72.590000  54.780000 ;
      RECT  72.465000  58.795000  72.635000  68.685000 ;
      RECT  72.480000  50.440000  79.050000  50.610000 ;
      RECT  72.565000  81.610000  73.375000  81.780000 ;
      RECT  72.620000  50.610000  78.910000  50.665000 ;
      RECT  72.640000  47.555000  73.170000  47.725000 ;
      RECT  72.725000  81.180000  73.255000  81.610000 ;
      RECT  72.740000 199.965000  72.910000 214.935000 ;
      RECT  72.755000  51.000000  77.505000  51.170000 ;
      RECT  72.760000  85.370000  76.760000  85.540000 ;
      RECT  72.760000  95.920000  76.760000  96.090000 ;
      RECT  72.760000 116.430000  76.760000 116.600000 ;
      RECT  72.760000 126.980000  76.760000 127.150000 ;
      RECT  72.810000  44.820000  72.980000  47.555000 ;
      RECT  72.810000  47.725000  72.980000  49.570000 ;
      RECT  72.815000  58.375000  73.485000  58.545000 ;
      RECT  72.815000  69.085000  73.485000  69.255000 ;
      RECT  72.875000  85.540000  76.645000  95.920000 ;
      RECT  72.875000 116.600000  76.645000 126.980000 ;
      RECT  72.935000 146.750000  73.105000 156.600000 ;
      RECT  72.990000 130.030000  73.950000 130.540000 ;
      RECT  72.990000 136.430000  73.950000 136.940000 ;
      RECT  73.110000  51.810000  73.640000  51.980000 ;
      RECT  73.130000  98.390000  87.790000  98.560000 ;
      RECT  73.130000 104.770000  87.780000 104.940000 ;
      RECT  73.130000 107.580000  87.780000 107.750000 ;
      RECT  73.130000 113.960000  87.790000 114.130000 ;
      RECT  73.160000 157.010000  77.160000 157.180000 ;
      RECT  73.170000  99.140000  73.340000 104.360000 ;
      RECT  73.170000 104.360000  74.395000 104.530000 ;
      RECT  73.170000 108.340000  73.340000 113.550000 ;
      RECT  73.170000 113.550000  74.395000 113.720000 ;
      RECT  73.300000  51.720000  73.470000  51.810000 ;
      RECT  73.300000  51.980000  73.470000  54.430000 ;
      RECT  73.315000 146.360000  77.045000 146.530000 ;
      RECT  73.350000   4.670000  78.510000   4.885000 ;
      RECT  73.350000   4.885000  73.520000  28.535000 ;
      RECT  73.350000  28.535000  78.510000  28.705000 ;
      RECT  73.520000 199.985000  74.710000 214.935000 ;
      RECT  73.550000  76.400000  73.720000  81.150000 ;
      RECT  73.620000 135.540000  74.580000 136.050000 ;
      RECT  73.620000 141.940000  74.580000 142.450000 ;
      RECT  73.635000 199.305000  74.595000 199.985000 ;
      RECT  73.635000 214.935000  74.595000 215.605000 ;
      RECT  73.645000  58.795000  73.815000  68.685000 ;
      RECT  73.690000  44.470000  73.860000  49.570000 ;
      RECT  73.780000 104.940000  73.950000 107.580000 ;
      RECT  73.845000  81.610000  74.655000  81.780000 ;
      RECT  73.850000  28.705000  78.510000  29.870000 ;
      RECT  73.850000  29.870000  74.990000  30.380000 ;
      RECT  73.980000   5.610000  74.150000  10.010000 ;
      RECT  73.980000  21.015000  74.150000  25.470000 ;
      RECT  73.980000  25.470000  75.380000  25.640000 ;
      RECT  73.995000  58.375000  74.665000  58.545000 ;
      RECT  73.995000  69.085000  74.665000  69.255000 ;
      RECT  74.005000  81.180000  74.535000  81.610000 ;
      RECT  74.180000  51.720000  74.350000  54.780000 ;
      RECT  74.250000 130.030000  75.210000 130.540000 ;
      RECT  74.250000 136.430000  75.210000 136.940000 ;
      RECT  74.360000 105.455000  74.530000 106.770000 ;
      RECT  74.370000   5.385000  75.380000   5.555000 ;
      RECT  74.370000   6.165000  75.380000   6.335000 ;
      RECT  74.370000   6.945000  75.380000   7.115000 ;
      RECT  74.370000   7.725000  75.380000   7.895000 ;
      RECT  74.370000   8.505000  75.380000   8.675000 ;
      RECT  74.370000   9.285000  75.380000   9.455000 ;
      RECT  74.370000  10.065000  75.380000  10.235000 ;
      RECT  74.370000  14.725000  75.380000  14.895000 ;
      RECT  74.370000  15.185000  75.380000  15.355000 ;
      RECT  74.370000  15.705000  75.380000  15.875000 ;
      RECT  74.370000  16.165000  75.380000  16.335000 ;
      RECT  74.370000  17.085000  75.380000  17.255000 ;
      RECT  74.370000  17.545000  75.380000  17.715000 ;
      RECT  74.370000  18.065000  75.380000  18.235000 ;
      RECT  74.370000  18.525000  75.380000  18.695000 ;
      RECT  74.370000  20.790000  75.380000  20.960000 ;
      RECT  74.370000  21.570000  75.380000  21.740000 ;
      RECT  74.370000  22.350000  75.380000  22.520000 ;
      RECT  74.370000  23.130000  75.380000  23.300000 ;
      RECT  74.370000  23.910000  75.380000  24.080000 ;
      RECT  74.370000  24.690000  75.380000  24.860000 ;
      RECT  74.400000  47.555000  74.930000  47.725000 ;
      RECT  74.445000 100.235000  74.620000 103.890000 ;
      RECT  74.445000 103.890000  74.615000 104.005000 ;
      RECT  74.450000  99.140000  74.620000 100.235000 ;
      RECT  74.450000 108.340000  74.620000 113.205000 ;
      RECT  74.460000  12.625000  75.590000  12.795000 ;
      RECT  74.460000  13.705000  75.130000  13.875000 ;
      RECT  74.460000  26.700000  75.130000  26.870000 ;
      RECT  74.460000  27.780000  75.590000  27.950000 ;
      RECT  74.570000  44.820000  74.740000  47.555000 ;
      RECT  74.570000  47.725000  74.740000  49.570000 ;
      RECT  74.700000 106.950000  75.370000 107.120000 ;
      RECT  74.765000 199.505000  77.605000 199.675000 ;
      RECT  74.765000 215.155000  77.605000 215.385000 ;
      RECT  74.825000  58.795000  74.995000  68.685000 ;
      RECT  74.830000  76.400000  75.000000  81.150000 ;
      RECT  74.840000 104.360000  84.470000 104.530000 ;
      RECT  74.840000 113.550000  84.470000 113.720000 ;
      RECT  74.875000  51.810000  75.405000  51.980000 ;
      RECT  74.880000 135.540000  75.840000 136.050000 ;
      RECT  74.880000 141.940000  75.840000 142.450000 ;
      RECT  75.060000  51.720000  75.230000  51.810000 ;
      RECT  75.060000  51.980000  75.230000  54.430000 ;
      RECT  75.125000  81.610000  75.935000  81.780000 ;
      RECT  75.285000  81.180000  75.815000  81.610000 ;
      RECT  75.320000 199.965000  75.490000 214.935000 ;
      RECT  75.420000  12.795000  75.590000  13.650000 ;
      RECT  75.420000  26.925000  75.590000  27.780000 ;
      RECT  75.450000  44.470000  75.620000  49.570000 ;
      RECT  75.510000 130.030000  76.470000 130.540000 ;
      RECT  75.510000 136.430000  76.470000 136.940000 ;
      RECT  75.530000  56.075000  77.280000  63.645000 ;
      RECT  75.530000  63.645000  78.330000  69.665000 ;
      RECT  75.540000 105.760000  75.710000 107.065000 ;
      RECT  75.615000 160.565000  76.145000 160.895000 ;
      RECT  75.615000 167.825000  76.145000 168.355000 ;
      RECT  75.615000 168.880000  76.145000 169.410000 ;
      RECT  75.730000  99.140000  75.900000 103.890000 ;
      RECT  75.730000 108.340000  75.900000 113.090000 ;
      RECT  75.780000  14.950000  75.950000  18.470000 ;
      RECT  75.780000 227.730000 136.095000 228.050000 ;
      RECT  75.780000 228.050000  76.630000 228.830000 ;
      RECT  75.940000  51.720000  76.110000  54.780000 ;
      RECT  76.100000 199.985000  76.270000 214.985000 ;
      RECT  76.110000  76.400000  76.280000  81.150000 ;
      RECT  76.140000 135.540000  77.100000 136.050000 ;
      RECT  76.140000 141.940000  77.100000 142.450000 ;
      RECT  76.160000  47.555000  76.690000  47.725000 ;
      RECT  76.200000   4.885000  78.510000  12.670000 ;
      RECT  76.200000  12.670000  76.370000  20.495000 ;
      RECT  76.200000  20.495000  78.510000  28.535000 ;
      RECT  76.330000  44.820000  76.500000  47.555000 ;
      RECT  76.330000  47.725000  76.500000  49.570000 ;
      RECT  76.330000 225.650000  77.310000 226.630000 ;
      RECT  76.330000 226.630000 136.095000 227.730000 ;
      RECT  76.330000 234.410000 136.095000 234.980000 ;
      RECT  76.330000 237.100000  77.310000 239.845000 ;
      RECT  76.405000  81.610000  77.215000  81.780000 ;
      RECT  76.565000  81.180000  77.095000  81.610000 ;
      RECT  76.630000  51.810000  77.160000  51.980000 ;
      RECT  76.715000 105.455000  76.885000 105.760000 ;
      RECT  76.715000 105.760000  76.890000 106.425000 ;
      RECT  76.720000 106.425000  76.890000 106.770000 ;
      RECT  76.720000 162.480000  86.720000 165.195000 ;
      RECT  76.720000 172.105000  86.720000 174.820000 ;
      RECT  76.770000 130.030000  77.730000 130.540000 ;
      RECT  76.770000 136.430000  77.730000 136.940000 ;
      RECT  76.800000 228.220000 136.095000 229.255000 ;
      RECT  76.800000 229.255000  77.650000 232.355000 ;
      RECT  76.800000 232.355000 136.095000 233.390000 ;
      RECT  76.815000  85.710000  77.665000  88.500000 ;
      RECT  76.815000  88.500000  77.705000  93.375000 ;
      RECT  76.815000  93.375000  77.665000  95.620000 ;
      RECT  76.815000 116.900000  77.665000 119.145000 ;
      RECT  76.815000 119.145000  77.705000 124.020000 ;
      RECT  76.815000 124.020000  77.665000 126.810000 ;
      RECT  76.820000  51.720000  76.990000  51.810000 ;
      RECT  76.820000  51.980000  76.990000  54.430000 ;
      RECT  76.850000  13.230000  77.180000  14.250000 ;
      RECT  76.850000  19.170000  77.180000  19.935000 ;
      RECT  76.880000 199.965000  77.050000 214.935000 ;
      RECT  77.010000  99.140000  77.180000 104.005000 ;
      RECT  77.010000 108.340000  77.180000 113.205000 ;
      RECT  77.140000 234.980000  77.310000 235.960000 ;
      RECT  77.210000  44.470000  77.380000  49.570000 ;
      RECT  77.215000 146.750000  77.385000 156.600000 ;
      RECT  77.300000 104.940000  87.780000 107.580000 ;
      RECT  77.390000  76.400000  77.560000  81.150000 ;
      RECT  77.400000 135.540000  78.360000 136.050000 ;
      RECT  77.400000 141.940000  78.360000 142.450000 ;
      RECT  77.495000  95.620000  77.665000  95.730000 ;
      RECT  77.495000 116.790000  77.665000 116.900000 ;
      RECT  77.555000 146.360000  81.320000 146.530000 ;
      RECT  77.570000 157.010000  85.720000 157.180000 ;
      RECT  77.660000  12.670000  78.510000  20.495000 ;
      RECT  77.660000 199.985000  79.190000 214.935000 ;
      RECT  77.685000  81.610000  78.495000  81.780000 ;
      RECT  77.700000  51.720000  77.870000  54.780000 ;
      RECT  77.845000  81.180000  78.375000  81.610000 ;
      RECT  77.880000 199.305000  79.190000 199.985000 ;
      RECT  77.880000 214.935000  79.190000 215.605000 ;
      RECT  77.920000  47.555000  78.450000  47.725000 ;
      RECT  78.005000  51.000000  82.755000  51.170000 ;
      RECT  78.030000 130.030000  78.990000 130.540000 ;
      RECT  78.030000 136.430000  78.990000 136.940000 ;
      RECT  78.080000 224.125000  88.080000 226.460000 ;
      RECT  78.080000 229.425000  88.080000 232.185000 ;
      RECT  78.080000 235.150000  88.080000 237.910000 ;
      RECT  78.080000 240.875000  88.080000 242.110000 ;
      RECT  78.090000  44.820000  78.260000  47.555000 ;
      RECT  78.090000  47.725000  78.260000  49.570000 ;
      RECT  78.290000  99.140000  78.460000 103.890000 ;
      RECT  78.290000 108.340000  78.460000 113.090000 ;
      RECT  78.385000  56.465000  78.555000  57.515000 ;
      RECT  78.385000  57.745000  78.555000  58.075000 ;
      RECT  78.385000  58.695000  78.555000  59.025000 ;
      RECT  78.385000  59.195000  78.555000  61.905000 ;
      RECT  78.390000  53.370000  78.920000  53.540000 ;
      RECT  78.410000 130.540000  78.580000 130.600000 ;
      RECT  78.410000 136.940000  78.580000 137.000000 ;
      RECT  78.580000  51.720000  78.750000  53.370000 ;
      RECT  78.580000  53.540000  78.750000  54.430000 ;
      RECT  78.655000  55.965000  79.165000  56.295000 ;
      RECT  78.655000  62.375000  79.165000  62.705000 ;
      RECT  78.660000 135.540000  79.620000 136.050000 ;
      RECT  78.660000 141.940000  79.620000 142.450000 ;
      RECT  78.670000  76.400000  78.840000  81.150000 ;
      RECT  78.725000  56.295000  79.095000  62.375000 ;
      RECT  78.880000 193.605000  79.410000 193.680000 ;
      RECT  78.880000 193.680000  79.415000 193.850000 ;
      RECT  78.880000 193.850000  79.410000 193.965000 ;
      RECT  78.965000  81.610000  79.775000  81.780000 ;
      RECT  78.970000  44.470000  79.140000  49.570000 ;
      RECT  79.005000  84.825000  79.175000  96.855000 ;
      RECT  79.005000 115.675000  79.175000 127.885000 ;
      RECT  79.125000  81.180000  79.655000  81.610000 ;
      RECT  79.265000  56.465000  79.435000  62.210000 ;
      RECT  79.275000  50.080000  83.385000  50.095000 ;
      RECT  79.275000  50.095000  83.465000  50.265000 ;
      RECT  79.275000  50.265000  80.805000  51.000000 ;
      RECT  79.280000   4.635000  86.510000   4.815000 ;
      RECT  79.280000   4.815000  79.460000   7.655000 ;
      RECT  79.280000   7.655000  81.850000   7.825000 ;
      RECT  79.280000   7.825000  80.280000   8.295000 ;
      RECT  79.280000   8.295000  79.460000  14.985000 ;
      RECT  79.280000  14.985000  80.280000  15.145000 ;
      RECT  79.280000  15.145000  81.850000  15.315000 ;
      RECT  79.280000  15.315000  79.460000  18.105000 ;
      RECT  79.280000  18.105000  80.280000  18.435000 ;
      RECT  79.280000  18.435000  79.460000  25.125000 ;
      RECT  79.280000  25.125000  80.280000  25.595000 ;
      RECT  79.280000  25.595000  81.850000  25.765000 ;
      RECT  79.280000  25.765000  79.460000  28.605000 ;
      RECT  79.280000  28.605000  86.510000  28.785000 ;
      RECT  79.290000 130.030000  80.250000 130.540000 ;
      RECT  79.290000 136.430000  80.250000 136.940000 ;
      RECT  79.460000  51.720000  79.630000  54.780000 ;
      RECT  79.520000  37.940000  80.190000  38.240000 ;
      RECT  79.520000  39.200000  80.190000  39.500000 ;
      RECT  79.520000  40.460000  80.190000  40.760000 ;
      RECT  79.520000  41.720000  80.190000  42.020000 ;
      RECT  79.535000  55.965000  80.925000  56.295000 ;
      RECT  79.535000  62.375000  80.925000  62.705000 ;
      RECT  79.570000  99.140000  79.740000 104.005000 ;
      RECT  79.570000 108.340000  79.740000 113.205000 ;
      RECT  79.605000  56.295000  79.975000  62.375000 ;
      RECT  79.605000 186.330000  79.775000 187.000000 ;
      RECT  79.605000 188.070000  79.775000 188.740000 ;
      RECT  79.605000 189.805000  79.775000 190.475000 ;
      RECT  79.605000 191.550000  79.775000 192.220000 ;
      RECT  79.630000  15.520000  80.280000  16.125000 ;
      RECT  79.720000  97.225000  87.790000  97.815000 ;
      RECT  79.720000 114.715000  87.790000 115.305000 ;
      RECT  79.750000  44.820000  79.920000  47.570000 ;
      RECT  79.750000  47.570000  80.280000  47.740000 ;
      RECT  79.750000  47.740000  79.920000  49.570000 ;
      RECT  79.920000 135.540000  80.880000 136.050000 ;
      RECT  79.920000 141.940000  80.880000 142.450000 ;
      RECT  79.950000  76.400000  80.120000  81.150000 ;
      RECT  79.960000 192.985000  80.130000 194.500000 ;
      RECT  80.130000 185.670000 121.065000 186.220000 ;
      RECT  80.130000 186.220000 101.370000 187.450000 ;
      RECT  80.130000 187.620000 101.370000 189.190000 ;
      RECT  80.130000 189.360000 101.370000 190.930000 ;
      RECT  80.130000 191.100000 101.370000 191.955000 ;
      RECT  80.145000  56.465000  80.315000  57.515000 ;
      RECT  80.145000  57.745000  80.315000  58.075000 ;
      RECT  80.145000  58.695000  80.315000  59.025000 ;
      RECT  80.145000  59.195000  80.315000  61.905000 ;
      RECT  80.155000  53.370000  80.685000  53.540000 ;
      RECT  80.190000 197.275000  81.040000 219.215000 ;
      RECT  80.245000  81.610000  81.055000  81.780000 ;
      RECT  80.330000  64.435000  81.895000  64.605000 ;
      RECT  80.330000  64.605000  80.840000  67.865000 ;
      RECT  80.340000  51.720000  80.510000  53.370000 ;
      RECT  80.340000  53.540000  80.510000  54.430000 ;
      RECT  80.405000  81.180000  80.935000  81.610000 ;
      RECT  80.420000  85.730000  80.590000  96.450000 ;
      RECT  80.420000  96.450000  87.790000  97.225000 ;
      RECT  80.420000  97.815000  87.790000  98.390000 ;
      RECT  80.420000 114.130000  87.790000 114.715000 ;
      RECT  80.420000 115.305000  87.790000 116.070000 ;
      RECT  80.420000 116.070000  80.590000 126.790000 ;
      RECT  80.485000  56.295000  80.855000  62.375000 ;
      RECT  80.500000   5.375000  81.850000   5.545000 ;
      RECT  80.500000   8.435000  81.850000   8.605000 ;
      RECT  80.500000   9.215000  81.850000   9.385000 ;
      RECT  80.500000   9.995000  81.850000  10.165000 ;
      RECT  80.500000  10.775000  81.850000  10.945000 ;
      RECT  80.500000  11.555000  81.850000  11.725000 ;
      RECT  80.500000  12.335000  81.850000  12.505000 ;
      RECT  80.500000  13.115000  81.850000  13.285000 ;
      RECT  80.500000  13.895000  81.850000  14.065000 ;
      RECT  80.500000  14.675000  81.850000  14.845000 ;
      RECT  80.500000  15.315000  81.850000  15.625000 ;
      RECT  80.500000  16.235000  81.850000  16.405000 ;
      RECT  80.500000  17.015000  81.850000  17.185000 ;
      RECT  80.500000  17.795000  81.850000  17.965000 ;
      RECT  80.500000  18.575000  81.850000  18.745000 ;
      RECT  80.500000  19.355000  81.850000  19.525000 ;
      RECT  80.500000  20.135000  81.850000  20.305000 ;
      RECT  80.500000  20.855000  81.850000  21.085000 ;
      RECT  80.500000  21.695000  81.850000  21.865000 ;
      RECT  80.500000  22.475000  81.850000  22.645000 ;
      RECT  80.500000  23.255000  81.850000  23.425000 ;
      RECT  80.500000  24.035000  81.850000  24.205000 ;
      RECT  80.500000  24.815000  81.850000  24.985000 ;
      RECT  80.500000  27.875000  81.850000  28.045000 ;
      RECT  80.530000  44.470000  80.700000  49.570000 ;
      RECT  80.540000  36.610000  80.710000  43.350000 ;
      RECT  80.550000 130.030000  81.510000 130.540000 ;
      RECT  80.550000 136.430000  81.510000 136.940000 ;
      RECT  80.850000  99.140000  81.020000 103.890000 ;
      RECT  80.850000 108.340000  81.020000 113.090000 ;
      RECT  81.000000  85.710000  81.170000  95.560000 ;
      RECT  81.000000 116.770000  81.170000 126.620000 ;
      RECT  81.015000  50.440000  89.000000  50.610000 ;
      RECT  81.025000  56.465000  81.195000  62.210000 ;
      RECT  81.130000  47.570000  81.660000  47.740000 ;
      RECT  81.180000 135.540000  82.140000 136.050000 ;
      RECT  81.180000 141.940000  82.140000 142.450000 ;
      RECT  81.220000  51.720000  81.390000  54.780000 ;
      RECT  81.225000  50.610000  88.955000  50.665000 ;
      RECT  81.225000  85.370000  85.225000  85.540000 ;
      RECT  81.225000  95.920000  85.225000  96.090000 ;
      RECT  81.225000 116.430000  85.225000 116.600000 ;
      RECT  81.225000 126.980000  85.225000 127.150000 ;
      RECT  81.230000  76.400000  81.400000  81.150000 ;
      RECT  81.255000 192.845000  81.425000 192.970000 ;
      RECT  81.255000 192.970000  85.155000 193.740000 ;
      RECT  81.255000 193.740000  81.425000 193.855000 ;
      RECT  81.295000  55.965000  81.805000  56.295000 ;
      RECT  81.295000  62.375000  81.805000  62.705000 ;
      RECT  81.310000  44.820000  81.480000  47.570000 ;
      RECT  81.310000  47.740000  81.480000  49.570000 ;
      RECT  81.320000  30.775000  83.340000  31.525000 ;
      RECT  81.320000  41.355000  83.340000  42.105000 ;
      RECT  81.340000  85.540000  85.110000  95.920000 ;
      RECT  81.340000 116.600000  85.110000 126.980000 ;
      RECT  81.365000  56.295000  81.735000  58.310000 ;
      RECT  81.365000  58.310000  82.370000  58.480000 ;
      RECT  81.365000  58.480000  81.735000  62.375000 ;
      RECT  81.495000 146.750000  81.665000 156.600000 ;
      RECT  81.525000  81.610000  82.335000  81.780000 ;
      RECT  81.685000  81.180000  82.215000  81.610000 ;
      RECT  81.810000 130.030000  82.770000 130.540000 ;
      RECT  81.810000 136.430000  82.770000 136.940000 ;
      RECT  81.835000 146.360000  85.605000 146.530000 ;
      RECT  81.900000 192.630000  84.685000 192.800000 ;
      RECT  81.900000 193.910000  84.685000 194.080000 ;
      RECT  81.905000  56.465000  82.075000  57.515000 ;
      RECT  81.905000  57.745000  82.075000  58.075000 ;
      RECT  81.905000  58.695000  82.075000  59.025000 ;
      RECT  81.905000  59.195000  82.075000  61.905000 ;
      RECT  81.910000  53.370000  82.440000  53.540000 ;
      RECT  81.950000  65.155000  82.120000  67.865000 ;
      RECT  81.975000 194.080000  84.685000 194.500000 ;
      RECT  82.040000 198.275000 157.330000 199.125000 ;
      RECT  82.040000 199.125000  85.950000 217.365000 ;
      RECT  82.040000 217.365000 157.330000 218.215000 ;
      RECT  82.090000  44.470000  82.260000  49.570000 ;
      RECT  82.100000  51.720000  82.270000  53.370000 ;
      RECT  82.100000  53.540000  82.270000  54.430000 ;
      RECT  82.130000  99.140000  82.300000 104.005000 ;
      RECT  82.130000 108.340000  82.300000 113.205000 ;
      RECT  82.175000  64.435000  92.135000  64.605000 ;
      RECT  82.260000   5.430000  82.430000  15.680000 ;
      RECT  82.260000  16.265000  82.430000  27.990000 ;
      RECT  82.440000 135.540000  83.400000 136.050000 ;
      RECT  82.440000 141.940000  83.400000 142.450000 ;
      RECT  82.510000  76.400000  82.680000  81.150000 ;
      RECT  82.585000  69.040000  97.970000  70.420000 ;
      RECT  82.690000  47.570000  83.220000  47.740000 ;
      RECT  82.805000  81.610000  83.615000  81.780000 ;
      RECT  82.870000  44.820000  83.040000  47.570000 ;
      RECT  82.870000  47.740000  83.040000  49.570000 ;
      RECT  82.965000  81.180000  83.495000  81.610000 ;
      RECT  82.980000   5.225000  85.690000   5.395000 ;
      RECT  82.980000   7.505000  85.690000   7.675000 ;
      RECT  82.980000   9.785000  85.690000   9.955000 ;
      RECT  82.980000  12.065000  85.690000  12.235000 ;
      RECT  82.980000  14.345000  85.690000  14.515000 ;
      RECT  82.980000  16.625000  85.690000  16.795000 ;
      RECT  82.980000  18.905000  85.690000  19.075000 ;
      RECT  82.980000  21.185000  85.690000  21.355000 ;
      RECT  82.980000  23.465000  85.690000  23.635000 ;
      RECT  82.980000  25.745000  85.690000  25.915000 ;
      RECT  82.980000  28.025000  85.690000  28.195000 ;
      RECT  82.980000  51.720000  83.150000  54.780000 ;
      RECT  83.025000  56.465000  83.195000  57.515000 ;
      RECT  83.025000  57.745000  83.195000  58.075000 ;
      RECT  83.025000  58.695000  83.195000  59.025000 ;
      RECT  83.025000  59.195000  83.195000  61.905000 ;
      RECT  83.070000 130.030000  84.030000 130.540000 ;
      RECT  83.070000 136.430000  84.030000 136.940000 ;
      RECT  83.230000  65.155000  83.400000  67.865000 ;
      RECT  83.295000  55.965000  83.805000  56.295000 ;
      RECT  83.295000  62.375000  83.805000  62.705000 ;
      RECT  83.365000  56.295000  83.735000  62.375000 ;
      RECT  83.410000  99.140000  83.580000 103.890000 ;
      RECT  83.410000 108.340000  83.580000 113.090000 ;
      RECT  83.530000  51.720000  83.700000  53.370000 ;
      RECT  83.530000  53.370000  84.060000  53.540000 ;
      RECT  83.530000  53.540000  83.700000  54.430000 ;
      RECT  83.650000  44.470000  83.820000  49.570000 ;
      RECT  83.700000 135.540000  84.660000 136.050000 ;
      RECT  83.700000 141.940000  84.660000 142.450000 ;
      RECT  83.790000  76.400000  83.960000  81.150000 ;
      RECT  83.810000  35.125000  88.170000  35.295000 ;
      RECT  83.810000  35.295000  83.980000  41.565000 ;
      RECT  83.810000  41.565000  88.170000  41.735000 ;
      RECT  83.810000  51.000000  85.160000  51.410000 ;
      RECT  83.895000  35.040000  88.085000  35.125000 ;
      RECT  83.905000  56.465000  84.075000  62.205000 ;
      RECT  83.995000  50.080000  89.050000  50.265000 ;
      RECT  84.085000  81.610000  84.895000  81.780000 ;
      RECT  84.120000  64.425000  91.375000  64.435000 ;
      RECT  84.175000  55.965000  84.685000  56.295000 ;
      RECT  84.175000  62.375000  84.685000  62.705000 ;
      RECT  84.210000  51.640000  84.740000  51.810000 ;
      RECT  84.225000  82.615000  84.755000  82.785000 ;
      RECT  84.240000  48.370000  84.770000  48.540000 ;
      RECT  84.245000  56.295000  84.615000  58.250000 ;
      RECT  84.245000  58.250000  85.545000  58.495000 ;
      RECT  84.245000  58.495000  84.615000  62.375000 ;
      RECT  84.330000 130.030000  85.290000 130.540000 ;
      RECT  84.330000 136.430000  85.290000 136.940000 ;
      RECT  84.410000  51.810000  84.580000  54.430000 ;
      RECT  84.430000  44.820000  84.600000  48.370000 ;
      RECT  84.430000  48.540000  84.600000  49.570000 ;
      RECT  84.510000  65.155000  84.680000  67.865000 ;
      RECT  84.660000  35.705000  87.370000  35.875000 ;
      RECT  84.660000  36.585000  87.370000  36.755000 ;
      RECT  84.660000  37.465000  87.370000  37.635000 ;
      RECT  84.660000  38.345000  87.370000  38.515000 ;
      RECT  84.660000  39.225000  87.370000  39.395000 ;
      RECT  84.660000  40.105000  87.370000  40.275000 ;
      RECT  84.660000  40.985000  87.370000  41.155000 ;
      RECT  84.690000  99.140000  84.860000 104.005000 ;
      RECT  84.690000 108.340000  84.860000 113.205000 ;
      RECT  84.785000  56.465000  84.955000  57.515000 ;
      RECT  84.785000  57.745000  84.955000  58.075000 ;
      RECT  84.785000  58.695000  84.955000  59.025000 ;
      RECT  84.785000  59.195000  84.955000  61.905000 ;
      RECT  84.825000 192.925000  85.155000 192.970000 ;
      RECT  84.825000 193.740000  85.155000 193.775000 ;
      RECT  84.915000 104.360000  85.640000 104.530000 ;
      RECT  84.915000 113.550000  85.640000 113.720000 ;
      RECT  84.960000 135.540000  85.920000 136.050000 ;
      RECT  84.960000 141.940000  85.920000 142.450000 ;
      RECT  85.070000  76.400000  85.240000  81.150000 ;
      RECT  85.100000  53.370000  85.630000  53.540000 ;
      RECT  85.210000  44.470000  85.380000  49.570000 ;
      RECT  85.280000  85.710000  85.450000  95.560000 ;
      RECT  85.280000 116.770000  85.450000 126.620000 ;
      RECT  85.290000  51.720000  85.460000  53.370000 ;
      RECT  85.290000  53.540000  85.460000  54.430000 ;
      RECT  85.375000  56.465000  85.545000  58.250000 ;
      RECT  85.375000  58.495000  85.545000  62.210000 ;
      RECT  85.470000  99.140000  85.640000 104.360000 ;
      RECT  85.470000 108.340000  85.640000 113.550000 ;
      RECT  85.545000  50.865000  86.895000  51.170000 ;
      RECT  85.590000 130.030000  86.550000 130.540000 ;
      RECT  85.590000 136.430000  86.550000 136.940000 ;
      RECT  85.645000  55.965000  93.190000  56.295000 ;
      RECT  85.645000  62.375000  86.155000  62.705000 ;
      RECT  85.650000  76.050000  85.820000  82.020000 ;
      RECT  85.705000  95.920000  86.235000  96.090000 ;
      RECT  85.715000  56.295000  86.085000  62.375000 ;
      RECT  85.720000 116.325000  86.250000 116.495000 ;
      RECT  85.775000 146.750000  85.945000 156.600000 ;
      RECT  85.790000  65.155000  85.960000  67.865000 ;
      RECT  85.800000  48.355000  86.330000  48.525000 ;
      RECT  85.890000  86.305000  86.060000  87.305000 ;
      RECT  85.910000   5.370000  86.090000  28.050000 ;
      RECT  85.990000  44.820000  86.160000  48.355000 ;
      RECT  85.990000  48.525000  86.160000  49.570000 ;
      RECT  85.995000  53.000000  86.525000  53.170000 ;
      RECT  86.020000  87.850000  86.190000  87.910000 ;
      RECT  86.020000  87.910000  87.790000  88.080000 ;
      RECT  86.020000  88.080000  86.190000  88.520000 ;
      RECT  86.020000  88.690000  87.150000  88.860000 ;
      RECT  86.020000  88.860000  86.190000  94.870000 ;
      RECT  86.020000  95.430000  86.190000  95.920000 ;
      RECT  86.020000  96.090000  86.190000  96.100000 ;
      RECT  86.020000  99.140000  86.190000 103.890000 ;
      RECT  86.020000 108.340000  86.190000 113.205000 ;
      RECT  86.020000 116.495000  86.190000 117.090000 ;
      RECT  86.020000 117.650000  86.190000 123.660000 ;
      RECT  86.020000 123.660000  87.150000 123.830000 ;
      RECT  86.020000 124.000000  86.190000 124.440000 ;
      RECT  86.020000 124.440000  87.790000 124.610000 ;
      RECT  86.020000 124.610000  86.190000 124.670000 ;
      RECT  86.115000 191.955000 101.370000 194.500000 ;
      RECT  86.170000  51.720000  86.340000  53.000000 ;
      RECT  86.170000  53.170000  86.340000  54.430000 ;
      RECT  86.220000 135.540000  87.180000 136.050000 ;
      RECT  86.220000 141.940000  87.180000 142.450000 ;
      RECT  86.255000  56.465000  86.425000  57.515000 ;
      RECT  86.255000  57.745000  86.425000  58.075000 ;
      RECT  86.255000  58.695000  86.425000  59.025000 ;
      RECT  86.255000  59.195000  86.425000  61.905000 ;
      RECT  86.260000  86.080000  87.280000  86.250000 ;
      RECT  86.260000  87.360000  87.790000  87.530000 ;
      RECT  86.325000 160.565000  86.855000 160.895000 ;
      RECT  86.330000   4.815000  86.510000  28.605000 ;
      RECT  86.355000 145.325000  86.525000 158.215000 ;
      RECT  86.370000  91.250000  87.260000  91.420000 ;
      RECT  86.370000  93.810000  87.260000  93.980000 ;
      RECT  86.370000 118.540000  87.260000 118.710000 ;
      RECT  86.370000 121.100000  87.260000 121.270000 ;
      RECT  86.380000 104.350000  87.390000 104.520000 ;
      RECT  86.380000 113.550000  87.455000 113.720000 ;
      RECT  86.430000  75.120000  87.720000  82.955000 ;
      RECT  86.460000 200.495000  86.990000 215.995000 ;
      RECT  86.480000  89.970000  87.790000  90.140000 ;
      RECT  86.480000  92.530000  87.370000  92.700000 ;
      RECT  86.480000  95.090000  87.425000  95.260000 ;
      RECT  86.480000  95.870000  87.150000  96.040000 ;
      RECT  86.480000 116.480000  87.150000 116.650000 ;
      RECT  86.480000 117.260000  87.300000 117.430000 ;
      RECT  86.480000 119.820000  87.370000 119.990000 ;
      RECT  86.480000 122.380000  87.790000 122.550000 ;
      RECT  86.495000  96.040000  87.025000  96.090000 ;
      RECT  86.690000  53.370000  87.220000  53.540000 ;
      RECT  86.770000  44.470000  86.940000  49.570000 ;
      RECT  86.800000  99.140000  86.970000 103.890000 ;
      RECT  86.800000 108.340000  86.970000 113.090000 ;
      RECT  86.850000 130.030000  87.180000 130.540000 ;
      RECT  86.850000 136.430000  87.180000 136.940000 ;
      RECT  86.930000 130.540000  87.100000 130.600000 ;
      RECT  86.930000 136.940000  87.100000 137.000000 ;
      RECT  87.050000  51.720000  87.220000  53.370000 ;
      RECT  87.050000  53.540000  87.220000  54.430000 ;
      RECT  87.070000  65.155000  87.240000  67.865000 ;
      RECT  87.130000 117.430000  87.300000 117.790000 ;
      RECT  87.175000  39.610000  87.760000  39.780000 ;
      RECT  87.185000 166.450000  87.355000 170.850000 ;
      RECT  87.225000  36.955000  87.760000  37.125000 ;
      RECT  87.255000  94.730000  87.425000  95.090000 ;
      RECT  87.275000   4.635000  90.020000   4.815000 ;
      RECT  87.275000   4.815000  87.455000  34.060000 ;
      RECT  87.275000  34.060000  90.020000  34.240000 ;
      RECT  87.290000 143.905000  90.225000 159.150000 ;
      RECT  87.380000  48.355000  87.910000  48.525000 ;
      RECT  87.420000 200.085000  88.355000 200.255000 ;
      RECT  87.550000  44.820000  87.720000  48.355000 ;
      RECT  87.550000  48.525000  87.720000  49.570000 ;
      RECT  87.580000  99.140000  87.750000 103.890000 ;
      RECT  87.580000 108.340000  87.750000 113.205000 ;
      RECT  87.590000  35.930000  87.760000  36.955000 ;
      RECT  87.590000  37.125000  87.760000  37.410000 ;
      RECT  87.590000  37.690000  87.760000  39.610000 ;
      RECT  87.590000  39.780000  87.760000  40.930000 ;
      RECT  87.595000 162.310000  88.445000 174.990000 ;
      RECT  87.600000  51.720000  87.770000  54.780000 ;
      RECT  87.620000  86.040000  87.790000  87.360000 ;
      RECT  87.620000  87.530000  87.790000  87.910000 ;
      RECT  87.620000  88.080000  87.790000  89.970000 ;
      RECT  87.620000  90.140000  87.790000  96.450000 ;
      RECT  87.620000 116.070000  87.790000 122.380000 ;
      RECT  87.620000 122.550000  87.790000 124.440000 ;
      RECT  87.620000 124.610000  87.790000 126.480000 ;
      RECT  87.620000 129.620000  87.790000 142.385000 ;
      RECT  87.750000  14.275000  87.920000  15.375000 ;
      RECT  87.750000  15.655000  87.920000  16.755000 ;
      RECT  87.750000  17.820000  89.160000  17.990000 ;
      RECT  87.750000  17.990000  87.920000  18.775000 ;
      RECT  87.930000  50.960000  90.980000  51.130000 ;
      RECT  88.000000  35.295000  88.170000  39.185000 ;
      RECT  88.000000  39.185000  88.560000  39.355000 ;
      RECT  88.000000  39.355000  88.170000  41.565000 ;
      RECT  88.085000   7.585000  89.160000   7.755000 ;
      RECT  88.150000   5.225000  89.160000   5.395000 ;
      RECT  88.150000   6.405000  89.160000   6.575000 ;
      RECT  88.150000   8.765000  89.160000   8.935000 ;
      RECT  88.150000   9.945000  89.160000  10.115000 ;
      RECT  88.150000  10.615000  89.160000  10.785000 ;
      RECT  88.150000  11.045000  89.160000  11.215000 ;
      RECT  88.150000  11.475000  89.160000  11.645000 ;
      RECT  88.150000  11.905000  89.160000  12.105000 ;
      RECT  88.150000  12.335000  89.160000  12.505000 ;
      RECT  88.150000  13.590000  89.160000  13.760000 ;
      RECT  88.150000  14.050000  89.160000  14.220000 ;
      RECT  88.150000  14.510000  89.160000  14.680000 ;
      RECT  88.150000  14.970000  89.160000  15.140000 ;
      RECT  88.150000  15.430000  89.160000  15.600000 ;
      RECT  88.150000  15.890000  89.160000  16.060000 ;
      RECT  88.150000  16.350000  89.160000  16.520000 ;
      RECT  88.150000  16.810000  89.160000  16.980000 ;
      RECT  88.150000  17.360000  89.160000  17.530000 ;
      RECT  88.150000  18.370000  89.160000  18.540000 ;
      RECT  88.150000  18.830000  89.160000  19.000000 ;
      RECT  88.150000  19.290000  89.160000  19.460000 ;
      RECT  88.150000  20.070000  89.160000  20.240000 ;
      RECT  88.150000  20.470000  89.040000  20.500000 ;
      RECT  88.150000  20.500000  89.160000  20.670000 ;
      RECT  88.150000  20.930000  89.160000  21.100000 ;
      RECT  88.150000  21.360000  89.160000  21.530000 ;
      RECT  88.150000  21.790000  89.160000  21.960000 ;
      RECT  88.150000  22.460000  89.160000  22.630000 ;
      RECT  88.150000  23.640000  89.160000  23.810000 ;
      RECT  88.150000  24.820000  89.160000  24.990000 ;
      RECT  88.150000  26.000000  89.160000  26.170000 ;
      RECT  88.150000  27.180000  89.160000  27.350000 ;
      RECT  88.150000  27.730000  88.820000  27.900000 ;
      RECT  88.150000  29.010000  88.820000  29.180000 ;
      RECT  88.150000  30.100000  88.820000  30.405000 ;
      RECT  88.150000  30.405000  89.590000  30.575000 ;
      RECT  88.150000  30.840000  89.160000  31.010000 ;
      RECT  88.150000  31.720000  89.160000  31.890000 ;
      RECT  88.150000  32.600000  89.160000  32.770000 ;
      RECT  88.150000  33.480000  89.160000  33.650000 ;
      RECT  88.190000  71.685000  90.210000  72.435000 ;
      RECT  88.190000  82.265000  90.210000  83.015000 ;
      RECT  88.250000 234.980000  89.855000 235.745000 ;
      RECT  88.330000  44.470000  88.500000  49.570000 ;
      RECT  88.350000  65.155000  88.520000  67.865000 ;
      RECT  88.480000  51.720000  88.650000  53.000000 ;
      RECT  88.480000  53.000000  89.010000  53.170000 ;
      RECT  88.480000  53.170000  88.650000  54.430000 ;
      RECT  88.520000 200.495000  89.050000 215.995000 ;
      RECT  88.745000 229.255000  89.595000 232.355000 ;
      RECT  88.745000 239.670000 136.095000 240.705000 ;
      RECT  88.745000 240.705000  89.595000 242.540000 ;
      RECT  88.875000 235.745000  89.855000 238.080000 ;
      RECT  88.875000 238.080000 136.095000 239.500000 ;
      RECT  88.880000  44.820000  89.050000  48.845000 ;
      RECT  88.880000  48.845000  89.410000  49.015000 ;
      RECT  88.880000  49.015000  89.050000  50.080000 ;
      RECT  88.930000  35.040000  95.400000  35.395000 ;
      RECT  88.930000  35.395000  89.100000  41.465000 ;
      RECT  88.930000  41.465000  99.560000  41.635000 ;
      RECT  88.985000 223.695000  89.595000 225.350000 ;
      RECT  89.035000  84.825000  89.205000 108.735000 ;
      RECT  89.035000 108.735000 190.325000 109.585000 ;
      RECT  89.035000 109.585000  90.225000 127.885000 ;
      RECT  89.035000 128.205000  90.225000 143.735000 ;
      RECT  89.050000  28.885000  89.220000  29.235000 ;
      RECT  89.050000  29.235000  89.405000  30.235000 ;
      RECT  89.060000  63.475000  93.915000  63.645000 ;
      RECT  89.085000 225.650000  89.255000 226.630000 ;
      RECT  89.100000  57.440000  89.270000  62.290000 ;
      RECT  89.250000  56.635000  89.920000  56.805000 ;
      RECT  89.340000  35.930000  89.510000  37.520000 ;
      RECT  89.340000  37.690000  89.510000  40.575000 ;
      RECT  89.340000  40.575000  89.910000  40.745000 ;
      RECT  89.340000  40.745000  89.510000  40.930000 ;
      RECT  89.355000  50.000000  89.525000  50.670000 ;
      RECT  89.360000  51.720000  89.530000  54.780000 ;
      RECT  89.375000 160.000000  90.225000 168.145000 ;
      RECT  89.375000 168.145000 190.325000 173.235000 ;
      RECT  89.375000 173.235000 162.890000 176.145000 ;
      RECT  89.375000 176.145000  90.225000 176.600000 ;
      RECT  89.390000  27.955000  89.590000  28.955000 ;
      RECT  89.420000   5.450000  89.590000   9.890000 ;
      RECT  89.420000  10.840000  89.590000  12.280000 ;
      RECT  89.420000  13.325000  89.590000  15.785000 ;
      RECT  89.420000  16.420000  89.590000  18.255000 ;
      RECT  89.420000  19.005000  89.960000  19.535000 ;
      RECT  89.420000  19.535000  89.590000  19.725000 ;
      RECT  89.420000  20.295000  89.590000  21.735000 ;
      RECT  89.420000  22.570000  89.590000  27.125000 ;
      RECT  89.420000  30.575000  89.590000  31.665000 ;
      RECT  89.420000  31.840000  89.590000  33.425000 ;
      RECT  89.480000 200.085000  90.150000 200.255000 ;
      RECT  89.630000  65.155000  89.800000  67.865000 ;
      RECT  89.660000  44.470000  89.830000  49.570000 ;
      RECT  89.840000   4.815000  90.020000  18.835000 ;
      RECT  89.840000  19.705000  90.020000  34.060000 ;
      RECT  89.880000  53.000000  90.410000  53.170000 ;
      RECT  89.880000  57.440000  90.050000  62.290000 ;
      RECT  90.025000 224.125000 100.025000 226.460000 ;
      RECT  90.025000 229.425000 100.025000 232.185000 ;
      RECT  90.025000 235.150000 100.025000 237.910000 ;
      RECT  90.025000 240.875000 100.025000 243.210000 ;
      RECT  90.050000  49.740000  92.290000  49.910000 ;
      RECT  90.050000  49.910000  90.220000  50.670000 ;
      RECT  90.060000  35.705000  92.770000  35.875000 ;
      RECT  90.060000  36.585000  92.770000  36.755000 ;
      RECT  90.060000  37.465000  92.770000  37.635000 ;
      RECT  90.060000  38.345000  92.770000  38.515000 ;
      RECT  90.060000  39.225000  92.770000  39.395000 ;
      RECT  90.060000  40.105000  92.770000  40.275000 ;
      RECT  90.060000  40.985000  92.770000  41.155000 ;
      RECT  90.240000  51.720000  90.410000  53.000000 ;
      RECT  90.240000  53.170000  90.410000  54.430000 ;
      RECT  90.250000  48.845000  90.780000  49.015000 ;
      RECT  90.375000   7.175000  90.965000   7.345000 ;
      RECT  90.435000  92.010000  98.825000  93.070000 ;
      RECT  90.435000  93.070000 299.570000  93.980000 ;
      RECT  90.440000  44.820000  90.610000  48.845000 ;
      RECT  90.440000  49.015000  90.610000  49.570000 ;
      RECT  90.450000  85.300000  98.820000  88.625000 ;
      RECT  90.450000  88.625000  98.825000  92.010000 ;
      RECT  90.450000  93.980000 299.555000  95.265000 ;
      RECT  90.450000  95.265000 153.450000 102.115000 ;
      RECT  90.450000 102.115000 116.880000 107.805000 ;
      RECT  90.470000  57.440000  90.640000  62.290000 ;
      RECT  90.580000 200.495000  91.110000 215.995000 ;
      RECT  90.780000  50.080000  90.950000  50.960000 ;
      RECT  90.785000   4.635000  93.605000   4.815000 ;
      RECT  90.785000   4.815000  90.965000   7.175000 ;
      RECT  90.785000   7.345000  90.965000  12.515000 ;
      RECT  90.785000  12.515000  93.605000  12.695000 ;
      RECT  90.785000  13.460000  93.605000  13.520000 ;
      RECT  90.785000  13.520000  93.685000  13.640000 ;
      RECT  90.785000  13.640000  90.965000  19.485000 ;
      RECT  90.785000  19.485000  93.605000  19.770000 ;
      RECT  90.785000  20.535000  93.605000  20.715000 ;
      RECT  90.785000  20.715000  90.965000  24.345000 ;
      RECT  90.785000  24.345000  93.605000  24.525000 ;
      RECT  90.785000  25.500000  93.605000  25.680000 ;
      RECT  90.785000  25.680000  90.965000  34.060000 ;
      RECT  90.785000  34.060000  93.605000  34.240000 ;
      RECT  90.860000  56.635000  92.810000  56.805000 ;
      RECT  90.910000  65.155000  91.080000  67.865000 ;
      RECT  91.120000  51.720000  91.290000  54.780000 ;
      RECT  91.155000 176.905000 160.800000 178.210000 ;
      RECT  91.215000  14.140000  92.645000  14.310000 ;
      RECT  91.215000  14.310000  91.385000  15.725000 ;
      RECT  91.215000  16.420000  91.385000  18.435000 ;
      RECT  91.215000  26.870000  91.385000  27.595000 ;
      RECT  91.215000  30.185000  91.385000  33.425000 ;
      RECT  91.220000  44.470000  91.390000  49.570000 ;
      RECT  91.300000  50.405000  91.830000  50.575000 ;
      RECT  91.540000 200.085000  92.210000 200.255000 ;
      RECT  91.630000  50.080000  91.800000  50.405000 ;
      RECT  91.630000  50.575000  91.800000  50.750000 ;
      RECT  91.635000  14.050000  92.645000  14.140000 ;
      RECT  91.635000  14.830000  92.645000  15.000000 ;
      RECT  91.635000  15.520000  93.035000  15.690000 ;
      RECT  91.635000  15.690000  92.645000  15.780000 ;
      RECT  91.635000  16.160000  92.645000  16.330000 ;
      RECT  91.635000  16.620000  92.645000  16.790000 ;
      RECT  91.635000  17.080000  92.645000  17.250000 ;
      RECT  91.635000  17.540000  92.645000  17.710000 ;
      RECT  91.635000  18.000000  93.105000  18.170000 ;
      RECT  91.635000  18.550000  92.645000  18.720000 ;
      RECT  91.635000  19.010000  92.645000  19.180000 ;
      RECT  91.695000   5.225000  92.705000   5.395000 ;
      RECT  91.695000   6.105000  92.705000   6.275000 ;
      RECT  91.695000   6.985000  92.705000   7.155000 ;
      RECT  91.695000   7.865000  92.705000   8.035000 ;
      RECT  91.695000   8.745000  92.705000   8.915000 ;
      RECT  91.695000   9.295000  92.705000   9.465000 ;
      RECT  91.695000  10.175000  92.705000  10.345000 ;
      RECT  91.695000  11.055000  92.705000  11.225000 ;
      RECT  91.695000  11.935000  92.705000  12.105000 ;
      RECT  91.695000  21.125000  92.705000  21.295000 ;
      RECT  91.695000  22.005000  92.705000  22.175000 ;
      RECT  91.695000  22.885000  92.705000  23.055000 ;
      RECT  91.695000  23.765000  92.705000  23.935000 ;
      RECT  91.695000  28.200000  92.705000  28.370000 ;
      RECT  91.695000  29.080000  92.705000  29.250000 ;
      RECT  91.695000  29.960000  92.705000  30.130000 ;
      RECT  91.695000  30.840000  92.705000  31.010000 ;
      RECT  91.695000  31.720000  92.705000  31.890000 ;
      RECT  91.695000  32.600000  92.705000  32.770000 ;
      RECT  91.695000  33.480000  92.705000  33.650000 ;
      RECT  91.750000  57.440000  91.920000  62.290000 ;
      RECT  91.760000  51.240000  92.290000  51.410000 ;
      RECT  91.795000 110.585000 187.905000 111.435000 ;
      RECT  91.795000 111.435000  92.645000 166.535000 ;
      RECT  91.795000 166.535000 187.905000 167.385000 ;
      RECT  91.915000  26.090000  92.585000  26.260000 ;
      RECT  91.915000  26.870000  92.585000  27.040000 ;
      RECT  91.915000  27.650000  92.585000  27.820000 ;
      RECT  92.000000  44.820000  92.290000  49.740000 ;
      RECT  92.000000  49.910000  92.290000  51.240000 ;
      RECT  92.000000  51.410000  92.290000  54.430000 ;
      RECT  92.190000  65.155000  92.360000  67.865000 ;
      RECT  92.415000  64.435000  93.980000  64.605000 ;
      RECT  92.550000  44.820000  92.820000  49.665000 ;
      RECT  92.550000  49.665000  93.080000  49.835000 ;
      RECT  92.550000  49.835000  92.820000  54.430000 ;
      RECT  92.625000  36.955000  93.160000  37.125000 ;
      RECT  92.625000  40.575000  93.160000  40.745000 ;
      RECT  92.640000 200.495000  93.170000 215.995000 ;
      RECT  92.865000  14.105000  93.035000  15.520000 ;
      RECT  92.865000  71.040000  97.970000  74.525000 ;
      RECT  92.865000  74.525000  99.865000  75.535000 ;
      RECT  92.865000  75.535000  98.820000  85.300000 ;
      RECT  92.925000  21.015000  94.780000  21.285000 ;
      RECT  92.925000  21.285000  93.095000  23.710000 ;
      RECT  92.935000   5.450000  93.105000   8.690000 ;
      RECT  92.935000   9.520000  93.105000  11.985000 ;
      RECT  92.935000  18.170000  93.105000  18.955000 ;
      RECT  92.990000  35.930000  93.160000  36.955000 ;
      RECT  92.990000  37.125000  93.160000  37.410000 ;
      RECT  92.990000  37.690000  93.160000  40.575000 ;
      RECT  92.990000  40.745000  93.160000  40.930000 ;
      RECT  92.990000  50.035000  93.520000  50.205000 ;
      RECT  93.005000  16.385000  93.175000  17.300000 ;
      RECT  93.005000  17.300000  93.605000  17.485000 ;
      RECT  93.005000  26.145000  93.175000  26.815000 ;
      RECT  93.005000  27.970000  93.175000  29.905000 ;
      RECT  93.020000  55.765000  93.190000  55.965000 ;
      RECT  93.030000  57.440000  93.200000  62.290000 ;
      RECT  93.050000  50.015000  93.220000  50.035000 ;
      RECT  93.050000  50.205000  93.220000  50.840000 ;
      RECT  93.050000  50.840000  94.480000  51.140000 ;
      RECT  93.250000 113.910000  96.250000 164.900000 ;
      RECT  93.425000   4.815000  93.605000  12.515000 ;
      RECT  93.425000  13.640000  93.685000  14.585000 ;
      RECT  93.425000  14.585000  93.605000  16.000000 ;
      RECT  93.425000  16.000000  93.685000  16.900000 ;
      RECT  93.425000  16.900000  93.605000  17.085000 ;
      RECT  93.425000  18.055000  93.605000  19.485000 ;
      RECT  93.425000  20.715000  93.605000  20.845000 ;
      RECT  93.425000  21.455000  93.605000  24.345000 ;
      RECT  93.425000  25.680000  93.605000  34.060000 ;
      RECT  93.430000  44.470000  93.600000  49.570000 ;
      RECT  93.430000  51.720000  93.600000  54.780000 ;
      RECT  93.435000  17.485000  93.605000  17.830000 ;
      RECT  93.470000  64.605000  93.980000  67.865000 ;
      RECT  93.600000 200.085000  94.270000 200.255000 ;
      RECT  93.710000  35.705000  96.420000  35.875000 ;
      RECT  93.710000  36.585000  96.420000  36.755000 ;
      RECT  93.710000  37.465000  96.420000  37.635000 ;
      RECT  93.710000  38.345000  96.420000  38.515000 ;
      RECT  93.710000  39.225000  96.420000  39.395000 ;
      RECT  93.710000  40.105000  96.420000  40.275000 ;
      RECT  93.710000  40.985000  96.420000  41.155000 ;
      RECT  93.745000  56.625000  93.915000  63.475000 ;
      RECT  93.750000  50.000000  94.040000  50.670000 ;
      RECT  93.770000  45.575000  94.040000  50.000000 ;
      RECT  94.210000  44.820000  94.480000  50.840000 ;
      RECT  94.210000  51.140000  94.480000  54.430000 ;
      RECT  94.610000  21.285000  94.780000  21.605000 ;
      RECT  94.700000 200.495000  95.230000 215.995000 ;
      RECT  94.790000  44.470000  94.960000  49.840000 ;
      RECT  94.890000  50.600000 113.595000  51.555000 ;
      RECT  94.890000  51.555000 113.590000  53.600000 ;
      RECT  94.890000  53.600000 110.720000  54.780000 ;
      RECT  95.230000  34.640000  99.560000  34.845000 ;
      RECT  95.230000  34.845000  95.400000  35.040000 ;
      RECT  95.380000  58.725000 110.720000  59.255000 ;
      RECT  95.415000  56.185000 110.720000  56.715000 ;
      RECT  95.490000  55.295000 110.720000  56.185000 ;
      RECT  95.490000  56.715000 110.720000  58.725000 ;
      RECT  95.490000  59.255000 110.720000  60.605000 ;
      RECT  95.490000  60.605000  99.865000  62.780000 ;
      RECT  95.505000  62.780000  99.865000  63.070000 ;
      RECT  95.660000 200.085000  96.330000 200.255000 ;
      RECT  95.705000 113.195000  96.375000 113.525000 ;
      RECT  95.720000  46.500000  99.970000  46.990000 ;
      RECT  95.760000  46.990000  99.890000  47.125000 ;
      RECT  95.775000 113.165000  96.305000 113.195000 ;
      RECT  96.120000  28.410000  99.460000  28.765000 ;
      RECT  96.120000  28.765000  96.290000  31.995000 ;
      RECT  96.120000  31.995000  99.460000  32.165000 ;
      RECT  96.485000 179.155000 158.850000 180.175000 ;
      RECT  96.485000 180.175000 122.340000 180.515000 ;
      RECT  96.485000 180.515000 121.065000 183.710000 ;
      RECT  96.530000  29.040000  96.720000  31.380000 ;
      RECT  96.570000  49.975000 113.910000  50.405000 ;
      RECT  96.570000  50.405000 113.595000  50.600000 ;
      RECT  96.715000  38.730000  97.250000  38.900000 ;
      RECT  96.715000  40.575000  97.250000  40.745000 ;
      RECT  96.760000 200.495000  97.290000 215.995000 ;
      RECT  96.830000  63.070000  97.970000  69.040000 ;
      RECT  96.950000  29.095000  97.640000  29.955000 ;
      RECT  96.950000  31.435000  97.640000  31.665000 ;
      RECT  97.080000  38.090000  97.250000  38.730000 ;
      RECT  97.080000  38.900000  97.250000  39.370000 ;
      RECT  97.080000  39.650000  97.250000  40.575000 ;
      RECT  97.080000  40.745000  97.250000  40.930000 ;
      RECT  97.240000   2.815000  99.760000   2.985000 ;
      RECT  97.240000   2.985000  97.670000   7.485000 ;
      RECT  97.240000   8.025000  97.670000  10.585000 ;
      RECT  97.240000  10.585000 100.195000  10.895000 ;
      RECT  97.355000  35.380000  97.525000  36.370000 ;
      RECT  97.420000  37.865000  99.110000  38.035000 ;
      RECT  97.420000  38.035000  97.590000  39.425000 ;
      RECT  97.420000  39.425000  99.110000  39.595000 ;
      RECT  97.420000  39.595000  97.590000  40.985000 ;
      RECT  97.420000  40.985000  99.110000  41.155000 ;
      RECT  97.500000   7.485000  97.670000   8.025000 ;
      RECT  97.500000  13.265000  99.760000  13.435000 ;
      RECT  97.500000  13.435000  97.670000  25.915000 ;
      RECT  97.500000  25.915000  99.760000  26.085000 ;
      RECT  97.680000  36.460000  97.930000  37.260000 ;
      RECT  97.720000 200.085000  98.390000 200.255000 ;
      RECT  97.760000  35.155000  99.110000  35.325000 ;
      RECT  97.760000  35.325000  97.930000  36.460000 ;
      RECT  97.760000  38.645000  99.110000  38.815000 ;
      RECT  97.760000  40.205000  99.110000  40.375000 ;
      RECT  97.760000 113.910000 100.760000 164.900000 ;
      RECT  97.855000  15.025000  98.930000  15.195000 ;
      RECT  97.920000   3.295000  98.930000   3.465000 ;
      RECT  97.920000   3.755000  98.930000   3.925000 ;
      RECT  97.920000   4.215000  98.930000   4.385000 ;
      RECT  97.920000   4.675000  98.930000   4.845000 ;
      RECT  97.920000   5.135000  98.930000   5.305000 ;
      RECT  97.920000   5.595000  98.930000   5.765000 ;
      RECT  97.920000   6.055000  98.930000   6.225000 ;
      RECT  97.920000   6.515000  98.930000   6.685000 ;
      RECT  97.920000   6.975000  98.930000   7.145000 ;
      RECT  97.920000   7.345000  98.880000   7.435000 ;
      RECT  97.920000   7.435000  98.930000   7.605000 ;
      RECT  97.920000   7.985000  98.930000   8.180000 ;
      RECT  97.920000   8.485000  98.930000   8.685000 ;
      RECT  97.920000   9.045000  98.930000   9.215000 ;
      RECT  97.920000   9.575000  98.930000   9.745000 ;
      RECT  97.920000  10.105000  98.930000  10.275000 ;
      RECT  97.920000  13.665000  98.950000  13.915000 ;
      RECT  97.920000  16.305000  98.950000  16.475000 ;
      RECT  97.920000  16.855000  99.350000  17.025000 ;
      RECT  97.920000  18.135000  98.930000  18.305000 ;
      RECT  97.920000  19.415000  98.930000  19.585000 ;
      RECT  97.920000  19.965000  99.350000  20.135000 ;
      RECT  97.920000  21.245000  98.930000  21.415000 ;
      RECT  97.920000  22.525000  98.930000  22.695000 ;
      RECT  97.920000  23.075000  98.930000  23.245000 ;
      RECT  97.920000  24.355000  98.930000  24.525000 ;
      RECT  97.920000  25.435000  98.930000  25.605000 ;
      RECT  97.970000  29.095000  98.660000  29.405000 ;
      RECT  97.970000  31.435000  98.660000  31.665000 ;
      RECT  98.100000  36.235000  99.110000  36.405000 ;
      RECT  98.100000  37.315000  99.110000  37.485000 ;
      RECT  98.465000  29.755000  99.050000  29.925000 ;
      RECT  98.590000  23.970000  99.350000  24.140000 ;
      RECT  98.610000  14.445000  99.350000  14.615000 ;
      RECT  98.820000  25.065000  99.350000  25.235000 ;
      RECT  98.820000 200.495000  99.350000 215.995000 ;
      RECT  98.880000  29.380000  99.050000  29.755000 ;
      RECT  98.880000  29.925000  99.050000  31.380000 ;
      RECT  99.050000  76.025000 101.480000  76.195000 ;
      RECT  99.050000  76.195000  99.220000  87.700000 ;
      RECT  99.050000  87.700000 175.800000  87.870000 ;
      RECT  99.050000  87.870000 100.935000  87.885000 ;
      RECT  99.100000   9.225000 101.250000   9.450000 ;
      RECT  99.180000   3.520000  99.350000   6.000000 ;
      RECT  99.180000   6.280000  99.350000   6.915000 ;
      RECT  99.180000   6.915000 101.250000   7.085000 ;
      RECT  99.180000   7.085000  99.350000   7.380000 ;
      RECT  99.180000   7.910000 101.250000   8.080000 ;
      RECT  99.180000   8.080000  99.350000   8.990000 ;
      RECT  99.180000   9.745000  99.350000  10.245000 ;
      RECT  99.180000  10.245000  99.715000  10.415000 ;
      RECT  99.180000  13.970000  99.350000  14.445000 ;
      RECT  99.180000  14.615000  99.350000  14.970000 ;
      RECT  99.180000  15.250000  99.350000  16.855000 ;
      RECT  99.180000  17.195000  99.350000  18.080000 ;
      RECT  99.180000  18.360000  99.350000  19.965000 ;
      RECT  99.180000  20.305000  99.350000  21.190000 ;
      RECT  99.180000  21.470000  99.350000  23.460000 ;
      RECT  99.180000  23.630000  99.350000  23.970000 ;
      RECT  99.180000  24.140000  99.350000  24.300000 ;
      RECT  99.180000  24.580000  99.350000  25.065000 ;
      RECT  99.180000  25.235000  99.350000  25.380000 ;
      RECT  99.205000  31.785000  99.460000  31.995000 ;
      RECT  99.290000  28.765000  99.460000  31.785000 ;
      RECT  99.390000  34.845000  99.560000  41.465000 ;
      RECT  99.425000  87.885000 100.225000  91.465000 ;
      RECT  99.425000  91.465000 145.515000  91.720000 ;
      RECT  99.425000  91.720000 125.530000  92.265000 ;
      RECT  99.575000   8.885000  99.760000   8.995000 ;
      RECT  99.575000   8.995000  99.745000   9.055000 ;
      RECT  99.590000   2.985000  99.760000   6.745000 ;
      RECT  99.590000   7.255000  99.760000   7.740000 ;
      RECT  99.590000   8.250000  99.760000   8.885000 ;
      RECT  99.590000   9.640000 100.195000  10.050000 ;
      RECT  99.590000  13.435000  99.760000  25.915000 ;
      RECT  99.605000  78.225000  99.935000  79.610000 ;
      RECT  99.605000  79.610000 101.600000  79.945000 ;
      RECT  99.685000  80.160000 101.835000  80.405000 ;
      RECT  99.685000  80.405000 100.100000  82.140000 ;
      RECT  99.685000  82.140000 100.715000  82.810000 ;
      RECT  99.685000  82.810000  99.950000  86.930000 ;
      RECT  99.685000  86.930000 101.650000  87.285000 ;
      RECT  99.780000 200.085000 100.650000 200.255000 ;
      RECT  99.780000 200.255000 100.450000 216.180000 ;
      RECT  99.780000 216.180000 100.970000 216.405000 ;
      RECT  99.800000  49.790000 113.910000  49.975000 ;
      RECT  99.885000  10.050000 100.195000  10.585000 ;
      RECT 100.130000  83.000000 100.300000  83.090000 ;
      RECT 100.130000  83.090000 100.305000  83.945000 ;
      RECT 100.130000  83.945000 100.300000  84.010000 ;
      RECT 100.230000  85.030000 100.815000  85.200000 ;
      RECT 100.295000   8.815000 100.840000   8.985000 ;
      RECT 100.440000  88.205000 102.660000  88.425000 ;
      RECT 100.455000 223.695000 101.305000 225.350000 ;
      RECT 100.455000 229.255000 101.305000 232.355000 ;
      RECT 100.455000 240.705000 101.305000 243.640000 ;
      RECT 100.630000  37.870000 100.800000  42.475000 ;
      RECT 100.630000  43.510000 100.800000  44.400000 ;
      RECT 100.630000  63.975000 102.070000  67.115000 ;
      RECT 100.630000  67.115000 101.375000  68.505000 ;
      RECT 100.630000  68.505000 101.480000  76.025000 ;
      RECT 100.645000  84.925000 100.815000  85.030000 ;
      RECT 100.645000  85.200000 100.815000  85.935000 ;
      RECT 100.670000   2.715000 108.535000   2.885000 ;
      RECT 100.670000   2.885000 100.840000   6.745000 ;
      RECT 100.670000   7.255000 100.840000   7.740000 ;
      RECT 100.670000   8.250000 100.840000   8.815000 ;
      RECT 100.670000   8.985000 100.840000   8.995000 ;
      RECT 100.670000   9.700000 100.840000  10.830000 ;
      RECT 100.670000  10.830000 102.455000  10.875000 ;
      RECT 100.670000  10.875000 102.460000  12.745000 ;
      RECT 100.670000  13.165000 102.460000  13.335000 ;
      RECT 100.670000  13.335000 100.840000  36.235000 ;
      RECT 100.670000  36.235000 103.000000  36.405000 ;
      RECT 100.685000  76.195000 101.480000  76.345000 ;
      RECT 100.685000  76.345000 101.375000  77.785000 ;
      RECT 100.740000  78.830000 100.910000  79.420000 ;
      RECT 100.775000  84.535000 101.445000  84.705000 ;
      RECT 100.795000 225.650000 100.965000 226.630000 ;
      RECT 100.795000 234.980000 100.965000 235.960000 ;
      RECT 100.795000 237.100000 100.965000 238.080000 ;
      RECT 100.880000 200.495000 101.410000 215.995000 ;
      RECT 100.915000  84.705000 101.445000  84.735000 ;
      RECT 100.935000  80.615000 101.255000  81.925000 ;
      RECT 101.010000  80.595000 101.180000  80.615000 ;
      RECT 101.010000  83.000000 101.180000  84.010000 ;
      RECT 101.060000 199.685000 101.590000 200.255000 ;
      RECT 101.080000   3.520000 101.250000   6.000000 ;
      RECT 101.080000   6.280000 101.250000   6.915000 ;
      RECT 101.080000   7.085000 101.250000   7.380000 ;
      RECT 101.080000   8.080000 101.250000   8.660000 ;
      RECT 101.080000   8.870000 101.250000   9.225000 ;
      RECT 101.080000   9.450000 101.250000   9.540000 ;
      RECT 101.080000   9.820000 101.250000  10.570000 ;
      RECT 101.080000  13.970000 101.250000  14.970000 ;
      RECT 101.080000  15.250000 101.250000  16.855000 ;
      RECT 101.080000  16.855000 102.480000  17.025000 ;
      RECT 101.080000  17.195000 101.250000  18.080000 ;
      RECT 101.080000  18.360000 101.250000  19.965000 ;
      RECT 101.080000  19.965000 102.480000  20.135000 ;
      RECT 101.080000  20.305000 101.250000  21.190000 ;
      RECT 101.080000  21.755000 101.250000  23.460000 ;
      RECT 101.080000  23.630000 101.665000  24.160000 ;
      RECT 101.080000  24.160000 101.250000  24.300000 ;
      RECT 101.080000  24.580000 101.250000  25.065000 ;
      RECT 101.080000  25.065000 101.610000  25.235000 ;
      RECT 101.080000  25.235000 101.250000  26.460000 ;
      RECT 101.080000  26.740000 101.250000  27.225000 ;
      RECT 101.080000  27.225000 101.610000  27.395000 ;
      RECT 101.080000  27.395000 101.250000  28.620000 ;
      RECT 101.080000  28.900000 101.250000  30.780000 ;
      RECT 101.080000  31.610000 101.250000  32.080000 ;
      RECT 101.080000  32.080000 101.720000  32.250000 ;
      RECT 101.080000  32.250000 101.250000  32.410000 ;
      RECT 101.080000  32.690000 101.250000  33.490000 ;
      RECT 101.080000  34.320000 101.250000  35.600000 ;
      RECT 101.205000  61.675000 101.375000  62.955000 ;
      RECT 101.205000  62.955000 102.070000  63.285000 ;
      RECT 101.205000  63.905000 102.070000  63.975000 ;
      RECT 101.425000  84.925000 101.595000  85.935000 ;
      RECT 101.470000   3.295000 102.480000   3.465000 ;
      RECT 101.470000   3.755000 102.480000   3.925000 ;
      RECT 101.470000   4.215000 102.480000   4.385000 ;
      RECT 101.470000   4.675000 102.480000   4.845000 ;
      RECT 101.470000   5.135000 102.480000   5.305000 ;
      RECT 101.470000   5.595000 102.480000   5.765000 ;
      RECT 101.470000   6.055000 102.480000   6.225000 ;
      RECT 101.470000   6.515000 102.480000   6.685000 ;
      RECT 101.470000   6.975000 102.480000   7.145000 ;
      RECT 101.470000   7.345000 102.480000   7.605000 ;
      RECT 101.470000   7.985000 102.480000   8.155000 ;
      RECT 101.470000   8.485000 102.480000   8.685000 ;
      RECT 101.470000   9.065000 102.480000   9.235000 ;
      RECT 101.470000   9.595000 102.480000   9.765000 ;
      RECT 101.470000  10.125000 102.480000  10.295000 ;
      RECT 101.470000  13.745000 102.480000  13.915000 ;
      RECT 101.470000  15.025000 102.480000  15.195000 ;
      RECT 101.470000  16.305000 102.480000  16.475000 ;
      RECT 101.470000  18.135000 102.480000  18.305000 ;
      RECT 101.470000  19.415000 102.480000  19.585000 ;
      RECT 101.470000  21.245000 102.480000  21.415000 ;
      RECT 101.470000  22.525000 102.480000  22.695000 ;
      RECT 101.470000  23.075000 102.480000  23.245000 ;
      RECT 101.470000  24.355000 102.480000  24.560000 ;
      RECT 101.470000  25.435000 102.480000  25.605000 ;
      RECT 101.470000  26.515000 102.480000  26.685000 ;
      RECT 101.470000  27.595000 102.480000  27.765000 ;
      RECT 101.470000  28.675000 102.480000  28.845000 ;
      RECT 101.470000  29.755000 102.480000  29.925000 ;
      RECT 101.470000  30.835000 102.480000  31.005000 ;
      RECT 101.470000  31.385000 102.480000  31.555000 ;
      RECT 101.470000  32.465000 102.480000  32.635000 ;
      RECT 101.470000  33.545000 102.480000  33.715000 ;
      RECT 101.470000  34.095000 102.480000  34.265000 ;
      RECT 101.470000  34.875000 102.480000  35.045000 ;
      RECT 101.470000  35.655000 102.480000  35.825000 ;
      RECT 101.475000  82.140000 102.440000  82.810000 ;
      RECT 101.505000   9.765000 102.035000   9.770000 ;
      RECT 101.520000  78.890000 102.380000  79.420000 ;
      RECT 101.735000 224.125000 111.735000 226.460000 ;
      RECT 101.735000 229.425000 111.735000 232.185000 ;
      RECT 101.735000 235.150000 111.735000 237.910000 ;
      RECT 101.735000 240.875000 111.735000 243.210000 ;
      RECT 101.805000  90.460000 123.885000  90.700000 ;
      RECT 101.820000  24.560000 102.480000  24.755000 ;
      RECT 101.840000 186.390000 105.860000 187.365000 ;
      RECT 101.840000 192.960000 105.860000 193.710000 ;
      RECT 101.840000 200.085000 102.510000 200.255000 ;
      RECT 101.840000 216.235000 102.510000 216.405000 ;
      RECT 101.850000  79.420000 102.380000  79.960000 ;
      RECT 101.890000  23.245000 102.480000  24.055000 ;
      RECT 101.890000  80.595000 102.060000  81.180000 ;
      RECT 101.890000  81.435000 102.060000  81.965000 ;
      RECT 101.890000  83.000000 102.060000  84.335000 ;
      RECT 101.900000  61.675000 102.070000  62.725000 ;
      RECT 102.060000  37.765000 102.670000  38.970000 ;
      RECT 102.060000  38.970000 102.910000  39.720000 ;
      RECT 102.060000  39.720000 102.670000  40.865000 ;
      RECT 102.060000  45.290000 102.230000  48.000000 ;
      RECT 102.060000  48.215000 103.670000  48.350000 ;
      RECT 102.060000  48.350000 103.830000  48.385000 ;
      RECT 102.145000  48.385000 103.830000  48.520000 ;
      RECT 102.165000 113.195000 102.835000 113.525000 ;
      RECT 102.170000  61.175000 102.680000  61.505000 ;
      RECT 102.170000  67.585000 102.680000  67.915000 ;
      RECT 102.240000  61.505000 102.610000  67.585000 ;
      RECT 102.240000  82.810000 102.440000  86.995000 ;
      RECT 102.255000  86.995000 102.425000  87.340000 ;
      RECT 102.270000 113.910000 105.270000 164.900000 ;
      RECT 102.285000  44.570000 103.400000  44.740000 ;
      RECT 102.350000  42.505000 102.880000  42.675000 ;
      RECT 102.350000  42.675000 102.520000  43.615000 ;
      RECT 102.510000  42.000000 103.180000  42.170000 ;
      RECT 102.545000  74.400000 102.715000  78.155000 ;
      RECT 102.545000  78.155000 117.835000  78.570000 ;
      RECT 102.560000  88.610000 102.730000  88.725000 ;
      RECT 102.560000  88.725000 103.115000  88.895000 ;
      RECT 102.560000  88.895000 102.730000  88.940000 ;
      RECT 102.560000  89.650000 102.730000  89.715000 ;
      RECT 102.560000  89.715000 103.115000  89.885000 ;
      RECT 102.560000  89.885000 102.730000  89.980000 ;
      RECT 102.580000  42.170000 103.110000  42.300000 ;
      RECT 102.620000  83.765000 102.790000  86.475000 ;
      RECT 102.765000  44.740000 103.400000  44.800000 ;
      RECT 102.780000  61.675000 102.950000  67.415000 ;
      RECT 102.780000  87.870000 110.985000  87.885000 ;
      RECT 102.785000  89.285000 122.600000  89.455000 ;
      RECT 102.815000  68.085000 115.865000  68.255000 ;
      RECT 102.815000  68.255000 102.985000  73.625000 ;
      RECT 102.830000  24.735000 105.415000  24.905000 ;
      RECT 102.830000  24.905000 103.000000  36.235000 ;
      RECT 102.840000  37.335000 105.095000  37.505000 ;
      RECT 102.840000  37.505000 104.980000  37.595000 ;
      RECT 102.840000  37.595000 103.220000  38.615000 ;
      RECT 102.840000  40.195000 103.010000  41.360000 ;
      RECT 102.840000  41.360000 103.760000  41.530000 ;
      RECT 102.840000  45.000000 103.010000  45.030000 ;
      RECT 102.840000  45.030000 103.385000  45.200000 ;
      RECT 102.840000  45.200000 103.010000  48.000000 ;
      RECT 102.845000  83.375000 104.125000  83.545000 ;
      RECT 102.910000  79.755000 103.080000  82.465000 ;
      RECT 102.940000 199.300000 103.470000 200.255000 ;
      RECT 102.940000 200.495000 103.470000 215.995000 ;
      RECT 103.015000   3.395000 104.485000   3.655000 ;
      RECT 103.015000  23.765000 103.395000  24.275000 ;
      RECT 103.050000  61.175000 103.560000  61.505000 ;
      RECT 103.050000  67.585000 103.560000  67.915000 ;
      RECT 103.120000  61.505000 103.490000  67.585000 ;
      RECT 103.125000  74.765000 103.295000  77.645000 ;
      RECT 103.125000  77.645000 106.815000  77.815000 ;
      RECT 103.135000  82.645000 107.495000  82.845000 ;
      RECT 103.135000  82.845000 106.375000  82.855000 ;
      RECT 103.225000  24.275000 103.395000  24.295000 ;
      RECT 103.230000  42.605000 103.400000  44.570000 ;
      RECT 103.350000  74.405000 104.700000  74.575000 ;
      RECT 103.390000  38.155000 103.560000  40.395000 ;
      RECT 103.390000  40.395000 104.100000  40.865000 ;
      RECT 103.395000  68.255000 103.565000  73.355000 ;
      RECT 103.400000  83.765000 103.570000  86.475000 ;
      RECT 103.435000  41.530000 103.760000  41.785000 ;
      RECT 103.435000  41.785000 104.055000  42.115000 ;
      RECT 103.620000  45.290000 103.790000  48.000000 ;
      RECT 103.660000  61.675000 103.830000  62.725000 ;
      RECT 103.660000  62.955000 103.830000  63.285000 ;
      RECT 103.660000  63.905000 103.830000  64.235000 ;
      RECT 103.660000  64.405000 103.830000  67.115000 ;
      RECT 103.665000   3.825000 103.835000  23.710000 ;
      RECT 103.665000  74.575000 103.835000  75.690000 ;
      RECT 103.785000  79.525000 103.955000  79.755000 ;
      RECT 103.785000  79.755000 103.960000  80.540000 ;
      RECT 103.790000  80.540000 103.960000  82.465000 ;
      RECT 103.900000 200.085000 104.570000 200.255000 ;
      RECT 103.900000 216.235000 104.570000 216.405000 ;
      RECT 103.930000  40.865000 104.100000  41.445000 ;
      RECT 103.930000  41.445000 104.395000  41.615000 ;
      RECT 103.930000  61.175000 104.440000  61.505000 ;
      RECT 103.930000  67.585000 104.440000  67.915000 ;
      RECT 104.000000  61.505000 104.370000  67.585000 ;
      RECT 104.005000  74.765000 104.175000  77.080000 ;
      RECT 104.005000  77.080000 104.535000  77.250000 ;
      RECT 104.005000  77.250000 104.175000  77.475000 ;
      RECT 104.065000  23.765000 104.485000  24.295000 ;
      RECT 104.110000  42.520000 104.395000  42.690000 ;
      RECT 104.110000  42.690000 104.280000  43.615000 ;
      RECT 104.180000  83.765000 104.350000  86.475000 ;
      RECT 104.225000  41.615000 104.395000  42.520000 ;
      RECT 104.270000  37.765000 104.440000  40.865000 ;
      RECT 104.275000  68.605000 104.445000  69.905000 ;
      RECT 104.275000  69.905000 104.810000  70.075000 ;
      RECT 104.275000  70.075000 104.445000  73.355000 ;
      RECT 104.345000  74.575000 104.515000  75.690000 ;
      RECT 104.425000  41.085000 105.095000  41.255000 ;
      RECT 104.450000  43.110000 104.980000  43.280000 ;
      RECT 104.500000  73.865000 105.850000  74.035000 ;
      RECT 104.540000  61.675000 104.710000  67.420000 ;
      RECT 104.550000  73.600000 105.800000  73.865000 ;
      RECT 104.565000  41.760000 105.095000  41.930000 ;
      RECT 104.565000  41.930000 104.875000  43.110000 ;
      RECT 104.590000  43.280000 104.760000  48.390000 ;
      RECT 104.610000  37.595000 104.980000  41.085000 ;
      RECT 104.610000  41.255000 105.095000  41.265000 ;
      RECT 104.610000  41.265000 105.575000  41.435000 ;
      RECT 104.670000  79.755000 104.840000  82.465000 ;
      RECT 104.725000 113.195000 105.395000 113.525000 ;
      RECT 104.780000  85.740000 104.950000  86.825000 ;
      RECT 104.835000   2.885000 105.245000  19.350000 ;
      RECT 104.835000  19.350000 130.720000  19.520000 ;
      RECT 104.835000  19.520000 105.415000  24.735000 ;
      RECT 104.835000  24.905000 105.415000  25.750000 ;
      RECT 104.850000  83.755000 105.020000  85.105000 ;
      RECT 104.885000  74.765000 105.055000  77.645000 ;
      RECT 105.000000 199.685000 105.530000 200.255000 ;
      RECT 105.000000 200.495000 105.530000 215.995000 ;
      RECT 105.005000  87.015000 106.925000  87.210000 ;
      RECT 105.005000  87.210000 106.005000  87.215000 ;
      RECT 105.045000  42.130000 105.575000  42.300000 ;
      RECT 105.075000  83.365000 106.075000  83.535000 ;
      RECT 105.090000  61.675000 105.260000  62.725000 ;
      RECT 105.090000  62.955000 105.260000  63.285000 ;
      RECT 105.090000  63.905000 105.260000  64.235000 ;
      RECT 105.090000  64.405000 105.260000  67.420000 ;
      RECT 105.135000  83.535000 106.015000  83.625000 ;
      RECT 105.150000  38.155000 105.435000  40.865000 ;
      RECT 105.155000  68.255000 105.325000  73.355000 ;
      RECT 105.170000  44.180000 106.730000  44.350000 ;
      RECT 105.170000  44.350000 105.340000  45.760000 ;
      RECT 105.170000  45.760000 107.700000  45.930000 ;
      RECT 105.170000  46.100000 105.340000  46.335000 ;
      RECT 105.170000  46.335000 105.700000  46.505000 ;
      RECT 105.170000  46.505000 105.340000  48.380000 ;
      RECT 105.230000  25.750000 105.415000  26.920000 ;
      RECT 105.230000  26.920000 124.675000  27.090000 ;
      RECT 105.265000  40.865000 105.435000  41.095000 ;
      RECT 105.265000  41.435000 105.575000  42.130000 ;
      RECT 105.270000  42.840000 105.440000  44.010000 ;
      RECT 105.430000  61.175000 105.940000  61.505000 ;
      RECT 105.430000  67.585000 105.940000  67.915000 ;
      RECT 105.500000  61.505000 105.870000  66.375000 ;
      RECT 105.500000  66.375000 106.030000  66.545000 ;
      RECT 105.500000  66.545000 105.870000  67.585000 ;
      RECT 105.505000   3.295000 108.555000   3.465000 ;
      RECT 105.505000   3.465000 105.675000   5.055000 ;
      RECT 105.505000   5.055000 108.555000   5.225000 ;
      RECT 105.545000  79.525000 105.715000  79.755000 ;
      RECT 105.545000  79.755000 105.720000  80.540000 ;
      RECT 105.550000  80.540000 105.720000  82.465000 ;
      RECT 105.555000  42.470000 106.905000  42.640000 ;
      RECT 105.655000  42.640000 106.905000  42.670000 ;
      RECT 105.700000  42.840000 105.870000  44.180000 ;
      RECT 105.730000  37.765000 105.900000  40.845000 ;
      RECT 105.765000  74.765000 106.205000  74.935000 ;
      RECT 105.765000  74.935000 105.935000  77.475000 ;
      RECT 105.830000  19.870000 106.000000  22.580000 ;
      RECT 105.830000  23.850000 106.000000  26.560000 ;
      RECT 105.845000   4.175000 108.555000   4.345000 ;
      RECT 105.845000   5.935000 108.555000   6.105000 ;
      RECT 105.855000  69.905000 106.385000  70.075000 ;
      RECT 105.960000  83.815000 106.360000  86.825000 ;
      RECT 105.960000 200.085000 106.630000 200.255000 ;
      RECT 105.960000 216.235000 106.630000 216.405000 ;
      RECT 105.995000  22.750000 111.055000  23.680000 ;
      RECT 106.000000   7.720000 106.230000   8.950000 ;
      RECT 106.000000  11.700000 106.230000  12.710000 ;
      RECT 106.030000   7.200000 109.970000   7.370000 ;
      RECT 106.030000   7.370000 106.200000   7.720000 ;
      RECT 106.030000   8.950000 106.200000  11.700000 ;
      RECT 106.030000  12.710000 106.200000  12.740000 ;
      RECT 106.030000  13.900000 106.200000  18.900000 ;
      RECT 106.035000  68.605000 106.205000  69.905000 ;
      RECT 106.035000  70.075000 106.205000  74.765000 ;
      RECT 106.040000  61.675000 106.210000  66.145000 ;
      RECT 106.130000  42.840000 106.300000  44.010000 ;
      RECT 106.130000  83.755000 106.300000  83.815000 ;
      RECT 106.310000  61.175000 106.820000  61.505000 ;
      RECT 106.310000  67.585000 106.820000  67.915000 ;
      RECT 106.330000 188.775000 121.065000 189.945000 ;
      RECT 106.335000 186.220000 121.065000 188.775000 ;
      RECT 106.335000 189.945000 121.065000 191.905000 ;
      RECT 106.335000 191.905000 143.505000 193.515000 ;
      RECT 106.335000 193.515000 158.850000 194.595000 ;
      RECT 106.350000  44.580000 106.520000  45.280000 ;
      RECT 106.350000  45.280000 107.025000  45.450000 ;
      RECT 106.350000  45.450000 106.520000  45.590000 ;
      RECT 106.350000  46.100000 106.520000  48.550000 ;
      RECT 106.350000  48.550000 109.240000  48.720000 ;
      RECT 106.380000  61.505000 106.750000  67.585000 ;
      RECT 106.430000  79.755000 106.600000  82.465000 ;
      RECT 106.560000  42.840000 106.730000  44.180000 ;
      RECT 106.590000  83.800000 107.180000  83.970000 ;
      RECT 106.590000  83.970000 106.925000  87.015000 ;
      RECT 106.610000   7.720000 106.780000  11.320000 ;
      RECT 106.610000  11.320000 107.140000  11.490000 ;
      RECT 106.610000  11.490000 106.780000  12.470000 ;
      RECT 106.610000  14.170000 106.780000  18.920000 ;
      RECT 106.645000  74.765000 106.815000  77.645000 ;
      RECT 106.710000  19.870000 106.880000  22.580000 ;
      RECT 106.710000  23.850000 106.880000  26.560000 ;
      RECT 106.780000 113.910000 109.780000 164.900000 ;
      RECT 106.850000  46.165000 107.180000  47.015000 ;
      RECT 106.915000  68.255000 107.085000  73.355000 ;
      RECT 106.930000  47.015000 107.100000  47.625000 ;
      RECT 106.990000  42.840000 107.160000  44.010000 ;
      RECT 106.990000  61.675000 107.160000  62.725000 ;
      RECT 106.990000  62.955000 107.160000  63.285000 ;
      RECT 106.990000  63.905000 107.160000  64.235000 ;
      RECT 106.990000  64.405000 107.160000  67.115000 ;
      RECT 107.015000   9.730000 107.660000   9.900000 ;
      RECT 107.060000 199.300000 107.590000 200.255000 ;
      RECT 107.060000 200.495000 107.590000 215.995000 ;
      RECT 107.075000  37.870000 107.245000  40.870000 ;
      RECT 107.195000  74.400000 107.365000  78.155000 ;
      RECT 107.195000  84.215000 107.365000  86.925000 ;
      RECT 107.260000  42.470000 108.610000  42.475000 ;
      RECT 107.260000  42.475000 109.920000  42.645000 ;
      RECT 107.295000  41.360000 107.825000  41.530000 ;
      RECT 107.295000  80.270000 107.495000  82.645000 ;
      RECT 107.310000  79.260000 107.480000  79.990000 ;
      RECT 107.330000  61.175000 107.860000  61.345000 ;
      RECT 107.330000  61.345000 107.840000  61.505000 ;
      RECT 107.330000  67.585000 107.840000  67.915000 ;
      RECT 107.400000  61.505000 107.770000  67.585000 ;
      RECT 107.420000  42.840000 107.590000  44.180000 ;
      RECT 107.420000  44.180000 109.240000  44.350000 ;
      RECT 107.435000  69.905000 107.965000  70.075000 ;
      RECT 107.490000   7.720000 107.660000   9.730000 ;
      RECT 107.490000   9.900000 107.660000  18.920000 ;
      RECT 107.530000  44.580000 107.700000  45.760000 ;
      RECT 107.530000  45.930000 107.700000  47.080000 ;
      RECT 107.530000  47.370000 108.400000  48.380000 ;
      RECT 107.530000  87.275000 109.560000  87.445000 ;
      RECT 107.590000  19.870000 107.760000  22.580000 ;
      RECT 107.590000  23.850000 107.760000  26.560000 ;
      RECT 107.590000  74.405000 108.600000  74.575000 ;
      RECT 107.590000  87.445000 109.500000  87.455000 ;
      RECT 107.650000  74.000000 108.540000  74.405000 ;
      RECT 107.655000  37.840000 111.895000  38.010000 ;
      RECT 107.655000  38.010000 107.825000  41.360000 ;
      RECT 107.775000  77.080000 108.305000  77.250000 ;
      RECT 107.795000  68.605000 107.965000  69.905000 ;
      RECT 107.795000  70.075000 107.965000  73.355000 ;
      RECT 107.830000  13.490000 108.500000  13.660000 ;
      RECT 107.850000  42.840000 108.020000  44.010000 ;
      RECT 107.860000  79.265000 110.760000  79.435000 ;
      RECT 107.860000  80.930000 110.760000  81.095000 ;
      RECT 107.860000  81.095000 109.070000  81.100000 ;
      RECT 107.870000  46.335000 108.400000  47.370000 ;
      RECT 107.880000  37.335000 109.910000  37.505000 ;
      RECT 107.880000  82.625000 110.530000  83.565000 ;
      RECT 107.940000  61.675000 108.110000  66.145000 ;
      RECT 108.020000 200.085000 108.690000 200.255000 ;
      RECT 108.020000 216.235000 108.690000 216.405000 ;
      RECT 108.040000   7.370000 108.210000  12.650000 ;
      RECT 108.050000  80.045000 110.760000  80.215000 ;
      RECT 108.050000  80.925000 110.760000  80.930000 ;
      RECT 108.050000  81.805000 110.760000  81.975000 ;
      RECT 108.055000  49.760000 113.910000  49.790000 ;
      RECT 108.075000  74.765000 108.245000  77.080000 ;
      RECT 108.075000  77.250000 108.245000  77.475000 ;
      RECT 108.210000  61.175000 108.720000  61.505000 ;
      RECT 108.210000  67.585000 108.720000  67.915000 ;
      RECT 108.280000  42.840000 108.450000  44.180000 ;
      RECT 108.280000  61.505000 108.650000  67.585000 ;
      RECT 108.290000  86.680000 108.820000  86.850000 ;
      RECT 108.330000  12.950000 110.635000  13.070000 ;
      RECT 108.330000  13.070000 110.625000  13.120000 ;
      RECT 108.350000  45.280000 108.880000  45.450000 ;
      RECT 108.370000  14.170000 108.540000  18.920000 ;
      RECT 108.390000  34.015000 111.390000  34.325000 ;
      RECT 108.395000  29.275000 111.105000  29.445000 ;
      RECT 108.395000  30.555000 111.305000  30.725000 ;
      RECT 108.470000  19.870000 108.640000  22.580000 ;
      RECT 108.470000  23.850000 108.640000  26.560000 ;
      RECT 108.475000  84.215000 108.645000  86.680000 ;
      RECT 108.475000  86.850000 108.645000  86.925000 ;
      RECT 108.535000  38.180000 108.795000  41.160000 ;
      RECT 108.560000  11.320000 109.090000  11.490000 ;
      RECT 108.675000  68.255000 108.845000  73.355000 ;
      RECT 108.700000  31.870000 111.410000  32.040000 ;
      RECT 108.700000  32.650000 111.410000  32.820000 ;
      RECT 108.700000  33.430000 111.410000  33.600000 ;
      RECT 108.710000  42.840000 108.880000  44.010000 ;
      RECT 108.710000  44.580000 108.880000  45.280000 ;
      RECT 108.710000  45.450000 108.880000  47.080000 ;
      RECT 108.710000  47.370000 109.240000  48.550000 ;
      RECT 108.745000   3.515000 108.915000   5.885000 ;
      RECT 108.890000  61.675000 109.610000  62.725000 ;
      RECT 108.890000  62.955000 109.610000  63.285000 ;
      RECT 108.890000  63.905000 109.610000  64.235000 ;
      RECT 108.890000  64.405000 109.060000  67.420000 ;
      RECT 108.920000   7.720000 109.090000  11.320000 ;
      RECT 108.920000  11.490000 109.090000  12.470000 ;
      RECT 108.920000  14.170000 109.090000  18.920000 ;
      RECT 108.955000  74.400000 109.125000  78.155000 ;
      RECT 108.995000  38.180000 109.255000  41.160000 ;
      RECT 109.050000  43.095000 109.580000  43.265000 ;
      RECT 109.050000  44.350000 109.240000  47.370000 ;
      RECT 109.120000 199.685000 109.650000 200.255000 ;
      RECT 109.120000 200.495000 109.650000 215.995000 ;
      RECT 109.140000  13.570000 114.020000  13.660000 ;
      RECT 109.140000  13.660000 111.470000  13.740000 ;
      RECT 109.170000  41.360000 109.700000  41.530000 ;
      RECT 109.255000  68.255000 109.425000  73.625000 ;
      RECT 109.270000  13.490000 114.020000  13.570000 ;
      RECT 109.315000   3.295000 110.325000   3.465000 ;
      RECT 109.315000   3.755000 110.325000   3.925000 ;
      RECT 109.315000   4.215000 110.325000   4.385000 ;
      RECT 109.350000  19.870000 109.520000  22.580000 ;
      RECT 109.350000  23.850000 109.520000  26.560000 ;
      RECT 109.350000  41.530000 109.520000  42.305000 ;
      RECT 109.385000  81.775000 110.645000  81.805000 ;
      RECT 109.410000  43.265000 109.580000  48.390000 ;
      RECT 109.440000  64.235000 109.610000  67.115000 ;
      RECT 109.450000  74.405000 110.460000  74.575000 ;
      RECT 109.495000  74.575000 109.665000  75.690000 ;
      RECT 109.555000  31.820000 110.195000  31.870000 ;
      RECT 109.555000  32.040000 110.195000  32.080000 ;
      RECT 109.555000  33.385000 110.195000  33.430000 ;
      RECT 109.555000  33.600000 110.195000  33.645000 ;
      RECT 109.620000  67.515000 110.150000  67.585000 ;
      RECT 109.620000  67.585000 110.220000  67.685000 ;
      RECT 109.655000  77.080000 110.185000  77.250000 ;
      RECT 109.710000  61.175000 110.220000  61.505000 ;
      RECT 109.710000  67.685000 110.220000  67.915000 ;
      RECT 109.750000  42.645000 109.920000  43.405000 ;
      RECT 109.750000  43.405000 110.400000  44.415000 ;
      RECT 109.755000  84.215000 109.925000  86.925000 ;
      RECT 109.780000  61.505000 110.150000  67.515000 ;
      RECT 109.800000   7.370000 109.970000  12.650000 ;
      RECT 109.800000  14.170000 109.970000  18.920000 ;
      RECT 109.835000  68.605000 110.005000  69.905000 ;
      RECT 109.835000  69.905000 110.365000  70.075000 ;
      RECT 109.835000  70.075000 110.005000  73.815000 ;
      RECT 109.835000  73.815000 113.525000  73.985000 ;
      RECT 109.835000  74.765000 110.005000  77.080000 ;
      RECT 109.835000  77.250000 110.005000  77.475000 ;
      RECT 109.870000  41.290000 110.540000  41.460000 ;
      RECT 109.870000  46.335000 110.400000  46.505000 ;
      RECT 109.890000  47.855000 110.060000  48.465000 ;
      RECT 109.890000  48.465000 115.420000  48.635000 ;
      RECT 109.930000  42.030000 110.460000  42.200000 ;
      RECT 109.965000  38.180000 110.135000  41.290000 ;
      RECT 109.965000  41.460000 110.460000  42.030000 ;
      RECT 110.080000 200.085000 110.750000 200.255000 ;
      RECT 110.080000 216.235000 110.750000 216.405000 ;
      RECT 110.090000  87.275000 112.120000  87.445000 ;
      RECT 110.105000  12.900000 110.635000  12.950000 ;
      RECT 110.120000  37.335000 112.385000  37.505000 ;
      RECT 110.150000  87.445000 112.060000  87.455000 ;
      RECT 110.175000  74.575000 110.345000  75.690000 ;
      RECT 110.215000   6.510000 110.745000   6.680000 ;
      RECT 110.230000  19.870000 110.400000  22.580000 ;
      RECT 110.230000  23.850000 110.400000  26.560000 ;
      RECT 110.230000  44.415000 110.400000  46.335000 ;
      RECT 110.230000  46.505000 110.400000  48.085000 ;
      RECT 110.320000  61.675000 110.490000  67.415000 ;
      RECT 110.500000  11.320000 111.030000  11.490000 ;
      RECT 110.525000   2.995000 110.695000   4.160000 ;
      RECT 110.525000   4.500000 110.695000   5.170000 ;
      RECT 110.550000   5.680000 110.720000   6.510000 ;
      RECT 110.570000  45.000000 111.100000  45.170000 ;
      RECT 110.590000  61.175000 111.100000  61.505000 ;
      RECT 110.590000  67.585000 111.100000  67.915000 ;
      RECT 110.630000  41.635000 110.880000  42.305000 ;
      RECT 110.660000  61.505000 111.030000  67.585000 ;
      RECT 110.665000  41.580000 110.880000  41.635000 ;
      RECT 110.665000  42.305000 110.835000  43.405000 ;
      RECT 110.665000  43.405000 110.860000  44.415000 ;
      RECT 110.680000   7.720000 110.850000  11.320000 ;
      RECT 110.680000  11.490000 110.850000  12.470000 ;
      RECT 110.680000  14.170000 110.850000  18.920000 ;
      RECT 110.680000  32.605000 111.320000  32.650000 ;
      RECT 110.680000  32.820000 111.320000  32.865000 ;
      RECT 110.690000  45.170000 110.860000  48.085000 ;
      RECT 110.705000  83.310000 111.235000  83.480000 ;
      RECT 110.710000  38.180000 111.015000  40.890000 ;
      RECT 110.710000  40.890000 110.880000  41.580000 ;
      RECT 110.715000  68.255000 110.885000  73.355000 ;
      RECT 110.715000  74.400000 110.885000  78.155000 ;
      RECT 110.720000   7.040000 111.390000   7.210000 ;
      RECT 110.860000   7.010000 111.390000   7.040000 ;
      RECT 110.865000   3.295000 116.005000   3.445000 ;
      RECT 110.865000   3.445000 115.955000   3.465000 ;
      RECT 110.865000   3.465000 111.035000   4.740000 ;
      RECT 110.865000   4.740000 116.005000   4.910000 ;
      RECT 110.875000  85.230000 111.405000  85.400000 ;
      RECT 110.905000  12.950000 111.935000  13.150000 ;
      RECT 110.975000   2.680000 135.050000   2.850000 ;
      RECT 111.010000  79.315000 111.575000  81.675000 ;
      RECT 111.010000  81.675000 111.235000  83.310000 ;
      RECT 111.030000   5.200000 115.955000   5.390000 ;
      RECT 111.030000   5.390000 111.200000   6.700000 ;
      RECT 111.030000  42.400000 111.560000  42.570000 ;
      RECT 111.030000  42.570000 111.440000  44.585000 ;
      RECT 111.030000  44.585000 111.520000  44.740000 ;
      RECT 111.030000  45.375000 111.520000  45.665000 ;
      RECT 111.030000  45.665000 111.320000  48.085000 ;
      RECT 111.035000  84.215000 111.205000  85.230000 ;
      RECT 111.035000  85.400000 111.205000  86.925000 ;
      RECT 111.050000  42.030000 112.080000  42.200000 ;
      RECT 111.055000  74.405000 112.185000  74.575000 ;
      RECT 111.055000  74.575000 111.225000  75.690000 ;
      RECT 111.110000  19.870000 111.280000  22.580000 ;
      RECT 111.110000  23.850000 111.280000  26.560000 ;
      RECT 111.140000  83.800000 111.730000  83.970000 ;
      RECT 111.150000  41.290000 111.895000  41.460000 ;
      RECT 111.180000 199.300000 111.710000 200.255000 ;
      RECT 111.180000 200.495000 111.710000 215.995000 ;
      RECT 111.185000 113.195000 111.855000 113.525000 ;
      RECT 111.200000  61.675000 111.370000  62.725000 ;
      RECT 111.200000  62.955000 112.180000  63.285000 ;
      RECT 111.200000  63.905000 112.180000  67.115000 ;
      RECT 111.205000   3.675000 115.695000   3.755000 ;
      RECT 111.205000   3.755000 115.955000   3.925000 ;
      RECT 111.205000   4.280000 115.955000   4.450000 ;
      RECT 111.220000  41.460000 111.750000  41.530000 ;
      RECT 111.270000  44.740000 111.520000  45.375000 ;
      RECT 111.290000 113.910000 114.290000 164.900000 ;
      RECT 111.335000  22.750000 123.980000  23.680000 ;
      RECT 111.380000   7.380000 111.910000   7.550000 ;
      RECT 111.400000   4.450000 115.890000   4.455000 ;
      RECT 111.405000  13.150000 111.935000  13.320000 ;
      RECT 111.405000  81.955000 111.730000  83.800000 ;
      RECT 111.415000  69.905000 111.945000  70.075000 ;
      RECT 111.415000  77.080000 111.945000  77.250000 ;
      RECT 111.490000  56.690000 111.660000  60.405000 ;
      RECT 111.500000  49.280000 113.680000  49.735000 ;
      RECT 111.500000  49.735000 113.910000  49.760000 ;
      RECT 111.520000  48.105000 112.275000  48.275000 ;
      RECT 111.560000   5.690000 111.730000   7.380000 ;
      RECT 111.560000   7.550000 111.730000  12.470000 ;
      RECT 111.560000  14.170000 111.730000  18.920000 ;
      RECT 111.595000  68.605000 111.765000  69.905000 ;
      RECT 111.595000  70.075000 111.765000  73.815000 ;
      RECT 111.595000  74.765000 111.765000  77.080000 ;
      RECT 111.595000  77.250000 111.765000  77.475000 ;
      RECT 111.610000  43.405000 111.900000  44.415000 ;
      RECT 111.630000  32.095000 111.800000  33.375000 ;
      RECT 111.655000  29.500000 111.830000  30.030000 ;
      RECT 111.655000  30.030000 111.825000  30.500000 ;
      RECT 111.725000  38.010000 111.895000  41.290000 ;
      RECT 111.730000  44.415000 111.900000  44.520000 ;
      RECT 111.730000  44.520000 111.935000  45.300000 ;
      RECT 111.745000  46.335000 112.275000  46.505000 ;
      RECT 111.765000  53.600000 113.590000  53.770000 ;
      RECT 111.765000  53.770000 113.770000  53.935000 ;
      RECT 111.765000  53.935000 114.730000  54.055000 ;
      RECT 111.765000  54.055000 115.890000  54.385000 ;
      RECT 111.765000  54.385000 111.935000  55.575000 ;
      RECT 111.805000  42.510000 112.340000  43.085000 ;
      RECT 111.910000  41.635000 112.080000  42.030000 ;
      RECT 111.910000  42.200000 112.080000  42.305000 ;
      RECT 111.915000  79.965000 115.685000  79.970000 ;
      RECT 111.915000  79.970000 116.805000  80.135000 ;
      RECT 111.915000  81.725000 115.550000  81.730000 ;
      RECT 111.915000  81.730000 116.805000  81.895000 ;
      RECT 111.930000   7.010000 112.460000   7.180000 ;
      RECT 111.930000   8.900000 112.460000   9.070000 ;
      RECT 111.935000  74.575000 112.105000  75.690000 ;
      RECT 111.985000  87.870000 175.800000  87.885000 ;
      RECT 112.010000  61.675000 112.180000  62.955000 ;
      RECT 112.010000  67.115000 112.180000  67.415000 ;
      RECT 112.055000  79.090000 116.805000  79.260000 ;
      RECT 112.055000  80.135000 116.805000  80.140000 ;
      RECT 112.055000  80.850000 116.805000  81.020000 ;
      RECT 112.055000  81.895000 116.805000  81.900000 ;
      RECT 112.055000  82.610000 116.805000  82.780000 ;
      RECT 112.070000  43.405000 112.275000  44.415000 ;
      RECT 112.070000  56.670000 112.240000  60.405000 ;
      RECT 112.105000  44.415000 112.275000  46.335000 ;
      RECT 112.105000  46.505000 112.275000  48.105000 ;
      RECT 112.110000   5.690000 112.280000   7.010000 ;
      RECT 112.110000   7.180000 112.280000   8.900000 ;
      RECT 112.110000   9.070000 112.280000  12.470000 ;
      RECT 112.140000 200.085000 112.810000 200.255000 ;
      RECT 112.140000 216.235000 112.810000 216.405000 ;
      RECT 112.165000 223.695000 113.015000 225.350000 ;
      RECT 112.165000 229.255000 113.015000 232.355000 ;
      RECT 112.165000 240.705000 113.015000 243.640000 ;
      RECT 112.215000  13.120000 112.745000  13.320000 ;
      RECT 112.215000  37.505000 112.385000  39.510000 ;
      RECT 112.265000  12.950000 112.935000  13.120000 ;
      RECT 112.315000  84.215000 112.485000  86.925000 ;
      RECT 112.360000  54.555000 112.530000  55.495000 ;
      RECT 112.360000  55.495000 112.890000  55.665000 ;
      RECT 112.390000  19.870000 112.560000  22.580000 ;
      RECT 112.390000  23.850000 112.560000  26.560000 ;
      RECT 112.410000  55.835000 113.080000  55.895000 ;
      RECT 112.410000  55.895000 113.125000  56.065000 ;
      RECT 112.410000  56.065000 113.080000  56.345000 ;
      RECT 112.410000  56.345000 112.680000  58.805000 ;
      RECT 112.410000  58.805000 113.020000  60.665000 ;
      RECT 112.410000  60.665000 115.175000  60.835000 ;
      RECT 112.440000  14.170000 112.610000  18.920000 ;
      RECT 112.475000  68.255000 112.645000  73.355000 ;
      RECT 112.475000  74.400000 112.645000  78.155000 ;
      RECT 112.505000 225.650000 112.675000 226.630000 ;
      RECT 112.505000 234.980000 112.675000 235.960000 ;
      RECT 112.505000 237.100000 112.675000 238.080000 ;
      RECT 112.570000  37.870000 113.005000  40.870000 ;
      RECT 112.570000  40.870000 112.740000  44.425000 ;
      RECT 112.570000  47.855000 112.740000  48.465000 ;
      RECT 112.595000  61.675000 112.765000  63.495000 ;
      RECT 112.595000  64.405000 112.765000  67.115000 ;
      RECT 112.620000   7.380000 116.060000   7.430000 ;
      RECT 112.620000   7.430000 113.150000   7.550000 ;
      RECT 112.630000   7.070000 114.085000   7.260000 ;
      RECT 112.630000   7.260000 116.060000   7.380000 ;
      RECT 112.640000   5.390000 112.810000   6.700000 ;
      RECT 112.810000  11.320000 113.340000  11.490000 ;
      RECT 112.850000  56.515000 114.055000  56.700000 ;
      RECT 112.850000  56.700000 113.020000  57.680000 ;
      RECT 112.865000  61.175000 113.440000  61.235000 ;
      RECT 112.865000  61.235000 113.375000  61.505000 ;
      RECT 112.865000  67.585000 113.375000  67.915000 ;
      RECT 112.865000  84.275000 113.035000  87.055000 ;
      RECT 112.910000  61.065000 113.440000  61.175000 ;
      RECT 112.935000  61.505000 113.305000  67.585000 ;
      RECT 112.970000  42.510000 113.505000  43.085000 ;
      RECT 112.980000   6.510000 113.510000   6.680000 ;
      RECT 112.990000   7.720000 113.160000  11.320000 ;
      RECT 112.990000  11.490000 113.160000  12.470000 ;
      RECT 113.025000  74.765000 113.195000  77.080000 ;
      RECT 113.025000  77.080000 113.555000  77.250000 ;
      RECT 113.025000  77.250000 113.195000  77.475000 ;
      RECT 113.035000  43.405000 113.240000  44.415000 ;
      RECT 113.035000  44.415000 113.205000  46.335000 ;
      RECT 113.035000  46.335000 113.565000  46.505000 ;
      RECT 113.035000  46.505000 113.205000  48.105000 ;
      RECT 113.035000  48.105000 113.790000  48.275000 ;
      RECT 113.120000   5.680000 113.290000   6.510000 ;
      RECT 113.175000  69.905000 113.705000  70.075000 ;
      RECT 113.200000  87.275000 115.770000  87.475000 ;
      RECT 113.215000  12.910000 113.745000  12.950000 ;
      RECT 113.215000  12.950000 113.885000  13.120000 ;
      RECT 113.230000  41.635000 113.400000  42.030000 ;
      RECT 113.230000  42.030000 114.260000  42.200000 ;
      RECT 113.230000  42.200000 113.400000  42.305000 ;
      RECT 113.240000  54.385000 113.770000  54.660000 ;
      RECT 113.240000  54.660000 113.410000  55.565000 ;
      RECT 113.240000 199.685000 113.770000 200.255000 ;
      RECT 113.240000 200.495000 113.770000 215.995000 ;
      RECT 113.320000  14.170000 113.490000  18.920000 ;
      RECT 113.355000  68.605000 113.525000  69.905000 ;
      RECT 113.355000  70.075000 113.525000  73.815000 ;
      RECT 113.355000  73.985000 113.525000  74.340000 ;
      RECT 113.355000  74.340000 115.835000  74.595000 ;
      RECT 113.375000  44.630000 113.545000  45.300000 ;
      RECT 113.415000  37.840000 117.655000  38.010000 ;
      RECT 113.415000  38.010000 113.585000  41.290000 ;
      RECT 113.415000  41.290000 114.160000  41.460000 ;
      RECT 113.445000 224.125000 123.445000 226.460000 ;
      RECT 113.445000 229.425000 123.445000 232.185000 ;
      RECT 113.445000 235.150000 123.445000 237.910000 ;
      RECT 113.445000 240.875000 123.445000 243.210000 ;
      RECT 113.475000  61.800000 113.645000  67.420000 ;
      RECT 113.485000  86.680000 114.015000  86.850000 ;
      RECT 113.500000  56.870000 114.395000  57.040000 ;
      RECT 113.500000  57.040000 113.670000  60.015000 ;
      RECT 113.525000  56.265000 114.055000  56.515000 ;
      RECT 113.530000  43.405000 113.700000  44.415000 ;
      RECT 113.545000  55.735000 114.055000  56.265000 ;
      RECT 113.560000  41.460000 114.090000  41.530000 ;
      RECT 113.570000  37.335000 114.240000  37.505000 ;
      RECT 113.645000  84.345000 113.815000  86.680000 ;
      RECT 113.645000  86.850000 113.815000  87.055000 ;
      RECT 113.655000  61.435000 114.255000  61.505000 ;
      RECT 113.655000  61.505000 114.185000  61.605000 ;
      RECT 113.670000  19.870000 113.840000  22.580000 ;
      RECT 113.670000  23.850000 113.840000  26.560000 ;
      RECT 113.740000  44.585000 114.280000  44.740000 ;
      RECT 113.740000  44.740000 114.040000  45.375000 ;
      RECT 113.740000  45.375000 114.280000  45.665000 ;
      RECT 113.745000  61.175000 114.255000  61.435000 ;
      RECT 113.745000  67.585000 114.255000  67.915000 ;
      RECT 113.745000 113.195000 114.415000 113.525000 ;
      RECT 113.750000  42.400000 114.280000  42.570000 ;
      RECT 113.815000  61.605000 114.185000  67.585000 ;
      RECT 113.815000  73.865000 114.825000  74.035000 ;
      RECT 113.850000  52.355000 114.360000  52.685000 ;
      RECT 113.870000   7.720000 114.040000  12.470000 ;
      RECT 113.870000  42.570000 114.280000  44.585000 ;
      RECT 113.875000  73.600000 114.765000  73.865000 ;
      RECT 113.905000  74.595000 114.075000  77.475000 ;
      RECT 113.915000   5.660000 114.085000   7.070000 ;
      RECT 113.970000  36.980000 114.140000  37.335000 ;
      RECT 113.970000  37.505000 114.140000  37.510000 ;
      RECT 113.990000  45.665000 114.280000  48.085000 ;
      RECT 114.060000  50.535000 115.150000  50.705000 ;
      RECT 114.060000  50.705000 114.230000  52.355000 ;
      RECT 114.060000  52.685000 114.230000  52.840000 ;
      RECT 114.120000  54.555000 114.395000  54.905000 ;
      RECT 114.120000  54.905000 114.650000  55.075000 ;
      RECT 114.120000  55.075000 114.395000  55.565000 ;
      RECT 114.200000  14.170000 114.370000  18.920000 ;
      RECT 114.200000 200.085000 114.870000 200.255000 ;
      RECT 114.200000 216.235000 114.870000 216.405000 ;
      RECT 114.210000  45.000000 114.740000  45.170000 ;
      RECT 114.220000   7.720000 114.750000   9.070000 ;
      RECT 114.225000  55.565000 114.395000  56.870000 ;
      RECT 114.235000  68.255000 114.405000  73.355000 ;
      RECT 114.255000  49.415000 114.925000  50.365000 ;
      RECT 114.280000  57.305000 114.450000  60.405000 ;
      RECT 114.295000  38.180000 114.600000  39.675000 ;
      RECT 114.295000  39.675000 114.825000  39.845000 ;
      RECT 114.295000  39.845000 114.600000  40.890000 ;
      RECT 114.320000   6.920000 114.990000   7.090000 ;
      RECT 114.355000  61.675000 114.525000  62.740000 ;
      RECT 114.355000  62.910000 114.525000  63.285000 ;
      RECT 114.355000  63.905000 114.525000  64.235000 ;
      RECT 114.355000  64.405000 114.525000  67.115000 ;
      RECT 114.425000  84.275000 114.595000  87.055000 ;
      RECT 114.430000  40.890000 114.600000  41.580000 ;
      RECT 114.430000  41.580000 114.645000  41.635000 ;
      RECT 114.430000  41.635000 114.680000  42.305000 ;
      RECT 114.450000   9.380000 114.620000   9.645000 ;
      RECT 114.450000   9.645000 120.800000  10.760000 ;
      RECT 114.450000  10.760000 125.745000  10.930000 ;
      RECT 114.450000  10.930000 119.090000  11.370000 ;
      RECT 114.450000  43.405000 114.645000  44.415000 ;
      RECT 114.450000  45.170000 114.620000  48.085000 ;
      RECT 114.475000  42.305000 114.645000  43.405000 ;
      RECT 114.480000  11.720000 114.650000  12.730000 ;
      RECT 114.520000  37.335000 115.190000  37.505000 ;
      RECT 114.520000  50.875000 114.730000  51.885000 ;
      RECT 114.520000  52.875000 114.730000  53.935000 ;
      RECT 114.530000  51.885000 114.730000  52.875000 ;
      RECT 114.565000  54.385000 115.890000  54.660000 ;
      RECT 114.565000  55.525000 115.095000  57.005000 ;
      RECT 114.565000  57.005000 115.230000  57.175000 ;
      RECT 114.605000  77.080000 115.135000  77.250000 ;
      RECT 114.625000  61.175000 115.135000  61.505000 ;
      RECT 114.625000  67.585000 115.135000  67.915000 ;
      RECT 114.695000  61.505000 115.065000  67.585000 ;
      RECT 114.755000  69.905000 115.285000  70.075000 ;
      RECT 114.770000  41.290000 115.440000  41.460000 ;
      RECT 114.780000  13.900000 114.950000  17.270000 ;
      RECT 114.780000  17.270000 118.750000  18.040000 ;
      RECT 114.780000  18.040000 128.285000  18.210000 ;
      RECT 114.785000  74.765000 114.955000  77.080000 ;
      RECT 114.785000  77.250000 114.955000  77.475000 ;
      RECT 114.850000  41.460000 115.345000  42.030000 ;
      RECT 114.850000  42.030000 115.380000  42.200000 ;
      RECT 114.910000  43.405000 115.560000  44.415000 ;
      RECT 114.910000  44.415000 115.080000  46.335000 ;
      RECT 114.910000  46.335000 115.440000  46.505000 ;
      RECT 114.910000  46.505000 115.080000  48.085000 ;
      RECT 114.950000  19.870000 115.120000  22.580000 ;
      RECT 114.950000  23.850000 115.120000  26.560000 ;
      RECT 114.980000  50.705000 115.150000  51.885000 ;
      RECT 114.980000  52.875000 115.150000  53.885000 ;
      RECT 115.000000   9.010000 115.715000   9.180000 ;
      RECT 115.000000   9.180000 115.530000   9.475000 ;
      RECT 115.005000  52.230000 115.535000  52.400000 ;
      RECT 115.025000  85.230000 115.555000  85.400000 ;
      RECT 115.060000  57.175000 115.230000  60.015000 ;
      RECT 115.065000  12.725000 115.530000  13.005000 ;
      RECT 115.065000  13.005000 115.345000  13.720000 ;
      RECT 115.065000  13.720000 116.745000  13.770000 ;
      RECT 115.100000  49.785000 115.955000  49.955000 ;
      RECT 115.115000  68.605000 115.285000  69.905000 ;
      RECT 115.115000  70.075000 115.285000  74.340000 ;
      RECT 115.120000  13.770000 116.745000  14.000000 ;
      RECT 115.120000  14.000000 115.530000  14.210000 ;
      RECT 115.175000  38.180000 115.345000  41.290000 ;
      RECT 115.195000   5.390000 115.365000   6.670000 ;
      RECT 115.205000  52.095000 115.535000  52.230000 ;
      RECT 115.205000  52.400000 115.535000  52.605000 ;
      RECT 115.205000  84.345000 115.375000  85.230000 ;
      RECT 115.205000  85.400000 115.375000  87.055000 ;
      RECT 115.235000  61.675000 115.405000  64.025000 ;
      RECT 115.235000  64.025000 116.495000  64.235000 ;
      RECT 115.235000  64.235000 115.405000  67.420000 ;
      RECT 115.250000  47.855000 115.420000  48.465000 ;
      RECT 115.300000 199.300000 115.830000 200.255000 ;
      RECT 115.300000 200.495000 115.830000 215.995000 ;
      RECT 115.360000  11.720000 115.530000  12.725000 ;
      RECT 115.360000  14.210000 115.530000  16.920000 ;
      RECT 115.360000  51.740000 115.890000  51.910000 ;
      RECT 115.360000  53.770000 115.890000  54.055000 ;
      RECT 115.390000   7.180000 116.060000   7.260000 ;
      RECT 115.390000  42.475000 118.050000  42.645000 ;
      RECT 115.390000  42.645000 115.560000  43.405000 ;
      RECT 115.400000  37.045000 117.430000  37.505000 ;
      RECT 115.425000  49.015000 115.955000  49.785000 ;
      RECT 115.440000  50.875000 115.890000  51.740000 ;
      RECT 115.440000  52.775000 115.890000  53.770000 ;
      RECT 115.475000   3.275000 116.005000   3.295000 ;
      RECT 115.515000  13.350000 116.185000  13.520000 ;
      RECT 115.610000  41.360000 116.140000  41.530000 ;
      RECT 115.655000   5.660000 115.825000   6.670000 ;
      RECT 115.655000   6.670000 115.830000   6.840000 ;
      RECT 115.655000   6.840000 116.400000   7.010000 ;
      RECT 115.665000  74.595000 115.835000  77.475000 ;
      RECT 115.695000  68.255000 115.865000  73.625000 ;
      RECT 115.700000  56.265000 116.230000  56.435000 ;
      RECT 115.705000  51.910000 115.890000  52.775000 ;
      RECT 115.730000  43.095000 116.260000  43.265000 ;
      RECT 115.730000  43.265000 115.900000  49.015000 ;
      RECT 115.740000  57.325000 115.910000  60.405000 ;
      RECT 115.770000   7.750000 115.940000   8.760000 ;
      RECT 115.785000  61.675000 115.955000  63.855000 ;
      RECT 115.785000  64.405000 115.955000  67.115000 ;
      RECT 115.790000  41.530000 115.960000  42.305000 ;
      RECT 115.800000 113.910000 118.800000 164.900000 ;
      RECT 115.985000  84.275000 116.155000  87.055000 ;
      RECT 116.055000  38.180000 116.315000  41.160000 ;
      RECT 116.055000  61.175000 116.565000  61.505000 ;
      RECT 116.055000  67.585000 116.565000  67.590000 ;
      RECT 116.055000  67.590000 117.445000  67.920000 ;
      RECT 116.060000  50.845000 116.230000  53.370000 ;
      RECT 116.060000  53.370000 116.590000  53.540000 ;
      RECT 116.060000  53.540000 116.230000  56.265000 ;
      RECT 116.070000  44.180000 117.890000  44.350000 ;
      RECT 116.070000  44.350000 116.260000  47.370000 ;
      RECT 116.070000  47.370000 116.600000  48.550000 ;
      RECT 116.070000  48.550000 118.960000  48.720000 ;
      RECT 116.115000   5.660000 116.285000   6.670000 ;
      RECT 116.125000  61.505000 116.495000  64.025000 ;
      RECT 116.125000  64.235000 116.495000  67.585000 ;
      RECT 116.175000   4.505000 116.380000   4.970000 ;
      RECT 116.175000   4.970000 116.345000   5.175000 ;
      RECT 116.185000  77.080000 116.715000  77.250000 ;
      RECT 116.210000   4.440000 116.380000   4.505000 ;
      RECT 116.210000   9.270000 120.800000   9.645000 ;
      RECT 116.215000  49.090000 116.885000  50.625000 ;
      RECT 116.230000   7.010000 116.400000   8.760000 ;
      RECT 116.230000  19.870000 116.400000  22.580000 ;
      RECT 116.230000  23.850000 116.400000  26.560000 ;
      RECT 116.240000  11.370000 116.410000  12.730000 ;
      RECT 116.240000  14.210000 116.410000  16.920000 ;
      RECT 116.260000 200.085000 116.930000 200.255000 ;
      RECT 116.260000 216.235000 116.930000 216.405000 ;
      RECT 116.420000  55.785000 116.750000  55.895000 ;
      RECT 116.420000  55.895000 116.950000  56.065000 ;
      RECT 116.420000  56.065000 116.750000  56.295000 ;
      RECT 116.430000  42.840000 116.600000  44.010000 ;
      RECT 116.430000  44.580000 116.600000  45.280000 ;
      RECT 116.430000  45.280000 116.960000  45.450000 ;
      RECT 116.430000  45.450000 116.600000  47.080000 ;
      RECT 116.430000  53.995000 116.760000  54.325000 ;
      RECT 116.465000  13.350000 117.475000  13.520000 ;
      RECT 116.465000  13.520000 116.745000  13.720000 ;
      RECT 116.465000  83.610000 116.635000  86.760000 ;
      RECT 116.515000  38.180000 116.775000  41.160000 ;
      RECT 116.545000  74.765000 116.715000  77.080000 ;
      RECT 116.545000  77.250000 116.715000  77.475000 ;
      RECT 116.635000   3.760000 116.805000   6.470000 ;
      RECT 116.665000  61.800000 116.835000  67.420000 ;
      RECT 116.690000   3.040000 117.360000   3.210000 ;
      RECT 116.700000  42.470000 118.050000  42.475000 ;
      RECT 116.750000   6.810000 118.760000   6.980000 ;
      RECT 116.750000   6.980000 116.920000   8.160000 ;
      RECT 116.750000   8.840000 120.800000   9.270000 ;
      RECT 116.860000  42.840000 117.030000  44.180000 ;
      RECT 116.910000  46.335000 117.440000  47.370000 ;
      RECT 116.910000  47.370000 117.780000  48.380000 ;
      RECT 116.935000  61.175000 117.445000  61.505000 ;
      RECT 116.935000  67.585000 117.445000  67.590000 ;
      RECT 116.940000  50.845000 117.110000  55.525000 ;
      RECT 116.945000  83.690000 119.995000  83.730000 ;
      RECT 116.945000  83.730000 120.235000  83.900000 ;
      RECT 116.945000  83.900000 117.115000  86.780000 ;
      RECT 116.950000  58.725000 117.840000  59.255000 ;
      RECT 116.975000   3.210000 117.245000   5.115000 ;
      RECT 116.990000  56.755000 117.840000  58.725000 ;
      RECT 116.990000  59.255000 117.840000  60.485000 ;
      RECT 117.005000  61.505000 117.375000  67.585000 ;
      RECT 117.120000  11.720000 117.290000  12.900000 ;
      RECT 117.120000  12.900000 119.050000  13.180000 ;
      RECT 117.120000  13.760000 117.925000  14.040000 ;
      RECT 117.120000  14.040000 117.650000  14.160000 ;
      RECT 117.120000  14.160000 117.290000  16.920000 ;
      RECT 117.120000  72.545000 117.835000  78.155000 ;
      RECT 117.120000  78.570000 117.835000  82.850000 ;
      RECT 117.165000  49.085000 117.835000  50.625000 ;
      RECT 117.165000  55.785000 117.495000  56.265000 ;
      RECT 117.165000  56.265000 117.695000  56.435000 ;
      RECT 117.180000 199.685000 117.710000 200.255000 ;
      RECT 117.210000   7.150000 117.380000   8.840000 ;
      RECT 117.235000  83.090000 120.625000  83.510000 ;
      RECT 117.240000  87.005000 119.955000  87.170000 ;
      RECT 117.240000  87.170000 119.930000  87.175000 ;
      RECT 117.245000  87.000000 119.955000  87.005000 ;
      RECT 117.280000  50.625000 117.650000  55.420000 ;
      RECT 117.290000  42.840000 117.460000  44.010000 ;
      RECT 117.360000 200.495000 117.890000 215.995000 ;
      RECT 117.415000   3.410000 118.690000   4.080000 ;
      RECT 117.415000   4.080000 117.995000   6.470000 ;
      RECT 117.415000   6.470000 118.955000   6.640000 ;
      RECT 117.485000  38.010000 117.655000  41.360000 ;
      RECT 117.485000  41.360000 118.015000  41.530000 ;
      RECT 117.510000  19.870000 117.680000  22.580000 ;
      RECT 117.510000  23.850000 117.680000  26.560000 ;
      RECT 117.545000  61.675000 117.715000  62.740000 ;
      RECT 117.545000  62.910000 117.715000  63.285000 ;
      RECT 117.545000  63.905000 117.715000  64.235000 ;
      RECT 117.545000  64.405000 117.715000  67.115000 ;
      RECT 117.555000  84.970000 118.085000  85.140000 ;
      RECT 117.610000  44.580000 117.780000  45.760000 ;
      RECT 117.610000  45.760000 120.140000  45.930000 ;
      RECT 117.610000  45.930000 117.780000  47.080000 ;
      RECT 117.645000  13.180000 117.925000  13.760000 ;
      RECT 117.670000   6.980000 117.840000   8.160000 ;
      RECT 117.670000  55.895000 118.200000  56.065000 ;
      RECT 117.720000  42.840000 117.890000  44.180000 ;
      RECT 117.725000  84.070000 117.895000  84.970000 ;
      RECT 117.725000  85.140000 117.895000  86.780000 ;
      RECT 117.815000  61.175000 118.325000  61.505000 ;
      RECT 117.815000  67.585000 118.325000  67.915000 ;
      RECT 117.820000  50.845000 118.655000  54.705000 ;
      RECT 117.820000  54.705000 117.990000  55.895000 ;
      RECT 117.885000  61.505000 118.255000  67.585000 ;
      RECT 117.975000  68.490000 118.145000  72.305000 ;
      RECT 118.000000  11.720000 118.170000  12.730000 ;
      RECT 118.000000  14.210000 118.170000  16.920000 ;
      RECT 118.035000 102.920000 166.055000 103.770000 ;
      RECT 118.035000 103.770000 121.145000 108.380000 ;
      RECT 118.035000 108.380000 166.055000 108.735000 ;
      RECT 118.065000  37.870000 118.235000  40.870000 ;
      RECT 118.130000   7.150000 118.300000   8.840000 ;
      RECT 118.130000  46.165000 118.460000  47.015000 ;
      RECT 118.150000  42.840000 118.320000  44.010000 ;
      RECT 118.210000  47.015000 118.380000  47.625000 ;
      RECT 118.235000  72.820000 118.525000  73.325000 ;
      RECT 118.235000  73.325000 118.765000  73.495000 ;
      RECT 118.235000  73.495000 118.525000  77.570000 ;
      RECT 118.235000  78.120000 118.405000  81.770000 ;
      RECT 118.235000  81.770000 118.765000  81.940000 ;
      RECT 118.235000  81.940000 118.405000  82.870000 ;
      RECT 118.285000  45.280000 118.960000  45.450000 ;
      RECT 118.315000  71.960000 118.920000  72.250000 ;
      RECT 118.315000  72.250000 118.525000  72.820000 ;
      RECT 118.320000 200.085000 118.990000 200.255000 ;
      RECT 118.320000 216.235000 118.990000 216.405000 ;
      RECT 118.390000 199.300000 118.920000 200.085000 ;
      RECT 118.405000  42.470000 119.755000  42.640000 ;
      RECT 118.405000  42.640000 119.655000  42.670000 ;
      RECT 118.425000  61.675000 118.595000  67.415000 ;
      RECT 118.450000  55.085000 120.980000  55.285000 ;
      RECT 118.450000  55.285000 118.620000  60.365000 ;
      RECT 118.485000  49.955000 118.655000  50.845000 ;
      RECT 118.505000  83.900000 118.675000  86.780000 ;
      RECT 118.570000   4.600000 143.990000   4.770000 ;
      RECT 118.570000   4.770000 118.740000   6.040000 ;
      RECT 118.580000  13.900000 118.750000  17.270000 ;
      RECT 118.580000  42.840000 118.750000  44.180000 ;
      RECT 118.580000  44.180000 120.140000  44.350000 ;
      RECT 118.590000   6.980000 118.760000   8.160000 ;
      RECT 118.630000  68.950000 118.920000  69.905000 ;
      RECT 118.630000  69.905000 119.200000  70.075000 ;
      RECT 118.630000  70.075000 118.920000  71.960000 ;
      RECT 118.695000  61.175000 119.205000  61.505000 ;
      RECT 118.695000  67.585000 119.205000  67.915000 ;
      RECT 118.715000  60.535000 122.445000  60.855000 ;
      RECT 118.720000  49.595000 120.750000  49.765000 ;
      RECT 118.765000  61.505000 119.135000  67.585000 ;
      RECT 118.790000  19.870000 118.960000  22.580000 ;
      RECT 118.790000  23.850000 118.960000  26.560000 ;
      RECT 118.790000  44.580000 118.960000  45.280000 ;
      RECT 118.790000  45.450000 118.960000  45.590000 ;
      RECT 118.790000  46.100000 118.960000  48.550000 ;
      RECT 118.880000  11.720000 119.050000  12.900000 ;
      RECT 118.910000   3.200000 124.100000   3.370000 ;
      RECT 118.910000   3.660000 123.760000   3.830000 ;
      RECT 118.910000   4.120000 124.100000   4.290000 ;
      RECT 118.965000  68.230000 121.680000  68.555000 ;
      RECT 119.010000  42.840000 119.180000  44.010000 ;
      RECT 119.045000  28.555000 168.425000  29.190000 ;
      RECT 119.045000  29.190000 160.450000  29.405000 ;
      RECT 119.050000   5.020000 119.220000   6.280000 ;
      RECT 119.050000   7.150000 119.220000   8.840000 ;
      RECT 119.115000  72.820000 119.285000  77.570000 ;
      RECT 119.115000  78.120000 119.285000  82.870000 ;
      RECT 119.115000  85.340000 119.645000  85.510000 ;
      RECT 119.120000  72.140000 120.810000  72.310000 ;
      RECT 119.265000  49.955000 119.435000  55.085000 ;
      RECT 119.280000  70.305000 119.810000  70.475000 ;
      RECT 119.285000  84.070000 119.455000  85.340000 ;
      RECT 119.285000  85.510000 119.455000  86.780000 ;
      RECT 119.305000  61.675000 119.475000  62.725000 ;
      RECT 119.305000  62.955000 120.870000  63.285000 ;
      RECT 119.305000  63.905000 120.870000  64.235000 ;
      RECT 119.305000  64.235000 120.285000  67.115000 ;
      RECT 119.410000  37.765000 119.580000  40.845000 ;
      RECT 119.420000 200.495000 119.950000 215.995000 ;
      RECT 119.440000  42.840000 119.610000  44.180000 ;
      RECT 119.450000  68.950000 119.620000  70.305000 ;
      RECT 119.450000  70.475000 119.620000  71.660000 ;
      RECT 119.455000  72.310000 119.825000  73.155000 ;
      RECT 119.610000  46.335000 120.140000  46.505000 ;
      RECT 119.630000  55.455000 119.800000  60.365000 ;
      RECT 119.735000  41.265000 120.700000  41.435000 ;
      RECT 119.735000  41.435000 120.045000  42.130000 ;
      RECT 119.735000  42.130000 120.265000  42.300000 ;
      RECT 119.750000  53.370000 120.280000  53.540000 ;
      RECT 119.780000  48.990000 120.310000  49.595000 ;
      RECT 119.805000  73.325000 120.335000  73.495000 ;
      RECT 119.805000  81.770000 120.335000  81.940000 ;
      RECT 119.870000  42.840000 120.040000  44.010000 ;
      RECT 119.875000  38.155000 120.160000  40.865000 ;
      RECT 119.875000  40.865000 120.045000  41.095000 ;
      RECT 119.970000  44.350000 120.140000  45.760000 ;
      RECT 119.970000  46.100000 120.140000  46.335000 ;
      RECT 119.970000  46.505000 120.140000  48.380000 ;
      RECT 119.995000  72.820000 120.165000  73.325000 ;
      RECT 119.995000  73.495000 120.165000  77.570000 ;
      RECT 119.995000  78.120000 120.165000  81.770000 ;
      RECT 119.995000  81.940000 120.165000  82.870000 ;
      RECT 120.030000  49.955000 120.200000  53.370000 ;
      RECT 120.030000  53.540000 120.200000  54.705000 ;
      RECT 120.045000  11.600000 120.215000  13.420000 ;
      RECT 120.045000  14.330000 120.215000  17.040000 ;
      RECT 120.055000  69.905000 120.585000  70.075000 ;
      RECT 120.065000  83.900000 120.235000  86.780000 ;
      RECT 120.070000  19.870000 120.240000  22.580000 ;
      RECT 120.070000  23.850000 120.240000  26.560000 ;
      RECT 120.115000  61.675000 120.285000  62.955000 ;
      RECT 120.115000  67.115000 120.285000  67.415000 ;
      RECT 120.150000   7.380000 120.680000   7.550000 ;
      RECT 120.205000 113.195000 120.875000 113.525000 ;
      RECT 120.215000  37.335000 122.470000  37.505000 ;
      RECT 120.215000  41.085000 120.885000  41.255000 ;
      RECT 120.215000  41.255000 120.700000  41.265000 ;
      RECT 120.215000  41.760000 120.745000  41.930000 ;
      RECT 120.230000  68.950000 120.400000  69.905000 ;
      RECT 120.230000  70.075000 120.400000  71.660000 ;
      RECT 120.305000  17.700000 120.835000  17.870000 ;
      RECT 120.310000 113.910000 123.310000 164.900000 ;
      RECT 120.315000  11.100000 120.825000  11.430000 ;
      RECT 120.315000  17.510000 120.825000  17.700000 ;
      RECT 120.330000   5.020000 120.500000   7.380000 ;
      RECT 120.330000   7.550000 120.500000   8.160000 ;
      RECT 120.330000  37.505000 122.470000  37.595000 ;
      RECT 120.330000  37.595000 120.700000  41.085000 ;
      RECT 120.330000  43.110000 120.860000  48.390000 ;
      RECT 120.335000  72.310000 120.705000  73.155000 ;
      RECT 120.355000  30.285000 120.525000  31.795000 ;
      RECT 120.355000  32.515000 120.525000  36.025000 ;
      RECT 120.380000 200.085000 121.050000 200.255000 ;
      RECT 120.380000 216.235000 121.050000 216.405000 ;
      RECT 120.385000  11.430000 120.755000  17.510000 ;
      RECT 120.435000  41.930000 120.745000  43.110000 ;
      RECT 120.615000  84.070000 120.785000  85.340000 ;
      RECT 120.615000  85.340000 121.145000  85.510000 ;
      RECT 120.615000  85.510000 120.785000  86.780000 ;
      RECT 120.670000   6.510000 122.700000   6.680000 ;
      RECT 120.700000  61.675000 120.870000  62.725000 ;
      RECT 120.700000  64.405000 120.870000  67.420000 ;
      RECT 120.810000  49.955000 121.600000  54.705000 ;
      RECT 120.810000  55.285000 120.980000  60.365000 ;
      RECT 120.830000  87.000000 121.840000  87.170000 ;
      RECT 120.840000  70.675000 121.370000  70.845000 ;
      RECT 120.870000  37.765000 121.040000  40.865000 ;
      RECT 120.875000  72.820000 121.045000  77.570000 ;
      RECT 120.875000  78.120000 121.045000  82.870000 ;
      RECT 120.915000  41.445000 121.380000  41.615000 ;
      RECT 120.915000  41.615000 121.085000  42.520000 ;
      RECT 120.915000  42.520000 121.200000  42.690000 ;
      RECT 120.925000  11.725000 121.095000  17.345000 ;
      RECT 121.010000  68.950000 121.180000  70.675000 ;
      RECT 121.010000  70.845000 121.180000  71.660000 ;
      RECT 121.020000  86.580000 121.670000  87.000000 ;
      RECT 121.030000  42.690000 121.200000  43.615000 ;
      RECT 121.040000  61.175000 121.550000  61.505000 ;
      RECT 121.040000  67.585000 122.430000  67.915000 ;
      RECT 121.050000  30.285000 121.220000  31.335000 ;
      RECT 121.050000  31.565000 121.220000  31.895000 ;
      RECT 121.050000  32.515000 121.220000  32.845000 ;
      RECT 121.050000  33.015000 121.220000  36.030000 ;
      RECT 121.100000  72.140000 121.770000  72.310000 ;
      RECT 121.100000  83.090000 121.770000  83.490000 ;
      RECT 121.110000  61.505000 121.480000  66.745000 ;
      RECT 121.110000  66.745000 121.640000  66.915000 ;
      RECT 121.110000  66.915000 121.480000  67.585000 ;
      RECT 121.140000  84.570000 121.670000  84.740000 ;
      RECT 121.185000  17.700000 121.715000  17.870000 ;
      RECT 121.195000  11.100000 121.705000  11.430000 ;
      RECT 121.195000  17.510000 121.705000  17.700000 ;
      RECT 121.210000  40.395000 121.920000  40.865000 ;
      RECT 121.210000  40.865000 121.380000  41.445000 ;
      RECT 121.215000  72.310000 121.585000  73.155000 ;
      RECT 121.235000 182.730000 139.290000 185.070000 ;
      RECT 121.235000 185.070000 122.525000 187.295000 ;
      RECT 121.235000 187.295000 139.290000 189.635000 ;
      RECT 121.235000 189.635000 121.920000 190.805000 ;
      RECT 121.255000  41.785000 121.875000  42.115000 ;
      RECT 121.265000  11.430000 121.635000  17.510000 ;
      RECT 121.315000  84.740000 121.670000  86.580000 ;
      RECT 121.350000  19.870000 121.520000  22.580000 ;
      RECT 121.350000  23.850000 121.520000  26.560000 ;
      RECT 121.385000  36.265000 121.915000  36.435000 ;
      RECT 121.390000  29.785000 121.900000  30.115000 ;
      RECT 121.390000  36.195000 121.900000  36.265000 ;
      RECT 121.390000  36.435000 121.900000  36.525000 ;
      RECT 121.395000  73.325000 121.925000  73.495000 ;
      RECT 121.395000  81.770000 121.925000  81.940000 ;
      RECT 121.405000  88.075000 124.800000  88.360000 ;
      RECT 121.405000  88.360000 122.110000  89.285000 ;
      RECT 121.430000  54.705000 121.600000  60.365000 ;
      RECT 121.440000  69.905000 121.970000  70.075000 ;
      RECT 121.460000  30.115000 121.830000  36.195000 ;
      RECT 121.480000  48.350000 124.850000  48.520000 ;
      RECT 121.480000 200.495000 122.010000 215.995000 ;
      RECT 121.520000  45.290000 121.690000  48.000000 ;
      RECT 121.550000  41.360000 122.470000  41.530000 ;
      RECT 121.550000  41.530000 121.875000  41.785000 ;
      RECT 121.610000   5.020000 121.780000   6.280000 ;
      RECT 121.610000   7.080000 121.780000   9.790000 ;
      RECT 121.640000  48.215000 124.690000  48.350000 ;
      RECT 121.650000  61.675000 121.820000  66.145000 ;
      RECT 121.750000  38.155000 121.920000  40.395000 ;
      RECT 121.755000  72.820000 121.925000  73.325000 ;
      RECT 121.755000  73.495000 121.925000  77.570000 ;
      RECT 121.755000  78.120000 121.925000  81.770000 ;
      RECT 121.755000  81.940000 121.925000  82.870000 ;
      RECT 121.770000  49.595000 122.440000  60.535000 ;
      RECT 121.790000  68.950000 121.960000  69.905000 ;
      RECT 121.790000  70.075000 121.960000  71.660000 ;
      RECT 121.805000  11.600000 121.975000  13.210000 ;
      RECT 121.805000  13.830000 121.975000  14.160000 ;
      RECT 121.805000  14.330000 121.975000  17.040000 ;
      RECT 121.895000  84.070000 122.065000  86.780000 ;
      RECT 121.910000  42.605000 122.080000  44.400000 ;
      RECT 121.910000 104.530000 139.430000 104.700000 ;
      RECT 121.910000 104.700000 122.080000 107.090000 ;
      RECT 121.910000 107.090000 139.430000 107.620000 ;
      RECT 121.920000  61.175000 122.430000  61.505000 ;
      RECT 121.925000  45.030000 122.470000  45.200000 ;
      RECT 121.990000  61.505000 122.360000  67.585000 ;
      RECT 122.000000  30.285000 122.170000  34.755000 ;
      RECT 122.005000  10.390000 122.615000  10.560000 ;
      RECT 122.015000  44.570000 123.025000  44.740000 ;
      RECT 122.015000  44.740000 122.545000  44.800000 ;
      RECT 122.075000  11.100000 122.585000  11.430000 ;
      RECT 122.075000  17.510000 122.585000  17.840000 ;
      RECT 122.090000  37.595000 122.470000  38.615000 ;
      RECT 122.090000 190.115000 122.600000 190.145000 ;
      RECT 122.090000 190.145000 124.650000 190.415000 ;
      RECT 122.090000 190.415000 122.600000 190.445000 ;
      RECT 122.090000 190.895000 122.600000 190.925000 ;
      RECT 122.090000 190.925000 126.800000 191.195000 ;
      RECT 122.090000 191.195000 122.600000 191.225000 ;
      RECT 122.105000  10.260000 122.615000  10.390000 ;
      RECT 122.105000  10.560000 122.615000  10.590000 ;
      RECT 122.120000  87.000000 123.130000  87.170000 ;
      RECT 122.130000  42.000000 122.800000  42.170000 ;
      RECT 122.130000  70.675000 122.660000  70.845000 ;
      RECT 122.130000  72.550000 122.695000  75.510000 ;
      RECT 122.130000  75.510000 122.795000  82.880000 ;
      RECT 122.145000  11.430000 122.515000  17.510000 ;
      RECT 122.200000  42.170000 122.730000  42.300000 ;
      RECT 122.270000  29.575000 122.800000  29.745000 ;
      RECT 122.270000  29.745000 122.780000  30.115000 ;
      RECT 122.270000  36.195000 122.780000  36.525000 ;
      RECT 122.300000  40.195000 122.470000  41.360000 ;
      RECT 122.300000  45.000000 122.470000  45.030000 ;
      RECT 122.300000  45.200000 122.470000  48.000000 ;
      RECT 122.305000  85.340000 122.955000  87.000000 ;
      RECT 122.320000 105.400000 122.490000 106.360000 ;
      RECT 122.320000 106.360000 122.850000 106.530000 ;
      RECT 122.320000 106.530000 122.490000 106.750000 ;
      RECT 122.340000  30.115000 122.710000  32.075000 ;
      RECT 122.340000  32.075000 122.930000  32.245000 ;
      RECT 122.340000  32.245000 122.710000  36.195000 ;
      RECT 122.340000  68.620000 122.510000  70.675000 ;
      RECT 122.340000  70.845000 122.510000  71.330000 ;
      RECT 122.400000  38.970000 123.930000  39.720000 ;
      RECT 122.420000 105.040000 138.910000 105.210000 ;
      RECT 122.430000  42.505000 122.960000  42.675000 ;
      RECT 122.440000 200.085000 123.110000 200.255000 ;
      RECT 122.440000 216.235000 123.110000 216.405000 ;
      RECT 122.555000  68.230000 124.855000  68.400000 ;
      RECT 122.600000  61.675000 122.770000  62.725000 ;
      RECT 122.600000  62.955000 122.770000  63.285000 ;
      RECT 122.600000  63.905000 122.770000  64.235000 ;
      RECT 122.600000  64.405000 122.770000  67.115000 ;
      RECT 122.610000  49.985000 122.780000  60.365000 ;
      RECT 122.630000  19.870000 122.800000  22.580000 ;
      RECT 122.630000  23.850000 122.800000  26.560000 ;
      RECT 122.640000  37.765000 123.690000  38.970000 ;
      RECT 122.640000  39.720000 123.690000  40.865000 ;
      RECT 122.685000  11.600000 122.925000  12.610000 ;
      RECT 122.685000  12.610000 122.855000  17.345000 ;
      RECT 122.710000   6.880000 123.240000   7.050000 ;
      RECT 122.720000  18.210000 127.210000  18.265000 ;
      RECT 122.755000  11.260000 123.285000  11.430000 ;
      RECT 122.755000  11.430000 122.925000  11.600000 ;
      RECT 122.765000 113.195000 123.435000 113.525000 ;
      RECT 122.790000  42.675000 122.960000  43.615000 ;
      RECT 122.815000  84.970000 123.345000  85.140000 ;
      RECT 122.820000 189.805000 137.770000 189.975000 ;
      RECT 122.820000 190.585000 137.770000 190.755000 ;
      RECT 122.820000 191.365000 137.770000 191.535000 ;
      RECT 122.840000  88.610000 123.635000  89.690000 ;
      RECT 122.840000  89.690000 133.305000  89.870000 ;
      RECT 122.840000  89.870000 143.765000  90.110000 ;
      RECT 122.840000  90.110000 123.885000  90.460000 ;
      RECT 122.870000  61.175000 123.380000  61.505000 ;
      RECT 122.870000  67.585000 123.380000  67.915000 ;
      RECT 122.890000   5.020000 123.060000   6.880000 ;
      RECT 122.890000   7.050000 123.060000   9.790000 ;
      RECT 122.900000  71.415000 124.740000  72.490000 ;
      RECT 122.900000  72.490000 124.795000  74.940000 ;
      RECT 122.910000 180.765000 137.860000 180.935000 ;
      RECT 122.910000 181.545000 137.860000 181.715000 ;
      RECT 122.910000 182.325000 137.860000 182.495000 ;
      RECT 122.910000 185.395000 137.860000 185.565000 ;
      RECT 122.910000 186.175000 137.860000 186.345000 ;
      RECT 122.910000 186.955000 137.860000 187.125000 ;
      RECT 122.940000  61.505000 123.310000  67.585000 ;
      RECT 122.950000  30.285000 123.120000  31.335000 ;
      RECT 122.950000  31.565000 123.120000  31.895000 ;
      RECT 122.950000  32.515000 123.120000  32.845000 ;
      RECT 122.950000  33.015000 123.120000  35.725000 ;
      RECT 122.950000 105.210000 127.700000 105.280000 ;
      RECT 122.950000 105.990000 127.700000 106.160000 ;
      RECT 122.950000 106.870000 127.770000 106.920000 ;
      RECT 122.950000 106.920000 138.910000 107.065000 ;
      RECT 122.950000 107.065000 139.430000 107.090000 ;
      RECT 122.960000  49.985000 123.400000  60.365000 ;
      RECT 123.080000  45.290000 123.250000  48.000000 ;
      RECT 123.175000  84.070000 123.345000  84.970000 ;
      RECT 123.175000  85.140000 123.345000  86.780000 ;
      RECT 123.235000  11.600000 123.405000  17.345000 ;
      RECT 123.260000   6.510000 123.790000   6.680000 ;
      RECT 123.305000  44.570000 124.315000  44.740000 ;
      RECT 123.370000  42.505000 123.900000  42.675000 ;
      RECT 123.370000  42.675000 123.540000  43.615000 ;
      RECT 123.410000  49.045000 124.080000  49.765000 ;
      RECT 123.410000  60.555000 124.080000  60.615000 ;
      RECT 123.410000  60.615000 125.470000  60.785000 ;
      RECT 123.440000   5.020000 123.610000   6.510000 ;
      RECT 123.440000   6.680000 123.610000   9.790000 ;
      RECT 123.480000  61.675000 123.650000  67.415000 ;
      RECT 123.505000  11.100000 124.015000  11.430000 ;
      RECT 123.505000  17.510000 124.015000  17.840000 ;
      RECT 123.515000  86.580000 124.045000  86.750000 ;
      RECT 123.530000  42.000000 124.200000  42.170000 ;
      RECT 123.540000 200.495000 124.070000 215.995000 ;
      RECT 123.570000  30.285000 123.740000  31.335000 ;
      RECT 123.570000  31.565000 123.740000  31.895000 ;
      RECT 123.570000  32.515000 123.740000  32.845000 ;
      RECT 123.570000  33.015000 123.740000  36.030000 ;
      RECT 123.575000  11.430000 123.945000  17.510000 ;
      RECT 123.600000  42.170000 124.130000  42.300000 ;
      RECT 123.620000  68.620000 123.790000  71.415000 ;
      RECT 123.660000  49.985000 123.830000  54.895000 ;
      RECT 123.660000  55.455000 123.830000  60.365000 ;
      RECT 123.725000  85.770000 123.895000  86.580000 ;
      RECT 123.725000  86.750000 123.895000  86.780000 ;
      RECT 123.750000  61.175000 124.260000  61.505000 ;
      RECT 123.750000  67.585000 124.260000  67.915000 ;
      RECT 123.785000  44.740000 124.315000  44.800000 ;
      RECT 123.820000  61.505000 124.190000  67.585000 ;
      RECT 123.860000  37.335000 126.115000  37.505000 ;
      RECT 123.860000  37.505000 126.000000  37.595000 ;
      RECT 123.860000  37.595000 124.240000  38.615000 ;
      RECT 123.860000  40.195000 124.030000  41.360000 ;
      RECT 123.860000  41.360000 124.780000  41.530000 ;
      RECT 123.860000  45.000000 124.030000  45.030000 ;
      RECT 123.860000  45.030000 124.405000  45.200000 ;
      RECT 123.860000  45.200000 124.030000  48.000000 ;
      RECT 123.865000  10.260000 124.375000  10.390000 ;
      RECT 123.865000  10.390000 124.395000  10.560000 ;
      RECT 123.865000  10.560000 124.375000  10.590000 ;
      RECT 123.875000 223.695000 124.725000 225.350000 ;
      RECT 123.875000 229.255000 124.725000 232.355000 ;
      RECT 123.875000 240.705000 124.725000 243.640000 ;
      RECT 123.895000  89.285000 143.690000  89.455000 ;
      RECT 123.910000  19.870000 124.080000  22.580000 ;
      RECT 123.910000  23.850000 124.080000  26.560000 ;
      RECT 123.910000  29.785000 124.420000  30.115000 ;
      RECT 123.910000  36.195000 124.420000  36.525000 ;
      RECT 123.930000   3.370000 124.100000   3.660000 ;
      RECT 123.930000   3.660000 129.130000   3.830000 ;
      RECT 123.930000   3.830000 124.100000   4.120000 ;
      RECT 123.960000  68.400000 124.370000  70.675000 ;
      RECT 123.960000  70.675000 124.550000  70.845000 ;
      RECT 123.975000  35.110000 124.505000  35.280000 ;
      RECT 123.980000  30.115000 124.350000  35.110000 ;
      RECT 123.980000  35.280000 124.350000  36.195000 ;
      RECT 124.070000  87.005000 127.840000  87.175000 ;
      RECT 124.090000  49.985000 131.700000  50.345000 ;
      RECT 124.090000  50.345000 126.655000  50.995000 ;
      RECT 124.090000  50.995000 124.840000  60.365000 ;
      RECT 124.110000  87.000000 127.840000  87.005000 ;
      RECT 124.115000  11.600000 124.285000  13.210000 ;
      RECT 124.115000  13.830000 124.285000  14.160000 ;
      RECT 124.115000  14.330000 124.285000  17.040000 ;
      RECT 124.135000  88.360000 124.800000  89.285000 ;
      RECT 124.140000   6.510000 125.830000   6.680000 ;
      RECT 124.215000 225.650000 124.385000 226.630000 ;
      RECT 124.215000 234.980000 124.385000 235.960000 ;
      RECT 124.215000 237.100000 124.385000 238.080000 ;
      RECT 124.250000  42.605000 124.420000  44.400000 ;
      RECT 124.360000  61.675000 124.530000  62.725000 ;
      RECT 124.360000  62.955000 124.530000  63.285000 ;
      RECT 124.360000  63.905000 124.530000  64.235000 ;
      RECT 124.360000  64.405000 124.530000  67.115000 ;
      RECT 124.375000  11.260000 124.905000  11.430000 ;
      RECT 124.380000   3.200000 129.470000   3.370000 ;
      RECT 124.380000   4.120000 129.470000   4.290000 ;
      RECT 124.385000  11.100000 124.895000  11.260000 ;
      RECT 124.385000  17.510000 124.895000  17.840000 ;
      RECT 124.410000  38.155000 124.580000  40.395000 ;
      RECT 124.410000  40.395000 125.120000  40.865000 ;
      RECT 124.410000 180.935000 133.710000 181.375000 ;
      RECT 124.410000 181.885000 133.710000 182.325000 ;
      RECT 124.410000 185.565000 133.710000 186.005000 ;
      RECT 124.410000 186.515000 133.710000 186.955000 ;
      RECT 124.455000  11.430000 124.825000  17.510000 ;
      RECT 124.455000  41.530000 124.780000  41.785000 ;
      RECT 124.455000  41.785000 125.075000  42.115000 ;
      RECT 124.490000  23.560000 124.660000  25.570000 ;
      RECT 124.490000  25.570000 130.755000  25.740000 ;
      RECT 124.490000  25.740000 124.675000  26.920000 ;
      RECT 124.500000 200.085000 125.170000 200.255000 ;
      RECT 124.500000 216.235000 125.170000 216.405000 ;
      RECT 124.520000  30.285000 124.690000  34.755000 ;
      RECT 124.540000  70.305000 125.070000  70.475000 ;
      RECT 124.555000  78.130000 124.725000  81.050000 ;
      RECT 124.555000  81.950000 124.725000  84.850000 ;
      RECT 124.630000  61.175000 125.140000  61.505000 ;
      RECT 124.630000  67.585000 125.140000  67.915000 ;
      RECT 124.640000  45.290000 124.810000  48.000000 ;
      RECT 124.670000  49.805000 131.120000  49.985000 ;
      RECT 124.670000  60.365000 124.840000  60.445000 ;
      RECT 124.700000  61.505000 125.070000  67.585000 ;
      RECT 124.720000   5.020000 124.890000   6.280000 ;
      RECT 124.720000   7.080000 124.890000   9.790000 ;
      RECT 124.730000  90.920000 145.515000  91.465000 ;
      RECT 124.790000  29.785000 125.300000  30.115000 ;
      RECT 124.790000  36.195000 125.300000  36.525000 ;
      RECT 124.820000 113.910000 127.820000 164.900000 ;
      RECT 124.840000  81.340000 125.790000  81.490000 ;
      RECT 124.840000  81.490000 125.730000  81.510000 ;
      RECT 124.860000  30.115000 125.230000  32.140000 ;
      RECT 124.860000  32.140000 125.390000  32.310000 ;
      RECT 124.860000  32.310000 125.230000  36.195000 ;
      RECT 124.865000  25.740000 125.245000  25.815000 ;
      RECT 124.900000  68.620000 125.070000  70.305000 ;
      RECT 124.900000  70.475000 125.070000  71.330000 ;
      RECT 124.950000  40.865000 125.120000  41.445000 ;
      RECT 124.950000  41.445000 125.415000  41.615000 ;
      RECT 124.995000  11.725000 125.165000  17.345000 ;
      RECT 125.060000  52.630000 125.590000  52.800000 ;
      RECT 125.070000  19.870000 125.240000  24.620000 ;
      RECT 125.070000  75.570000 125.600000  75.740000 ;
      RECT 125.080000  51.955000 125.470000  52.630000 ;
      RECT 125.080000  52.800000 125.470000  54.985000 ;
      RECT 125.080000  54.985000 125.590000  55.315000 ;
      RECT 125.085000  82.220000 125.255000  84.070000 ;
      RECT 125.085000  84.070000 125.615000  84.240000 ;
      RECT 125.085000  84.240000 125.255000  84.930000 ;
      RECT 125.105000  51.235000 125.775000  51.785000 ;
      RECT 125.120000  81.320000 125.790000  81.340000 ;
      RECT 125.130000  42.520000 125.415000  42.690000 ;
      RECT 125.130000  42.690000 125.300000  43.615000 ;
      RECT 125.145000  78.070000 125.315000  79.055000 ;
      RECT 125.145000  79.055000 125.845000  79.225000 ;
      RECT 125.145000  79.225000 125.315000  80.780000 ;
      RECT 125.155000 224.125000 135.155000 226.460000 ;
      RECT 125.155000 229.425000 135.155000 232.185000 ;
      RECT 125.155000 235.150000 135.155000 237.910000 ;
      RECT 125.155000 240.875000 135.155000 243.210000 ;
      RECT 125.240000  61.675000 125.410000  67.415000 ;
      RECT 125.245000  41.615000 125.415000  42.520000 ;
      RECT 125.265000  11.100000 125.775000  11.430000 ;
      RECT 125.265000  17.510000 125.775000  17.840000 ;
      RECT 125.290000  37.765000 125.460000  40.865000 ;
      RECT 125.300000  55.785000 125.470000  60.615000 ;
      RECT 125.335000  11.430000 125.705000  13.590000 ;
      RECT 125.335000  13.590000 126.595000  13.850000 ;
      RECT 125.335000  13.850000 125.705000  17.510000 ;
      RECT 125.355000  72.250000 125.525000  75.570000 ;
      RECT 125.355000  75.740000 125.525000  77.230000 ;
      RECT 125.435000  77.680000 126.785000  77.850000 ;
      RECT 125.445000  41.085000 126.115000  41.255000 ;
      RECT 125.450000  68.620000 125.620000  68.725000 ;
      RECT 125.450000  68.725000 126.380000  69.905000 ;
      RECT 125.450000  70.120000 125.620000  71.945000 ;
      RECT 125.470000  30.285000 125.640000  31.335000 ;
      RECT 125.470000  31.565000 125.640000  31.895000 ;
      RECT 125.470000  32.515000 125.640000  32.845000 ;
      RECT 125.470000  33.015000 125.640000  35.725000 ;
      RECT 125.470000  43.110000 126.000000  48.390000 ;
      RECT 125.475000  21.220000 126.020000  23.410000 ;
      RECT 125.475000  26.060000 126.005000  27.100000 ;
      RECT 125.490000  21.120000 126.020000  21.220000 ;
      RECT 125.510000  61.175000 126.020000  61.505000 ;
      RECT 125.510000  67.585000 126.020000  67.915000 ;
      RECT 125.575000   8.840000 129.030000   9.010000 ;
      RECT 125.575000   9.010000 125.745000  10.760000 ;
      RECT 125.580000  61.505000 125.950000  67.585000 ;
      RECT 125.585000  41.760000 126.115000  41.930000 ;
      RECT 125.585000  41.930000 125.895000  43.110000 ;
      RECT 125.600000 200.495000 126.130000 215.995000 ;
      RECT 125.630000  37.595000 126.000000  41.085000 ;
      RECT 125.630000  41.255000 126.115000  41.265000 ;
      RECT 125.630000  41.265000 126.595000  41.435000 ;
      RECT 125.640000  59.125000 130.150000  60.315000 ;
      RECT 125.740000  29.785000 128.890000  30.115000 ;
      RECT 125.740000  36.195000 126.250000  36.220000 ;
      RECT 125.740000  36.220000 128.890000  36.525000 ;
      RECT 125.750000  68.230000 129.520000  68.385000 ;
      RECT 125.750000  68.385000 129.560000  68.400000 ;
      RECT 125.760000  51.955000 125.930000  58.495000 ;
      RECT 125.785000  59.115000 129.915000  59.125000 ;
      RECT 125.790000  68.400000 129.560000  68.555000 ;
      RECT 125.810000  30.115000 126.180000  36.195000 ;
      RECT 125.820000   7.365000 126.350000   7.535000 ;
      RECT 125.835000  70.985000 129.560000  71.350000 ;
      RECT 125.835000  71.350000 129.565000  71.520000 ;
      RECT 125.850000  69.905000 126.380000  70.075000 ;
      RECT 125.850000  75.180000 126.180000  75.880000 ;
      RECT 125.850000  75.880000 128.375000  76.050000 ;
      RECT 125.865000  82.200000 126.035000  84.930000 ;
      RECT 125.875000  11.600000 126.115000  13.420000 ;
      RECT 125.875000  14.330000 126.045000  17.040000 ;
      RECT 125.945000  11.260000 126.475000  11.430000 ;
      RECT 125.945000  11.430000 126.115000  11.600000 ;
      RECT 125.985000  51.235000 126.655000  51.405000 ;
      RECT 125.985000  58.715000 127.335000  58.885000 ;
      RECT 126.000000   5.020000 126.170000   7.365000 ;
      RECT 126.000000   7.535000 126.170000   8.160000 ;
      RECT 126.010000  25.130000 129.915000  25.300000 ;
      RECT 126.025000  78.070000 126.195000  80.780000 ;
      RECT 126.060000  27.350000 126.960000  27.520000 ;
      RECT 126.065000  42.130000 126.595000  42.300000 ;
      RECT 126.075000  25.740000 130.720000  25.815000 ;
      RECT 126.100000  51.405000 126.370000  58.715000 ;
      RECT 126.120000  61.675000 126.290000  62.725000 ;
      RECT 126.120000  62.955000 126.290000  63.285000 ;
      RECT 126.120000  63.905000 126.290000  64.235000 ;
      RECT 126.120000  64.405000 126.290000  67.115000 ;
      RECT 126.170000  38.155000 126.455000  40.865000 ;
      RECT 126.190000  44.180000 127.750000  44.350000 ;
      RECT 126.190000  44.350000 126.360000  45.760000 ;
      RECT 126.190000  45.760000 128.720000  45.930000 ;
      RECT 126.190000  46.100000 126.360000  46.335000 ;
      RECT 126.190000  46.335000 126.720000  46.505000 ;
      RECT 126.190000  46.505000 126.360000  48.380000 ;
      RECT 126.270000  85.150000 127.960000  85.320000 ;
      RECT 126.285000  40.865000 126.455000  41.095000 ;
      RECT 126.285000  41.435000 126.595000  42.130000 ;
      RECT 126.290000  42.840000 126.460000  44.010000 ;
      RECT 126.305000  71.775000 126.475000  74.960000 ;
      RECT 126.305000  76.220000 126.475000  77.360000 ;
      RECT 126.350000  19.870000 126.520000  24.620000 ;
      RECT 126.350000  30.285000 126.520000  36.030000 ;
      RECT 126.425000  11.600000 126.595000  13.590000 ;
      RECT 126.425000  13.850000 126.595000  17.345000 ;
      RECT 126.460000  61.175000 126.970000  61.505000 ;
      RECT 126.460000  67.585000 127.850000  67.885000 ;
      RECT 126.460000  67.885000 127.865000  67.915000 ;
      RECT 126.515000  84.070000 127.045000  84.240000 ;
      RECT 126.530000  26.780000 127.185000  27.040000 ;
      RECT 126.530000  61.505000 126.900000  67.585000 ;
      RECT 126.540000  51.765000 126.995000  51.935000 ;
      RECT 126.540000  51.935000 126.710000  58.495000 ;
      RECT 126.560000 200.085000 127.230000 200.255000 ;
      RECT 126.560000 216.235000 127.230000 216.405000 ;
      RECT 126.575000  42.470000 127.925000  42.640000 ;
      RECT 126.620000  36.195000 128.010000  36.220000 ;
      RECT 126.640000  75.160000 127.170000  75.330000 ;
      RECT 126.645000  80.950000 127.955000  81.165000 ;
      RECT 126.645000  81.165000 126.815000  84.070000 ;
      RECT 126.645000  84.240000 126.815000  84.930000 ;
      RECT 126.675000  42.640000 127.925000  42.670000 ;
      RECT 126.690000  30.115000 127.060000  36.195000 ;
      RECT 126.695000  11.100000 127.205000  11.430000 ;
      RECT 126.695000  17.510000 127.205000  17.840000 ;
      RECT 126.715000  79.055000 127.245000  79.225000 ;
      RECT 126.720000  42.840000 126.890000  44.180000 ;
      RECT 126.735000  75.330000 127.065000  75.690000 ;
      RECT 126.750000  37.765000 126.920000  40.845000 ;
      RECT 126.765000  11.430000 127.135000  17.510000 ;
      RECT 126.825000  50.515000 126.995000  51.765000 ;
      RECT 126.880000  52.210000 127.150000  58.715000 ;
      RECT 126.905000  78.070000 127.075000  79.055000 ;
      RECT 126.905000  79.225000 127.075000  80.780000 ;
      RECT 126.970000 189.975000 136.270000 190.415000 ;
      RECT 126.970000 190.925000 136.270000 191.365000 ;
      RECT 127.015000  26.090000 127.185000  26.780000 ;
      RECT 127.015000  27.040000 127.185000  27.100000 ;
      RECT 127.070000  61.675000 127.240000  66.145000 ;
      RECT 127.150000  42.840000 127.320000  44.010000 ;
      RECT 127.165000  50.345000 128.625000  50.995000 ;
      RECT 127.195000  77.680000 128.545000  77.850000 ;
      RECT 127.195000  81.335000 128.545000  81.805000 ;
      RECT 127.195000  81.805000 128.515000  81.940000 ;
      RECT 127.230000  30.285000 127.400000  31.335000 ;
      RECT 127.230000  31.565000 127.400000  31.895000 ;
      RECT 127.230000  32.515000 127.400000  32.845000 ;
      RECT 127.230000  33.015000 127.400000  35.725000 ;
      RECT 127.240000  27.350000 131.680000  27.520000 ;
      RECT 127.255000  76.050000 127.425000  77.230000 ;
      RECT 127.280000   5.020000 127.450000   6.280000 ;
      RECT 127.280000   7.150000 127.450000   8.840000 ;
      RECT 127.305000  11.600000 127.475000  13.210000 ;
      RECT 127.305000  13.830000 127.475000  14.160000 ;
      RECT 127.305000  14.330000 127.475000  17.040000 ;
      RECT 127.320000  51.955000 127.490000  58.495000 ;
      RECT 127.335000  67.915000 127.865000  68.055000 ;
      RECT 127.340000  61.175000 127.850000  61.505000 ;
      RECT 127.370000  44.580000 127.540000  45.280000 ;
      RECT 127.370000  45.280000 128.045000  45.450000 ;
      RECT 127.370000  45.450000 127.540000  45.590000 ;
      RECT 127.370000  46.100000 127.540000  48.550000 ;
      RECT 127.370000  48.550000 130.260000  48.720000 ;
      RECT 127.410000  61.505000 127.780000  67.585000 ;
      RECT 127.425000  82.200000 127.595000  84.930000 ;
      RECT 127.435000  26.315000 127.965000  27.350000 ;
      RECT 127.505000  75.160000 128.035000  75.330000 ;
      RECT 127.565000  17.700000 128.095000  17.870000 ;
      RECT 127.570000  30.115000 127.940000  36.195000 ;
      RECT 127.575000  11.100000 128.085000  11.430000 ;
      RECT 127.575000  17.510000 128.085000  17.700000 ;
      RECT 127.580000  42.840000 127.750000  44.180000 ;
      RECT 127.615000  75.330000 127.945000  75.690000 ;
      RECT 127.630000  19.870000 127.800000  24.620000 ;
      RECT 127.645000  11.430000 128.015000  17.510000 ;
      RECT 127.660000 200.495000 128.190000 215.995000 ;
      RECT 127.785000  78.070000 127.955000  80.950000 ;
      RECT 127.810000  51.665000 127.980000  58.425000 ;
      RECT 127.815000 106.360000 128.345000 106.530000 ;
      RECT 127.845000  74.000000 128.375000  74.170000 ;
      RECT 127.845000  84.070000 128.375000  84.240000 ;
      RECT 127.870000  46.165000 128.200000  47.015000 ;
      RECT 127.895000 105.400000 128.065000 106.360000 ;
      RECT 127.895000 106.530000 128.065000 106.750000 ;
      RECT 127.950000  47.015000 128.120000  47.625000 ;
      RECT 128.005000  85.770000 128.175000  86.780000 ;
      RECT 128.010000  42.840000 128.180000  44.010000 ;
      RECT 128.020000  61.675000 128.740000  62.725000 ;
      RECT 128.020000  62.955000 128.740000  63.285000 ;
      RECT 128.020000  63.905000 128.740000  64.235000 ;
      RECT 128.020000  64.405000 128.190000  67.420000 ;
      RECT 128.095000  37.870000 128.265000  40.870000 ;
      RECT 128.110000  30.285000 128.280000  36.030000 ;
      RECT 128.135000  79.055000 128.835000  79.225000 ;
      RECT 128.185000  11.725000 128.355000  17.345000 ;
      RECT 128.190000 106.870000 133.375000 106.920000 ;
      RECT 128.195000  26.090000 128.365000  26.145000 ;
      RECT 128.195000  26.145000 128.895000  26.405000 ;
      RECT 128.195000  26.405000 128.365000  27.100000 ;
      RECT 128.205000  72.250000 128.375000  74.000000 ;
      RECT 128.205000  74.170000 128.375000  75.880000 ;
      RECT 128.205000  76.220000 128.375000  77.360000 ;
      RECT 128.205000  82.220000 128.375000  84.070000 ;
      RECT 128.205000  84.240000 128.375000  84.930000 ;
      RECT 128.280000  42.470000 129.630000  42.475000 ;
      RECT 128.280000  42.475000 130.940000  42.645000 ;
      RECT 128.290000  87.005000 132.060000  87.175000 ;
      RECT 128.300000  51.955000 128.470000  58.495000 ;
      RECT 128.305000  87.000000 132.035000  87.005000 ;
      RECT 128.315000  41.360000 128.845000  41.530000 ;
      RECT 128.380000  36.195000 128.890000  36.220000 ;
      RECT 128.410000  19.870000 128.580000  24.620000 ;
      RECT 128.430000  18.465000 128.965000  18.635000 ;
      RECT 128.440000  42.840000 128.610000  44.180000 ;
      RECT 128.440000  44.180000 130.260000  44.350000 ;
      RECT 128.450000  30.115000 128.820000  32.140000 ;
      RECT 128.450000  32.140000 129.085000  32.310000 ;
      RECT 128.450000  32.310000 128.820000  36.195000 ;
      RECT 128.455000  11.100000 128.965000  11.430000 ;
      RECT 128.455000  17.510000 128.965000  18.465000 ;
      RECT 128.455000  58.715000 129.805000  58.885000 ;
      RECT 128.525000  11.430000 128.895000  17.510000 ;
      RECT 128.550000  44.580000 128.720000  45.760000 ;
      RECT 128.550000  45.930000 128.720000  47.080000 ;
      RECT 128.550000  47.370000 129.420000  48.380000 ;
      RECT 128.555000 105.210000 133.305000 105.280000 ;
      RECT 128.555000 105.990000 133.305000 106.160000 ;
      RECT 128.560000   5.020000 128.730000   8.160000 ;
      RECT 128.570000  64.405000 128.740000  67.420000 ;
      RECT 128.620000 200.085000 129.290000 200.255000 ;
      RECT 128.620000 216.235000 129.290000 216.405000 ;
      RECT 128.640000  52.210000 128.910000  58.715000 ;
      RECT 128.665000  78.070000 128.835000  79.055000 ;
      RECT 128.665000  79.225000 128.835000  80.780000 ;
      RECT 128.675000  37.840000 132.915000  38.010000 ;
      RECT 128.675000  38.010000 128.845000  41.360000 ;
      RECT 128.695000  81.950000 128.865000  84.850000 ;
      RECT 128.785000  71.775000 128.955000  74.940000 ;
      RECT 128.795000  50.515000 128.965000  51.765000 ;
      RECT 128.795000  51.765000 129.250000  51.935000 ;
      RECT 128.860000   9.010000 129.030000  10.760000 ;
      RECT 128.860000  10.760000 133.975000  10.930000 ;
      RECT 128.870000  42.840000 129.040000  44.010000 ;
      RECT 128.890000  46.335000 129.420000  47.370000 ;
      RECT 128.900000   6.510000 130.930000   6.680000 ;
      RECT 128.900000  37.335000 130.930000  37.505000 ;
      RECT 128.910000  61.175000 129.420000  61.505000 ;
      RECT 128.910000  67.585000 129.420000  67.915000 ;
      RECT 128.980000  61.505000 129.350000  67.585000 ;
      RECT 128.990000  30.285000 129.160000  31.335000 ;
      RECT 128.990000  31.565000 129.160000  31.895000 ;
      RECT 128.990000  32.515000 129.160000  32.845000 ;
      RECT 128.990000  33.015000 129.160000  35.725000 ;
      RECT 128.995000  76.420000 132.395000  76.590000 ;
      RECT 128.995000  76.590000 129.165000  77.155000 ;
      RECT 129.065000  11.600000 129.235000  13.420000 ;
      RECT 129.065000  14.330000 129.235000  17.040000 ;
      RECT 129.080000  51.935000 129.250000  58.495000 ;
      RECT 129.135000  18.040000 130.275000  18.210000 ;
      RECT 129.135000  50.345000 131.700000  50.995000 ;
      RECT 129.135000  51.235000 129.805000  51.405000 ;
      RECT 129.140000  26.780000 129.780000  27.040000 ;
      RECT 129.190000  19.870000 129.360000  24.620000 ;
      RECT 129.225000 113.195000 129.895000 113.525000 ;
      RECT 129.260000  29.785000 129.770000  30.115000 ;
      RECT 129.260000  36.195000 129.770000  36.525000 ;
      RECT 129.300000   3.370000 129.470000   4.120000 ;
      RECT 129.300000  42.840000 129.470000  44.180000 ;
      RECT 129.310000  18.210000 130.200000  18.270000 ;
      RECT 129.310000  78.090000 129.860000  81.090000 ;
      RECT 129.330000  30.115000 129.700000  36.195000 ;
      RECT 129.330000 113.910000 132.330000 164.900000 ;
      RECT 129.370000  45.280000 129.900000  45.450000 ;
      RECT 129.375000  26.090000 129.545000  26.780000 ;
      RECT 129.375000  27.040000 129.545000  27.100000 ;
      RECT 129.385000  81.335000 130.055000  81.570000 ;
      RECT 129.420000  51.405000 129.690000  58.715000 ;
      RECT 129.445000  82.220000 129.615000  83.290000 ;
      RECT 129.445000  83.290000 130.055000  83.460000 ;
      RECT 129.445000  83.460000 129.615000  84.930000 ;
      RECT 129.520000  61.675000 129.690000  66.145000 ;
      RECT 129.555000  38.180000 129.815000  41.160000 ;
      RECT 129.610000  72.450000 131.450000  73.365000 ;
      RECT 129.615000  11.600000 129.785000  13.210000 ;
      RECT 129.615000  13.830000 129.785000  14.160000 ;
      RECT 129.615000  14.330000 129.785000  17.040000 ;
      RECT 129.640000   3.430000 129.810000   4.430000 ;
      RECT 129.685000  77.200000 132.395000  77.370000 ;
      RECT 129.720000 200.495000 130.250000 215.995000 ;
      RECT 129.730000  42.840000 129.900000  44.010000 ;
      RECT 129.730000  44.580000 129.900000  45.280000 ;
      RECT 129.730000  45.450000 129.900000  47.080000 ;
      RECT 129.730000  47.370000 130.260000  48.550000 ;
      RECT 129.730000  68.620000 129.900000  71.130000 ;
      RECT 129.755000  74.760000 129.925000  74.790000 ;
      RECT 129.755000  74.790000 130.345000  74.960000 ;
      RECT 129.755000  74.960000 129.925000  75.770000 ;
      RECT 129.765000  76.370000 132.095000  76.420000 ;
      RECT 129.765000  77.080000 132.095000  77.200000 ;
      RECT 129.790000  61.175000 130.300000  61.505000 ;
      RECT 129.790000  67.585000 130.300000  67.915000 ;
      RECT 129.840000   5.020000 130.010000   6.280000 ;
      RECT 129.840000   7.080000 130.010000   9.790000 ;
      RECT 129.860000  51.955000 130.030000  58.495000 ;
      RECT 129.860000  61.505000 130.230000  67.585000 ;
      RECT 129.865000  85.150000 130.875000  85.320000 ;
      RECT 129.870000  30.285000 130.040000  32.140000 ;
      RECT 129.870000  32.140000 130.400000  32.310000 ;
      RECT 129.870000  32.310000 130.040000  36.030000 ;
      RECT 129.885000  11.100000 130.395000  11.430000 ;
      RECT 129.885000  17.510000 130.395000  17.840000 ;
      RECT 129.955000  11.430000 130.325000  17.510000 ;
      RECT 129.970000  19.870000 130.140000  24.620000 ;
      RECT 129.980000   3.200000 135.070000   3.370000 ;
      RECT 129.980000   3.370000 130.150000   4.120000 ;
      RECT 129.980000   4.120000 135.070000   4.290000 ;
      RECT 130.015000  38.180000 130.275000  41.160000 ;
      RECT 130.015000  51.235000 130.685000  51.785000 ;
      RECT 130.025000  74.000000 134.225000  74.540000 ;
      RECT 130.035000  84.280000 130.565000  84.450000 ;
      RECT 130.070000  43.095000 130.600000  43.265000 ;
      RECT 130.070000  44.350000 130.260000  47.370000 ;
      RECT 130.190000  41.360000 130.720000  41.530000 ;
      RECT 130.200000  52.630000 130.730000  52.800000 ;
      RECT 130.200000  54.985000 130.710000  55.315000 ;
      RECT 130.225000  80.950000 131.390000  81.120000 ;
      RECT 130.225000  81.120000 130.395000  84.280000 ;
      RECT 130.225000  84.450000 130.395000  84.930000 ;
      RECT 130.320000   3.660000 135.070000   3.830000 ;
      RECT 130.320000  26.145000 131.460000  26.405000 ;
      RECT 130.320000  51.955000 130.710000  52.630000 ;
      RECT 130.320000  52.800000 130.710000  54.985000 ;
      RECT 130.320000  55.785000 130.490000  60.615000 ;
      RECT 130.320000  60.615000 132.380000  60.785000 ;
      RECT 130.325000  10.390000 130.855000  10.560000 ;
      RECT 130.335000  10.260000 130.845000  10.390000 ;
      RECT 130.335000  10.560000 130.845000  10.590000 ;
      RECT 130.340000  78.070000 130.510000  80.780000 ;
      RECT 130.370000  41.530000 130.540000  42.305000 ;
      RECT 130.430000  43.265000 130.600000  48.390000 ;
      RECT 130.440000  18.875000 130.970000  19.045000 ;
      RECT 130.470000  61.675000 130.640000  62.740000 ;
      RECT 130.470000  62.910000 130.640000  63.285000 ;
      RECT 130.470000  63.905000 130.640000  64.235000 ;
      RECT 130.470000  64.405000 130.640000  67.115000 ;
      RECT 130.475000  77.680000 131.145000  77.850000 ;
      RECT 130.490000  30.285000 130.660000  31.335000 ;
      RECT 130.490000  33.015000 130.660000  35.725000 ;
      RECT 130.495000  11.600000 130.665000  17.345000 ;
      RECT 130.550000  19.520000 130.720000  20.525000 ;
      RECT 130.550000  24.090000 130.720000  25.130000 ;
      RECT 130.550000  25.130000 130.755000  25.570000 ;
      RECT 130.555000  26.090000 130.725000  26.145000 ;
      RECT 130.555000  26.405000 130.725000  27.100000 ;
      RECT 130.565000  17.515000 131.825000  17.840000 ;
      RECT 130.565000  17.840000 130.970000  18.875000 ;
      RECT 130.600000  68.460000 131.450000  71.440000 ;
      RECT 130.600000  71.440000 131.490000  72.330000 ;
      RECT 130.600000  72.330000 131.450000  72.450000 ;
      RECT 130.665000  75.180000 131.205000  75.350000 ;
      RECT 130.680000  36.195000 134.790000  36.525000 ;
      RECT 130.680000 200.085000 131.350000 200.255000 ;
      RECT 130.680000 216.235000 131.350000 216.405000 ;
      RECT 130.740000  61.175000 131.250000  61.505000 ;
      RECT 130.740000  67.585000 131.250000  67.915000 ;
      RECT 130.765000  29.785000 132.295000  30.115000 ;
      RECT 130.770000  42.645000 130.940000  43.405000 ;
      RECT 130.770000  43.405000 131.420000  44.415000 ;
      RECT 130.810000  61.505000 131.180000  67.585000 ;
      RECT 130.825000  83.290000 131.355000  83.460000 ;
      RECT 130.830000  30.115000 131.200000  36.195000 ;
      RECT 130.890000  41.290000 131.560000  41.460000 ;
      RECT 130.890000  46.335000 131.420000  46.505000 ;
      RECT 130.910000  47.855000 131.080000  48.465000 ;
      RECT 130.910000  48.465000 136.440000  48.635000 ;
      RECT 130.940000   6.880000 131.470000   7.050000 ;
      RECT 130.950000  42.030000 131.480000  42.200000 ;
      RECT 130.950000  50.995000 131.700000  60.365000 ;
      RECT 130.950000  60.365000 131.120000  60.445000 ;
      RECT 130.985000  38.180000 131.155000  41.290000 ;
      RECT 130.985000  41.460000 131.480000  42.030000 ;
      RECT 131.005000  82.220000 131.175000  83.290000 ;
      RECT 131.005000  83.460000 131.175000  84.930000 ;
      RECT 131.035000  74.760000 131.205000  75.180000 ;
      RECT 131.035000  75.350000 131.205000  75.770000 ;
      RECT 131.045000  11.600000 131.215000  13.420000 ;
      RECT 131.045000  14.330000 131.215000  17.040000 ;
      RECT 131.095000  19.745000 131.355000  20.385000 ;
      RECT 131.120000   5.020000 131.290000   6.880000 ;
      RECT 131.120000   7.050000 131.290000   9.790000 ;
      RECT 131.140000  18.945000 131.340000  19.745000 ;
      RECT 131.140000  20.385000 131.310000  21.025000 ;
      RECT 131.140000  37.335000 131.810000  37.505000 ;
      RECT 131.180000  21.610000 131.350000  24.645000 ;
      RECT 131.200000  24.955000 132.130000  25.215000 ;
      RECT 131.200000  25.215000 131.460000  26.145000 ;
      RECT 131.220000  78.070000 131.390000  80.950000 ;
      RECT 131.250000  44.415000 131.420000  46.335000 ;
      RECT 131.250000  46.505000 131.420000  48.085000 ;
      RECT 131.265000  26.780000 131.905000  27.040000 ;
      RECT 131.315000  11.100000 131.825000  11.430000 ;
      RECT 131.315000  17.510000 131.825000  17.515000 ;
      RECT 131.330000  85.150000 132.340000  85.320000 ;
      RECT 131.350000  61.800000 131.520000  67.420000 ;
      RECT 131.370000  30.285000 131.540000  35.725000 ;
      RECT 131.385000  11.430000 131.755000  17.510000 ;
      RECT 131.405000  18.040000 139.275000  18.210000 ;
      RECT 131.465000  81.335000 132.475000  81.505000 ;
      RECT 131.475000  77.680000 132.145000  77.850000 ;
      RECT 131.490000   6.510000 132.020000   6.680000 ;
      RECT 131.525000  19.625000 132.205000  19.795000 ;
      RECT 131.530000  21.225000 132.205000  21.395000 ;
      RECT 131.590000  19.795000 132.205000  21.225000 ;
      RECT 131.590000  45.000000 132.120000  45.170000 ;
      RECT 131.620000  61.175000 132.130000  61.505000 ;
      RECT 131.620000  67.585000 132.130000  67.915000 ;
      RECT 131.650000  41.635000 131.900000  42.305000 ;
      RECT 131.670000   5.020000 131.840000   6.510000 ;
      RECT 131.670000   6.680000 131.840000   9.790000 ;
      RECT 131.685000  41.580000 131.900000  41.635000 ;
      RECT 131.685000  42.305000 131.855000  43.405000 ;
      RECT 131.685000  43.405000 131.880000  44.415000 ;
      RECT 131.690000  61.505000 132.060000  67.585000 ;
      RECT 131.710000  30.115000 132.080000  36.195000 ;
      RECT 131.710000  45.170000 131.880000  48.085000 ;
      RECT 131.710000  49.045000 132.380000  49.765000 ;
      RECT 131.710000  60.555000 132.380000  60.615000 ;
      RECT 131.730000  38.180000 132.035000  40.890000 ;
      RECT 131.730000  40.890000 131.900000  41.580000 ;
      RECT 131.735000  26.090000 131.905000  26.780000 ;
      RECT 131.735000  27.040000 131.905000  27.100000 ;
      RECT 131.780000 200.495000 132.310000 215.995000 ;
      RECT 131.785000  82.140000 131.955000  84.930000 ;
      RECT 131.785000 113.195000 132.455000 113.525000 ;
      RECT 131.890000  81.020000 132.420000  81.190000 ;
      RECT 131.890000  81.190000 132.475000  81.335000 ;
      RECT 131.925000  11.725000 132.095000  17.345000 ;
      RECT 131.960000  49.985000 132.130000  54.895000 ;
      RECT 131.960000  55.455000 132.130000  60.365000 ;
      RECT 131.995000  18.210000 132.885000  18.300000 ;
      RECT 132.050000  42.400000 132.580000  42.570000 ;
      RECT 132.050000  42.570000 132.460000  44.585000 ;
      RECT 132.050000  44.585000 132.590000  44.740000 ;
      RECT 132.050000  45.375000 132.590000  45.665000 ;
      RECT 132.050000  45.665000 132.340000  48.085000 ;
      RECT 132.070000  42.030000 133.100000  42.200000 ;
      RECT 132.090000  37.335000 132.760000  37.505000 ;
      RECT 132.095000   9.215000 132.625000  10.590000 ;
      RECT 132.100000  78.070000 132.270000  80.780000 ;
      RECT 132.125000  83.290000 132.735000  83.460000 ;
      RECT 132.145000  74.790000 132.675000  74.960000 ;
      RECT 132.150000  68.810000 133.400000  69.700000 ;
      RECT 132.170000  41.290000 132.915000  41.460000 ;
      RECT 132.195000  11.100000 132.705000  11.430000 ;
      RECT 132.195000  17.510000 132.705000  17.840000 ;
      RECT 132.210000  69.700000 133.400000  73.365000 ;
      RECT 132.230000  61.675000 132.400000  63.495000 ;
      RECT 132.230000  64.405000 132.400000  67.115000 ;
      RECT 132.240000  25.360000 132.780000  28.030000 ;
      RECT 132.240000  41.460000 132.770000  41.530000 ;
      RECT 132.250000  28.030000 132.780000  28.200000 ;
      RECT 132.250000  30.285000 132.420000  31.335000 ;
      RECT 132.250000  33.015000 132.420000  35.725000 ;
      RECT 132.265000  11.430000 132.635000  17.510000 ;
      RECT 132.285000  85.770000 132.935000  86.780000 ;
      RECT 132.290000  44.740000 132.590000  45.375000 ;
      RECT 132.315000  74.760000 132.485000  74.790000 ;
      RECT 132.315000  74.960000 132.485000  75.770000 ;
      RECT 132.350000  24.795000 135.430000  25.310000 ;
      RECT 132.350000  25.310000 132.780000  25.360000 ;
      RECT 132.355000  75.990000 132.885000  76.160000 ;
      RECT 132.370000   6.510000 134.060000   6.680000 ;
      RECT 132.390000  49.985000 132.830000  60.365000 ;
      RECT 132.410000  18.940000 132.700000  21.330000 ;
      RECT 132.410000  21.330000 132.705000  22.705000 ;
      RECT 132.460000  22.705000 132.630000  24.320000 ;
      RECT 132.540000  48.105000 133.295000  48.275000 ;
      RECT 132.565000  82.220000 132.735000  83.290000 ;
      RECT 132.565000  83.460000 132.735000  84.930000 ;
      RECT 132.630000  43.405000 132.800000  44.415000 ;
      RECT 132.715000  76.160000 132.885000  80.820000 ;
      RECT 132.740000 200.085000 133.410000 200.255000 ;
      RECT 132.740000 216.235000 133.410000 216.405000 ;
      RECT 132.745000  38.010000 132.915000  41.290000 ;
      RECT 132.765000  46.335000 133.295000  46.505000 ;
      RECT 132.765000  85.760000 132.935000  85.770000 ;
      RECT 132.780000  61.675000 132.950000  67.420000 ;
      RECT 132.785000  44.630000 132.955000  45.300000 ;
      RECT 132.805000  11.600000 132.975000  13.210000 ;
      RECT 132.805000  13.830000 132.975000  14.160000 ;
      RECT 132.805000  14.330000 132.975000  17.040000 ;
      RECT 132.825000  42.510000 133.360000  43.085000 ;
      RECT 132.870000  81.330000 133.540000  81.500000 ;
      RECT 132.925000  21.225000 133.470000  21.395000 ;
      RECT 132.930000  41.635000 133.100000  42.030000 ;
      RECT 132.930000  42.200000 133.100000  42.305000 ;
      RECT 132.950000   5.020000 133.120000   6.280000 ;
      RECT 132.950000   7.080000 133.120000   9.790000 ;
      RECT 133.010000  49.985000 133.180000  60.365000 ;
      RECT 133.035000  26.165000 133.205000  26.835000 ;
      RECT 133.050000  61.175000 133.560000  61.505000 ;
      RECT 133.050000  67.585000 133.560000  67.915000 ;
      RECT 133.055000  81.950000 133.225000  84.850000 ;
      RECT 133.065000  17.700000 133.595000  17.870000 ;
      RECT 133.075000  11.100000 133.585000  11.430000 ;
      RECT 133.075000  17.510000 133.585000  17.700000 ;
      RECT 133.090000  43.405000 133.295000  44.415000 ;
      RECT 133.120000  61.505000 133.490000  67.585000 ;
      RECT 133.125000  44.415000 133.295000  46.335000 ;
      RECT 133.125000  46.505000 133.295000  48.105000 ;
      RECT 133.130000  33.015000 133.300000  35.725000 ;
      RECT 133.145000  11.430000 133.515000  17.510000 ;
      RECT 133.235000  75.160000 133.765000  75.330000 ;
      RECT 133.255000  27.175000 134.535000  28.305000 ;
      RECT 133.345000  60.535000 137.075000  60.855000 ;
      RECT 133.350000  49.595000 134.020000  60.535000 ;
      RECT 133.420000 106.360000 133.950000 106.530000 ;
      RECT 133.440000  85.785000 136.550000  86.315000 ;
      RECT 133.500000 105.400000 133.670000 106.360000 ;
      RECT 133.500000 106.530000 133.670000 106.750000 ;
      RECT 133.545000  82.220000 133.715000  83.300000 ;
      RECT 133.545000  83.300000 134.245000  83.470000 ;
      RECT 133.545000  83.470000 133.715000  84.930000 ;
      RECT 133.555000  77.300000 138.835000  77.480000 ;
      RECT 133.555000  77.480000 134.085000  78.010000 ;
      RECT 133.565000  25.730000 134.145000  26.865000 ;
      RECT 133.570000  70.200000 134.100000  70.370000 ;
      RECT 133.575000  85.555000 136.550000  85.785000 ;
      RECT 133.575000  86.315000 136.550000  87.700000 ;
      RECT 133.590000  37.870000 133.760000  44.425000 ;
      RECT 133.590000  45.065000 133.760000  48.465000 ;
      RECT 133.595000  74.760000 133.765000  75.160000 ;
      RECT 133.595000  75.330000 133.765000  75.770000 ;
      RECT 133.595000  76.070000 133.765000  77.300000 ;
      RECT 133.595000  78.010000 133.765000  80.820000 ;
      RECT 133.660000  61.675000 133.830000  62.725000 ;
      RECT 133.660000  62.955000 133.830000  63.285000 ;
      RECT 133.660000  63.905000 133.830000  64.235000 ;
      RECT 133.660000  64.405000 133.830000  67.115000 ;
      RECT 133.685000  11.725000 133.855000  17.345000 ;
      RECT 133.695000  19.960000 134.205000  24.415000 ;
      RECT 133.790000  81.030000 134.800000  81.545000 ;
      RECT 133.795000 106.870000 138.910000 106.920000 ;
      RECT 133.805000   8.840000 137.260000   9.010000 ;
      RECT 133.805000   9.010000 133.975000  10.760000 ;
      RECT 133.835000  69.485000 134.005000  70.200000 ;
      RECT 133.835000  70.370000 134.005000  73.215000 ;
      RECT 133.835000  85.150000 135.185000  85.320000 ;
      RECT 133.840000 113.910000 136.840000 164.900000 ;
      RECT 133.840000 200.495000 134.370000 215.995000 ;
      RECT 133.880000 181.885000 138.590000 182.155000 ;
      RECT 133.880000 185.735000 138.590000 186.005000 ;
      RECT 133.935000  74.540000 134.225000  76.420000 ;
      RECT 133.935000  76.420000 138.835000  76.590000 ;
      RECT 133.955000  11.100000 134.465000  11.430000 ;
      RECT 133.955000  17.510000 134.465000  17.840000 ;
      RECT 133.990000  42.510000 134.525000  43.085000 ;
      RECT 134.010000  30.285000 134.180000  31.350000 ;
      RECT 134.010000  31.520000 134.180000  31.895000 ;
      RECT 134.010000  32.515000 134.180000  35.725000 ;
      RECT 134.025000  11.430000 134.395000  13.590000 ;
      RECT 134.025000  13.590000 135.285000  13.850000 ;
      RECT 134.025000  13.850000 134.395000  17.510000 ;
      RECT 134.050000   4.990000 134.580000   5.160000 ;
      RECT 134.055000  43.405000 134.260000  44.415000 ;
      RECT 134.055000  44.415000 134.225000  46.335000 ;
      RECT 134.055000  46.335000 134.585000  46.505000 ;
      RECT 134.055000  46.505000 134.225000  48.105000 ;
      RECT 134.055000  48.105000 134.810000  48.275000 ;
      RECT 134.070000  18.210000 139.275000  18.880000 ;
      RECT 134.070000  18.880000 144.775000  18.920000 ;
      RECT 134.160000 105.210000 138.910000 105.280000 ;
      RECT 134.160000 105.990000 138.910000 106.160000 ;
      RECT 134.185000  18.920000 144.775000  19.030000 ;
      RECT 134.190000  49.045000 134.720000  49.595000 ;
      RECT 134.190000  49.595000 137.070000  49.765000 ;
      RECT 134.190000  49.955000 134.980000  54.705000 ;
      RECT 134.190000  54.705000 134.360000  60.365000 ;
      RECT 134.230000   5.160000 134.400000   8.160000 ;
      RECT 134.250000  41.635000 134.420000  42.030000 ;
      RECT 134.250000  42.030000 135.280000  42.200000 ;
      RECT 134.250000  42.200000 134.420000  42.305000 ;
      RECT 134.255000  78.070000 134.425000  80.780000 ;
      RECT 134.280000  29.785000 134.790000  30.115000 ;
      RECT 134.350000  30.115000 134.720000  36.195000 ;
      RECT 134.355000  69.125000 135.405000  69.295000 ;
      RECT 134.355000  73.405000 134.725000  73.575000 ;
      RECT 134.375000  19.550000 135.895000  21.085000 ;
      RECT 134.375000  21.085000 134.545000  24.200000 ;
      RECT 134.390000  77.700000 135.060000  77.870000 ;
      RECT 134.395000  44.630000 134.565000  45.300000 ;
      RECT 134.395000  73.575000 134.725000  74.760000 ;
      RECT 134.395000  74.760000 135.045000  74.930000 ;
      RECT 134.425000  82.140000 134.595000  84.930000 ;
      RECT 134.435000  37.840000 138.675000  38.010000 ;
      RECT 134.435000  38.010000 134.605000  41.290000 ;
      RECT 134.435000  41.290000 135.180000  41.460000 ;
      RECT 134.550000  43.405000 134.720000  44.415000 ;
      RECT 134.565000  11.600000 134.735000  13.420000 ;
      RECT 134.565000  14.330000 134.735000  17.040000 ;
      RECT 134.580000  41.460000 135.110000  41.530000 ;
      RECT 134.590000  37.335000 135.260000  37.505000 ;
      RECT 134.595000  26.165000 134.765000  26.835000 ;
      RECT 134.760000  44.585000 135.300000  44.740000 ;
      RECT 134.760000  44.740000 135.060000  45.375000 ;
      RECT 134.760000  45.375000 135.300000  45.665000 ;
      RECT 134.770000  42.400000 135.300000  42.570000 ;
      RECT 134.775000  83.300000 135.475000  83.470000 ;
      RECT 134.800000 200.085000 135.470000 200.255000 ;
      RECT 134.800000 216.235000 135.470000 216.405000 ;
      RECT 134.810000  55.085000 137.340000  55.285000 ;
      RECT 134.810000  55.285000 134.980000  60.365000 ;
      RECT 134.875000  74.930000 135.045000  75.770000 ;
      RECT 134.890000  30.410000 135.060000  36.045000 ;
      RECT 134.890000  42.570000 135.300000  44.585000 ;
      RECT 134.915000  73.405000 135.445000  73.575000 ;
      RECT 134.940000  22.850000 136.390000  23.360000 ;
      RECT 134.940000  23.360000 135.430000  24.795000 ;
      RECT 135.010000  45.665000 135.300000  48.085000 ;
      RECT 135.100000  74.370000 139.220000  74.540000 ;
      RECT 135.115000  11.600000 135.285000  13.590000 ;
      RECT 135.115000  13.850000 135.285000  17.345000 ;
      RECT 135.135000  78.070000 135.305000  81.810000 ;
      RECT 135.135000  81.810000 136.355000  81.980000 ;
      RECT 135.150000  36.195000 135.680000  36.845000 ;
      RECT 135.160000  29.785000 135.670000  30.115000 ;
      RECT 135.225000  74.760000 135.925000  75.770000 ;
      RECT 135.225000  75.770000 135.755000  76.250000 ;
      RECT 135.230000  30.115000 135.600000  36.195000 ;
      RECT 135.230000  45.000000 135.760000  45.170000 ;
      RECT 135.305000  82.220000 135.475000  83.300000 ;
      RECT 135.305000  83.470000 135.475000  84.930000 ;
      RECT 135.315000  38.180000 135.620000  40.890000 ;
      RECT 135.385000  11.100000 135.895000  11.430000 ;
      RECT 135.385000  17.510000 135.895000  17.840000 ;
      RECT 135.390000  77.700000 136.060000  77.870000 ;
      RECT 135.450000  40.890000 135.620000  41.580000 ;
      RECT 135.450000  41.580000 135.665000  41.635000 ;
      RECT 135.450000  41.635000 135.700000  42.305000 ;
      RECT 135.455000  11.430000 135.825000  17.510000 ;
      RECT 135.470000  43.405000 135.665000  44.415000 ;
      RECT 135.470000  45.170000 135.640000  48.085000 ;
      RECT 135.495000  42.305000 135.665000  43.405000 ;
      RECT 135.510000   5.020000 135.680000   6.280000 ;
      RECT 135.510000   7.150000 135.680000   8.840000 ;
      RECT 135.510000  53.370000 136.040000  53.540000 ;
      RECT 135.540000  37.335000 136.210000  37.505000 ;
      RECT 135.585000 223.695000 136.195000 225.350000 ;
      RECT 135.590000  49.955000 135.760000  53.370000 ;
      RECT 135.590000  53.540000 135.760000  54.705000 ;
      RECT 135.620000  81.325000 136.290000  81.570000 ;
      RECT 135.690000  23.610000 135.860000  26.080000 ;
      RECT 135.770000  30.285000 135.940000  32.105000 ;
      RECT 135.770000  33.015000 135.940000  35.725000 ;
      RECT 135.790000  41.290000 136.460000  41.460000 ;
      RECT 135.825000  84.280000 136.355000  84.450000 ;
      RECT 135.870000  41.460000 136.365000  42.030000 ;
      RECT 135.870000  42.030000 136.400000  42.200000 ;
      RECT 135.890000  29.945000 136.420000  30.115000 ;
      RECT 135.900000 200.495000 136.430000 215.995000 ;
      RECT 135.925000  76.020000 136.595000  76.190000 ;
      RECT 135.925000 225.650000 136.095000 226.630000 ;
      RECT 135.925000 234.980000 136.095000 235.960000 ;
      RECT 135.925000 237.100000 136.095000 238.080000 ;
      RECT 135.930000  43.405000 136.580000  44.415000 ;
      RECT 135.930000  44.415000 136.100000  46.335000 ;
      RECT 135.930000  46.335000 136.460000  46.505000 ;
      RECT 135.930000  46.505000 136.100000  48.085000 ;
      RECT 135.970000  61.675000 136.140000  62.740000 ;
      RECT 135.970000  62.910000 136.140000  63.285000 ;
      RECT 135.970000  63.905000 136.140000  64.235000 ;
      RECT 135.970000  64.405000 136.140000  67.115000 ;
      RECT 135.980000  21.340000 136.390000  22.850000 ;
      RECT 135.980000  23.360000 136.390000  23.375000 ;
      RECT 135.990000  55.455000 136.160000  60.365000 ;
      RECT 135.995000  11.600000 136.165000  13.210000 ;
      RECT 135.995000  13.830000 136.165000  14.160000 ;
      RECT 135.995000  14.330000 136.165000  17.040000 ;
      RECT 136.015000  78.070000 136.185000  80.780000 ;
      RECT 136.030000 181.105000 138.590000 181.375000 ;
      RECT 136.030000 186.515000 138.590000 186.785000 ;
      RECT 136.090000   4.970000 136.620000   6.680000 ;
      RECT 136.110000  30.115000 136.420000  30.260000 ;
      RECT 136.110000  30.260000 136.490000  36.030000 ;
      RECT 136.155000  68.635000 136.325000  71.415000 ;
      RECT 136.155000  71.415000 137.045000  72.305000 ;
      RECT 136.155000  72.305000 136.325000  73.575000 ;
      RECT 136.185000  81.980000 136.355000  84.280000 ;
      RECT 136.185000  84.450000 136.355000  84.930000 ;
      RECT 136.195000  38.180000 136.365000  41.290000 ;
      RECT 136.240000  61.175000 136.750000  61.505000 ;
      RECT 136.240000  67.585000 136.750000  67.915000 ;
      RECT 136.255000  17.700000 136.785000  17.870000 ;
      RECT 136.265000  11.100000 136.775000  11.430000 ;
      RECT 136.265000  17.510000 136.775000  17.700000 ;
      RECT 136.270000  47.855000 136.440000  48.465000 ;
      RECT 136.275000  74.790000 136.805000  74.960000 ;
      RECT 136.280000  77.480000 137.170000  77.620000 ;
      RECT 136.310000  61.505000 136.680000  67.585000 ;
      RECT 136.335000  11.430000 136.705000  17.510000 ;
      RECT 136.355000  49.955000 136.525000  55.085000 ;
      RECT 136.410000  42.475000 139.070000  42.645000 ;
      RECT 136.410000  42.645000 136.580000  43.405000 ;
      RECT 136.420000  37.335000 138.450000  37.505000 ;
      RECT 136.495000  73.120000 137.025000  73.405000 ;
      RECT 136.495000  73.405000 137.045000  73.575000 ;
      RECT 136.515000  69.125000 137.045000  71.415000 ;
      RECT 136.515000  72.305000 137.045000  72.365000 ;
      RECT 136.570000  20.410000 136.740000  25.940000 ;
      RECT 136.590000  29.575000 137.120000  30.115000 ;
      RECT 136.590000  36.195000 137.100000  36.525000 ;
      RECT 136.630000  41.360000 137.160000  41.530000 ;
      RECT 136.635000  74.760000 136.805000  74.790000 ;
      RECT 136.635000  74.960000 136.805000  75.770000 ;
      RECT 136.660000  30.115000 137.030000  36.195000 ;
      RECT 136.675000  78.130000 136.845000  81.050000 ;
      RECT 136.675000  81.950000 136.845000  84.850000 ;
      RECT 136.680000  19.030000 144.775000  19.135000 ;
      RECT 136.680000  19.135000 142.810000  19.500000 ;
      RECT 136.750000  43.095000 137.280000  43.265000 ;
      RECT 136.750000  43.265000 136.920000  48.390000 ;
      RECT 136.790000   5.020000 136.960000   8.160000 ;
      RECT 136.810000  41.530000 136.980000  42.305000 ;
      RECT 136.820000 223.695000 137.670000 243.640000 ;
      RECT 136.850000  61.800000 137.020000  67.420000 ;
      RECT 136.860000 200.085000 137.530000 200.255000 ;
      RECT 136.860000 216.235000 137.530000 216.405000 ;
      RECT 136.875000  11.725000 137.045000  17.345000 ;
      RECT 136.975000  74.760000 137.685000  75.770000 ;
      RECT 136.975000  75.770000 137.515000  76.420000 ;
      RECT 137.025000  74.000000 137.615000  74.170000 ;
      RECT 137.075000  38.180000 137.335000  41.160000 ;
      RECT 137.090000   9.010000 137.260000  10.760000 ;
      RECT 137.090000  10.760000 146.035000  10.930000 ;
      RECT 137.090000  44.180000 138.910000  44.350000 ;
      RECT 137.090000  44.350000 137.280000  47.370000 ;
      RECT 137.090000  47.370000 137.620000  48.550000 ;
      RECT 137.090000  48.550000 139.980000  48.720000 ;
      RECT 137.120000  61.175000 137.630000  61.505000 ;
      RECT 137.120000  67.585000 137.630000  67.915000 ;
      RECT 137.130000   6.510000 139.160000   6.680000 ;
      RECT 137.135000  17.700000 137.665000  17.870000 ;
      RECT 137.135000  49.955000 137.305000  50.845000 ;
      RECT 137.135000  50.845000 137.970000  54.705000 ;
      RECT 137.145000  11.100000 137.655000  11.430000 ;
      RECT 137.145000  17.510000 137.655000  17.700000 ;
      RECT 137.165000  26.945000 144.190000  27.115000 ;
      RECT 137.170000  55.285000 137.340000  60.365000 ;
      RECT 137.180000  19.775000 142.890000  19.945000 ;
      RECT 137.190000  61.505000 137.560000  67.585000 ;
      RECT 137.200000  30.285000 137.370000  31.895000 ;
      RECT 137.200000  32.515000 137.370000  35.725000 ;
      RECT 137.215000  11.430000 137.585000  17.510000 ;
      RECT 137.220000  20.300000 137.390000  21.570000 ;
      RECT 137.220000  23.670000 137.390000  26.595000 ;
      RECT 137.235000  82.180000 137.405000  83.690000 ;
      RECT 137.235000  83.690000 137.765000  83.860000 ;
      RECT 137.235000  83.860000 137.405000  86.930000 ;
      RECT 137.265000  68.925000 137.615000  74.000000 ;
      RECT 137.335000  78.075000 137.505000  80.785000 ;
      RECT 137.355000  81.430000 138.025000  81.600000 ;
      RECT 137.415000  68.205000 138.085000  68.545000 ;
      RECT 137.425000  49.005000 138.625000  49.175000 ;
      RECT 137.450000  42.840000 137.620000  44.010000 ;
      RECT 137.450000  44.580000 137.620000  45.280000 ;
      RECT 137.450000  45.280000 137.980000  45.450000 ;
      RECT 137.450000  45.450000 137.620000  47.080000 ;
      RECT 137.470000  29.785000 137.980000  29.945000 ;
      RECT 137.470000  29.945000 138.000000  30.115000 ;
      RECT 137.470000  36.195000 137.980000  36.525000 ;
      RECT 137.470000  77.700000 138.140000  77.870000 ;
      RECT 137.495000  81.400000 138.025000  81.430000 ;
      RECT 137.535000  38.180000 137.795000  41.160000 ;
      RECT 137.540000  30.115000 137.910000  36.195000 ;
      RECT 137.590000  55.895000 138.120000  56.065000 ;
      RECT 137.625000  22.080000 139.505000  22.670000 ;
      RECT 137.685000  76.020000 138.355000  76.065000 ;
      RECT 137.685000  76.065000 138.735000  76.190000 ;
      RECT 137.720000  42.470000 139.070000  42.475000 ;
      RECT 137.730000  61.675000 137.900000  63.495000 ;
      RECT 137.730000  64.405000 137.900000  67.115000 ;
      RECT 137.755000  11.600000 137.925000  13.420000 ;
      RECT 137.755000  14.330000 137.925000  17.040000 ;
      RECT 137.800000  54.705000 137.970000  55.895000 ;
      RECT 137.815000  73.830000 139.135000  74.370000 ;
      RECT 137.845000  76.190000 138.735000  76.235000 ;
      RECT 137.880000  42.840000 138.050000  44.180000 ;
      RECT 137.930000  46.335000 138.460000  47.370000 ;
      RECT 137.930000  47.370000 138.800000  48.380000 ;
      RECT 137.950000  56.755000 138.800000  58.725000 ;
      RECT 137.950000  58.725000 138.840000  59.255000 ;
      RECT 137.950000  59.255000 138.800000  60.485000 ;
      RECT 137.955000  20.240000 138.215000  21.310000 ;
      RECT 137.955000  25.675000 138.215000  26.655000 ;
      RECT 137.955000  49.175000 138.625000  50.625000 ;
      RECT 137.960000 200.495000 138.490000 215.995000 ;
      RECT 138.000000  23.885000 138.170000  25.675000 ;
      RECT 138.010000  70.655000 138.885000  71.185000 ;
      RECT 138.035000  71.380000 138.205000  72.600000 ;
      RECT 138.035000  72.600000 138.255000  73.610000 ;
      RECT 138.070000   5.020000 138.240000   6.280000 ;
      RECT 138.070000   7.080000 138.240000   9.790000 ;
      RECT 138.080000  30.285000 138.250000  36.030000 ;
      RECT 138.080000 181.075000 138.590000 181.105000 ;
      RECT 138.080000 181.375000 138.590000 181.405000 ;
      RECT 138.080000 181.855000 138.590000 181.885000 ;
      RECT 138.080000 182.155000 138.590000 182.185000 ;
      RECT 138.080000 185.705000 138.590000 185.735000 ;
      RECT 138.080000 186.005000 138.590000 186.035000 ;
      RECT 138.080000 186.485000 138.590000 186.515000 ;
      RECT 138.080000 186.785000 138.590000 186.815000 ;
      RECT 138.095000  56.265000 138.625000  56.435000 ;
      RECT 138.115000  82.180000 138.285000  86.930000 ;
      RECT 138.215000  78.075000 138.385000  80.785000 ;
      RECT 138.225000  74.790000 138.755000  74.960000 ;
      RECT 138.245000 113.195000 138.915000 113.525000 ;
      RECT 138.280000  61.675000 138.450000  62.725000 ;
      RECT 138.280000  62.955000 138.450000  63.285000 ;
      RECT 138.280000  63.905000 138.450000  64.235000 ;
      RECT 138.280000  64.405000 138.450000  67.115000 ;
      RECT 138.295000  55.785000 138.625000  56.265000 ;
      RECT 138.305000  11.600000 138.475000  13.420000 ;
      RECT 138.305000  14.330000 138.475000  17.040000 ;
      RECT 138.310000  42.840000 138.480000  44.010000 ;
      RECT 138.350000  29.785000 139.740000  30.115000 ;
      RECT 138.350000  36.195000 139.740000  36.525000 ;
      RECT 138.350000 113.910000 141.350000 164.900000 ;
      RECT 138.375000  71.185000 138.885000  72.250000 ;
      RECT 138.395000  74.760000 138.565000  74.790000 ;
      RECT 138.395000  74.960000 138.565000  75.770000 ;
      RECT 138.405000  87.150000 139.755000  87.320000 ;
      RECT 138.420000  30.115000 138.790000  36.195000 ;
      RECT 138.435000 222.080000 139.285000 245.255000 ;
      RECT 138.470000  77.700000 139.140000  77.870000 ;
      RECT 138.505000  38.010000 138.675000  41.360000 ;
      RECT 138.505000  41.360000 139.035000  41.530000 ;
      RECT 138.505000  72.935000 139.035000  73.105000 ;
      RECT 138.550000  61.175000 139.060000  61.505000 ;
      RECT 138.550000  67.585000 139.060000  67.915000 ;
      RECT 138.565000   9.990000 139.095000  10.590000 ;
      RECT 138.565000  11.260000 139.095000  11.430000 ;
      RECT 138.575000  11.100000 139.085000  11.260000 ;
      RECT 138.575000  17.510000 139.085000  17.840000 ;
      RECT 138.620000  61.505000 138.990000  67.585000 ;
      RECT 138.630000  44.580000 138.800000  45.760000 ;
      RECT 138.630000  45.760000 141.160000  45.930000 ;
      RECT 138.630000  45.930000 138.800000  47.080000 ;
      RECT 138.645000  11.430000 139.015000  17.510000 ;
      RECT 138.680000  50.845000 138.850000  55.525000 ;
      RECT 138.740000  42.840000 138.910000  44.180000 ;
      RECT 138.760000 181.235000 138.930000 181.560000 ;
      RECT 138.760000 181.560000 139.290000 182.730000 ;
      RECT 138.760000 185.070000 139.290000 187.295000 ;
      RECT 138.760000 189.635000 139.290000 190.805000 ;
      RECT 138.780000  20.300000 138.950000  21.570000 ;
      RECT 138.780000  23.670000 138.950000  26.595000 ;
      RECT 138.805000  83.690000 139.335000  83.860000 ;
      RECT 138.840000  55.895000 139.370000  56.065000 ;
      RECT 138.865000  72.600000 139.035000  72.935000 ;
      RECT 138.865000  73.105000 139.035000  73.490000 ;
      RECT 138.865000  73.490000 139.475000  73.660000 ;
      RECT 138.905000  49.090000 139.575000  50.625000 ;
      RECT 138.920000 200.085000 139.590000 200.255000 ;
      RECT 138.920000 216.235000 139.590000 216.405000 ;
      RECT 138.960000  30.285000 139.130000  31.895000 ;
      RECT 138.960000  32.515000 139.130000  35.725000 ;
      RECT 138.995000  81.430000 139.265000  81.600000 ;
      RECT 138.995000  81.600000 139.165000  83.690000 ;
      RECT 138.995000  83.860000 139.165000  86.930000 ;
      RECT 139.005000  77.080000 139.535000  77.250000 ;
      RECT 139.040000  55.785000 139.370000  55.895000 ;
      RECT 139.040000  56.065000 139.370000  56.295000 ;
      RECT 139.045000  53.995000 139.375000  54.325000 ;
      RECT 139.085000  37.870000 139.255000  40.870000 ;
      RECT 139.095000  68.375000 139.845000  68.545000 ;
      RECT 139.095000  78.075000 139.265000  81.430000 ;
      RECT 139.120000 181.235000 139.290000 181.560000 ;
      RECT 139.150000  46.165000 139.480000  47.015000 ;
      RECT 139.160000  61.675000 139.330000  67.415000 ;
      RECT 139.170000   6.880000 139.700000   7.050000 ;
      RECT 139.170000  42.840000 139.340000  44.010000 ;
      RECT 139.175000  68.205000 139.845000  68.375000 ;
      RECT 139.185000  11.725000 139.355000  17.345000 ;
      RECT 139.200000  53.370000 139.730000  53.540000 ;
      RECT 139.230000  47.015000 139.400000  47.625000 ;
      RECT 139.260000 104.700000 139.430000 107.065000 ;
      RECT 139.275000  74.760000 139.560000  75.770000 ;
      RECT 139.300000  30.115000 139.670000  36.195000 ;
      RECT 139.305000  45.280000 139.980000  45.450000 ;
      RECT 139.305000  73.660000 139.475000  73.930000 ;
      RECT 139.305000  73.930000 139.560000  74.000000 ;
      RECT 139.305000  74.000000 139.980000  74.170000 ;
      RECT 139.305000  74.170000 139.560000  74.200000 ;
      RECT 139.345000  76.575000 139.515000  77.080000 ;
      RECT 139.350000   5.020000 139.520000   6.880000 ;
      RECT 139.350000   7.050000 139.520000   9.790000 ;
      RECT 139.390000  74.200000 139.560000  74.760000 ;
      RECT 139.425000  42.470000 140.775000  42.640000 ;
      RECT 139.425000  42.640000 140.675000  42.670000 ;
      RECT 139.430000  61.175000 139.940000  61.505000 ;
      RECT 139.430000  67.585000 139.940000  67.915000 ;
      RECT 139.435000  81.450000 140.105000  81.940000 ;
      RECT 139.445000  17.510000 139.975000  18.670000 ;
      RECT 139.455000  11.100000 139.965000  11.430000 ;
      RECT 139.460000 181.075000 139.970000 181.105000 ;
      RECT 139.460000 181.105000 142.020000 181.375000 ;
      RECT 139.460000 181.375000 139.970000 181.405000 ;
      RECT 139.460000 181.855000 139.970000 181.885000 ;
      RECT 139.460000 181.885000 144.170000 182.155000 ;
      RECT 139.460000 182.155000 139.970000 182.185000 ;
      RECT 139.460000 185.705000 139.970000 185.735000 ;
      RECT 139.460000 185.735000 144.170000 186.005000 ;
      RECT 139.460000 186.005000 139.970000 186.035000 ;
      RECT 139.460000 186.485000 139.970000 186.515000 ;
      RECT 139.460000 186.515000 142.020000 186.785000 ;
      RECT 139.460000 186.785000 139.970000 186.815000 ;
      RECT 139.460000 190.115000 139.970000 190.145000 ;
      RECT 139.460000 190.145000 142.020000 190.415000 ;
      RECT 139.460000 190.415000 139.970000 190.445000 ;
      RECT 139.460000 190.895000 139.970000 190.925000 ;
      RECT 139.460000 190.925000 144.170000 191.195000 ;
      RECT 139.460000 191.195000 139.970000 191.225000 ;
      RECT 139.500000  61.505000 139.870000  63.455000 ;
      RECT 139.500000  63.455000 140.120000  63.625000 ;
      RECT 139.500000  63.625000 139.870000  67.585000 ;
      RECT 139.515000  20.240000 139.775000  21.310000 ;
      RECT 139.515000  25.675000 139.775000  26.655000 ;
      RECT 139.525000  11.430000 139.895000  17.510000 ;
      RECT 139.560000  23.885000 139.730000  25.675000 ;
      RECT 139.560000  50.845000 139.730000  53.370000 ;
      RECT 139.560000  53.540000 139.730000  56.265000 ;
      RECT 139.560000  56.265000 140.090000  56.435000 ;
      RECT 139.565000  71.415000 140.455000  72.305000 ;
      RECT 139.600000  42.840000 139.770000  44.180000 ;
      RECT 139.600000  44.180000 141.160000  44.350000 ;
      RECT 139.645000  68.925000 140.305000  70.860000 ;
      RECT 139.645000  70.860000 140.455000  71.415000 ;
      RECT 139.645000  72.305000 140.455000  72.365000 ;
      RECT 139.645000  72.365000 140.305000  73.610000 ;
      RECT 139.720000   6.510000 140.250000   6.680000 ;
      RECT 139.785000  22.080000 141.065000  22.670000 ;
      RECT 139.810000  44.580000 139.980000  45.280000 ;
      RECT 139.810000  45.450000 139.980000  45.590000 ;
      RECT 139.810000  46.100000 139.980000  48.550000 ;
      RECT 139.840000  30.285000 140.010000  36.045000 ;
      RECT 139.875000  82.180000 140.045000  86.930000 ;
      RECT 139.880000  57.325000 140.050000  60.405000 ;
      RECT 139.900000   5.020000 140.070000   6.510000 ;
      RECT 139.900000   6.680000 140.070000   9.790000 ;
      RECT 139.900000  50.875000 140.350000  51.740000 ;
      RECT 139.900000  51.740000 140.430000  51.910000 ;
      RECT 139.900000  51.910000 140.085000  52.775000 ;
      RECT 139.900000  52.775000 140.350000  53.770000 ;
      RECT 139.900000  53.770000 140.430000  54.055000 ;
      RECT 139.900000  54.055000 142.550000  54.385000 ;
      RECT 139.900000  54.385000 141.225000  54.660000 ;
      RECT 140.020000 200.495000 140.550000 215.995000 ;
      RECT 140.030000  42.840000 140.200000  44.010000 ;
      RECT 140.040000  61.675000 140.210000  62.740000 ;
      RECT 140.040000  62.910000 140.210000  63.285000 ;
      RECT 140.040000  63.905000 140.210000  64.235000 ;
      RECT 140.040000  64.405000 140.210000  67.115000 ;
      RECT 140.050000 220.085000 140.900000 247.105000 ;
      RECT 140.065000  11.600000 140.235000  13.210000 ;
      RECT 140.065000  13.830000 140.235000  14.160000 ;
      RECT 140.065000  14.330000 140.235000  17.040000 ;
      RECT 140.110000  29.785000 140.620000  30.115000 ;
      RECT 140.110000  36.195000 140.620000  36.525000 ;
      RECT 140.135000  68.635000 140.305000  68.925000 ;
      RECT 140.145000  18.040000 143.345000  18.855000 ;
      RECT 140.145000  18.855000 144.775000  18.880000 ;
      RECT 140.180000  30.115000 140.550000  36.195000 ;
      RECT 140.190000 180.765000 155.140000 180.935000 ;
      RECT 140.190000 181.545000 155.140000 181.715000 ;
      RECT 140.190000 182.325000 155.140000 182.495000 ;
      RECT 140.190000 185.395000 155.140000 185.565000 ;
      RECT 140.190000 186.175000 155.140000 186.345000 ;
      RECT 140.190000 186.955000 155.140000 187.125000 ;
      RECT 140.190000 189.805000 155.140000 189.975000 ;
      RECT 140.190000 190.585000 155.140000 190.755000 ;
      RECT 140.190000 191.365000 155.140000 191.535000 ;
      RECT 140.195000 103.770000 140.365000 108.380000 ;
      RECT 140.250000 183.525000 158.850000 184.375000 ;
      RECT 140.250000 188.010000 158.850000 188.860000 ;
      RECT 140.255000  52.095000 140.585000  52.230000 ;
      RECT 140.255000  52.230000 140.785000  52.400000 ;
      RECT 140.255000  52.400000 140.585000  52.605000 ;
      RECT 140.265000  74.400000 140.435000  81.020000 ;
      RECT 140.310000  61.175000 140.820000  61.505000 ;
      RECT 140.310000  67.585000 140.820000  67.590000 ;
      RECT 140.310000  67.590000 141.700000  67.915000 ;
      RECT 140.325000  10.260000 140.835000  10.390000 ;
      RECT 140.325000  10.390000 140.855000  10.560000 ;
      RECT 140.325000  10.560000 140.835000  10.590000 ;
      RECT 140.335000  11.100000 140.845000  11.430000 ;
      RECT 140.335000  17.510000 140.845000  17.840000 ;
      RECT 140.340000  20.300000 140.510000  21.655000 ;
      RECT 140.340000  23.670000 140.510000  26.595000 ;
      RECT 140.355000  85.820000 140.535000  86.350000 ;
      RECT 140.365000  81.950000 140.535000  85.820000 ;
      RECT 140.365000  86.350000 140.535000  86.765000 ;
      RECT 140.380000  61.505000 140.750000  67.585000 ;
      RECT 140.405000  11.430000 140.775000  17.510000 ;
      RECT 140.430000  37.765000 140.600000  40.845000 ;
      RECT 140.460000  42.840000 140.630000  44.180000 ;
      RECT 140.560000  57.005000 141.225000  57.175000 ;
      RECT 140.560000  57.175000 141.195000  57.205000 ;
      RECT 140.560000  57.205000 140.730000  60.015000 ;
      RECT 140.600000   6.510000 142.290000   6.680000 ;
      RECT 140.605000  77.400000 141.025000  78.240000 ;
      RECT 140.605000  78.240000 141.445000  78.410000 ;
      RECT 140.605000  78.410000 141.025000  78.750000 ;
      RECT 140.605000  78.750000 140.775000  79.730000 ;
      RECT 140.605000  79.730000 141.025000  81.080000 ;
      RECT 140.615000  60.665000 143.380000  60.835000 ;
      RECT 140.625000  68.885000 140.795000  73.635000 ;
      RECT 140.630000  46.335000 141.160000  46.505000 ;
      RECT 140.640000  50.535000 141.730000  50.705000 ;
      RECT 140.640000  50.705000 140.810000  51.885000 ;
      RECT 140.640000  52.875000 140.810000  53.885000 ;
      RECT 140.680000  68.205000 141.350000  68.555000 ;
      RECT 140.695000  55.525000 141.225000  57.005000 ;
      RECT 140.720000  30.285000 140.890000  31.895000 ;
      RECT 140.720000  32.515000 140.890000  35.725000 ;
      RECT 140.755000  41.265000 141.720000  41.435000 ;
      RECT 140.755000  41.435000 141.065000  42.130000 ;
      RECT 140.755000  42.130000 141.285000  42.300000 ;
      RECT 140.805000 113.195000 141.475000 113.525000 ;
      RECT 140.855000  74.420000 141.025000  76.020000 ;
      RECT 140.855000  81.890000 141.025000  83.290000 ;
      RECT 140.855000  83.290000 141.385000  83.460000 ;
      RECT 140.855000  83.460000 141.025000  86.640000 ;
      RECT 140.865000  49.415000 141.535000  50.365000 ;
      RECT 140.890000  42.840000 141.060000  44.010000 ;
      RECT 140.895000  38.155000 141.180000  40.865000 ;
      RECT 140.895000  40.865000 141.065000  41.095000 ;
      RECT 140.920000  61.800000 141.090000  67.420000 ;
      RECT 140.945000  11.600000 141.185000  17.345000 ;
      RECT 140.980000 200.085000 141.650000 200.255000 ;
      RECT 140.980000 216.235000 141.650000 216.405000 ;
      RECT 140.990000  29.785000 141.500000  30.115000 ;
      RECT 140.990000  36.195000 141.500000  36.525000 ;
      RECT 140.990000  44.350000 141.160000  45.760000 ;
      RECT 140.990000  46.100000 141.160000  46.335000 ;
      RECT 140.990000  46.505000 141.160000  48.380000 ;
      RECT 140.990000  79.075000 141.500000  79.120000 ;
      RECT 140.990000  79.120000 141.555000  79.290000 ;
      RECT 140.990000  79.290000 141.500000  79.405000 ;
      RECT 141.015000  11.260000 141.545000  11.430000 ;
      RECT 141.015000  11.430000 141.185000  11.600000 ;
      RECT 141.060000  30.115000 141.430000  36.195000 ;
      RECT 141.060000  50.875000 141.270000  51.885000 ;
      RECT 141.060000  51.885000 141.260000  52.875000 ;
      RECT 141.060000  52.875000 141.270000  53.935000 ;
      RECT 141.060000  53.935000 142.550000  54.055000 ;
      RECT 141.075000  20.240000 141.335000  21.310000 ;
      RECT 141.075000  25.675000 141.335000  26.655000 ;
      RECT 141.100000  76.370000 144.830000  76.540000 ;
      RECT 141.120000  23.885000 141.290000  25.675000 ;
      RECT 141.130000 104.530000 153.065000 104.700000 ;
      RECT 141.130000 104.700000 141.300000 107.450000 ;
      RECT 141.130000 107.450000 153.065000 107.620000 ;
      RECT 141.140000  54.920000 141.670000  55.090000 ;
      RECT 141.145000  87.150000 143.175000  87.320000 ;
      RECT 141.180000   5.020000 141.350000   6.280000 ;
      RECT 141.180000   7.080000 141.350000   9.790000 ;
      RECT 141.190000  61.175000 141.700000  61.505000 ;
      RECT 141.190000  67.585000 141.700000  67.590000 ;
      RECT 141.230000 239.550000 146.095000 241.240000 ;
      RECT 141.230000 242.025000 146.425000 243.720000 ;
      RECT 141.235000  37.335000 143.490000  37.505000 ;
      RECT 141.235000  41.085000 141.905000  41.255000 ;
      RECT 141.235000  41.255000 141.720000  41.265000 ;
      RECT 141.235000  41.760000 141.765000  41.930000 ;
      RECT 141.260000  61.505000 141.630000  63.695000 ;
      RECT 141.260000  63.695000 142.520000  63.865000 ;
      RECT 141.260000  63.865000 141.630000  67.585000 ;
      RECT 141.310000 243.890000 143.665000 244.175000 ;
      RECT 141.310000 244.175000 141.680000 244.345000 ;
      RECT 141.310000 244.345000 142.060000 246.365000 ;
      RECT 141.310000 246.365000 141.680000 246.535000 ;
      RECT 141.310000 246.535000 143.665000 246.935000 ;
      RECT 141.340000  57.305000 141.510000  60.405000 ;
      RECT 141.345000  22.080000 143.990000  22.670000 ;
      RECT 141.350000  37.505000 143.490000  37.595000 ;
      RECT 141.350000  37.595000 141.720000  41.085000 ;
      RECT 141.350000  43.110000 141.880000  48.390000 ;
      RECT 141.395000  54.555000 141.670000  54.920000 ;
      RECT 141.395000  55.090000 141.670000  55.565000 ;
      RECT 141.395000  55.565000 141.565000  56.870000 ;
      RECT 141.395000  56.870000 142.290000  57.040000 ;
      RECT 141.405000  68.885000 141.575000  73.635000 ;
      RECT 141.430000  52.355000 141.940000  52.685000 ;
      RECT 141.455000  41.930000 141.765000  43.110000 ;
      RECT 141.495000  11.600000 141.665000  17.345000 ;
      RECT 141.545000  75.100000 144.935000  75.270000 ;
      RECT 141.560000  50.705000 141.730000  52.355000 ;
      RECT 141.560000  52.685000 141.730000  52.840000 ;
      RECT 141.600000  30.285000 141.770000  36.025000 ;
      RECT 141.650000 105.035000 152.555000 105.205000 ;
      RECT 141.650000 105.205000 146.400000 105.280000 ;
      RECT 141.650000 105.990000 146.400000 106.160000 ;
      RECT 141.650000 106.870000 146.400000 106.940000 ;
      RECT 141.650000 106.940000 152.555000 107.110000 ;
      RECT 141.660000 221.045000 170.470000 221.215000 ;
      RECT 141.660000 221.215000 141.830000 231.605000 ;
      RECT 141.660000 231.605000 163.760000 232.050000 ;
      RECT 141.660000 232.050000 141.830000 238.575000 ;
      RECT 141.660000 238.575000 164.550000 239.105000 ;
      RECT 141.715000  68.205000 148.770000  68.385000 ;
      RECT 141.715000  68.385000 147.485000  68.555000 ;
      RECT 141.735000  55.735000 142.245000  56.265000 ;
      RECT 141.735000  56.265000 142.265000  56.515000 ;
      RECT 141.735000  56.515000 142.940000  56.700000 ;
      RECT 141.735000  81.890000 141.905000  86.640000 ;
      RECT 141.765000  11.100000 142.275000  11.430000 ;
      RECT 141.765000  17.510000 142.275000  17.840000 ;
      RECT 141.790000  77.010000 142.800000  77.180000 ;
      RECT 141.790000  81.300000 142.800000  81.470000 ;
      RECT 141.800000  61.675000 141.970000  63.495000 ;
      RECT 141.800000  64.405000 141.970000  67.115000 ;
      RECT 141.835000  11.430000 142.205000  17.510000 ;
      RECT 141.855000  21.125000 142.115000  21.765000 ;
      RECT 141.855000  23.495000 142.115000  26.595000 ;
      RECT 141.870000  29.785000 143.260000  30.085000 ;
      RECT 141.870000  30.085000 142.380000  30.115000 ;
      RECT 141.870000  36.195000 142.380000  36.225000 ;
      RECT 141.870000  36.225000 143.260000  36.525000 ;
      RECT 141.890000  37.765000 142.060000  40.865000 ;
      RECT 141.900000  20.300000 142.070000  21.125000 ;
      RECT 141.935000  41.445000 142.400000  41.615000 ;
      RECT 141.935000  41.615000 142.105000  42.520000 ;
      RECT 141.935000  42.520000 142.220000  42.690000 ;
      RECT 141.940000  30.115000 142.310000  36.195000 ;
      RECT 142.020000  53.770000 142.550000  53.935000 ;
      RECT 142.020000  54.385000 142.550000  54.660000 ;
      RECT 142.020000  80.875000 142.550000  81.300000 ;
      RECT 142.035000   8.840000 146.035000  10.760000 ;
      RECT 142.050000  42.690000 142.220000  43.615000 ;
      RECT 142.080000 200.495000 142.610000 215.995000 ;
      RECT 142.100000   4.970000 142.630000   5.140000 ;
      RECT 142.120000  57.040000 142.290000  60.015000 ;
      RECT 142.185000  68.555000 142.355000  73.635000 ;
      RECT 142.190000  76.895000 142.720000  77.010000 ;
      RECT 142.200000  50.865000 142.370000  53.770000 ;
      RECT 142.230000  40.395000 142.940000  40.865000 ;
      RECT 142.230000  40.865000 142.400000  41.445000 ;
      RECT 142.230000 244.175000 143.665000 246.535000 ;
      RECT 142.240000 221.465000 161.950000 222.075000 ;
      RECT 142.240000 222.245000 161.950000 222.855000 ;
      RECT 142.240000 223.025000 161.950000 223.635000 ;
      RECT 142.240000 223.805000 161.950000 224.415000 ;
      RECT 142.240000 224.585000 161.950000 225.195000 ;
      RECT 142.240000 225.365000 161.950000 225.975000 ;
      RECT 142.240000 226.145000 161.950000 226.755000 ;
      RECT 142.240000 226.925000 161.950000 227.535000 ;
      RECT 142.240000 227.705000 161.950000 228.315000 ;
      RECT 142.240000 228.485000 161.950000 229.095000 ;
      RECT 142.240000 229.265000 161.950000 229.875000 ;
      RECT 142.240000 230.045000 161.950000 230.655000 ;
      RECT 142.240000 230.825000 161.950000 231.435000 ;
      RECT 142.240000 232.220000 161.950000 232.715000 ;
      RECT 142.240000 232.885000 161.965000 233.495000 ;
      RECT 142.240000 233.665000 161.950000 234.160000 ;
      RECT 142.240000 234.330000 161.950000 234.825000 ;
      RECT 142.240000 234.995000 161.950000 235.605000 ;
      RECT 142.240000 235.775000 161.950000 236.270000 ;
      RECT 142.240000 236.465000 161.950000 236.960000 ;
      RECT 142.240000 237.130000 161.950000 237.740000 ;
      RECT 142.240000 237.910000 161.950000 238.405000 ;
      RECT 142.275000  41.785000 142.895000  42.115000 ;
      RECT 142.325000  22.670000 142.585000  23.405000 ;
      RECT 142.325000  23.405000 143.515000  23.710000 ;
      RECT 142.350000  61.675000 142.520000  63.695000 ;
      RECT 142.350000  63.865000 142.520000  67.420000 ;
      RECT 142.375000  11.600000 142.545000  13.210000 ;
      RECT 142.375000  13.830000 142.545000  14.160000 ;
      RECT 142.375000  14.330000 142.545000  17.040000 ;
      RECT 142.380000  54.660000 142.550000  55.565000 ;
      RECT 142.445000  83.290000 142.975000  83.460000 ;
      RECT 142.460000   5.140000 142.630000   8.160000 ;
      RECT 142.475000  25.675000 142.735000  26.655000 ;
      RECT 142.480000  30.285000 142.650000  31.895000 ;
      RECT 142.480000  32.515000 142.650000  35.725000 ;
      RECT 142.500000  48.350000 145.870000  48.520000 ;
      RECT 142.520000  23.885000 142.690000  25.675000 ;
      RECT 142.540000  45.290000 142.710000  48.000000 ;
      RECT 142.570000  41.360000 143.490000  41.530000 ;
      RECT 142.570000  41.530000 142.895000  41.785000 ;
      RECT 142.615000  81.890000 142.785000  83.290000 ;
      RECT 142.615000  83.460000 142.785000  86.640000 ;
      RECT 142.620000  61.175000 143.130000  61.505000 ;
      RECT 142.620000  67.585000 143.130000  67.915000 ;
      RECT 142.635000  20.240000 142.895000  21.310000 ;
      RECT 142.645000  11.100000 143.155000  11.430000 ;
      RECT 142.645000  17.510000 143.155000  17.840000 ;
      RECT 142.660000  48.215000 145.710000  48.350000 ;
      RECT 142.665000  55.895000 143.380000  56.065000 ;
      RECT 142.690000  61.505000 143.060000  63.455000 ;
      RECT 142.690000  63.455000 143.220000  63.625000 ;
      RECT 142.690000  63.625000 143.060000  67.585000 ;
      RECT 142.710000  55.835000 143.380000  55.895000 ;
      RECT 142.710000  56.065000 143.380000  56.345000 ;
      RECT 142.715000  11.430000 143.085000  17.510000 ;
      RECT 142.750000  30.085000 143.260000  30.115000 ;
      RECT 142.750000  36.195000 143.260000  36.225000 ;
      RECT 142.755000  22.840000 144.700000  23.235000 ;
      RECT 142.770000  38.155000 142.940000  40.395000 ;
      RECT 142.770000  56.700000 142.940000  57.680000 ;
      RECT 142.770000  58.805000 143.380000  60.665000 ;
      RECT 142.820000  30.115000 143.190000  36.195000 ;
      RECT 142.845000  77.400000 143.015000  78.750000 ;
      RECT 142.845000  79.540000 143.015000  81.080000 ;
      RECT 142.860000 113.910000 145.860000 164.900000 ;
      RECT 142.900000  55.495000 143.430000  55.665000 ;
      RECT 142.930000  42.605000 143.100000  44.400000 ;
      RECT 142.945000  45.030000 143.490000  45.200000 ;
      RECT 142.965000  68.885000 143.135000  73.635000 ;
      RECT 143.035000  44.570000 144.045000  44.740000 ;
      RECT 143.035000  44.740000 143.565000  44.800000 ;
      RECT 143.040000 200.085000 143.710000 200.255000 ;
      RECT 143.040000 216.235000 143.710000 216.405000 ;
      RECT 143.070000  77.010000 144.080000  77.180000 ;
      RECT 143.070000  81.300000 144.080000  81.470000 ;
      RECT 143.110000  37.595000 143.490000  38.615000 ;
      RECT 143.110000  56.345000 143.380000  58.805000 ;
      RECT 143.150000  42.000000 143.820000  42.170000 ;
      RECT 143.220000  42.170000 143.750000  42.300000 ;
      RECT 143.230000  61.675000 143.400000  62.740000 ;
      RECT 143.230000  62.910000 143.400000  63.285000 ;
      RECT 143.230000  63.905000 143.400000  64.235000 ;
      RECT 143.230000  64.405000 143.400000  67.115000 ;
      RECT 143.255000  11.725000 143.425000  17.345000 ;
      RECT 143.255000  23.710000 143.515000  26.595000 ;
      RECT 143.260000  54.555000 143.430000  55.495000 ;
      RECT 143.300000  80.875000 143.830000  81.300000 ;
      RECT 143.315000  20.815000 143.990000  21.145000 ;
      RECT 143.320000  40.195000 143.490000  41.360000 ;
      RECT 143.320000  45.000000 143.490000  45.030000 ;
      RECT 143.320000  45.200000 143.490000  48.000000 ;
      RECT 143.360000  30.285000 143.530000  36.025000 ;
      RECT 143.385000  88.895000 143.915000  89.065000 ;
      RECT 143.400000  19.325000 143.990000  20.815000 ;
      RECT 143.400000  21.145000 143.990000  22.080000 ;
      RECT 143.420000  38.970000 144.950000  39.720000 ;
      RECT 143.450000  42.505000 143.980000  42.675000 ;
      RECT 143.470000  76.895000 144.000000  77.010000 ;
      RECT 143.495000  81.890000 143.665000  86.640000 ;
      RECT 143.500000  61.175000 144.175000  61.345000 ;
      RECT 143.500000  61.345000 144.010000  61.505000 ;
      RECT 143.500000  67.585000 144.010000  67.915000 ;
      RECT 143.515000  17.510000 144.045000  18.670000 ;
      RECT 143.525000  11.100000 144.035000  11.430000 ;
      RECT 143.550000  56.670000 143.720000  60.405000 ;
      RECT 143.570000  61.505000 143.940000  67.585000 ;
      RECT 143.595000  11.430000 143.965000  17.510000 ;
      RECT 143.630000  29.785000 145.020000  30.085000 ;
      RECT 143.630000  30.085000 144.140000  30.115000 ;
      RECT 143.630000  36.195000 144.140000  36.225000 ;
      RECT 143.630000  36.225000 145.020000  36.525000 ;
      RECT 143.660000  37.765000 144.710000  38.970000 ;
      RECT 143.660000  39.720000 144.710000  40.865000 ;
      RECT 143.700000  30.115000 144.070000  36.195000 ;
      RECT 143.740000   5.020000 143.910000   6.280000 ;
      RECT 143.740000   7.150000 143.910000   8.840000 ;
      RECT 143.740000  87.150000 144.410000  87.320000 ;
      RECT 143.745000  68.555000 143.915000  73.635000 ;
      RECT 143.745000  88.610000 143.915000  88.895000 ;
      RECT 143.810000  42.675000 143.980000  43.615000 ;
      RECT 143.995000  83.290000 144.545000  83.460000 ;
      RECT 144.020000 192.700000 144.560000 192.870000 ;
      RECT 144.035000  25.675000 144.295000  26.655000 ;
      RECT 144.050000 192.620000 144.560000 192.700000 ;
      RECT 144.050000 192.870000 144.560000 192.950000 ;
      RECT 144.080000  23.885000 144.250000  25.675000 ;
      RECT 144.100000  45.290000 144.270000  48.000000 ;
      RECT 144.110000  61.800000 144.280000  67.420000 ;
      RECT 144.135000  11.600000 144.305000  13.420000 ;
      RECT 144.135000  14.330000 144.305000  17.040000 ;
      RECT 144.140000 200.495000 144.670000 215.995000 ;
      RECT 144.215000  18.040000 146.535000  18.440000 ;
      RECT 144.215000  18.440000 148.190000  18.660000 ;
      RECT 144.240000  30.285000 144.410000  31.895000 ;
      RECT 144.240000  32.515000 144.410000  35.725000 ;
      RECT 144.310000  22.190000 144.700000  22.840000 ;
      RECT 144.325000  44.570000 145.335000  44.740000 ;
      RECT 144.340000 180.935000 153.640000 181.375000 ;
      RECT 144.340000 181.885000 153.640000 182.325000 ;
      RECT 144.340000 185.565000 153.640000 186.005000 ;
      RECT 144.340000 186.515000 153.640000 186.955000 ;
      RECT 144.340000 189.975000 153.640000 190.415000 ;
      RECT 144.340000 190.925000 153.640000 191.365000 ;
      RECT 144.360000  75.270000 144.890000  75.330000 ;
      RECT 144.360000  79.110000 144.890000  79.280000 ;
      RECT 144.370000  79.075000 144.880000  79.110000 ;
      RECT 144.370000  79.280000 144.880000  79.405000 ;
      RECT 144.375000  81.890000 144.545000  83.290000 ;
      RECT 144.375000  83.460000 144.545000  86.640000 ;
      RECT 144.380000  61.175000 144.890000  61.505000 ;
      RECT 144.380000  67.585000 144.890000  67.915000 ;
      RECT 144.390000  42.505000 144.920000  42.675000 ;
      RECT 144.390000  42.675000 144.560000  43.615000 ;
      RECT 144.395000  18.660000 144.775000  18.855000 ;
      RECT 144.395000  19.135000 144.775000  21.150000 ;
      RECT 144.415000  78.240000 145.320000  78.410000 ;
      RECT 144.450000  61.505000 144.820000  67.585000 ;
      RECT 144.510000  30.085000 145.020000  30.115000 ;
      RECT 144.510000  36.195000 145.020000  36.225000 ;
      RECT 144.525000  68.885000 144.695000  73.635000 ;
      RECT 144.550000  42.000000 145.220000  42.170000 ;
      RECT 144.580000  30.115000 144.950000  36.195000 ;
      RECT 144.620000  42.170000 145.150000  42.300000 ;
      RECT 144.640000   4.515000 146.035000   8.840000 ;
      RECT 144.650000  61.075000 144.820000  61.175000 ;
      RECT 144.685000  11.600000 144.855000  13.420000 ;
      RECT 144.685000  14.330000 144.855000  17.040000 ;
      RECT 144.715000  87.885000 145.515000  90.920000 ;
      RECT 144.795000  50.330000 153.885000  59.670000 ;
      RECT 144.805000  44.740000 145.335000  44.800000 ;
      RECT 144.845000  77.400000 145.320000  78.240000 ;
      RECT 144.845000  78.410000 145.320000  78.750000 ;
      RECT 144.845000  79.730000 145.320000  81.080000 ;
      RECT 144.865000  17.295000 145.395000  17.465000 ;
      RECT 144.880000  37.335000 147.135000  37.505000 ;
      RECT 144.880000  37.505000 147.020000  37.595000 ;
      RECT 144.880000  37.595000 145.260000  38.615000 ;
      RECT 144.880000  40.195000 145.050000  41.360000 ;
      RECT 144.880000  41.360000 145.800000  41.530000 ;
      RECT 144.880000  45.000000 145.050000  45.030000 ;
      RECT 144.880000  45.030000 145.425000  45.200000 ;
      RECT 144.880000  45.200000 145.050000  48.000000 ;
      RECT 144.945000  19.565000 145.205000  24.340000 ;
      RECT 144.955000  11.100000 145.465000  11.430000 ;
      RECT 144.955000  17.465000 145.395000  17.510000 ;
      RECT 144.955000  17.510000 145.465000  17.840000 ;
      RECT 144.970000  25.390000 149.720000  25.560000 ;
      RECT 144.970000  26.470000 149.720000  26.640000 ;
      RECT 144.970000  27.550000 149.720000  27.720000 ;
      RECT 144.975000  83.290000 146.205000  83.460000 ;
      RECT 144.990000  19.530000 145.160000  19.565000 ;
      RECT 144.990000  61.675000 145.160000  63.495000 ;
      RECT 144.990000  64.405000 145.160000  67.115000 ;
      RECT 145.025000  11.430000 145.395000  17.295000 ;
      RECT 145.065000  81.920000 145.395000  83.290000 ;
      RECT 145.065000  86.430000 146.225000  86.940000 ;
      RECT 145.100000 200.085000 145.770000 200.255000 ;
      RECT 145.100000 216.235000 145.770000 216.405000 ;
      RECT 145.110000  61.260000 145.640000  61.430000 ;
      RECT 145.120000  30.285000 145.290000  36.025000 ;
      RECT 145.135000  74.400000 145.305000  74.930000 ;
      RECT 145.135000  75.430000 145.305000  76.020000 ;
      RECT 145.150000  78.750000 145.320000  79.730000 ;
      RECT 145.160000  24.800000 150.850000  24.970000 ;
      RECT 145.215000  18.850000 150.235000  19.020000 ;
      RECT 145.270000  42.605000 145.440000  44.400000 ;
      RECT 145.305000  68.555000 145.475000  73.635000 ;
      RECT 145.330000  61.430000 145.500000  61.645000 ;
      RECT 145.330000  61.645000 145.710000  61.815000 ;
      RECT 145.385000  36.195000 145.895000  36.225000 ;
      RECT 145.385000  36.225000 146.780000  36.525000 ;
      RECT 145.390000  29.785000 146.780000  30.085000 ;
      RECT 145.390000  30.085000 145.900000  30.115000 ;
      RECT 145.430000  38.155000 145.600000  40.395000 ;
      RECT 145.430000  40.395000 146.140000  40.865000 ;
      RECT 145.460000  30.115000 145.830000  36.195000 ;
      RECT 145.475000  41.530000 145.800000  41.785000 ;
      RECT 145.475000  41.785000 146.095000  42.115000 ;
      RECT 145.540000  61.815000 145.710000  63.495000 ;
      RECT 145.540000  64.405000 145.710000  67.115000 ;
      RECT 145.565000  11.725000 145.735000  17.345000 ;
      RECT 145.615000  78.240000 146.205000  78.410000 ;
      RECT 145.615000  78.950000 146.205000  79.120000 ;
      RECT 145.660000  45.290000 145.830000  48.000000 ;
      RECT 145.720000  63.695000 146.250000  63.865000 ;
      RECT 145.725000  22.700000 145.985000  23.340000 ;
      RECT 145.770000  19.530000 145.940000  22.700000 ;
      RECT 145.770000  23.340000 145.940000  24.280000 ;
      RECT 145.810000  61.175000 146.320000  61.505000 ;
      RECT 145.810000  67.585000 146.320000  67.590000 ;
      RECT 145.810000  67.590000 147.200000  67.915000 ;
      RECT 145.825000  11.260000 146.355000  11.430000 ;
      RECT 145.835000  11.100000 146.345000  11.260000 ;
      RECT 145.835000  17.510000 146.345000  17.840000 ;
      RECT 145.875000  74.920000 146.205000  78.240000 ;
      RECT 145.875000  78.410000 146.205000  78.440000 ;
      RECT 145.875000  79.120000 146.205000  83.290000 ;
      RECT 145.875000  83.460000 146.205000  83.830000 ;
      RECT 145.880000  61.505000 146.250000  63.695000 ;
      RECT 145.880000  63.865000 146.250000  67.585000 ;
      RECT 145.905000  11.430000 146.275000  17.510000 ;
      RECT 145.970000  40.865000 146.140000  41.445000 ;
      RECT 145.970000  41.445000 146.435000  41.615000 ;
      RECT 146.000000  30.285000 146.170000  31.895000 ;
      RECT 146.000000  32.515000 146.170000  35.725000 ;
      RECT 146.085000  68.885000 146.255000  73.635000 ;
      RECT 146.150000  42.520000 146.435000  42.690000 ;
      RECT 146.150000  42.690000 146.320000  43.615000 ;
      RECT 146.200000 200.495000 146.730000 215.995000 ;
      RECT 146.265000  41.615000 146.435000  42.520000 ;
      RECT 146.270000  30.085000 146.780000  30.115000 ;
      RECT 146.270000  36.195000 146.780000  36.225000 ;
      RECT 146.310000  37.765000 146.480000  40.865000 ;
      RECT 146.340000  30.115000 146.710000  36.195000 ;
      RECT 146.420000  61.800000 146.590000  67.420000 ;
      RECT 146.445000  11.600000 146.615000  13.210000 ;
      RECT 146.445000  13.830000 146.615000  14.160000 ;
      RECT 146.445000  14.330000 146.615000  17.040000 ;
      RECT 146.465000  41.085000 147.135000  41.255000 ;
      RECT 146.490000  43.110000 147.020000  48.390000 ;
      RECT 146.505000  19.565000 146.765000  24.340000 ;
      RECT 146.550000  19.530000 146.720000  19.565000 ;
      RECT 146.580000   4.515000 154.900000   4.685000 ;
      RECT 146.580000   4.685000 146.750000   9.785000 ;
      RECT 146.605000  41.760000 147.135000  41.930000 ;
      RECT 146.605000  41.930000 146.915000  43.110000 ;
      RECT 146.610000 106.360000 147.140000 106.530000 ;
      RECT 146.615000 239.550000 152.280000 241.240000 ;
      RECT 146.650000  37.595000 147.020000  41.085000 ;
      RECT 146.650000  41.255000 147.135000  41.265000 ;
      RECT 146.650000  41.265000 147.615000  41.435000 ;
      RECT 146.665000  86.430000 147.825000  86.940000 ;
      RECT 146.685000  74.920000 147.015000  78.240000 ;
      RECT 146.685000  78.240000 147.275000  78.410000 ;
      RECT 146.685000  78.410000 147.015000  78.440000 ;
      RECT 146.685000  78.950000 147.275000  79.120000 ;
      RECT 146.685000  79.120000 147.015000  83.290000 ;
      RECT 146.685000  83.290000 147.915000  83.460000 ;
      RECT 146.685000  83.460000 147.015000  83.830000 ;
      RECT 146.690000  61.175000 147.200000  61.505000 ;
      RECT 146.690000  67.585000 147.200000  67.590000 ;
      RECT 146.705000  17.510000 147.235000  18.270000 ;
      RECT 146.715000  11.100000 147.225000  11.430000 ;
      RECT 146.760000  61.505000 147.130000  67.585000 ;
      RECT 146.785000  11.430000 147.155000  17.510000 ;
      RECT 146.790000  88.630000 243.215000  93.070000 ;
      RECT 146.865000  68.555000 147.035000  73.635000 ;
      RECT 146.880000  10.295000 149.590000  10.465000 ;
      RECT 146.880000  30.285000 147.050000  36.025000 ;
      RECT 146.880000 105.400000 147.050000 106.360000 ;
      RECT 146.880000 106.530000 147.050000 106.750000 ;
      RECT 146.920000   8.830000 147.190000  10.295000 ;
      RECT 146.955000 242.030000 152.180000 243.720000 ;
      RECT 147.085000  42.130000 147.615000  42.300000 ;
      RECT 147.125000  22.015000 147.385000  22.655000 ;
      RECT 147.150000  29.785000 147.660000  30.115000 ;
      RECT 147.150000  36.195000 147.660000  36.525000 ;
      RECT 147.160000 200.085000 147.830000 200.255000 ;
      RECT 147.160000 216.235000 147.830000 216.405000 ;
      RECT 147.170000  19.530000 147.340000  22.015000 ;
      RECT 147.170000  22.655000 147.340000  24.280000 ;
      RECT 147.190000  38.155000 147.475000  40.865000 ;
      RECT 147.210000  44.180000 148.770000  44.350000 ;
      RECT 147.210000  44.350000 147.380000  45.760000 ;
      RECT 147.210000  45.760000 149.740000  45.930000 ;
      RECT 147.210000  46.100000 147.380000  46.335000 ;
      RECT 147.210000  46.335000 147.740000  46.505000 ;
      RECT 147.210000  46.505000 147.380000  48.380000 ;
      RECT 147.220000  30.115000 147.590000  36.195000 ;
      RECT 147.255000 105.205000 152.005000 105.280000 ;
      RECT 147.255000 105.990000 152.005000 106.160000 ;
      RECT 147.255000 106.870000 152.005000 106.940000 ;
      RECT 147.265000 113.195000 147.935000 113.525000 ;
      RECT 147.300000  61.675000 147.470000  62.740000 ;
      RECT 147.300000  62.910000 147.470000  63.285000 ;
      RECT 147.300000  63.905000 147.470000  64.235000 ;
      RECT 147.300000  64.405000 147.470000  67.115000 ;
      RECT 147.305000  40.865000 147.475000  41.095000 ;
      RECT 147.305000  41.435000 147.615000  42.130000 ;
      RECT 147.310000  42.840000 147.480000  44.010000 ;
      RECT 147.315000  71.040000 148.305000  71.240000 ;
      RECT 147.325000  11.600000 147.495000  17.345000 ;
      RECT 147.360000   5.035000 147.530000   8.850000 ;
      RECT 147.360000   8.850000 147.890000   9.020000 ;
      RECT 147.360000   9.020000 147.530000   9.785000 ;
      RECT 147.370000 113.910000 150.370000 164.900000 ;
      RECT 147.385000  71.240000 148.305000  72.305000 ;
      RECT 147.405000  18.040000 148.190000  18.440000 ;
      RECT 147.495000  81.920000 147.825000  83.290000 ;
      RECT 147.565000  61.260000 148.095000  61.430000 ;
      RECT 147.570000  61.175000 148.080000  61.260000 ;
      RECT 147.570000  61.430000 148.080000  61.505000 ;
      RECT 147.570000  67.585000 148.080000  67.915000 ;
      RECT 147.570000  77.400000 148.045000  78.240000 ;
      RECT 147.570000  78.240000 148.475000  78.410000 ;
      RECT 147.570000  78.410000 148.045000  78.750000 ;
      RECT 147.570000  78.750000 147.740000  79.730000 ;
      RECT 147.570000  79.730000 148.045000  81.080000 ;
      RECT 147.585000  74.400000 147.755000  74.930000 ;
      RECT 147.585000  75.430000 147.755000  76.020000 ;
      RECT 147.595000  42.470000 148.945000  42.640000 ;
      RECT 147.640000  61.505000 148.010000  67.585000 ;
      RECT 147.645000  68.635000 148.305000  71.040000 ;
      RECT 147.645000  72.305000 148.305000  73.635000 ;
      RECT 147.695000  42.640000 148.945000  42.670000 ;
      RECT 147.740000  42.840000 147.910000  44.180000 ;
      RECT 147.760000  30.285000 147.930000  31.895000 ;
      RECT 147.760000  32.515000 147.930000  35.725000 ;
      RECT 147.770000  37.765000 147.940000  40.845000 ;
      RECT 147.905000  20.875000 148.165000  21.515000 ;
      RECT 147.950000  19.530000 148.120000  20.875000 ;
      RECT 147.950000  21.515000 148.120000  24.280000 ;
      RECT 147.955000  75.100000 151.345000  75.270000 ;
      RECT 148.000000  75.270000 148.530000  75.330000 ;
      RECT 148.000000  79.110000 148.530000  79.280000 ;
      RECT 148.010000  79.075000 148.520000  79.110000 ;
      RECT 148.010000  79.280000 148.520000  79.405000 ;
      RECT 148.020000  11.600000 148.190000  13.410000 ;
      RECT 148.020000  13.830000 148.190000  18.040000 ;
      RECT 148.030000  29.785000 148.540000  30.115000 ;
      RECT 148.030000  36.195000 148.540000  36.525000 ;
      RECT 148.060000  76.370000 151.790000  76.540000 ;
      RECT 148.100000  30.115000 148.470000  36.195000 ;
      RECT 148.140000   4.685000 148.310000   9.785000 ;
      RECT 148.170000  42.840000 148.340000  44.010000 ;
      RECT 148.180000  61.675000 148.350000  67.415000 ;
      RECT 148.260000 200.495000 148.790000 215.995000 ;
      RECT 148.345000  81.890000 148.515000  83.290000 ;
      RECT 148.345000  83.290000 148.895000  83.460000 ;
      RECT 148.345000  83.460000 148.515000  86.640000 ;
      RECT 148.390000  44.580000 148.560000  45.280000 ;
      RECT 148.390000  45.280000 149.065000  45.450000 ;
      RECT 148.390000  45.450000 148.560000  45.590000 ;
      RECT 148.390000  46.100000 148.560000  48.550000 ;
      RECT 148.390000  48.550000 151.280000  48.720000 ;
      RECT 148.450000  61.175000 148.960000  61.505000 ;
      RECT 148.450000  67.585000 148.960000  67.915000 ;
      RECT 148.480000  87.150000 149.150000  87.320000 ;
      RECT 148.520000  61.505000 148.890000  67.585000 ;
      RECT 148.560000   8.850000 149.090000   9.020000 ;
      RECT 148.600000  42.840000 148.770000  44.180000 ;
      RECT 148.600000  68.385000 148.770000  68.885000 ;
      RECT 148.600000  68.885000 148.795000  71.015000 ;
      RECT 148.600000  71.015000 149.160000  71.185000 ;
      RECT 148.600000  71.185000 148.795000  73.345000 ;
      RECT 148.625000  73.345000 148.795000  73.635000 ;
      RECT 148.625000 112.085000 149.155000 112.255000 ;
      RECT 148.635000 112.000000 149.145000 112.085000 ;
      RECT 148.635000 112.255000 149.145000 112.330000 ;
      RECT 148.640000  30.285000 148.810000  36.025000 ;
      RECT 148.685000  22.015000 148.945000  22.655000 ;
      RECT 148.730000  19.530000 148.900000  22.015000 ;
      RECT 148.730000  22.655000 148.900000  24.280000 ;
      RECT 148.755000  17.235000 149.645000  17.615000 ;
      RECT 148.810000  77.010000 151.100000  77.180000 ;
      RECT 148.810000  77.180000 149.705000  79.150000 ;
      RECT 148.810000  79.150000 151.040000  79.320000 ;
      RECT 148.810000  79.320000 149.705000  81.250000 ;
      RECT 148.810000  81.250000 151.040000  81.300000 ;
      RECT 148.810000  81.300000 151.100000  81.470000 ;
      RECT 148.875000  15.140000 149.545000  15.310000 ;
      RECT 148.890000  46.165000 149.220000  47.015000 ;
      RECT 148.910000  29.785000 150.300000  30.085000 ;
      RECT 148.910000  30.085000 149.420000  30.115000 ;
      RECT 148.910000  36.195000 149.420000  36.225000 ;
      RECT 148.910000  36.225000 150.300000  36.525000 ;
      RECT 148.920000   5.035000 149.090000   8.850000 ;
      RECT 148.920000   9.020000 149.090000   9.785000 ;
      RECT 148.940000  68.205000 154.710000  68.555000 ;
      RECT 148.970000  47.015000 149.140000  47.625000 ;
      RECT 148.980000  30.115000 149.350000  36.195000 ;
      RECT 149.030000  42.840000 149.200000  44.010000 ;
      RECT 149.060000  61.675000 149.230000  62.725000 ;
      RECT 149.060000  62.955000 149.230000  63.285000 ;
      RECT 149.060000  63.905000 149.230000  64.235000 ;
      RECT 149.060000  64.405000 149.230000  67.115000 ;
      RECT 149.115000  37.870000 149.285000  40.870000 ;
      RECT 149.220000 200.085000 149.890000 200.255000 ;
      RECT 149.220000 216.235000 149.890000 216.405000 ;
      RECT 149.225000  81.890000 149.395000  86.640000 ;
      RECT 149.235000  72.535000 149.765000  72.705000 ;
      RECT 149.300000  42.470000 150.650000  42.475000 ;
      RECT 149.300000  42.475000 151.960000  42.645000 ;
      RECT 149.335000  41.360000 149.865000  41.530000 ;
      RECT 149.400000  61.175000 149.910000  61.285000 ;
      RECT 149.400000  61.285000 149.930000  61.455000 ;
      RECT 149.400000  61.455000 149.910000  61.505000 ;
      RECT 149.400000  67.585000 149.910000  67.915000 ;
      RECT 149.405000  68.555000 149.575000  72.535000 ;
      RECT 149.405000  72.705000 149.575000  73.635000 ;
      RECT 149.460000  42.840000 149.630000  44.180000 ;
      RECT 149.460000  44.180000 151.280000  44.350000 ;
      RECT 149.465000  20.875000 149.725000  21.515000 ;
      RECT 149.470000  61.505000 149.840000  67.585000 ;
      RECT 149.510000  19.530000 149.680000  20.875000 ;
      RECT 149.510000  21.515000 149.680000  24.280000 ;
      RECT 149.520000  30.285000 149.690000  31.895000 ;
      RECT 149.520000  32.515000 149.690000  35.725000 ;
      RECT 149.545000 243.890000 152.640000 244.175000 ;
      RECT 149.545000 244.175000 151.720000 246.535000 ;
      RECT 149.545000 246.535000 152.640000 246.935000 ;
      RECT 149.570000  44.580000 149.740000  45.760000 ;
      RECT 149.570000  45.930000 149.740000  47.080000 ;
      RECT 149.570000  47.370000 150.440000  48.380000 ;
      RECT 149.695000  37.840000 153.935000  38.010000 ;
      RECT 149.695000  38.010000 149.865000  41.360000 ;
      RECT 149.700000   4.685000 149.870000   9.785000 ;
      RECT 149.715000  87.150000 151.745000  87.320000 ;
      RECT 149.780000   9.960000 150.310000  10.130000 ;
      RECT 149.780000  10.130000 150.300000  10.965000 ;
      RECT 149.790000  30.085000 150.300000  30.115000 ;
      RECT 149.790000  36.195000 150.300000  36.225000 ;
      RECT 149.825000 113.195000 150.495000 113.525000 ;
      RECT 149.860000  30.115000 150.230000  36.195000 ;
      RECT 149.870000  15.350000 152.430000  18.455000 ;
      RECT 149.875000  77.400000 150.045000  78.750000 ;
      RECT 149.875000  79.540000 150.045000  81.080000 ;
      RECT 149.890000  42.840000 150.060000  44.010000 ;
      RECT 149.910000  46.335000 150.440000  47.370000 ;
      RECT 149.915000  83.290000 150.445000  83.460000 ;
      RECT 149.920000  37.335000 151.950000  37.505000 ;
      RECT 149.920000  60.665000 151.890000  60.835000 ;
      RECT 150.010000  61.675000 150.180000  66.135000 ;
      RECT 150.020000  71.015000 150.550000  71.185000 ;
      RECT 150.060000  14.655000 155.270000  14.825000 ;
      RECT 150.105000  81.890000 150.275000  83.290000 ;
      RECT 150.105000  83.460000 150.275000  86.640000 ;
      RECT 150.185000  68.885000 150.355000  71.015000 ;
      RECT 150.185000  71.185000 150.355000  73.635000 ;
      RECT 150.215000  77.180000 151.040000  79.150000 ;
      RECT 150.215000  79.320000 151.040000  81.250000 ;
      RECT 150.230000  25.475000 150.400000  27.495000 ;
      RECT 150.245000  22.015000 150.505000  22.655000 ;
      RECT 150.260000  67.115000 150.790000  67.285000 ;
      RECT 150.280000  61.175000 150.790000  61.505000 ;
      RECT 150.280000  67.585000 150.790000  67.915000 ;
      RECT 150.290000  19.530000 150.460000  22.015000 ;
      RECT 150.290000  22.655000 150.460000  24.280000 ;
      RECT 150.320000  42.840000 150.490000  44.180000 ;
      RECT 150.320000 200.495000 150.850000 215.995000 ;
      RECT 150.350000  61.505000 150.720000  67.115000 ;
      RECT 150.350000  67.285000 150.720000  67.585000 ;
      RECT 150.390000  45.280000 150.920000  45.450000 ;
      RECT 150.400000  30.285000 150.570000  36.025000 ;
      RECT 150.470000  10.860000 151.000000  11.030000 ;
      RECT 150.480000   5.035000 150.650000  10.295000 ;
      RECT 150.480000  10.295000 152.500000  10.465000 ;
      RECT 150.575000  38.180000 150.835000  41.160000 ;
      RECT 150.650000  10.855000 150.820000  10.860000 ;
      RECT 150.650000  11.030000 150.820000  14.185000 ;
      RECT 150.650000  14.185000 154.320000  14.355000 ;
      RECT 150.670000  29.785000 152.060000  30.085000 ;
      RECT 150.670000  30.085000 151.180000  30.115000 ;
      RECT 150.670000  36.195000 151.180000  36.225000 ;
      RECT 150.670000  36.225000 152.060000  36.525000 ;
      RECT 150.670000 239.105000 159.120000 239.275000 ;
      RECT 150.680000  24.970000 150.850000  26.470000 ;
      RECT 150.680000  26.470000 156.430000  26.640000 ;
      RECT 150.740000  30.115000 151.110000  36.195000 ;
      RECT 150.750000  42.840000 150.920000  44.010000 ;
      RECT 150.750000  44.580000 150.920000  45.280000 ;
      RECT 150.750000  45.450000 150.920000  47.080000 ;
      RECT 150.750000  47.370000 151.280000  48.550000 ;
      RECT 150.795000  72.535000 151.325000  72.705000 ;
      RECT 150.960000  61.675000 151.130000  62.725000 ;
      RECT 150.960000  62.955000 151.130000  63.285000 ;
      RECT 150.960000  63.905000 151.130000  64.235000 ;
      RECT 150.960000  64.405000 151.130000  67.420000 ;
      RECT 150.965000  68.555000 151.135000  72.535000 ;
      RECT 150.965000  72.705000 151.135000  73.635000 ;
      RECT 150.985000  81.890000 151.155000  86.640000 ;
      RECT 151.030000   5.035000 151.200000   8.850000 ;
      RECT 151.030000   8.850000 151.560000   9.020000 ;
      RECT 151.030000   9.020000 151.200000   9.785000 ;
      RECT 151.035000  38.180000 151.295000  41.160000 ;
      RECT 151.090000  43.095000 151.620000  43.265000 ;
      RECT 151.090000  44.350000 151.280000  47.370000 ;
      RECT 151.210000  41.360000 151.740000  41.530000 ;
      RECT 151.230000  10.795000 151.400000  11.360000 ;
      RECT 151.230000  11.360000 151.760000  11.530000 ;
      RECT 151.230000  11.530000 151.400000  13.505000 ;
      RECT 151.280000  30.285000 151.450000  31.895000 ;
      RECT 151.280000  32.515000 151.450000  35.725000 ;
      RECT 151.280000 200.085000 151.950000 200.255000 ;
      RECT 151.280000 216.235000 151.950000 216.405000 ;
      RECT 151.290000 199.685000 151.950000 200.085000 ;
      RECT 151.300000  19.565000 151.560000  20.600000 ;
      RECT 151.335000  79.120000 151.900000  79.290000 ;
      RECT 151.345000  19.080000 151.515000  19.565000 ;
      RECT 151.345000  20.600000 151.515000  25.870000 ;
      RECT 151.390000  41.530000 151.560000  42.305000 ;
      RECT 151.390000  79.075000 151.900000  79.120000 ;
      RECT 151.390000  79.290000 151.900000  79.405000 ;
      RECT 151.445000  78.240000 152.285000  78.410000 ;
      RECT 151.450000  43.265000 151.620000  48.390000 ;
      RECT 151.505000  83.290000 152.035000  83.460000 ;
      RECT 151.510000  61.675000 151.680000  63.695000 ;
      RECT 151.510000  63.695000 152.040000  63.865000 ;
      RECT 151.510000  63.865000 151.680000  67.115000 ;
      RECT 151.550000  30.085000 152.060000  30.115000 ;
      RECT 151.550000  36.195000 152.060000  36.225000 ;
      RECT 151.570000  18.650000 155.515000  18.820000 ;
      RECT 151.580000  71.015000 152.110000  71.185000 ;
      RECT 151.620000  30.115000 151.990000  36.195000 ;
      RECT 151.725000  22.940000 152.255000  23.110000 ;
      RECT 151.745000  68.885000 151.915000  71.015000 ;
      RECT 151.745000  71.185000 151.915000  73.635000 ;
      RECT 151.760000  61.255000 152.290000  61.425000 ;
      RECT 151.765000  18.820000 152.190000  22.940000 ;
      RECT 151.765000  23.110000 152.190000  26.185000 ;
      RECT 151.780000  61.175000 152.290000  61.255000 ;
      RECT 151.780000  61.425000 152.290000  61.505000 ;
      RECT 151.790000  42.645000 151.960000  43.405000 ;
      RECT 151.790000  43.405000 152.440000  44.415000 ;
      RECT 151.810000   5.035000 151.980000   9.220000 ;
      RECT 151.810000   9.220000 152.340000   9.390000 ;
      RECT 151.810000   9.390000 151.980000   9.785000 ;
      RECT 151.850000  61.505000 152.220000  61.885000 ;
      RECT 151.865000  74.420000 152.035000  76.020000 ;
      RECT 151.865000  77.400000 152.285000  78.240000 ;
      RECT 151.865000  78.410000 152.285000  78.750000 ;
      RECT 151.865000  79.730000 152.285000  81.080000 ;
      RECT 151.865000  81.890000 152.035000  83.290000 ;
      RECT 151.865000  83.460000 152.035000  86.640000 ;
      RECT 151.880000 113.910000 154.880000 164.900000 ;
      RECT 151.890000 244.345000 152.640000 246.365000 ;
      RECT 151.910000  41.290000 152.580000  41.460000 ;
      RECT 151.910000  46.335000 152.440000  46.505000 ;
      RECT 151.930000  47.855000 152.100000  48.465000 ;
      RECT 151.930000  48.465000 157.460000  48.635000 ;
      RECT 151.970000  42.030000 152.500000  42.200000 ;
      RECT 152.005000  38.180000 152.175000  41.290000 ;
      RECT 152.005000  41.460000 152.500000  42.030000 ;
      RECT 152.010000  10.795000 152.180000  14.185000 ;
      RECT 152.115000  78.750000 152.285000  79.730000 ;
      RECT 152.125000 106.360000 152.655000 106.530000 ;
      RECT 152.150000   9.590000 152.420000  10.295000 ;
      RECT 152.160000  30.285000 152.330000  36.025000 ;
      RECT 152.160000  37.335000 152.830000  37.505000 ;
      RECT 152.215000  60.665000 152.745000  60.835000 ;
      RECT 152.230000   8.850000 152.760000   9.020000 ;
      RECT 152.250000  36.975000 152.420000  37.335000 ;
      RECT 152.270000  44.415000 152.440000  46.335000 ;
      RECT 152.270000  46.505000 152.440000  48.085000 ;
      RECT 152.270000 244.175000 152.640000 244.345000 ;
      RECT 152.270000 246.365000 152.640000 246.535000 ;
      RECT 152.345000  87.070000 175.800000  87.700000 ;
      RECT 152.355000  72.535000 152.885000  72.705000 ;
      RECT 152.355000  81.950000 152.525000  87.070000 ;
      RECT 152.380000  23.495000 152.640000  25.000000 ;
      RECT 152.380000 200.495000 152.910000 215.995000 ;
      RECT 152.390000  61.675000 152.560000  62.685000 ;
      RECT 152.390000  62.955000 152.560000  63.285000 ;
      RECT 152.390000  63.905000 152.560000  64.235000 ;
      RECT 152.390000  64.405000 152.560000  67.115000 ;
      RECT 152.425000  19.080000 152.595000  23.495000 ;
      RECT 152.425000  25.000000 152.595000  25.870000 ;
      RECT 152.425000  36.195000 152.935000  36.225000 ;
      RECT 152.425000  36.225000 153.820000  36.525000 ;
      RECT 152.430000  11.360000 152.960000  11.530000 ;
      RECT 152.430000  29.785000 153.820000  30.085000 ;
      RECT 152.430000  30.085000 152.940000  30.115000 ;
      RECT 152.455000  74.400000 152.625000  81.020000 ;
      RECT 152.470000  67.515000 153.100000  67.585000 ;
      RECT 152.470000  67.585000 153.155000  67.685000 ;
      RECT 152.485000 105.375000 152.655000 106.360000 ;
      RECT 152.485000 106.530000 152.655000 106.725000 ;
      RECT 152.500000  30.115000 152.870000  36.195000 ;
      RECT 152.525000  68.555000 152.695000  72.535000 ;
      RECT 152.525000  72.705000 152.695000  73.635000 ;
      RECT 152.590000   5.035000 152.760000   8.850000 ;
      RECT 152.590000   9.020000 152.760000   9.785000 ;
      RECT 152.610000  45.000000 153.140000  45.170000 ;
      RECT 152.645000  67.685000 153.155000  67.915000 ;
      RECT 152.650000  61.255000 153.180000  61.425000 ;
      RECT 152.670000  41.635000 152.920000  42.305000 ;
      RECT 152.705000  41.580000 152.920000  41.635000 ;
      RECT 152.705000  42.305000 152.875000  43.405000 ;
      RECT 152.705000  43.405000 152.900000  44.415000 ;
      RECT 152.730000  45.170000 152.900000  48.085000 ;
      RECT 152.730000  61.175000 153.100000  61.255000 ;
      RECT 152.730000  61.425000 153.100000  67.515000 ;
      RECT 152.750000  38.180000 153.055000  40.890000 ;
      RECT 152.750000  40.890000 152.920000  41.580000 ;
      RECT 152.790000  10.015000 153.540000  10.185000 ;
      RECT 152.790000  10.185000 152.960000  11.360000 ;
      RECT 152.790000  11.530000 152.960000  13.505000 ;
      RECT 152.800000 239.550000 161.420000 241.240000 ;
      RECT 152.810000  15.225000 157.660000  15.395000 ;
      RECT 152.820000 242.090000 158.990000 243.700000 ;
      RECT 152.845000  18.820000 153.270000  26.185000 ;
      RECT 152.895000 104.700000 153.065000 107.450000 ;
      RECT 152.910000  16.505000 157.660000  16.675000 ;
      RECT 152.940000 242.030000 158.990000 242.090000 ;
      RECT 152.940000 243.700000 158.990000 243.720000 ;
      RECT 153.005000   9.220000 153.540000   9.390000 ;
      RECT 153.040000  30.285000 153.210000  31.895000 ;
      RECT 153.040000  32.515000 153.210000  35.725000 ;
      RECT 153.060000 244.355000 165.290000 247.105000 ;
      RECT 153.070000  42.400000 153.600000  42.570000 ;
      RECT 153.070000  42.570000 153.480000  44.585000 ;
      RECT 153.070000  44.585000 153.610000  44.740000 ;
      RECT 153.070000  45.375000 153.610000  45.665000 ;
      RECT 153.070000  45.665000 153.360000  48.085000 ;
      RECT 153.090000  42.030000 154.120000  42.200000 ;
      RECT 153.110000  37.335000 153.780000  37.505000 ;
      RECT 153.140000  71.015000 153.670000  71.185000 ;
      RECT 153.170000  60.665000 156.280000  60.835000 ;
      RECT 153.190000  41.290000 153.935000  41.460000 ;
      RECT 153.205000  75.275000 170.475000  75.525000 ;
      RECT 153.205000  75.525000 153.375000  79.145000 ;
      RECT 153.260000  41.460000 153.790000  41.530000 ;
      RECT 153.270000  64.405000 153.440000  67.115000 ;
      RECT 153.305000  68.885000 153.475000  71.015000 ;
      RECT 153.305000  71.185000 153.475000  73.635000 ;
      RECT 153.310000  30.085000 153.820000  30.115000 ;
      RECT 153.310000  36.195000 153.820000  36.225000 ;
      RECT 153.310000  44.740000 153.610000  45.375000 ;
      RECT 153.370000   5.035000 153.540000   9.220000 ;
      RECT 153.370000   9.390000 153.540000  10.015000 ;
      RECT 153.375000  80.895000 154.045000  81.065000 ;
      RECT 153.380000  30.115000 153.750000  36.195000 ;
      RECT 153.395000  74.255000 159.835000  74.505000 ;
      RECT 153.420000 199.125000 157.330000 217.365000 ;
      RECT 153.435000  80.800000 153.965000  80.895000 ;
      RECT 153.435000  81.285000 153.605000  86.270000 ;
      RECT 153.440000  80.145000 153.745000  80.475000 ;
      RECT 153.450000  63.415000 153.980000  63.585000 ;
      RECT 153.460000  19.565000 153.720000  20.600000 ;
      RECT 153.505000  19.080000 153.675000  19.565000 ;
      RECT 153.505000  20.600000 153.675000  25.870000 ;
      RECT 153.535000  67.585000 154.045000  67.915000 ;
      RECT 153.545000  79.140000 154.745000  79.370000 ;
      RECT 153.545000  79.370000 153.745000  80.145000 ;
      RECT 153.560000  48.105000 154.315000  48.275000 ;
      RECT 153.570000  10.795000 153.740000  14.185000 ;
      RECT 153.610000  63.585000 153.980000  67.585000 ;
      RECT 153.650000  43.405000 153.820000  44.415000 ;
      RECT 153.765000  38.010000 153.935000  41.290000 ;
      RECT 153.785000  46.335000 154.315000  46.505000 ;
      RECT 153.790000   8.850000 154.320000   9.020000 ;
      RECT 153.795000  75.775000 155.200000  75.945000 ;
      RECT 153.795000  75.945000 153.965000  78.350000 ;
      RECT 153.795000  78.350000 154.325000  78.520000 ;
      RECT 153.795000  78.520000 153.965000  78.875000 ;
      RECT 153.805000  44.630000 153.975000  45.300000 ;
      RECT 153.830000 103.770000 166.055000 108.380000 ;
      RECT 153.845000  42.510000 154.380000  43.085000 ;
      RECT 153.910000  10.860000 154.440000  11.030000 ;
      RECT 153.915000  72.535000 154.445000  72.705000 ;
      RECT 153.920000  30.285000 154.090000  36.025000 ;
      RECT 153.950000  41.635000 154.120000  42.030000 ;
      RECT 153.950000  42.200000 154.120000  42.305000 ;
      RECT 154.085000  68.555000 154.255000  72.535000 ;
      RECT 154.085000  72.705000 154.255000  73.635000 ;
      RECT 154.110000  43.405000 154.315000  44.415000 ;
      RECT 154.145000  44.415000 154.315000  46.335000 ;
      RECT 154.145000  46.505000 154.315000  48.105000 ;
      RECT 154.150000   5.035000 154.320000   8.850000 ;
      RECT 154.150000   9.020000 154.320000   9.785000 ;
      RECT 154.150000  10.855000 154.320000  10.860000 ;
      RECT 154.150000  11.030000 154.320000  14.185000 ;
      RECT 154.150000  61.675000 154.320000  65.585000 ;
      RECT 154.150000  65.585000 154.680000  65.755000 ;
      RECT 154.150000  65.755000 154.320000  67.420000 ;
      RECT 154.190000  29.785000 154.700000  30.115000 ;
      RECT 154.190000  36.195000 154.700000  36.525000 ;
      RECT 154.215000  79.620000 156.305000  79.790000 ;
      RECT 154.215000  79.790000 154.385000  86.035000 ;
      RECT 154.260000  30.115000 154.630000  36.195000 ;
      RECT 154.280000  96.030000 190.275000  96.880000 ;
      RECT 154.280000  96.880000 190.270000  97.045000 ;
      RECT 154.280000  97.045000 166.055000 102.920000 ;
      RECT 154.410000  61.255000 154.940000  61.425000 ;
      RECT 154.420000  61.175000 154.930000  61.255000 ;
      RECT 154.420000  61.425000 154.930000  61.505000 ;
      RECT 154.490000  61.505000 154.860000  61.880000 ;
      RECT 154.490000  63.455000 154.820000  63.695000 ;
      RECT 154.490000  63.695000 155.020000  63.865000 ;
      RECT 154.490000  63.865000 154.820000  63.965000 ;
      RECT 154.510000  71.015000 155.040000  71.185000 ;
      RECT 154.540000  23.495000 154.800000  25.000000 ;
      RECT 154.555000  80.895000 155.225000  81.065000 ;
      RECT 154.575000  76.165000 154.745000  79.140000 ;
      RECT 154.585000  19.080000 154.755000  23.495000 ;
      RECT 154.585000  25.000000 154.755000  25.870000 ;
      RECT 154.595000  58.725000 154.780000  59.255000 ;
      RECT 154.610000  37.870000 154.780000  44.425000 ;
      RECT 154.610000  45.065000 154.780000  48.465000 ;
      RECT 154.610000  49.535000 157.460000  49.705000 ;
      RECT 154.610000  49.705000 154.780000  52.000000 ;
      RECT 154.610000  52.610000 154.780000  58.725000 ;
      RECT 154.610000  59.255000 154.780000  60.320000 ;
      RECT 154.635000  80.800000 155.165000  80.895000 ;
      RECT 154.730000   4.685000 154.900000  10.055000 ;
      RECT 154.760000 192.620000 158.850000 192.950000 ;
      RECT 154.800000  30.285000 155.665000  31.565000 ;
      RECT 154.800000  31.565000 156.025000  31.735000 ;
      RECT 154.800000  31.735000 155.665000  31.795000 ;
      RECT 154.800000  31.795000 154.970000  31.895000 ;
      RECT 154.800000  32.515000 155.665000  35.725000 ;
      RECT 154.865000  68.885000 155.035000  71.015000 ;
      RECT 154.865000  71.185000 155.035000  73.635000 ;
      RECT 154.995000  81.285000 155.165000  86.270000 ;
      RECT 155.010000  42.510000 155.545000  43.085000 ;
      RECT 155.010000  55.085000 155.545000  55.660000 ;
      RECT 155.030000  64.405000 155.200000  67.115000 ;
      RECT 155.075000  43.405000 155.280000  44.415000 ;
      RECT 155.075000  44.415000 155.245000  46.335000 ;
      RECT 155.075000  46.335000 155.605000  46.505000 ;
      RECT 155.075000  46.505000 155.245000  48.105000 ;
      RECT 155.075000  48.105000 155.830000  48.275000 ;
      RECT 155.075000  49.895000 155.830000  50.065000 ;
      RECT 155.075000  50.065000 155.245000  51.665000 ;
      RECT 155.075000  51.665000 155.605000  51.835000 ;
      RECT 155.075000  51.835000 155.245000  53.755000 ;
      RECT 155.075000  53.755000 155.280000  54.765000 ;
      RECT 155.170000  78.350000 155.700000  78.520000 ;
      RECT 155.270000  41.635000 155.440000  42.030000 ;
      RECT 155.270000  42.030000 156.300000  42.200000 ;
      RECT 155.270000  42.200000 155.440000  42.305000 ;
      RECT 155.270000  55.865000 155.440000  55.970000 ;
      RECT 155.270000  55.970000 156.300000  56.140000 ;
      RECT 155.270000  56.140000 155.440000  56.535000 ;
      RECT 155.300000  61.175000 155.810000  61.285000 ;
      RECT 155.300000  61.285000 155.835000  61.455000 ;
      RECT 155.300000  61.455000 155.810000  61.505000 ;
      RECT 155.315000  67.585000 155.825000  67.915000 ;
      RECT 155.355000  68.635000 156.015000  71.415000 ;
      RECT 155.355000  71.415000 156.250000  72.305000 ;
      RECT 155.355000  72.305000 156.015000  74.255000 ;
      RECT 155.355000  76.165000 155.525000  78.350000 ;
      RECT 155.355000  78.520000 155.525000  78.875000 ;
      RECT 155.370000  61.505000 155.740000  67.585000 ;
      RECT 155.415000  44.630000 155.585000  45.300000 ;
      RECT 155.415000  52.870000 155.585000  53.540000 ;
      RECT 155.455000  37.840000 159.695000  38.010000 ;
      RECT 155.455000  38.010000 155.625000  41.290000 ;
      RECT 155.455000  41.290000 156.200000  41.460000 ;
      RECT 155.455000  56.710000 156.200000  56.880000 ;
      RECT 155.455000  56.880000 155.625000  60.160000 ;
      RECT 155.455000  60.160000 159.695000  60.330000 ;
      RECT 155.495000  35.725000 155.665000  36.025000 ;
      RECT 155.530000  84.545000 159.070000  84.560000 ;
      RECT 155.530000  84.560000 158.240000  84.715000 ;
      RECT 155.545000  84.380000 159.070000  84.545000 ;
      RECT 155.570000  43.405000 155.740000  44.415000 ;
      RECT 155.570000  53.755000 155.740000  54.765000 ;
      RECT 155.600000  41.460000 156.130000  41.530000 ;
      RECT 155.600000  56.640000 156.130000  56.710000 ;
      RECT 155.610000  37.335000 156.280000  37.505000 ;
      RECT 155.620000  22.010000 155.880000  22.655000 ;
      RECT 155.665000  19.080000 155.835000  22.010000 ;
      RECT 155.665000  22.655000 155.835000  25.870000 ;
      RECT 155.725000  86.210000 170.705000  86.320000 ;
      RECT 155.725000  86.320000 170.730000  86.375000 ;
      RECT 155.725000  86.375000 175.800000  86.380000 ;
      RECT 155.740000  86.380000 175.800000  87.070000 ;
      RECT 155.750000  75.775000 156.760000  75.945000 ;
      RECT 155.780000  44.585000 156.320000  44.740000 ;
      RECT 155.780000  44.740000 156.080000  45.375000 ;
      RECT 155.780000  45.375000 156.320000  45.665000 ;
      RECT 155.780000  52.505000 156.320000  52.795000 ;
      RECT 155.780000  52.795000 156.080000  53.430000 ;
      RECT 155.780000  53.430000 156.320000  53.585000 ;
      RECT 155.780000  85.025000 158.150000  86.210000 ;
      RECT 155.790000  42.400000 156.320000  42.570000 ;
      RECT 155.790000  55.600000 156.320000  55.770000 ;
      RECT 155.895000 180.175000 158.850000 183.525000 ;
      RECT 155.895000 184.375000 158.850000 188.010000 ;
      RECT 155.895000 188.860000 158.850000 192.620000 ;
      RECT 155.895000 192.950000 158.850000 193.515000 ;
      RECT 155.910000  42.570000 156.320000  44.585000 ;
      RECT 155.910000  53.585000 156.320000  55.600000 ;
      RECT 155.910000  61.675000 156.080000  62.725000 ;
      RECT 155.910000  62.955000 156.080000  63.285000 ;
      RECT 155.910000  63.905000 156.080000  64.235000 ;
      RECT 155.910000  64.405000 156.080000  67.115000 ;
      RECT 156.010000  80.770000 156.540000  80.940000 ;
      RECT 156.010000  80.940000 156.180000  83.995000 ;
      RECT 156.030000  45.665000 156.320000  48.085000 ;
      RECT 156.030000  50.085000 156.320000  52.505000 ;
      RECT 156.135000  75.945000 156.305000  79.620000 ;
      RECT 156.160000  68.205000 161.930000  68.525000 ;
      RECT 156.250000  45.000000 156.780000  45.170000 ;
      RECT 156.250000  53.000000 156.780000  53.170000 ;
      RECT 156.260000  19.055000 156.430000  26.470000 ;
      RECT 156.285000 113.195000 156.955000 113.525000 ;
      RECT 156.335000  38.180000 156.640000  40.890000 ;
      RECT 156.335000  57.280000 156.640000  59.990000 ;
      RECT 156.390000 113.910000 159.390000 164.900000 ;
      RECT 156.430000  63.415000 156.960000  63.585000 ;
      RECT 156.460000  71.015000 156.990000  71.185000 ;
      RECT 156.470000  40.890000 156.640000  41.580000 ;
      RECT 156.470000  41.580000 156.685000  41.635000 ;
      RECT 156.470000  41.635000 156.720000  42.305000 ;
      RECT 156.470000  55.865000 156.720000  56.535000 ;
      RECT 156.470000  56.535000 156.685000  56.590000 ;
      RECT 156.470000  56.590000 156.640000  57.280000 ;
      RECT 156.490000  43.405000 156.685000  44.415000 ;
      RECT 156.490000  45.170000 156.660000  48.085000 ;
      RECT 156.490000  50.085000 156.660000  53.000000 ;
      RECT 156.490000  53.755000 156.685000  54.765000 ;
      RECT 156.515000  42.305000 156.685000  43.405000 ;
      RECT 156.515000  54.765000 156.685000  55.865000 ;
      RECT 156.555000  78.350000 157.085000  78.520000 ;
      RECT 156.560000  37.335000 157.230000  37.505000 ;
      RECT 156.560000  60.665000 157.230000  60.835000 ;
      RECT 156.625000  68.885000 156.795000  71.015000 ;
      RECT 156.625000  71.185000 156.795000  73.635000 ;
      RECT 156.790000  61.675000 156.960000  63.415000 ;
      RECT 156.790000  63.585000 156.960000  67.115000 ;
      RECT 156.790000  81.285000 156.960000  83.995000 ;
      RECT 156.810000  41.290000 157.480000  41.460000 ;
      RECT 156.810000  56.710000 157.480000  56.880000 ;
      RECT 156.890000  41.460000 157.385000  42.030000 ;
      RECT 156.890000  42.030000 157.420000  42.200000 ;
      RECT 156.890000  55.970000 157.420000  56.140000 ;
      RECT 156.890000  56.140000 157.385000  56.710000 ;
      RECT 156.915000  76.165000 157.085000  78.350000 ;
      RECT 156.915000  78.520000 157.085000  78.875000 ;
      RECT 156.950000  43.405000 157.600000  44.415000 ;
      RECT 156.950000  44.415000 157.120000  46.335000 ;
      RECT 156.950000  46.335000 157.480000  46.505000 ;
      RECT 156.950000  46.505000 157.120000  48.085000 ;
      RECT 156.950000  50.085000 157.120000  51.665000 ;
      RECT 156.950000  51.665000 157.480000  51.835000 ;
      RECT 156.950000  51.835000 157.120000  53.755000 ;
      RECT 156.950000  53.755000 157.600000  54.765000 ;
      RECT 157.060000  29.405000 160.450000  30.145000 ;
      RECT 157.060000  30.145000 161.030000  31.535000 ;
      RECT 157.060000  31.535000 159.170000  31.735000 ;
      RECT 157.060000  31.735000 158.470000  32.785000 ;
      RECT 157.060000  32.785000 157.570000  35.945000 ;
      RECT 157.060000  35.945000 168.445000  36.455000 ;
      RECT 157.060000  79.140000 157.635000  79.310000 ;
      RECT 157.215000  38.180000 157.385000  41.290000 ;
      RECT 157.215000  56.880000 157.385000  59.990000 ;
      RECT 157.290000  47.855000 157.460000  48.465000 ;
      RECT 157.290000  49.705000 157.460000  50.315000 ;
      RECT 157.340000  61.675000 157.510000  63.415000 ;
      RECT 157.340000  63.415000 157.870000  63.585000 ;
      RECT 157.340000  63.585000 157.510000  67.115000 ;
      RECT 157.385000  80.770000 157.915000  80.940000 ;
      RECT 157.405000  68.885000 157.575000  74.255000 ;
      RECT 157.430000  42.475000 160.090000  42.645000 ;
      RECT 157.430000  42.645000 157.600000  43.405000 ;
      RECT 157.430000  54.765000 157.600000  55.525000 ;
      RECT 157.430000  55.525000 160.090000  55.695000 ;
      RECT 157.440000  37.335000 159.470000  37.505000 ;
      RECT 157.440000  60.665000 159.470000  60.835000 ;
      RECT 157.465000  76.165000 157.635000  79.140000 ;
      RECT 157.570000  80.940000 157.740000  83.995000 ;
      RECT 157.650000  41.360000 158.180000  41.530000 ;
      RECT 157.650000  56.640000 158.180000  56.810000 ;
      RECT 157.770000  43.095000 158.300000  43.265000 ;
      RECT 157.770000  43.265000 157.940000  48.390000 ;
      RECT 157.770000  49.780000 157.940000  54.905000 ;
      RECT 157.770000  54.905000 158.300000  55.075000 ;
      RECT 157.830000  41.530000 158.000000  42.305000 ;
      RECT 157.830000  55.865000 158.000000  56.640000 ;
      RECT 157.845000  75.775000 158.855000  75.945000 ;
      RECT 158.015000  71.015000 158.545000  71.185000 ;
      RECT 158.075000   3.840000 160.095000   4.590000 ;
      RECT 158.075000  14.420000 160.095000  15.170000 ;
      RECT 158.095000  38.180000 158.355000  41.160000 ;
      RECT 158.095000  57.010000 158.355000  59.990000 ;
      RECT 158.110000  44.180000 159.930000  44.350000 ;
      RECT 158.110000  44.350000 158.300000  47.370000 ;
      RECT 158.110000  47.370000 158.640000  48.550000 ;
      RECT 158.110000  48.550000 161.000000  48.720000 ;
      RECT 158.110000  49.450000 161.000000  49.620000 ;
      RECT 158.110000  49.620000 158.640000  50.800000 ;
      RECT 158.110000  50.800000 158.300000  53.820000 ;
      RECT 158.110000  53.820000 159.930000  53.990000 ;
      RECT 158.185000  68.885000 158.355000  71.015000 ;
      RECT 158.185000  71.185000 158.355000  73.635000 ;
      RECT 158.220000  35.165000 166.795000  35.335000 ;
      RECT 158.220000  61.675000 158.390000  62.725000 ;
      RECT 158.220000  62.955000 158.390000  63.285000 ;
      RECT 158.220000  63.905000 158.390000  64.235000 ;
      RECT 158.220000  64.405000 158.390000  67.115000 ;
      RECT 158.245000  76.165000 158.415000  78.875000 ;
      RECT 158.300000  33.860000 158.470000  34.915000 ;
      RECT 158.330000 197.275000 159.180000 209.275000 ;
      RECT 158.330000 209.275000 159.930000 214.785000 ;
      RECT 158.330000 214.785000 164.210000 218.740000 ;
      RECT 158.330000 218.740000 172.950000 219.215000 ;
      RECT 158.350000  80.695000 161.400000  80.865000 ;
      RECT 158.350000  80.865000 158.520000  83.995000 ;
      RECT 158.470000  42.840000 158.640000  44.010000 ;
      RECT 158.470000  44.580000 158.640000  45.280000 ;
      RECT 158.470000  45.280000 159.000000  45.450000 ;
      RECT 158.470000  45.450000 158.640000  47.080000 ;
      RECT 158.470000  51.090000 158.640000  52.720000 ;
      RECT 158.470000  52.720000 159.000000  52.890000 ;
      RECT 158.470000  52.890000 158.640000  53.590000 ;
      RECT 158.470000  54.160000 158.640000  55.330000 ;
      RECT 158.470000  61.285000 159.000000  61.455000 ;
      RECT 158.475000  67.585000 158.985000  67.915000 ;
      RECT 158.480000  84.780000 159.070000  84.950000 ;
      RECT 158.490000  61.175000 159.000000  61.285000 ;
      RECT 158.490000  61.455000 159.000000  61.505000 ;
      RECT 158.555000  38.180000 158.815000  41.160000 ;
      RECT 158.555000  57.010000 158.815000  59.990000 ;
      RECT 158.560000  61.505000 158.930000  67.585000 ;
      RECT 158.585000  78.265000 159.195000  78.435000 ;
      RECT 158.740000  42.470000 160.090000  42.475000 ;
      RECT 158.740000  55.695000 160.090000  55.700000 ;
      RECT 158.845000 113.195000 159.515000 113.525000 ;
      RECT 158.900000  42.840000 159.070000  44.180000 ;
      RECT 158.900000  53.990000 159.070000  55.330000 ;
      RECT 158.900000  81.285000 159.070000  84.380000 ;
      RECT 158.900000  84.950000 159.070000  85.465000 ;
      RECT 158.950000  46.335000 159.480000  47.370000 ;
      RECT 158.950000  47.370000 159.820000  48.380000 ;
      RECT 158.950000  49.790000 159.820000  50.800000 ;
      RECT 158.950000  50.800000 159.480000  51.835000 ;
      RECT 158.965000  68.885000 159.135000  74.255000 ;
      RECT 159.025000  76.165000 159.195000  78.265000 ;
      RECT 159.025000  78.435000 159.195000  78.875000 ;
      RECT 159.100000  64.405000 159.270000  67.115000 ;
      RECT 159.105000  75.785000 159.835000  75.870000 ;
      RECT 159.105000  75.870000 159.635000  75.955000 ;
      RECT 159.165000  75.700000 159.835000  75.785000 ;
      RECT 159.240000  84.465000 159.850000  84.795000 ;
      RECT 159.280000  63.695000 159.810000  63.865000 ;
      RECT 159.330000  42.840000 159.500000  44.010000 ;
      RECT 159.330000  54.160000 159.500000  55.330000 ;
      RECT 159.335000 112.085000 159.865000 112.255000 ;
      RECT 159.345000 112.000000 159.855000 112.085000 ;
      RECT 159.345000 112.255000 159.855000 112.330000 ;
      RECT 159.350000 208.205000 160.075000 208.735000 ;
      RECT 159.360000  61.255000 159.890000  61.425000 ;
      RECT 159.370000  61.175000 159.880000  61.255000 ;
      RECT 159.370000  61.425000 159.880000  61.505000 ;
      RECT 159.440000  61.505000 159.810000  61.880000 ;
      RECT 159.480000  63.455000 159.810000  63.695000 ;
      RECT 159.480000  63.865000 159.810000  63.965000 ;
      RECT 159.525000  38.010000 159.695000  41.360000 ;
      RECT 159.525000  41.360000 160.055000  41.530000 ;
      RECT 159.525000  56.640000 160.055000  56.810000 ;
      RECT 159.525000  56.810000 159.695000  60.160000 ;
      RECT 159.545000  71.015000 160.075000  71.185000 ;
      RECT 159.580000  31.775000 159.750000  34.915000 ;
      RECT 159.620000  65.585000 160.150000  65.755000 ;
      RECT 159.650000  44.580000 159.820000  45.760000 ;
      RECT 159.650000  45.760000 162.180000  45.930000 ;
      RECT 159.650000  45.930000 159.820000  47.080000 ;
      RECT 159.650000  51.090000 159.820000  52.240000 ;
      RECT 159.650000  52.240000 162.180000  52.410000 ;
      RECT 159.650000  52.410000 159.820000  53.590000 ;
      RECT 159.680000  81.285000 159.850000  84.010000 ;
      RECT 159.680000  84.010000 160.210000  84.180000 ;
      RECT 159.680000  84.180000 159.850000  84.465000 ;
      RECT 159.745000  68.885000 159.915000  71.015000 ;
      RECT 159.745000  71.185000 159.915000  73.635000 ;
      RECT 159.745000 197.515000 160.075000 198.485000 ;
      RECT 159.745000 198.485000 160.860000 198.655000 ;
      RECT 159.760000  42.840000 159.930000  44.180000 ;
      RECT 159.760000  53.990000 159.930000  55.330000 ;
      RECT 159.805000  76.165000 159.975000  78.875000 ;
      RECT 159.920000  31.535000 161.030000  31.735000 ;
      RECT 159.920000  33.255000 161.950000  33.425000 ;
      RECT 159.950000 178.905000 160.800000 196.425000 ;
      RECT 159.980000  61.675000 160.150000  65.585000 ;
      RECT 159.980000  65.755000 160.150000  67.420000 ;
      RECT 160.090000  79.250000 162.800000  79.595000 ;
      RECT 160.105000  37.870000 160.275000  40.870000 ;
      RECT 160.105000  57.300000 160.275000  60.300000 ;
      RECT 160.105000  79.140000 162.795000  79.250000 ;
      RECT 160.170000  46.165000 160.500000  47.015000 ;
      RECT 160.170000  51.155000 160.500000  52.005000 ;
      RECT 160.190000  42.840000 160.360000  44.010000 ;
      RECT 160.190000  54.160000 160.360000  55.330000 ;
      RECT 160.230000  80.865000 160.760000  83.070000 ;
      RECT 160.245000  68.885000 160.695000  71.415000 ;
      RECT 160.245000  71.415000 160.805000  72.305000 ;
      RECT 160.245000  72.305000 160.695000  74.515000 ;
      RECT 160.245000  74.515000 160.415000  74.525000 ;
      RECT 160.250000  47.015000 160.420000  47.625000 ;
      RECT 160.250000  50.545000 160.420000  51.155000 ;
      RECT 160.255000  67.585000 160.765000  67.915000 ;
      RECT 160.315000  84.745000 167.105000  84.915000 ;
      RECT 160.320000  63.415000 160.850000  63.585000 ;
      RECT 160.320000  63.585000 160.690000  67.585000 ;
      RECT 160.325000  45.280000 161.000000  45.450000 ;
      RECT 160.325000  52.720000 161.000000  52.890000 ;
      RECT 160.395000  78.340000 160.925000  78.510000 ;
      RECT 160.445000  42.470000 161.795000  42.640000 ;
      RECT 160.445000  42.640000 161.695000  42.670000 ;
      RECT 160.445000  55.500000 161.695000  55.530000 ;
      RECT 160.445000  55.530000 161.795000  55.700000 ;
      RECT 160.585000  76.165000 160.755000  78.340000 ;
      RECT 160.585000  78.510000 160.755000  78.875000 ;
      RECT 160.590000  74.745000 168.400000  74.915000 ;
      RECT 160.620000  42.840000 160.790000  44.180000 ;
      RECT 160.620000  44.180000 162.180000  44.350000 ;
      RECT 160.620000  53.820000 162.180000  53.990000 ;
      RECT 160.620000  53.990000 160.790000  55.330000 ;
      RECT 160.690000 198.065000 171.340000 198.235000 ;
      RECT 160.690000 198.235000 160.860000 198.485000 ;
      RECT 160.690000 198.655000 160.860000 213.855000 ;
      RECT 160.690000 213.855000 165.140000 214.025000 ;
      RECT 160.695000  83.290000 163.025000  83.460000 ;
      RECT 160.755000  83.460000 163.025000  84.745000 ;
      RECT 160.830000  44.580000 161.000000  45.280000 ;
      RECT 160.830000  45.450000 161.000000  45.590000 ;
      RECT 160.830000  46.100000 161.000000  48.550000 ;
      RECT 160.830000  49.620000 161.000000  52.070000 ;
      RECT 160.830000  52.580000 161.000000  52.720000 ;
      RECT 160.830000  52.890000 161.000000  53.590000 ;
      RECT 160.860000  31.735000 161.030000  32.855000 ;
      RECT 160.860000  33.860000 161.030000  34.915000 ;
      RECT 160.860000  64.405000 161.030000  67.115000 ;
      RECT 160.900000 113.910000 163.900000 164.900000 ;
      RECT 161.020000   5.035000 174.910000   5.735000 ;
      RECT 161.020000   5.735000 161.720000  15.795000 ;
      RECT 161.020000  15.795000 174.910000  16.495000 ;
      RECT 161.020000  16.495000 161.720000  26.555000 ;
      RECT 161.020000  26.555000 174.910000  27.255000 ;
      RECT 161.050000  42.840000 161.220000  44.010000 ;
      RECT 161.050000  54.160000 161.220000  55.330000 ;
      RECT 161.120000  61.255000 161.650000  61.425000 ;
      RECT 161.135000  71.015000 161.665000  71.185000 ;
      RECT 161.145000  67.585000 161.655000  67.915000 ;
      RECT 161.200000  61.175000 161.570000  61.255000 ;
      RECT 161.200000  61.425000 161.570000  67.585000 ;
      RECT 161.270000 198.815000 161.440000 205.605000 ;
      RECT 161.270000 206.465000 161.440000 213.255000 ;
      RECT 161.275000  29.420000 161.945000  29.590000 ;
      RECT 161.305000  68.885000 161.475000  71.015000 ;
      RECT 161.305000  71.185000 161.475000  73.635000 ;
      RECT 161.310000  81.770000 161.840000  81.940000 ;
      RECT 161.310000  81.940000 161.480000  83.060000 ;
      RECT 161.335000  29.590000 161.865000  30.115000 ;
      RECT 161.365000  76.165000 161.535000  78.875000 ;
      RECT 161.385000 242.030000 163.790000 243.720000 ;
      RECT 161.450000  37.765000 161.620000  40.845000 ;
      RECT 161.450000  57.325000 161.620000  60.405000 ;
      RECT 161.480000  42.840000 161.650000  44.180000 ;
      RECT 161.480000  53.990000 161.650000  55.330000 ;
      RECT 161.560000 198.425000 164.270000 198.595000 ;
      RECT 161.560000 205.815000 164.270000 206.245000 ;
      RECT 161.610000 198.595000 161.880000 205.815000 ;
      RECT 161.650000  46.335000 162.180000  46.505000 ;
      RECT 161.650000  51.665000 162.180000  51.835000 ;
      RECT 161.720000  79.900000 161.890000  80.475000 ;
      RECT 161.740000  61.675000 161.910000  62.685000 ;
      RECT 161.740000  62.955000 161.910000  63.285000 ;
      RECT 161.740000  63.905000 161.910000  64.235000 ;
      RECT 161.740000  64.405000 161.910000  67.115000 ;
      RECT 161.775000  41.265000 162.740000  41.435000 ;
      RECT 161.775000  41.435000 162.085000  42.130000 ;
      RECT 161.775000  42.130000 162.305000  42.300000 ;
      RECT 161.775000  55.870000 162.305000  56.040000 ;
      RECT 161.775000  56.040000 162.085000  56.735000 ;
      RECT 161.775000  56.735000 162.740000  56.905000 ;
      RECT 161.840000   0.710000 168.030000   0.880000 ;
      RECT 161.840000   0.880000 162.010000   5.035000 ;
      RECT 161.855000  71.415000 162.745000  72.305000 ;
      RECT 161.910000  42.840000 162.080000  44.010000 ;
      RECT 161.910000  54.160000 162.080000  55.330000 ;
      RECT 161.915000  38.155000 162.200000  40.865000 ;
      RECT 161.915000  40.865000 162.085000  41.095000 ;
      RECT 161.915000  57.075000 162.085000  57.305000 ;
      RECT 161.915000  57.305000 162.200000  60.015000 ;
      RECT 161.965000 239.550000 163.790000 241.160000 ;
      RECT 161.990000  32.885000 162.520000  33.055000 ;
      RECT 162.010000  44.350000 162.180000  45.760000 ;
      RECT 162.010000  46.100000 162.180000  46.335000 ;
      RECT 162.010000  46.505000 162.180000  48.380000 ;
      RECT 162.010000  49.790000 162.180000  51.665000 ;
      RECT 162.010000  51.835000 162.180000  52.070000 ;
      RECT 162.010000  52.410000 162.180000  53.820000 ;
      RECT 162.010000  61.175000 162.520000  61.255000 ;
      RECT 162.010000  61.255000 162.540000  61.425000 ;
      RECT 162.010000  61.425000 162.520000  61.505000 ;
      RECT 162.025000  67.885000 162.555000  68.055000 ;
      RECT 162.040000 176.145000 162.890000 194.305000 ;
      RECT 162.040000 194.305000 175.920000 195.155000 ;
      RECT 162.050000 198.815000 162.220000 205.605000 ;
      RECT 162.050000 206.465000 162.220000 213.255000 ;
      RECT 162.080000  61.505000 162.450000  61.885000 ;
      RECT 162.080000  66.015000 162.450000  67.885000 ;
      RECT 162.085000  68.885000 162.255000  71.415000 ;
      RECT 162.085000  72.305000 162.255000  73.635000 ;
      RECT 162.130000  80.695000 165.520000  80.790000 ;
      RECT 162.130000  80.790000 166.720000  80.960000 ;
      RECT 162.130000  80.960000 165.520000  81.205000 ;
      RECT 162.130000  81.430000 164.840000  81.600000 ;
      RECT 162.135000 241.160000 163.790000 241.240000 ;
      RECT 162.140000  30.145000 162.310000  32.885000 ;
      RECT 162.140000  33.055000 162.310000  34.915000 ;
      RECT 162.145000  76.165000 162.315000  78.340000 ;
      RECT 162.145000  78.340000 162.675000  78.510000 ;
      RECT 162.145000  78.510000 162.315000  78.875000 ;
      RECT 162.255000  37.335000 164.510000  37.505000 ;
      RECT 162.255000  41.085000 162.925000  41.255000 ;
      RECT 162.255000  41.255000 162.740000  41.265000 ;
      RECT 162.255000  41.760000 162.785000  41.930000 ;
      RECT 162.255000  56.240000 162.785000  56.410000 ;
      RECT 162.255000  56.905000 162.740000  56.915000 ;
      RECT 162.255000  56.915000 162.925000  57.085000 ;
      RECT 162.255000  60.665000 164.510000  60.835000 ;
      RECT 162.260000  63.695000 162.790000  63.865000 ;
      RECT 162.370000  37.505000 164.510000  37.595000 ;
      RECT 162.370000  37.595000 162.740000  41.085000 ;
      RECT 162.370000  43.110000 162.900000  48.390000 ;
      RECT 162.370000  54.890000 162.900000  55.060000 ;
      RECT 162.370000  57.085000 162.740000  60.575000 ;
      RECT 162.370000  60.575000 164.510000  60.665000 ;
      RECT 162.390000  82.050000 162.560000  83.060000 ;
      RECT 162.390000 198.595000 162.660000 205.815000 ;
      RECT 162.400000 232.550000 162.765000 238.030000 ;
      RECT 162.475000  41.930000 162.785000  43.110000 ;
      RECT 162.475000  55.060000 162.785000  56.240000 ;
      RECT 162.480000   6.495000 166.855000   7.195000 ;
      RECT 162.480000   7.195000 163.180000  14.325000 ;
      RECT 162.480000  14.325000 166.855000  15.035000 ;
      RECT 162.480000  17.255000 166.855000  17.965000 ;
      RECT 162.480000  17.965000 163.180000  25.095000 ;
      RECT 162.480000  25.095000 166.855000  25.795000 ;
      RECT 162.500000 221.910000 162.755000 230.710000 ;
      RECT 162.500000 230.710000 165.500000 230.990000 ;
      RECT 162.500000 238.030000 162.670000 238.050000 ;
      RECT 162.510000  33.255000 163.040000  33.425000 ;
      RECT 162.575000  68.635000 162.745000  71.415000 ;
      RECT 162.575000  72.305000 162.745000  73.575000 ;
      RECT 162.590000  49.780000 162.760000  54.890000 ;
      RECT 162.620000  61.675000 162.790000  63.695000 ;
      RECT 162.620000  63.865000 162.790000  67.115000 ;
      RECT 162.690000  30.145000 162.860000  33.255000 ;
      RECT 162.690000  33.425000 162.860000  34.915000 ;
      RECT 162.770000   1.640000 167.100000   1.810000 ;
      RECT 162.770000   1.810000 162.940000   4.080000 ;
      RECT 162.770000   4.080000 167.100000   4.250000 ;
      RECT 162.830000 198.815000 163.000000 205.605000 ;
      RECT 162.830000 206.465000 163.000000 213.255000 ;
      RECT 162.910000  37.765000 163.080000  40.865000 ;
      RECT 162.910000  57.305000 163.080000  60.405000 ;
      RECT 162.925000  76.165000 163.095000  78.875000 ;
      RECT 162.925000 221.215000 165.025000 230.235000 ;
      RECT 162.935000 231.160000 163.760000 231.605000 ;
      RECT 162.935000 232.050000 163.760000 238.575000 ;
      RECT 162.955000  41.445000 163.420000  41.615000 ;
      RECT 162.955000  41.615000 163.125000  42.520000 ;
      RECT 162.955000  42.520000 163.240000  42.690000 ;
      RECT 162.955000  55.480000 163.240000  55.650000 ;
      RECT 162.955000  55.650000 163.125000  56.555000 ;
      RECT 162.955000  56.555000 163.420000  56.725000 ;
      RECT 163.035000  29.425000 163.705000  29.595000 ;
      RECT 163.065000  68.885000 163.235000  71.015000 ;
      RECT 163.065000  71.015000 163.595000  71.185000 ;
      RECT 163.065000  71.185000 163.235000  73.635000 ;
      RECT 163.070000  42.690000 163.240000  43.615000 ;
      RECT 163.070000  52.095000 163.240000  55.480000 ;
      RECT 163.095000  29.595000 163.625000  29.745000 ;
      RECT 163.170000  61.675000 163.340000  63.495000 ;
      RECT 163.170000  64.405000 163.340000  67.115000 ;
      RECT 163.170000 198.595000 163.440000 205.815000 ;
      RECT 163.210000  75.775000 165.920000  75.945000 ;
      RECT 163.225000  83.310000 163.895000  83.480000 ;
      RECT 163.240000   2.220000 166.000000   2.390000 ;
      RECT 163.250000  40.395000 163.960000  40.865000 ;
      RECT 163.250000  40.865000 163.420000  41.445000 ;
      RECT 163.250000  56.725000 163.420000  57.305000 ;
      RECT 163.250000  57.305000 163.960000  57.775000 ;
      RECT 163.280000  81.770000 163.810000  81.940000 ;
      RECT 163.290000   3.500000 166.000000   3.670000 ;
      RECT 163.295000  41.785000 163.915000  42.115000 ;
      RECT 163.295000  56.055000 163.915000  56.385000 ;
      RECT 163.350000  67.515000 163.880000  67.585000 ;
      RECT 163.350000  67.585000 163.950000  67.685000 ;
      RECT 163.360000  68.205000 166.070000  68.375000 ;
      RECT 163.390000  33.255000 165.080000  33.425000 ;
      RECT 163.435000 192.285000 164.105000 193.605000 ;
      RECT 163.435000 193.605000 169.140000 194.135000 ;
      RECT 163.440000  61.175000 163.950000  61.505000 ;
      RECT 163.440000  67.685000 163.950000  67.915000 ;
      RECT 163.465000  83.895000 166.940000  84.405000 ;
      RECT 163.470000  81.940000 163.640000  83.060000 ;
      RECT 163.510000  61.505000 163.880000  67.515000 ;
      RECT 163.515000  78.340000 164.045000  78.510000 ;
      RECT 163.520000  48.350000 166.890000  48.520000 ;
      RECT 163.520000  49.650000 166.890000  49.820000 ;
      RECT 163.560000  45.290000 163.730000  48.000000 ;
      RECT 163.560000  50.170000 163.730000  52.880000 ;
      RECT 163.590000  41.360000 164.510000  41.530000 ;
      RECT 163.590000  41.530000 163.915000  41.785000 ;
      RECT 163.590000  56.385000 163.915000  56.640000 ;
      RECT 163.590000  56.640000 164.510000  56.810000 ;
      RECT 163.610000 198.815000 163.780000 205.605000 ;
      RECT 163.610000 206.465000 163.780000 213.255000 ;
      RECT 163.665000   8.065000 164.205000  13.460000 ;
      RECT 163.665000  18.830000 164.205000  24.225000 ;
      RECT 163.675000  70.335000 164.205000  70.505000 ;
      RECT 163.680000  48.215000 166.730000  48.350000 ;
      RECT 163.680000  49.820000 166.730000  49.955000 ;
      RECT 163.705000  75.945000 163.875000  78.340000 ;
      RECT 163.705000  78.510000 163.875000  78.875000 ;
      RECT 163.790000  38.155000 163.960000  40.395000 ;
      RECT 163.790000  57.775000 163.960000  60.015000 ;
      RECT 163.845000  68.375000 164.015000  70.335000 ;
      RECT 163.845000  70.505000 164.015000  73.635000 ;
      RECT 163.930000 230.990000 164.820000 238.295000 ;
      RECT 163.950000  42.605000 164.120000  44.400000 ;
      RECT 163.950000  53.770000 164.120000  55.565000 ;
      RECT 163.950000 198.595000 164.220000 205.815000 ;
      RECT 163.965000  45.030000 164.510000  45.200000 ;
      RECT 163.965000  52.970000 164.510000  53.140000 ;
      RECT 163.970000  30.145000 168.425000  31.485000 ;
      RECT 163.970000  31.485000 165.080000  31.735000 ;
      RECT 163.970000  31.735000 164.140000  32.855000 ;
      RECT 163.970000  33.860000 164.140000  34.915000 ;
      RECT 164.010000  13.630000 165.335000  14.040000 ;
      RECT 164.010000  18.250000 165.335000  18.660000 ;
      RECT 164.050000  61.800000 164.220000  67.420000 ;
      RECT 164.055000  44.570000 165.065000  44.740000 ;
      RECT 164.055000  44.740000 164.585000  44.800000 ;
      RECT 164.055000  53.370000 164.585000  53.430000 ;
      RECT 164.055000  53.430000 165.065000  53.600000 ;
      RECT 164.095000  82.050000 164.880000  83.895000 ;
      RECT 164.130000  37.595000 164.510000  38.615000 ;
      RECT 164.130000  59.555000 164.510000  60.575000 ;
      RECT 164.170000  42.000000 164.840000  42.170000 ;
      RECT 164.170000  56.000000 164.840000  56.170000 ;
      RECT 164.240000  42.170000 164.770000  42.300000 ;
      RECT 164.240000  55.870000 164.770000  56.000000 ;
      RECT 164.320000  61.175000 164.830000  61.505000 ;
      RECT 164.320000  67.585000 164.830000  67.915000 ;
      RECT 164.340000  40.195000 164.510000  41.360000 ;
      RECT 164.340000  45.000000 164.510000  45.030000 ;
      RECT 164.340000  45.200000 164.510000  48.000000 ;
      RECT 164.340000  50.170000 164.510000  52.970000 ;
      RECT 164.340000  53.140000 164.510000  53.170000 ;
      RECT 164.340000  56.810000 164.510000  57.975000 ;
      RECT 164.380000 239.105000 164.550000 240.355000 ;
      RECT 164.380000 240.355000 171.340000 240.525000 ;
      RECT 164.390000  61.505000 164.760000  67.585000 ;
      RECT 164.390000 198.815000 164.560000 205.605000 ;
      RECT 164.390000 206.465000 164.560000 213.315000 ;
      RECT 164.440000  38.970000 165.970000  39.720000 ;
      RECT 164.440000  58.450000 165.970000  59.200000 ;
      RECT 164.440000 241.585000 172.950000 242.435000 ;
      RECT 164.440000 242.435000 165.290000 244.355000 ;
      RECT 164.455000  71.015000 164.985000  71.185000 ;
      RECT 164.470000  42.505000 165.000000  42.675000 ;
      RECT 164.470000  55.495000 165.000000  55.665000 ;
      RECT 164.485000  76.165000 164.655000  78.875000 ;
      RECT 164.550000  29.190000 168.425000  30.145000 ;
      RECT 164.625000  68.885000 164.795000  71.015000 ;
      RECT 164.625000  71.185000 164.795000  73.635000 ;
      RECT 164.680000  37.765000 165.730000  38.970000 ;
      RECT 164.680000  39.720000 165.730000  40.865000 ;
      RECT 164.680000  57.305000 165.730000  58.450000 ;
      RECT 164.680000  59.200000 165.730000  60.405000 ;
      RECT 164.830000  42.675000 165.000000  43.615000 ;
      RECT 164.830000  54.555000 165.000000  55.495000 ;
      RECT 164.930000  61.675000 165.100000  62.740000 ;
      RECT 164.930000  62.910000 165.100000  63.285000 ;
      RECT 164.930000  63.905000 165.100000  64.235000 ;
      RECT 164.930000  64.405000 165.100000  67.115000 ;
      RECT 164.970000 198.235000 165.140000 206.440000 ;
      RECT 164.970000 206.440000 171.340000 206.610000 ;
      RECT 164.970000 206.610000 165.140000 213.855000 ;
      RECT 164.970000 214.025000 165.140000 217.810000 ;
      RECT 164.970000 217.810000 169.420000 217.980000 ;
      RECT 164.990000 231.315000 166.520000 235.420000 ;
      RECT 165.020000  63.455000 165.640000  63.625000 ;
      RECT 165.050000  83.310000 166.400000  83.480000 ;
      RECT 165.080000  78.340000 165.610000  78.510000 ;
      RECT 165.120000  45.290000 165.290000  48.000000 ;
      RECT 165.120000  50.170000 165.290000  52.880000 ;
      RECT 165.140000   8.065000 165.680000  13.460000 ;
      RECT 165.140000  18.830000 165.680000  24.225000 ;
      RECT 165.195000 221.910000 165.500000 230.710000 ;
      RECT 165.200000  61.175000 165.710000  61.505000 ;
      RECT 165.200000  67.585000 165.710000  67.915000 ;
      RECT 165.210000  81.395000 165.800000  81.940000 ;
      RECT 165.230000  70.335000 165.760000  70.505000 ;
      RECT 165.250000  31.775000 165.420000  32.165000 ;
      RECT 165.250000  32.165000 165.830000  32.335000 ;
      RECT 165.250000  32.335000 165.420000  34.915000 ;
      RECT 165.265000  75.945000 165.435000  78.340000 ;
      RECT 165.265000  78.510000 165.435000  78.875000 ;
      RECT 165.270000  61.505000 165.640000  63.455000 ;
      RECT 165.270000  63.625000 165.640000  67.585000 ;
      RECT 165.305000 113.195000 165.975000 113.525000 ;
      RECT 165.330000 236.270000 165.500000 236.485000 ;
      RECT 165.330000 236.485000 170.885000 236.655000 ;
      RECT 165.330000 236.655000 165.500000 239.660000 ;
      RECT 165.345000  44.570000 166.355000  44.740000 ;
      RECT 165.345000  53.430000 166.355000  53.600000 ;
      RECT 165.365000  79.140000 166.170000  79.310000 ;
      RECT 165.405000  68.375000 165.575000  70.335000 ;
      RECT 165.405000  70.505000 165.575000  73.635000 ;
      RECT 165.410000  42.505000 165.940000  42.675000 ;
      RECT 165.410000  42.675000 165.580000  43.615000 ;
      RECT 165.410000  54.555000 165.580000  55.495000 ;
      RECT 165.410000  55.495000 165.940000  55.665000 ;
      RECT 165.410000 113.910000 168.410000 164.900000 ;
      RECT 165.550000 198.705000 170.425000 198.875000 ;
      RECT 165.550000 199.485000 170.425000 199.655000 ;
      RECT 165.550000 200.265000 170.425000 200.435000 ;
      RECT 165.550000 200.815000 170.425000 200.985000 ;
      RECT 165.550000 201.595000 170.425000 201.765000 ;
      RECT 165.550000 202.375000 170.425000 202.545000 ;
      RECT 165.550000 202.925000 170.425000 203.095000 ;
      RECT 165.550000 203.705000 170.425000 203.875000 ;
      RECT 165.550000 204.255000 170.420000 204.425000 ;
      RECT 165.550000 205.035000 170.425000 205.205000 ;
      RECT 165.550000 205.815000 170.420000 205.985000 ;
      RECT 165.550000 207.380000 165.720000 217.230000 ;
      RECT 165.570000  42.000000 166.240000  42.170000 ;
      RECT 165.570000  56.000000 166.240000  56.170000 ;
      RECT 165.630000  81.940000 165.800000  83.060000 ;
      RECT 165.640000  42.170000 166.170000  42.300000 ;
      RECT 165.640000  55.870000 166.170000  56.000000 ;
      RECT 165.670000 228.585000 166.520000 231.315000 ;
      RECT 165.720000 221.465000 170.470000 222.075000 ;
      RECT 165.720000 222.245000 170.470000 222.855000 ;
      RECT 165.720000 223.025000 170.470000 223.635000 ;
      RECT 165.720000 223.805000 170.470000 224.415000 ;
      RECT 165.720000 224.585000 170.470000 225.195000 ;
      RECT 165.720000 225.365000 170.470000 225.975000 ;
      RECT 165.720000 226.145000 170.470000 226.755000 ;
      RECT 165.720000 226.925000 170.470000 227.535000 ;
      RECT 165.720000 227.705000 170.470000 228.200000 ;
      RECT 165.720000 235.940000 170.470000 236.215000 ;
      RECT 165.720000 236.825000 170.470000 237.215000 ;
      RECT 165.720000 237.385000 170.470000 237.880000 ;
      RECT 165.720000 238.050000 170.470000 238.545000 ;
      RECT 165.720000 238.715000 170.470000 239.325000 ;
      RECT 165.720000 239.495000 170.470000 239.990000 ;
      RECT 165.810000  61.800000 165.980000  67.420000 ;
      RECT 165.825000  44.740000 166.355000  44.800000 ;
      RECT 165.825000  53.370000 166.355000  53.430000 ;
      RECT 165.830000  31.485000 168.425000  31.595000 ;
      RECT 165.830000  31.595000 168.445000  31.765000 ;
      RECT 165.840000 206.800000 168.550000 206.980000 ;
      RECT 165.840000 217.440000 168.550000 217.620000 ;
      RECT 165.885000 236.215000 170.375000 236.315000 ;
      RECT 165.890000 206.980000 166.160000 217.440000 ;
      RECT 165.900000  37.335000 168.155000  37.505000 ;
      RECT 165.900000  37.505000 168.040000  37.595000 ;
      RECT 165.900000  37.595000 166.280000  38.615000 ;
      RECT 165.900000  40.195000 166.070000  41.360000 ;
      RECT 165.900000  41.360000 166.820000  41.530000 ;
      RECT 165.900000  45.000000 166.070000  45.030000 ;
      RECT 165.900000  45.030000 166.445000  45.200000 ;
      RECT 165.900000  45.200000 166.070000  48.000000 ;
      RECT 165.900000  50.170000 166.070000  52.970000 ;
      RECT 165.900000  52.970000 166.445000  53.140000 ;
      RECT 165.900000  53.140000 166.070000  53.170000 ;
      RECT 165.900000  56.640000 166.820000  56.810000 ;
      RECT 165.900000  56.810000 166.070000  57.975000 ;
      RECT 165.900000  59.555000 166.280000  60.575000 ;
      RECT 165.900000  60.575000 168.040000  60.665000 ;
      RECT 165.900000  60.665000 168.155000  60.835000 ;
      RECT 166.000000  79.310000 166.170000  80.475000 ;
      RECT 166.015000  71.015000 166.545000  71.185000 ;
      RECT 166.045000  76.165000 166.215000  78.875000 ;
      RECT 166.050000 243.195000 175.920000 244.045000 ;
      RECT 166.050000 244.045000 166.900000 252.535000 ;
      RECT 166.080000  61.175000 166.590000  61.505000 ;
      RECT 166.080000  67.585000 166.590000  67.915000 ;
      RECT 166.150000  61.505000 166.520000  63.695000 ;
      RECT 166.150000  63.695000 166.680000  63.865000 ;
      RECT 166.150000  63.865000 166.520000  67.585000 ;
      RECT 166.155000   7.195000 166.855000  14.325000 ;
      RECT 166.155000  17.965000 166.855000  25.095000 ;
      RECT 166.185000  68.885000 166.410000  71.015000 ;
      RECT 166.185000  71.185000 166.410000  73.345000 ;
      RECT 166.185000  73.345000 166.355000  73.635000 ;
      RECT 166.240000  68.205000 169.475000  68.375000 ;
      RECT 166.240000  68.375000 166.410000  68.885000 ;
      RECT 166.290000  42.605000 166.460000  44.400000 ;
      RECT 166.290000  53.770000 166.460000  55.565000 ;
      RECT 166.330000 207.380000 166.500000 217.230000 ;
      RECT 166.450000  38.155000 166.620000  40.395000 ;
      RECT 166.450000  40.395000 167.160000  40.865000 ;
      RECT 166.450000  57.305000 167.160000  57.775000 ;
      RECT 166.450000  57.775000 166.620000  60.015000 ;
      RECT 166.495000  41.530000 166.820000  41.785000 ;
      RECT 166.495000  41.785000 167.115000  42.115000 ;
      RECT 166.495000  56.055000 167.115000  56.385000 ;
      RECT 166.495000  56.385000 166.820000  56.640000 ;
      RECT 166.520000   2.435000 166.690000   3.445000 ;
      RECT 166.530000  31.765000 168.425000  32.710000 ;
      RECT 166.530000  32.710000 168.445000  32.785000 ;
      RECT 166.530000  33.860000 166.700000  34.915000 ;
      RECT 166.550000  79.635000 166.720000  80.790000 ;
      RECT 166.550000  80.960000 166.720000  80.985000 ;
      RECT 166.570000  82.050000 166.940000  83.895000 ;
      RECT 166.580000  81.395000 167.250000  81.565000 ;
      RECT 166.590000  75.775000 169.590000  75.945000 ;
      RECT 166.595000  76.165000 166.765000  78.340000 ;
      RECT 166.595000  78.340000 167.125000  78.510000 ;
      RECT 166.595000  78.510000 166.765000  78.875000 ;
      RECT 166.670000 206.980000 166.940000 217.440000 ;
      RECT 166.680000  45.290000 166.850000  48.000000 ;
      RECT 166.680000  50.170000 166.850000  52.880000 ;
      RECT 166.690000  61.675000 166.860000  63.495000 ;
      RECT 166.690000  64.405000 166.860000  67.115000 ;
      RECT 166.690000 228.700000 167.010000 235.275000 ;
      RECT 166.690000 235.275000 170.155000 235.770000 ;
      RECT 166.795000  69.905000 167.325000  70.075000 ;
      RECT 166.820000  97.825000 173.070000  98.675000 ;
      RECT 166.820000  98.675000 167.670000 106.775000 ;
      RECT 166.820000 106.775000 173.070000 107.625000 ;
      RECT 166.930000   1.810000 167.100000   4.080000 ;
      RECT 166.965000  68.885000 167.135000  69.905000 ;
      RECT 166.965000  70.075000 167.135000  73.635000 ;
      RECT 166.990000  40.865000 167.160000  41.445000 ;
      RECT 166.990000  41.445000 167.455000  41.615000 ;
      RECT 166.990000  56.555000 167.455000  56.725000 ;
      RECT 166.990000  56.725000 167.160000  57.305000 ;
      RECT 167.110000 207.380000 167.280000 217.230000 ;
      RECT 167.130000  95.995000 173.880000  96.030000 ;
      RECT 167.170000  42.520000 167.455000  42.690000 ;
      RECT 167.170000  42.690000 167.340000  43.615000 ;
      RECT 167.170000  54.555000 167.340000  55.480000 ;
      RECT 167.170000  55.480000 167.455000  55.650000 ;
      RECT 167.180000 228.370000 170.155000 228.865000 ;
      RECT 167.180000 229.035000 169.890000 229.645000 ;
      RECT 167.180000 229.815000 170.155000 230.425000 ;
      RECT 167.180000 230.595000 169.890000 231.205000 ;
      RECT 167.180000 231.375000 170.155000 231.985000 ;
      RECT 167.180000 232.155000 169.890000 232.765000 ;
      RECT 167.180000 232.935000 170.155000 233.545000 ;
      RECT 167.180000 233.715000 169.890000 234.325000 ;
      RECT 167.180000 234.495000 170.155000 234.990000 ;
      RECT 167.240000  61.675000 167.410000  62.725000 ;
      RECT 167.240000  62.955000 167.410000  63.285000 ;
      RECT 167.240000  63.905000 167.410000  64.235000 ;
      RECT 167.240000  64.405000 167.410000  67.420000 ;
      RECT 167.275000 192.395000 167.945000 192.875000 ;
      RECT 167.275000 192.875000 169.140000 193.405000 ;
      RECT 167.285000  41.615000 167.455000  42.520000 ;
      RECT 167.285000  55.650000 167.455000  56.555000 ;
      RECT 167.325000  83.310000 168.675000  83.480000 ;
      RECT 167.330000  37.765000 167.500000  40.865000 ;
      RECT 167.330000  57.305000 167.500000  60.405000 ;
      RECT 167.375000  75.945000 167.545000  78.875000 ;
      RECT 167.415000  84.555000 167.585000  86.210000 ;
      RECT 167.430000  81.820000 167.960000  81.990000 ;
      RECT 167.450000 206.980000 167.720000 217.440000 ;
      RECT 167.460000  81.480000 168.130000  81.650000 ;
      RECT 167.485000  41.085000 168.155000  41.255000 ;
      RECT 167.485000  56.915000 168.155000  57.085000 ;
      RECT 167.510000  43.110000 168.040000  43.280000 ;
      RECT 167.510000  54.890000 168.040000  55.060000 ;
      RECT 167.520000  81.395000 168.050000  81.480000 ;
      RECT 167.555000  32.785000 168.445000  33.600000 ;
      RECT 167.555000  35.565000 168.445000  35.945000 ;
      RECT 167.560000  84.070000 168.450000  84.240000 ;
      RECT 167.575000  33.600000 168.425000  35.565000 ;
      RECT 167.575000  71.015000 168.105000  71.185000 ;
      RECT 167.580000  61.175000 168.090000  61.505000 ;
      RECT 167.580000  67.115000 168.110000  67.285000 ;
      RECT 167.580000  67.585000 168.090000  67.915000 ;
      RECT 167.615000   5.735000 168.315000  15.795000 ;
      RECT 167.615000  16.495000 168.315000  26.555000 ;
      RECT 167.625000  41.760000 168.155000  41.930000 ;
      RECT 167.625000  41.930000 167.935000  43.110000 ;
      RECT 167.625000  55.060000 167.935000  56.240000 ;
      RECT 167.625000  56.240000 168.155000  56.410000 ;
      RECT 167.650000  43.280000 167.820000  48.390000 ;
      RECT 167.650000  49.780000 167.820000  54.890000 ;
      RECT 167.650000  61.505000 168.020000  67.115000 ;
      RECT 167.650000  67.285000 168.020000  67.585000 ;
      RECT 167.660000 244.805000 173.410000 245.655000 ;
      RECT 167.660000 245.655000 168.510000 250.435000 ;
      RECT 167.660000 250.435000 173.410000 251.715000 ;
      RECT 167.670000  37.595000 168.040000  41.085000 ;
      RECT 167.670000  41.255000 168.155000  41.265000 ;
      RECT 167.670000  41.265000 168.635000  41.435000 ;
      RECT 167.670000  56.735000 168.635000  56.905000 ;
      RECT 167.670000  56.905000 168.155000  56.915000 ;
      RECT 167.670000  57.085000 168.040000  60.575000 ;
      RECT 167.745000  68.375000 167.915000  71.015000 ;
      RECT 167.745000  71.185000 167.915000  73.635000 ;
      RECT 167.755000  84.595000 168.365000  84.765000 ;
      RECT 167.790000  81.990000 167.960000  83.060000 ;
      RECT 167.850000 251.715000 173.220000 251.845000 ;
      RECT 167.860000   0.880000 168.030000   5.035000 ;
      RECT 167.865000 113.195000 168.535000 113.525000 ;
      RECT 167.890000 207.380000 168.060000 217.230000 ;
      RECT 167.920000  83.735000 168.450000  84.070000 ;
      RECT 167.965000  78.340000 168.495000  78.510000 ;
      RECT 168.105000  42.130000 168.635000  42.300000 ;
      RECT 168.105000  55.870000 168.635000  56.040000 ;
      RECT 168.155000  76.165000 168.325000  78.340000 ;
      RECT 168.155000  78.510000 168.325000  78.875000 ;
      RECT 168.190000  61.675000 168.360000  66.145000 ;
      RECT 168.195000  84.555000 168.365000  84.595000 ;
      RECT 168.195000  84.765000 168.365000  85.565000 ;
      RECT 168.210000  38.155000 168.495000  40.865000 ;
      RECT 168.210000  57.305000 168.495000  60.015000 ;
      RECT 168.230000  44.180000 169.790000  44.350000 ;
      RECT 168.230000  44.350000 168.400000  45.760000 ;
      RECT 168.230000  45.760000 170.760000  45.930000 ;
      RECT 168.230000  46.100000 168.400000  46.335000 ;
      RECT 168.230000  46.335000 168.760000  46.505000 ;
      RECT 168.230000  46.505000 168.400000  48.380000 ;
      RECT 168.230000  49.790000 168.400000  51.665000 ;
      RECT 168.230000  51.665000 168.760000  51.835000 ;
      RECT 168.230000  51.835000 168.400000  52.070000 ;
      RECT 168.230000  52.240000 170.760000  52.410000 ;
      RECT 168.230000  52.410000 168.400000  53.820000 ;
      RECT 168.230000  53.820000 169.790000  53.990000 ;
      RECT 168.230000 206.980000 168.500000 217.440000 ;
      RECT 168.325000  40.865000 168.495000  41.095000 ;
      RECT 168.325000  41.435000 168.635000  42.130000 ;
      RECT 168.325000  56.040000 168.635000  56.735000 ;
      RECT 168.325000  57.075000 168.495000  57.305000 ;
      RECT 168.330000  42.840000 168.500000  44.010000 ;
      RECT 168.330000  54.160000 168.500000  55.330000 ;
      RECT 168.335000  85.870000 169.005000  86.040000 ;
      RECT 168.340000  81.395000 169.530000  81.565000 ;
      RECT 168.350000  69.905000 168.880000  70.075000 ;
      RECT 168.460000  61.175000 168.970000  61.385000 ;
      RECT 168.460000  61.385000 169.015000  61.505000 ;
      RECT 168.460000  67.585000 168.970000  67.915000 ;
      RECT 168.485000  61.505000 169.015000  61.555000 ;
      RECT 168.525000  68.885000 168.695000  69.905000 ;
      RECT 168.525000  70.075000 168.695000  74.525000 ;
      RECT 168.530000  61.555000 168.900000  67.585000 ;
      RECT 168.555000 173.755000 169.225000 173.925000 ;
      RECT 168.555000 174.115000 169.225000 174.285000 ;
      RECT 168.555000 175.785000 169.225000 175.955000 ;
      RECT 168.555000 176.325000 169.225000 176.495000 ;
      RECT 168.555000 177.995000 169.225000 178.165000 ;
      RECT 168.555000 178.535000 169.225000 178.705000 ;
      RECT 168.555000 180.205000 169.225000 180.375000 ;
      RECT 168.555000 180.745000 169.225000 180.915000 ;
      RECT 168.555000 182.415000 169.225000 188.785000 ;
      RECT 168.555000 189.915000 169.225000 192.565000 ;
      RECT 168.585000  84.485000 168.755000  85.870000 ;
      RECT 168.600000  99.085000 171.490000  99.255000 ;
      RECT 168.600000  99.865000 171.490000 100.035000 ;
      RECT 168.600000 100.415000 171.520000 100.585000 ;
      RECT 168.600000 101.195000 171.525000 101.365000 ;
      RECT 168.600000 101.975000 171.490000 102.145000 ;
      RECT 168.600000 102.525000 171.465000 102.695000 ;
      RECT 168.600000 103.305000 171.465000 103.475000 ;
      RECT 168.600000 104.085000 171.465000 104.255000 ;
      RECT 168.600000 104.635000 171.465000 104.805000 ;
      RECT 168.600000 105.415000 171.465000 105.585000 ;
      RECT 168.600000 106.195000 171.465000 106.365000 ;
      RECT 168.615000  42.470000 169.965000  42.640000 ;
      RECT 168.615000  55.530000 169.965000  55.700000 ;
      RECT 168.625000 173.705000 169.155000 173.755000 ;
      RECT 168.670000 207.380000 168.840000 217.230000 ;
      RECT 168.715000  42.640000 169.965000  42.670000 ;
      RECT 168.715000  55.500000 169.965000  55.530000 ;
      RECT 168.760000  42.840000 168.930000  44.180000 ;
      RECT 168.760000  53.990000 168.930000  55.330000 ;
      RECT 168.790000  37.765000 168.960000  40.845000 ;
      RECT 168.790000  57.325000 168.960000  60.405000 ;
      RECT 168.820000  35.165000 169.350000  35.335000 ;
      RECT 168.870000  79.540000 169.040000  80.985000 ;
      RECT 168.870000  82.050000 169.145000  83.060000 ;
      RECT 168.925000  83.060000 169.145000  84.615000 ;
      RECT 168.925000  84.615000 169.585000  85.575000 ;
      RECT 168.935000  75.945000 169.105000  78.875000 ;
      RECT 168.945000  71.015000 169.475000  71.185000 ;
      RECT 169.075000   6.495000 173.450000   7.195000 ;
      RECT 169.075000   7.195000 169.775000  14.325000 ;
      RECT 169.075000  14.325000 173.450000  15.035000 ;
      RECT 169.075000  17.255000 173.450000  17.965000 ;
      RECT 169.075000  17.965000 169.775000  25.095000 ;
      RECT 169.075000  25.095000 173.450000  25.795000 ;
      RECT 169.140000  61.675000 169.310000  62.740000 ;
      RECT 169.140000  62.910000 169.310000  63.285000 ;
      RECT 169.140000  63.905000 169.310000  64.235000 ;
      RECT 169.140000  64.405000 169.310000  67.115000 ;
      RECT 169.175000  85.575000 169.585000  85.850000 ;
      RECT 169.175000  85.850000 169.705000  86.020000 ;
      RECT 169.180000  32.125000 169.350000  32.135000 ;
      RECT 169.180000  32.135000 169.900000  33.645000 ;
      RECT 169.180000  33.815000 169.900000  34.145000 ;
      RECT 169.180000  34.145000 169.350000  35.165000 ;
      RECT 169.190000  42.840000 169.360000  44.010000 ;
      RECT 169.190000  54.160000 169.360000  55.330000 ;
      RECT 169.245000  79.140000 170.135000  79.240000 ;
      RECT 169.245000  79.240000 170.155000  79.310000 ;
      RECT 169.250000 206.610000 169.420000 217.810000 ;
      RECT 169.250000 246.125000 171.960000 246.295000 ;
      RECT 169.250000 246.905000 171.960000 247.075000 ;
      RECT 169.250000 247.685000 171.960000 247.855000 ;
      RECT 169.250000 248.235000 171.960000 248.405000 ;
      RECT 169.250000 249.015000 171.960000 249.185000 ;
      RECT 169.250000 249.795000 171.960000 249.965000 ;
      RECT 169.260000 220.235000 171.000000 220.765000 ;
      RECT 169.305000  68.375000 169.475000  71.015000 ;
      RECT 169.305000  71.185000 169.475000  73.635000 ;
      RECT 169.355000  78.340000 169.885000  78.510000 ;
      RECT 169.360000  81.565000 169.530000  84.030000 ;
      RECT 169.360000  84.030000 169.950000  84.200000 ;
      RECT 169.360000  84.200000 169.530000  84.415000 ;
      RECT 169.410000  44.580000 169.580000  45.280000 ;
      RECT 169.410000  45.280000 170.085000  45.450000 ;
      RECT 169.410000  45.450000 169.580000  45.590000 ;
      RECT 169.410000  46.100000 169.580000  48.550000 ;
      RECT 169.410000  48.550000 172.300000  48.720000 ;
      RECT 169.410000  49.450000 172.300000  49.620000 ;
      RECT 169.410000  49.620000 169.580000  52.070000 ;
      RECT 169.410000  52.580000 169.580000  52.720000 ;
      RECT 169.410000  52.720000 170.085000  52.890000 ;
      RECT 169.410000  52.890000 169.580000  53.590000 ;
      RECT 169.410000  61.175000 169.920000  61.505000 ;
      RECT 169.410000  67.585000 169.920000  67.915000 ;
      RECT 169.480000  61.505000 169.850000  67.585000 ;
      RECT 169.620000  42.840000 169.790000  44.180000 ;
      RECT 169.620000  53.990000 169.790000  55.330000 ;
      RECT 169.715000  76.165000 169.885000  78.340000 ;
      RECT 169.715000  78.510000 169.885000  78.875000 ;
      RECT 169.730000  34.315000 169.900000  35.325000 ;
      RECT 169.755000  79.310000 170.155000  83.060000 ;
      RECT 169.755000  84.555000 169.925000  85.565000 ;
      RECT 169.760000 173.655000 171.780000 174.405000 ;
      RECT 169.760000 184.235000 171.780000 184.985000 ;
      RECT 169.780000  83.660000 170.310000  83.830000 ;
      RECT 169.845000 186.225000 170.515000 188.785000 ;
      RECT 169.845000 189.915000 170.515000 192.565000 ;
      RECT 169.855000  68.885000 170.025000  69.905000 ;
      RECT 169.855000  69.905000 170.385000  70.075000 ;
      RECT 169.855000  70.075000 170.025000  73.635000 ;
      RECT 169.910000  46.165000 170.240000  47.015000 ;
      RECT 169.910000  51.155000 170.240000  52.005000 ;
      RECT 169.920000 113.910000 172.920000 164.900000 ;
      RECT 169.990000  47.015000 170.160000  47.625000 ;
      RECT 169.990000  50.545000 170.160000  51.155000 ;
      RECT 169.990000  73.855000 171.340000  74.170000 ;
      RECT 170.020000  61.800000 170.190000  67.420000 ;
      RECT 170.050000  42.840000 170.220000  44.010000 ;
      RECT 170.050000  54.160000 170.220000  55.330000 ;
      RECT 170.070000  31.635000 170.240000  35.825000 ;
      RECT 170.135000  37.870000 170.305000  40.870000 ;
      RECT 170.135000  57.300000 170.305000  60.300000 ;
      RECT 170.140000  83.405000 170.310000  83.660000 ;
      RECT 170.140000  83.830000 170.310000  84.415000 ;
      RECT 170.180000 207.370000 172.950000 218.740000 ;
      RECT 170.250000   8.065000 170.790000  13.460000 ;
      RECT 170.250000  18.830000 170.790000  24.225000 ;
      RECT 170.290000  61.175000 170.800000  61.505000 ;
      RECT 170.290000  67.585000 170.800000  67.915000 ;
      RECT 170.305000  75.525000 170.475000  79.145000 ;
      RECT 170.320000  42.470000 171.670000  42.475000 ;
      RECT 170.320000  42.475000 172.980000  42.645000 ;
      RECT 170.320000  55.525000 172.980000  55.695000 ;
      RECT 170.320000  55.695000 171.670000  55.700000 ;
      RECT 170.355000  41.360000 170.885000  41.530000 ;
      RECT 170.355000  56.640000 170.885000  56.810000 ;
      RECT 170.360000  61.505000 170.730000  67.585000 ;
      RECT 170.440000  31.635000 170.610000  35.995000 ;
      RECT 170.440000  35.995000 172.060000  36.165000 ;
      RECT 170.480000  42.840000 170.650000  44.180000 ;
      RECT 170.480000  44.180000 172.300000  44.350000 ;
      RECT 170.480000  53.820000 172.300000  53.990000 ;
      RECT 170.480000  53.990000 170.650000  55.330000 ;
      RECT 170.535000  82.050000 170.705000  86.210000 ;
      RECT 170.590000  44.580000 170.760000  45.760000 ;
      RECT 170.590000  45.930000 170.760000  47.080000 ;
      RECT 170.590000  47.370000 171.460000  48.380000 ;
      RECT 170.590000  49.790000 171.460000  50.800000 ;
      RECT 170.590000  51.090000 170.760000  52.240000 ;
      RECT 170.590000  52.410000 170.760000  53.590000 ;
      RECT 170.595000  13.630000 171.920000  14.040000 ;
      RECT 170.595000  18.250000 171.920000  18.660000 ;
      RECT 170.635000  68.885000 170.805000  70.685000 ;
      RECT 170.635000  70.685000 170.860000  71.225000 ;
      RECT 170.635000  71.225000 170.805000  73.635000 ;
      RECT 170.640000 220.765000 171.000000 222.010000 ;
      RECT 170.640000 234.695000 170.885000 236.485000 ;
      RECT 170.665000  77.480000 173.715000  78.010000 ;
      RECT 170.675000 203.150000 170.980000 203.820000 ;
      RECT 170.675000 204.480000 170.980000 205.760000 ;
      RECT 170.685000 199.005000 170.980000 200.255000 ;
      RECT 170.685000 201.020000 170.980000 202.270000 ;
      RECT 170.705000 204.205000 170.875000 204.480000 ;
      RECT 170.715000  37.840000 174.955000  38.010000 ;
      RECT 170.715000  38.010000 170.885000  41.360000 ;
      RECT 170.715000  56.810000 170.885000  60.160000 ;
      RECT 170.715000  60.160000 174.955000  60.330000 ;
      RECT 170.785000  75.265000 173.675000  77.480000 ;
      RECT 170.785000  78.010000 173.675000  79.185000 ;
      RECT 170.810000  31.635000 171.660000  31.965000 ;
      RECT 170.810000  31.965000 170.980000  35.495000 ;
      RECT 170.810000  35.495000 171.660000  35.825000 ;
      RECT 170.810000 198.930000 170.980000 199.005000 ;
      RECT 170.810000 200.255000 170.980000 200.280000 ;
      RECT 170.810000 200.970000 170.980000 201.020000 ;
      RECT 170.810000 202.270000 170.980000 202.320000 ;
      RECT 170.900000  61.675000 171.070000  63.495000 ;
      RECT 170.900000  64.405000 171.070000  67.115000 ;
      RECT 170.910000  42.840000 171.080000  44.010000 ;
      RECT 170.910000  54.160000 171.080000  55.330000 ;
      RECT 170.930000  46.335000 171.460000  47.370000 ;
      RECT 170.930000  50.800000 171.460000  51.835000 ;
      RECT 170.935000  80.165000 171.155000  81.175000 ;
      RECT 170.935000  81.175000 171.105000  82.380000 ;
      RECT 170.935000  82.380000 171.255000  85.090000 ;
      RECT 170.940000  37.335000 172.970000  37.505000 ;
      RECT 170.940000  60.665000 172.970000  60.835000 ;
      RECT 171.055000  72.535000 171.585000  72.705000 ;
      RECT 171.125000 192.395000 171.795000 192.565000 ;
      RECT 171.150000  32.135000 171.320000  33.645000 ;
      RECT 171.150000  33.815000 171.320000  34.145000 ;
      RECT 171.150000  34.315000 171.320000  35.325000 ;
      RECT 171.170000 198.235000 171.340000 206.440000 ;
      RECT 171.170000 221.045000 171.340000 240.355000 ;
      RECT 171.275000  81.370000 171.785000  81.700000 ;
      RECT 171.325000  80.660000 171.695000  81.370000 ;
      RECT 171.340000  42.840000 171.510000  44.180000 ;
      RECT 171.340000  53.990000 171.510000  55.330000 ;
      RECT 171.410000  45.280000 171.940000  45.450000 ;
      RECT 171.410000  52.720000 171.940000  52.890000 ;
      RECT 171.415000  68.885000 171.585000  72.535000 ;
      RECT 171.415000  72.705000 171.585000  73.635000 ;
      RECT 171.450000  61.675000 171.620000  63.495000 ;
      RECT 171.450000  64.405000 171.620000  67.115000 ;
      RECT 171.490000  31.965000 171.660000  35.495000 ;
      RECT 171.595000  38.180000 171.855000  41.160000 ;
      RECT 171.595000  57.010000 171.855000  59.990000 ;
      RECT 171.630000  63.695000 172.160000  63.865000 ;
      RECT 171.660000  85.650000 175.800000  86.375000 ;
      RECT 171.720000  61.175000 172.230000  61.505000 ;
      RECT 171.720000  67.585000 172.230000  67.915000 ;
      RECT 171.725000   8.065000 172.265000  13.460000 ;
      RECT 171.725000  18.830000 172.265000  24.225000 ;
      RECT 171.735000  99.215000 172.040000 106.140000 ;
      RECT 171.770000  42.840000 171.940000  44.010000 ;
      RECT 171.770000  44.580000 171.940000  45.280000 ;
      RECT 171.770000  45.450000 171.940000  47.080000 ;
      RECT 171.770000  47.370000 172.300000  48.550000 ;
      RECT 171.770000  49.620000 172.300000  50.800000 ;
      RECT 171.770000  51.090000 171.940000  52.720000 ;
      RECT 171.770000  52.890000 171.940000  53.590000 ;
      RECT 171.770000  54.160000 171.940000  55.330000 ;
      RECT 171.790000  61.505000 172.160000  63.695000 ;
      RECT 171.790000  63.865000 172.160000  67.585000 ;
      RECT 171.860000  31.635000 172.030000  35.995000 ;
      RECT 171.865000  79.540000 172.035000  81.175000 ;
      RECT 171.880000  70.285000 175.800000  71.225000 ;
      RECT 171.895000  68.615000 175.800000  70.285000 ;
      RECT 171.895000  71.225000 175.800000  73.615000 ;
      RECT 171.965000  82.170000 172.135000  85.650000 ;
      RECT 172.055000  38.180000 172.315000  41.160000 ;
      RECT 172.055000  57.010000 172.315000  59.990000 ;
      RECT 172.100000 197.275000 172.950000 207.370000 ;
      RECT 172.100000 220.065000 172.950000 241.585000 ;
      RECT 172.110000  43.095000 172.640000  43.265000 ;
      RECT 172.110000  44.350000 172.300000  47.370000 ;
      RECT 172.110000  50.800000 172.300000  53.820000 ;
      RECT 172.110000  54.905000 172.640000  55.075000 ;
      RECT 172.150000 246.350000 172.320000 249.820000 ;
      RECT 172.165000  81.285000 172.675000  81.615000 ;
      RECT 172.220000  98.675000 173.070000 106.775000 ;
      RECT 172.230000  31.635000 172.400000  35.825000 ;
      RECT 172.230000  41.360000 172.760000  41.530000 ;
      RECT 172.230000  56.640000 172.760000  56.810000 ;
      RECT 172.305000  81.615000 172.675000  84.930000 ;
      RECT 172.330000  61.800000 172.500000  67.420000 ;
      RECT 172.405000 173.755000 174.095000 173.925000 ;
      RECT 172.405000 173.925000 174.090000 174.150000 ;
      RECT 172.405000 174.150000 174.095000 174.320000 ;
      RECT 172.405000 174.320000 174.090000 174.355000 ;
      RECT 172.405000 181.435000 174.095000 184.885000 ;
      RECT 172.405000 192.395000 173.075000 192.565000 ;
      RECT 172.410000  41.530000 172.580000  42.305000 ;
      RECT 172.410000  55.865000 172.580000  56.640000 ;
      RECT 172.470000  43.265000 172.640000  48.390000 ;
      RECT 172.470000  49.780000 172.640000  54.905000 ;
      RECT 172.560000 245.655000 173.410000 250.435000 ;
      RECT 172.570000  32.135000 173.290000  33.645000 ;
      RECT 172.570000  33.815000 173.290000  34.145000 ;
      RECT 172.570000  34.315000 172.740000  35.325000 ;
      RECT 172.600000  61.175000 173.110000  61.505000 ;
      RECT 172.600000  67.585000 173.110000  67.915000 ;
      RECT 172.670000  61.505000 173.040000  67.585000 ;
      RECT 172.750000   7.195000 173.450000  14.325000 ;
      RECT 172.750000  17.965000 173.450000  25.095000 ;
      RECT 172.810000  42.645000 172.980000  43.405000 ;
      RECT 172.810000  43.405000 173.460000  44.415000 ;
      RECT 172.810000  53.755000 173.460000  54.765000 ;
      RECT 172.810000  54.765000 172.980000  55.525000 ;
      RECT 172.845000  80.660000 173.795000  81.175000 ;
      RECT 172.845000  81.175000 173.015000  85.090000 ;
      RECT 172.910000  35.165000 173.440000  35.335000 ;
      RECT 172.930000  41.290000 173.600000  41.460000 ;
      RECT 172.930000  46.335000 173.460000  46.505000 ;
      RECT 172.930000  51.665000 173.460000  51.835000 ;
      RECT 172.930000  56.710000 173.600000  56.880000 ;
      RECT 172.950000  47.855000 173.120000  48.465000 ;
      RECT 172.950000  48.465000 175.800000  48.635000 ;
      RECT 172.950000  49.535000 175.800000  49.705000 ;
      RECT 172.950000  49.705000 173.120000  50.315000 ;
      RECT 172.990000  42.030000 173.520000  42.200000 ;
      RECT 172.990000  55.970000 173.520000  56.140000 ;
      RECT 173.025000  38.180000 173.195000  41.290000 ;
      RECT 173.025000  41.460000 173.520000  42.030000 ;
      RECT 173.025000  56.140000 173.520000  56.710000 ;
      RECT 173.025000  56.880000 173.195000  59.990000 ;
      RECT 173.120000  32.125000 173.290000  32.135000 ;
      RECT 173.120000  34.145000 173.290000  35.165000 ;
      RECT 173.180000  37.335000 173.850000  37.505000 ;
      RECT 173.180000  60.665000 173.850000  60.835000 ;
      RECT 173.185000  81.370000 173.715000  81.940000 ;
      RECT 173.210000  61.675000 173.380000  62.740000 ;
      RECT 173.210000  62.910000 173.380000  63.285000 ;
      RECT 173.210000  63.905000 173.380000  64.235000 ;
      RECT 173.210000  64.405000 173.380000  67.115000 ;
      RECT 173.250000  48.635000 174.420000  48.655000 ;
      RECT 173.250000  60.835000 173.780000  60.885000 ;
      RECT 173.270000  36.975000 173.440000  37.335000 ;
      RECT 173.290000  44.415000 173.460000  46.335000 ;
      RECT 173.290000  46.505000 173.460000  48.085000 ;
      RECT 173.290000  50.085000 173.460000  51.665000 ;
      RECT 173.290000  51.835000 173.460000  53.755000 ;
      RECT 173.480000  61.175000 173.990000  61.415000 ;
      RECT 173.480000  61.415000 174.080000  61.505000 ;
      RECT 173.480000  67.585000 173.990000  67.915000 ;
      RECT 173.550000  61.505000 174.080000  61.585000 ;
      RECT 173.550000  61.585000 173.920000  67.585000 ;
      RECT 173.625000  80.165000 173.795000  80.660000 ;
      RECT 173.630000  45.000000 174.160000  45.170000 ;
      RECT 173.630000  53.000000 174.160000  53.170000 ;
      RECT 173.690000  41.635000 173.940000  42.305000 ;
      RECT 173.690000  55.865000 173.940000  56.535000 ;
      RECT 173.725000  41.580000 173.940000  41.635000 ;
      RECT 173.725000  42.305000 173.895000  43.405000 ;
      RECT 173.725000  43.405000 173.920000  44.415000 ;
      RECT 173.725000  53.755000 173.920000  54.765000 ;
      RECT 173.725000  54.765000 173.895000  55.865000 ;
      RECT 173.725000  56.535000 173.940000  56.590000 ;
      RECT 173.725000  82.170000 173.895000  85.650000 ;
      RECT 173.750000  45.170000 173.920000  48.085000 ;
      RECT 173.750000  50.085000 173.920000  53.000000 ;
      RECT 173.770000  38.180000 174.075000  40.890000 ;
      RECT 173.770000  40.890000 173.940000  41.580000 ;
      RECT 173.770000  56.590000 173.940000  57.280000 ;
      RECT 173.770000  57.280000 174.075000  59.990000 ;
      RECT 173.880000  97.045000 190.270000  97.095000 ;
      RECT 173.880000  97.095000 190.275000 101.900000 ;
      RECT 173.880000 101.900000 174.730000 108.735000 ;
      RECT 174.000000 195.155000 175.920000 243.195000 ;
      RECT 174.090000  42.400000 174.620000  42.570000 ;
      RECT 174.090000  42.570000 174.500000  44.585000 ;
      RECT 174.090000  44.585000 174.630000  44.740000 ;
      RECT 174.090000  45.375000 174.630000  45.665000 ;
      RECT 174.090000  45.665000 174.380000  48.085000 ;
      RECT 174.090000  50.085000 174.380000  52.505000 ;
      RECT 174.090000  52.505000 174.630000  52.795000 ;
      RECT 174.090000  53.430000 174.630000  53.585000 ;
      RECT 174.090000  53.585000 174.500000  55.600000 ;
      RECT 174.090000  55.600000 174.620000  55.770000 ;
      RECT 174.090000  61.800000 174.260000  67.420000 ;
      RECT 174.110000  42.030000 175.140000  42.200000 ;
      RECT 174.110000  55.970000 175.140000  56.140000 ;
      RECT 174.130000  37.335000 174.800000  37.505000 ;
      RECT 174.130000  60.665000 174.800000  60.835000 ;
      RECT 174.160000 244.045000 175.920000 252.535000 ;
      RECT 174.180000  95.995000 190.270000  96.030000 ;
      RECT 174.210000   5.735000 174.910000  15.795000 ;
      RECT 174.210000  16.495000 174.910000  26.555000 ;
      RECT 174.210000  41.290000 174.955000  41.460000 ;
      RECT 174.210000  56.710000 174.955000  56.880000 ;
      RECT 174.280000  41.460000 174.810000  41.530000 ;
      RECT 174.280000  56.640000 174.810000  56.710000 ;
      RECT 174.305000  95.985000 190.270000  95.995000 ;
      RECT 174.325000 113.195000 174.995000 113.525000 ;
      RECT 174.330000  44.740000 174.630000  45.375000 ;
      RECT 174.330000  52.795000 174.630000  53.430000 ;
      RECT 174.360000  61.175000 174.870000  61.505000 ;
      RECT 174.360000  67.585000 174.870000  67.915000 ;
      RECT 174.430000  61.505000 174.800000  67.585000 ;
      RECT 174.430000 113.910000 177.430000 164.900000 ;
      RECT 174.580000  48.105000 175.335000  48.275000 ;
      RECT 174.580000  49.895000 175.335000  50.065000 ;
      RECT 174.670000  43.405000 174.840000  44.415000 ;
      RECT 174.670000  53.755000 174.840000  54.765000 ;
      RECT 174.730000  73.615000 175.800000  85.650000 ;
      RECT 174.785000  38.010000 174.955000  41.290000 ;
      RECT 174.785000  56.880000 174.955000  60.160000 ;
      RECT 174.805000  46.335000 175.335000  46.505000 ;
      RECT 174.805000  51.665000 175.335000  51.835000 ;
      RECT 174.825000  44.630000 174.995000  45.300000 ;
      RECT 174.825000  52.870000 174.995000  53.540000 ;
      RECT 174.865000  42.510000 175.400000  43.085000 ;
      RECT 174.865000  55.085000 175.400000  55.660000 ;
      RECT 174.970000  41.635000 175.140000  42.030000 ;
      RECT 174.970000  42.200000 175.140000  42.305000 ;
      RECT 174.970000  55.865000 175.140000  55.970000 ;
      RECT 174.970000  56.140000 175.140000  56.535000 ;
      RECT 174.970000  61.675000 175.140000  63.855000 ;
      RECT 174.970000  64.405000 175.140000  67.115000 ;
      RECT 175.020000 173.235000 190.325000 174.305000 ;
      RECT 175.020000 174.305000 175.920000 194.305000 ;
      RECT 175.130000  43.405000 175.335000  44.415000 ;
      RECT 175.130000  53.755000 175.335000  54.765000 ;
      RECT 175.165000  44.415000 175.335000  46.335000 ;
      RECT 175.165000  46.505000 175.335000  48.105000 ;
      RECT 175.165000  50.065000 175.335000  51.665000 ;
      RECT 175.165000  51.835000 175.335000  53.755000 ;
      RECT 175.270000  64.065000 175.800000  64.235000 ;
      RECT 175.345000  48.635000 175.800000  48.655000 ;
      RECT 175.630000  37.870000 175.800000  44.425000 ;
      RECT 175.630000  45.065000 175.800000  48.465000 ;
      RECT 175.630000  49.705000 175.800000  52.000000 ;
      RECT 175.630000  52.610000 175.800000  63.485000 ;
      RECT 175.630000  63.905000 175.800000  64.065000 ;
      RECT 175.630000  64.235000 175.800000  68.615000 ;
      RECT 175.995000 105.870000 176.465000 105.900000 ;
      RECT 175.995000 105.900000 176.545000 106.070000 ;
      RECT 175.995000 106.070000 176.465000 106.545000 ;
      RECT 176.050000 102.445000 176.380000 102.615000 ;
      RECT 176.050000 102.785000 176.380000 102.955000 ;
      RECT 176.130000 102.425000 176.300000 102.445000 ;
      RECT 176.130000 102.615000 176.300000 102.785000 ;
      RECT 176.755000 175.100000 213.250000 253.240000 ;
      RECT 176.885000 113.195000 177.555000 113.525000 ;
      RECT 176.975000  23.665000 178.995000  24.415000 ;
      RECT 176.975000  34.245000 178.995000  34.995000 ;
      RECT 177.320000  37.110000 212.685000  88.630000 ;
      RECT 177.595000 101.900000 190.275000 108.735000 ;
      RECT 178.940000 113.910000 181.940000 164.900000 ;
      RECT 183.345000 113.195000 184.015000 113.525000 ;
      RECT 183.415000 113.165000 183.945000 113.195000 ;
      RECT 183.450000 113.910000 186.450000 164.900000 ;
      RECT 183.940000   0.330000 205.860000  37.110000 ;
      RECT 187.055000 111.435000 187.905000 166.535000 ;
      RECT 189.475000 109.585000 190.325000 168.145000 ;
      RECT 191.735000  95.265000 198.365000 175.100000 ;
      RECT 199.680000 108.735000 300.970000 109.585000 ;
      RECT 199.680000 109.585000 200.530000 168.145000 ;
      RECT 199.680000 168.145000 300.630000 173.235000 ;
      RECT 199.680000 173.235000 214.985000 174.305000 ;
      RECT 199.730000  96.030000 235.725000  96.880000 ;
      RECT 199.730000  97.095000 216.125000 101.900000 ;
      RECT 199.730000 101.900000 212.410000 108.735000 ;
      RECT 199.735000  95.985000 215.700000  95.995000 ;
      RECT 199.735000  95.995000 215.825000  96.030000 ;
      RECT 199.735000  96.880000 235.725000  97.045000 ;
      RECT 199.735000  97.045000 216.125000  97.095000 ;
      RECT 202.100000 110.585000 298.210000 111.435000 ;
      RECT 202.100000 111.435000 202.950000 166.535000 ;
      RECT 202.100000 166.535000 298.210000 167.385000 ;
      RECT 203.555000 113.910000 206.555000 164.900000 ;
      RECT 205.990000 113.195000 206.660000 113.525000 ;
      RECT 206.060000 113.165000 206.590000 113.195000 ;
      RECT 208.065000 113.910000 211.065000 164.900000 ;
      RECT 211.010000  23.665000 213.030000  24.415000 ;
      RECT 211.010000  34.245000 213.030000  34.995000 ;
      RECT 212.450000 113.195000 213.120000 113.525000 ;
      RECT 212.575000 113.910000 215.575000 164.900000 ;
      RECT 213.460000 105.900000 214.010000 106.070000 ;
      RECT 213.540000 105.870000 214.010000 105.900000 ;
      RECT 213.540000 106.070000 214.010000 106.545000 ;
      RECT 213.625000 102.445000 213.955000 102.615000 ;
      RECT 213.625000 102.785000 213.955000 102.955000 ;
      RECT 213.705000 102.425000 213.875000 102.445000 ;
      RECT 213.705000 102.615000 213.875000 102.785000 ;
      RECT 214.085000 174.305000 214.985000 194.305000 ;
      RECT 214.085000 194.305000 227.965000 195.155000 ;
      RECT 214.085000 195.155000 216.005000 243.195000 ;
      RECT 214.085000 243.195000 223.955000 244.045000 ;
      RECT 214.085000 244.045000 215.845000 252.535000 ;
      RECT 214.085000 252.535000 348.425000 253.385000 ;
      RECT 214.205000  37.870000 214.375000  44.425000 ;
      RECT 214.205000  45.065000 214.375000  48.465000 ;
      RECT 214.205000  48.465000 217.055000  48.635000 ;
      RECT 214.205000  48.635000 214.660000  48.655000 ;
      RECT 214.205000  49.535000 217.055000  49.705000 ;
      RECT 214.205000  49.705000 214.375000  52.000000 ;
      RECT 214.205000  52.610000 214.375000  63.485000 ;
      RECT 214.205000  63.905000 214.375000  64.065000 ;
      RECT 214.205000  64.065000 214.735000  64.235000 ;
      RECT 214.205000  64.235000 214.375000  68.615000 ;
      RECT 214.205000  68.615000 218.110000  70.285000 ;
      RECT 214.205000  70.285000 218.125000  71.225000 ;
      RECT 214.205000  71.225000 218.110000  73.615000 ;
      RECT 214.205000  73.615000 215.275000  85.650000 ;
      RECT 214.205000  85.650000 218.345000  86.375000 ;
      RECT 214.205000  86.375000 234.280000  86.380000 ;
      RECT 214.205000  86.380000 234.265000  87.070000 ;
      RECT 214.205000  87.070000 237.660000  87.700000 ;
      RECT 214.205000  87.700000 290.955000  87.870000 ;
      RECT 214.205000  87.870000 278.020000  87.885000 ;
      RECT 214.605000  42.510000 215.140000  43.085000 ;
      RECT 214.605000  55.085000 215.140000  55.660000 ;
      RECT 214.670000  43.405000 214.875000  44.415000 ;
      RECT 214.670000  44.415000 214.840000  46.335000 ;
      RECT 214.670000  46.335000 215.200000  46.505000 ;
      RECT 214.670000  46.505000 214.840000  48.105000 ;
      RECT 214.670000  48.105000 215.425000  48.275000 ;
      RECT 214.670000  49.895000 215.425000  50.065000 ;
      RECT 214.670000  50.065000 214.840000  51.665000 ;
      RECT 214.670000  51.665000 215.200000  51.835000 ;
      RECT 214.670000  51.835000 214.840000  53.755000 ;
      RECT 214.670000  53.755000 214.875000  54.765000 ;
      RECT 214.865000  41.635000 215.035000  42.030000 ;
      RECT 214.865000  42.030000 215.895000  42.200000 ;
      RECT 214.865000  42.200000 215.035000  42.305000 ;
      RECT 214.865000  55.865000 215.035000  55.970000 ;
      RECT 214.865000  55.970000 215.895000  56.140000 ;
      RECT 214.865000  56.140000 215.035000  56.535000 ;
      RECT 214.865000  61.675000 215.035000  63.855000 ;
      RECT 214.865000  64.405000 215.035000  67.115000 ;
      RECT 215.010000  44.630000 215.180000  45.300000 ;
      RECT 215.010000  52.870000 215.180000  53.540000 ;
      RECT 215.010000 113.195000 215.680000 113.525000 ;
      RECT 215.050000  37.840000 219.290000  38.010000 ;
      RECT 215.050000  38.010000 215.220000  41.290000 ;
      RECT 215.050000  41.290000 215.795000  41.460000 ;
      RECT 215.050000  56.710000 215.795000  56.880000 ;
      RECT 215.050000  56.880000 215.220000  60.160000 ;
      RECT 215.050000  60.160000 219.290000  60.330000 ;
      RECT 215.095000   5.035000 228.985000   5.735000 ;
      RECT 215.095000   5.735000 215.795000  15.795000 ;
      RECT 215.095000  15.795000 228.985000  16.495000 ;
      RECT 215.095000  16.495000 215.795000  26.555000 ;
      RECT 215.095000  26.555000 228.985000  27.255000 ;
      RECT 215.135000  61.175000 215.645000  61.505000 ;
      RECT 215.135000  67.585000 215.645000  67.915000 ;
      RECT 215.165000  43.405000 215.335000  44.415000 ;
      RECT 215.165000  53.755000 215.335000  54.765000 ;
      RECT 215.195000  41.460000 215.725000  41.530000 ;
      RECT 215.195000  56.640000 215.725000  56.710000 ;
      RECT 215.205000  37.335000 215.875000  37.505000 ;
      RECT 215.205000  60.665000 215.875000  60.835000 ;
      RECT 215.205000  61.505000 215.575000  67.585000 ;
      RECT 215.275000 101.900000 216.125000 108.735000 ;
      RECT 215.375000  44.585000 215.915000  44.740000 ;
      RECT 215.375000  44.740000 215.675000  45.375000 ;
      RECT 215.375000  45.375000 215.915000  45.665000 ;
      RECT 215.375000  52.505000 215.915000  52.795000 ;
      RECT 215.375000  52.795000 215.675000  53.430000 ;
      RECT 215.375000  53.430000 215.915000  53.585000 ;
      RECT 215.385000  42.400000 215.915000  42.570000 ;
      RECT 215.385000  55.600000 215.915000  55.770000 ;
      RECT 215.505000  42.570000 215.915000  44.585000 ;
      RECT 215.505000  53.585000 215.915000  55.600000 ;
      RECT 215.585000  48.635000 216.755000  48.655000 ;
      RECT 215.625000  45.665000 215.915000  48.085000 ;
      RECT 215.625000  50.085000 215.915000  52.505000 ;
      RECT 215.745000  61.800000 215.915000  67.420000 ;
      RECT 215.845000  45.000000 216.375000  45.170000 ;
      RECT 215.845000  53.000000 216.375000  53.170000 ;
      RECT 215.910000 173.755000 217.600000 173.925000 ;
      RECT 215.910000 174.150000 217.600000 174.320000 ;
      RECT 215.910000 181.435000 217.600000 184.885000 ;
      RECT 215.915000 173.925000 217.600000 174.150000 ;
      RECT 215.915000 174.320000 217.600000 174.355000 ;
      RECT 215.925000  61.415000 216.525000  61.505000 ;
      RECT 215.925000  61.505000 216.455000  61.585000 ;
      RECT 215.930000  38.180000 216.235000  40.890000 ;
      RECT 215.930000  57.280000 216.235000  59.990000 ;
      RECT 216.015000  61.175000 216.525000  61.415000 ;
      RECT 216.015000  67.585000 216.525000  67.915000 ;
      RECT 216.065000  40.890000 216.235000  41.580000 ;
      RECT 216.065000  41.580000 216.280000  41.635000 ;
      RECT 216.065000  41.635000 216.315000  42.305000 ;
      RECT 216.065000  55.865000 216.315000  56.535000 ;
      RECT 216.065000  56.535000 216.280000  56.590000 ;
      RECT 216.065000  56.590000 216.235000  57.280000 ;
      RECT 216.085000  43.405000 216.280000  44.415000 ;
      RECT 216.085000  45.170000 216.255000  48.085000 ;
      RECT 216.085000  50.085000 216.255000  53.000000 ;
      RECT 216.085000  53.755000 216.280000  54.765000 ;
      RECT 216.085000  61.585000 216.455000  67.585000 ;
      RECT 216.110000  42.305000 216.280000  43.405000 ;
      RECT 216.110000  54.765000 216.280000  55.865000 ;
      RECT 216.110000  82.170000 216.280000  85.650000 ;
      RECT 216.125000  95.995000 222.875000  96.030000 ;
      RECT 216.155000  37.335000 216.825000  37.505000 ;
      RECT 216.155000  60.665000 216.825000  60.835000 ;
      RECT 216.210000  80.165000 216.380000  80.660000 ;
      RECT 216.210000  80.660000 217.160000  81.175000 ;
      RECT 216.225000  60.835000 216.755000  60.885000 ;
      RECT 216.290000  77.480000 219.340000  78.010000 ;
      RECT 216.290000  81.370000 216.820000  81.940000 ;
      RECT 216.330000  75.265000 219.220000  77.480000 ;
      RECT 216.330000  78.010000 219.220000  79.185000 ;
      RECT 216.405000  41.290000 217.075000  41.460000 ;
      RECT 216.405000  56.710000 217.075000  56.880000 ;
      RECT 216.485000  41.460000 216.980000  42.030000 ;
      RECT 216.485000  42.030000 217.015000  42.200000 ;
      RECT 216.485000  55.970000 217.015000  56.140000 ;
      RECT 216.485000  56.140000 216.980000  56.710000 ;
      RECT 216.545000  43.405000 217.195000  44.415000 ;
      RECT 216.545000  44.415000 216.715000  46.335000 ;
      RECT 216.545000  46.335000 217.075000  46.505000 ;
      RECT 216.545000  46.505000 216.715000  48.085000 ;
      RECT 216.545000  50.085000 216.715000  51.665000 ;
      RECT 216.545000  51.665000 217.075000  51.835000 ;
      RECT 216.545000  51.835000 216.715000  53.755000 ;
      RECT 216.545000  53.755000 217.195000  54.765000 ;
      RECT 216.555000   6.495000 220.930000   7.195000 ;
      RECT 216.555000   7.195000 217.255000  14.325000 ;
      RECT 216.555000  14.325000 220.930000  15.035000 ;
      RECT 216.555000  17.255000 220.930000  17.965000 ;
      RECT 216.555000  17.965000 217.255000  25.095000 ;
      RECT 216.555000  25.095000 220.930000  25.795000 ;
      RECT 216.565000  35.165000 217.095000  35.335000 ;
      RECT 216.565000  36.975000 216.735000  37.335000 ;
      RECT 216.595000 244.805000 222.345000 245.655000 ;
      RECT 216.595000 245.655000 217.445000 250.435000 ;
      RECT 216.595000 250.435000 222.345000 251.715000 ;
      RECT 216.625000  61.675000 216.795000  62.740000 ;
      RECT 216.625000  62.910000 216.795000  63.285000 ;
      RECT 216.625000  63.905000 216.795000  64.235000 ;
      RECT 216.625000  64.405000 216.795000  67.115000 ;
      RECT 216.715000  32.125000 216.885000  32.135000 ;
      RECT 216.715000  32.135000 217.435000  33.645000 ;
      RECT 216.715000  33.815000 217.435000  34.145000 ;
      RECT 216.715000  34.145000 216.885000  35.165000 ;
      RECT 216.785000 251.715000 222.155000 251.845000 ;
      RECT 216.810000  38.180000 216.980000  41.290000 ;
      RECT 216.810000  56.880000 216.980000  59.990000 ;
      RECT 216.885000  47.855000 217.055000  48.465000 ;
      RECT 216.885000  49.705000 217.055000  50.315000 ;
      RECT 216.895000  61.175000 217.405000  61.505000 ;
      RECT 216.895000  67.585000 217.405000  67.915000 ;
      RECT 216.930000 192.395000 217.600000 192.565000 ;
      RECT 216.935000  97.825000 223.185000  98.675000 ;
      RECT 216.935000  98.675000 217.785000 106.775000 ;
      RECT 216.935000 106.775000 223.185000 107.625000 ;
      RECT 216.965000  61.505000 217.335000  67.585000 ;
      RECT 216.990000  81.175000 217.160000  85.090000 ;
      RECT 217.025000  42.475000 219.685000  42.645000 ;
      RECT 217.025000  42.645000 217.195000  43.405000 ;
      RECT 217.025000  54.765000 217.195000  55.525000 ;
      RECT 217.025000  55.525000 219.685000  55.695000 ;
      RECT 217.035000  37.335000 219.065000  37.505000 ;
      RECT 217.035000  60.665000 219.065000  60.835000 ;
      RECT 217.055000 196.425000 344.705000 197.275000 ;
      RECT 217.055000 197.275000 217.905000 207.370000 ;
      RECT 217.055000 207.370000 219.825000 218.740000 ;
      RECT 217.055000 218.740000 231.675000 219.215000 ;
      RECT 217.055000 219.215000 346.520000 220.065000 ;
      RECT 217.055000 220.065000 217.905000 241.585000 ;
      RECT 217.055000 241.585000 225.565000 242.435000 ;
      RECT 217.085000 113.910000 220.085000 164.900000 ;
      RECT 217.245000  41.360000 217.775000  41.530000 ;
      RECT 217.245000  56.640000 217.775000  56.810000 ;
      RECT 217.265000  34.315000 217.435000  35.325000 ;
      RECT 217.330000  81.285000 217.840000  81.615000 ;
      RECT 217.330000  81.615000 217.700000  84.930000 ;
      RECT 217.365000  43.095000 217.895000  43.265000 ;
      RECT 217.365000  43.265000 217.535000  48.390000 ;
      RECT 217.365000  49.780000 217.535000  54.905000 ;
      RECT 217.365000  54.905000 217.895000  55.075000 ;
      RECT 217.425000  41.530000 217.595000  42.305000 ;
      RECT 217.425000  55.865000 217.595000  56.640000 ;
      RECT 217.505000  61.800000 217.675000  67.420000 ;
      RECT 217.605000  31.635000 217.775000  35.825000 ;
      RECT 217.685000 246.350000 217.855000 249.820000 ;
      RECT 217.690000  38.180000 217.950000  41.160000 ;
      RECT 217.690000  57.010000 217.950000  59.990000 ;
      RECT 217.705000  44.180000 219.525000  44.350000 ;
      RECT 217.705000  44.350000 217.895000  47.370000 ;
      RECT 217.705000  47.370000 218.235000  48.550000 ;
      RECT 217.705000  48.550000 220.595000  48.720000 ;
      RECT 217.705000  49.450000 220.595000  49.620000 ;
      RECT 217.705000  49.620000 218.235000  50.800000 ;
      RECT 217.705000  50.800000 217.895000  53.820000 ;
      RECT 217.705000  53.820000 219.525000  53.990000 ;
      RECT 217.740000   8.065000 218.280000  13.460000 ;
      RECT 217.740000  18.830000 218.280000  24.225000 ;
      RECT 217.775000  61.175000 218.285000  61.505000 ;
      RECT 217.775000  67.585000 218.285000  67.915000 ;
      RECT 217.845000  61.505000 218.215000  63.695000 ;
      RECT 217.845000  63.695000 218.375000  63.865000 ;
      RECT 217.845000  63.865000 218.215000  67.585000 ;
      RECT 217.870000  82.170000 218.040000  85.650000 ;
      RECT 217.945000  35.995000 219.565000  36.165000 ;
      RECT 217.965000  99.215000 218.270000 106.140000 ;
      RECT 217.970000  79.540000 218.140000  81.175000 ;
      RECT 217.975000  31.635000 218.145000  35.995000 ;
      RECT 218.045000 246.125000 220.755000 246.295000 ;
      RECT 218.045000 246.905000 220.755000 247.075000 ;
      RECT 218.045000 247.685000 220.755000 247.855000 ;
      RECT 218.045000 248.235000 220.755000 248.405000 ;
      RECT 218.045000 249.015000 220.755000 249.185000 ;
      RECT 218.045000 249.795000 220.755000 249.965000 ;
      RECT 218.065000  42.840000 218.235000  44.010000 ;
      RECT 218.065000  44.580000 218.235000  45.280000 ;
      RECT 218.065000  45.280000 218.595000  45.450000 ;
      RECT 218.065000  45.450000 218.235000  47.080000 ;
      RECT 218.065000  51.090000 218.235000  52.720000 ;
      RECT 218.065000  52.720000 218.595000  52.890000 ;
      RECT 218.065000  52.890000 218.235000  53.590000 ;
      RECT 218.065000  54.160000 218.235000  55.330000 ;
      RECT 218.085000  13.630000 219.410000  14.040000 ;
      RECT 218.085000  18.250000 219.410000  18.660000 ;
      RECT 218.150000  38.180000 218.410000  41.160000 ;
      RECT 218.150000  57.010000 218.410000  59.990000 ;
      RECT 218.210000 192.395000 218.880000 192.565000 ;
      RECT 218.220000  81.370000 218.730000  81.700000 ;
      RECT 218.225000 173.655000 220.245000 174.405000 ;
      RECT 218.225000 184.235000 220.245000 184.985000 ;
      RECT 218.310000  80.660000 218.680000  81.370000 ;
      RECT 218.335000  42.470000 219.685000  42.475000 ;
      RECT 218.335000  55.695000 219.685000  55.700000 ;
      RECT 218.345000  31.635000 219.195000  31.965000 ;
      RECT 218.345000  31.965000 218.515000  35.495000 ;
      RECT 218.345000  35.495000 219.195000  35.825000 ;
      RECT 218.385000  61.675000 218.555000  63.495000 ;
      RECT 218.385000  64.405000 218.555000  67.115000 ;
      RECT 218.420000  68.885000 218.590000  72.535000 ;
      RECT 218.420000  72.535000 218.950000  72.705000 ;
      RECT 218.420000  72.705000 218.590000  73.635000 ;
      RECT 218.480000 101.195000 221.405000 101.365000 ;
      RECT 218.485000 100.415000 221.405000 100.585000 ;
      RECT 218.495000  42.840000 218.665000  44.180000 ;
      RECT 218.495000  53.990000 218.665000  55.330000 ;
      RECT 218.515000  99.085000 221.405000  99.255000 ;
      RECT 218.515000  99.865000 221.405000 100.035000 ;
      RECT 218.515000 101.975000 221.405000 102.145000 ;
      RECT 218.540000 102.525000 221.405000 102.695000 ;
      RECT 218.540000 103.305000 221.405000 103.475000 ;
      RECT 218.540000 104.085000 221.405000 104.255000 ;
      RECT 218.540000 104.635000 221.405000 104.805000 ;
      RECT 218.540000 105.415000 221.405000 105.585000 ;
      RECT 218.540000 106.195000 221.405000 106.365000 ;
      RECT 218.545000  46.335000 219.075000  47.370000 ;
      RECT 218.545000  47.370000 219.415000  48.380000 ;
      RECT 218.545000  49.790000 219.415000  50.800000 ;
      RECT 218.545000  50.800000 219.075000  51.835000 ;
      RECT 218.665000  73.855000 220.015000  74.170000 ;
      RECT 218.665000 198.065000 229.315000 198.235000 ;
      RECT 218.665000 198.235000 218.835000 206.440000 ;
      RECT 218.665000 206.440000 225.035000 206.610000 ;
      RECT 218.665000 221.045000 218.835000 240.355000 ;
      RECT 218.665000 240.355000 225.625000 240.525000 ;
      RECT 218.685000  32.135000 218.855000  33.645000 ;
      RECT 218.685000  33.815000 218.855000  34.145000 ;
      RECT 218.685000  34.315000 218.855000  35.325000 ;
      RECT 218.750000  82.380000 219.070000  85.090000 ;
      RECT 218.850000  80.165000 219.070000  81.175000 ;
      RECT 218.900000  81.175000 219.070000  82.380000 ;
      RECT 218.925000  42.840000 219.095000  44.010000 ;
      RECT 218.925000  54.160000 219.095000  55.330000 ;
      RECT 218.935000  61.675000 219.105000  63.495000 ;
      RECT 218.935000  64.405000 219.105000  67.115000 ;
      RECT 219.005000 220.235000 220.745000 220.765000 ;
      RECT 219.005000 220.765000 219.365000 222.010000 ;
      RECT 219.025000  31.965000 219.195000  35.495000 ;
      RECT 219.025000 198.930000 219.195000 199.005000 ;
      RECT 219.025000 199.005000 219.320000 200.255000 ;
      RECT 219.025000 200.255000 219.195000 200.280000 ;
      RECT 219.025000 200.970000 219.195000 201.020000 ;
      RECT 219.025000 201.020000 219.320000 202.270000 ;
      RECT 219.025000 202.270000 219.195000 202.320000 ;
      RECT 219.025000 203.150000 219.330000 203.820000 ;
      RECT 219.025000 204.480000 219.330000 205.760000 ;
      RECT 219.120000  38.010000 219.290000  41.360000 ;
      RECT 219.120000  41.360000 219.650000  41.530000 ;
      RECT 219.120000  56.640000 219.650000  56.810000 ;
      RECT 219.120000  56.810000 219.290000  60.160000 ;
      RECT 219.120000 234.695000 219.365000 236.485000 ;
      RECT 219.120000 236.485000 224.675000 236.655000 ;
      RECT 219.130000 204.205000 219.300000 204.480000 ;
      RECT 219.145000  70.685000 219.370000  71.225000 ;
      RECT 219.200000  68.885000 219.370000  70.685000 ;
      RECT 219.200000  71.225000 219.370000  73.635000 ;
      RECT 219.205000  61.175000 219.715000  61.505000 ;
      RECT 219.205000  67.585000 219.715000  67.915000 ;
      RECT 219.215000   8.065000 219.755000  13.460000 ;
      RECT 219.215000  18.830000 219.755000  24.225000 ;
      RECT 219.245000  44.580000 219.415000  45.760000 ;
      RECT 219.245000  45.760000 221.775000  45.930000 ;
      RECT 219.245000  45.930000 219.415000  47.080000 ;
      RECT 219.245000  51.090000 219.415000  52.240000 ;
      RECT 219.245000  52.240000 221.775000  52.410000 ;
      RECT 219.245000  52.410000 219.415000  53.590000 ;
      RECT 219.275000  61.505000 219.645000  67.585000 ;
      RECT 219.275000  86.320000 234.280000  86.375000 ;
      RECT 219.300000  82.050000 219.470000  86.210000 ;
      RECT 219.300000  86.210000 234.280000  86.320000 ;
      RECT 219.355000  42.840000 219.525000  44.180000 ;
      RECT 219.355000  53.990000 219.525000  55.330000 ;
      RECT 219.395000  31.635000 219.565000  35.995000 ;
      RECT 219.490000 186.225000 220.160000 188.785000 ;
      RECT 219.490000 189.915000 220.160000 192.565000 ;
      RECT 219.530000  75.275000 236.800000  75.525000 ;
      RECT 219.530000  75.525000 219.700000  79.145000 ;
      RECT 219.535000 221.045000 248.345000 221.215000 ;
      RECT 219.535000 221.465000 224.285000 222.075000 ;
      RECT 219.535000 222.245000 224.285000 222.855000 ;
      RECT 219.535000 223.025000 224.285000 223.635000 ;
      RECT 219.535000 223.805000 224.285000 224.415000 ;
      RECT 219.535000 224.585000 224.285000 225.195000 ;
      RECT 219.535000 225.365000 224.285000 225.975000 ;
      RECT 219.535000 226.145000 224.285000 226.755000 ;
      RECT 219.535000 226.925000 224.285000 227.535000 ;
      RECT 219.535000 227.705000 224.285000 228.200000 ;
      RECT 219.535000 235.940000 224.285000 236.215000 ;
      RECT 219.535000 236.825000 224.285000 237.215000 ;
      RECT 219.535000 237.385000 224.285000 237.880000 ;
      RECT 219.535000 238.050000 224.285000 238.545000 ;
      RECT 219.535000 238.715000 224.285000 239.325000 ;
      RECT 219.535000 239.495000 224.285000 239.990000 ;
      RECT 219.580000 198.705000 224.455000 198.875000 ;
      RECT 219.580000 199.485000 224.455000 199.655000 ;
      RECT 219.580000 200.265000 224.455000 200.435000 ;
      RECT 219.580000 200.815000 224.455000 200.985000 ;
      RECT 219.580000 201.595000 224.455000 201.765000 ;
      RECT 219.580000 202.375000 224.455000 202.545000 ;
      RECT 219.580000 202.925000 224.455000 203.095000 ;
      RECT 219.580000 203.705000 224.455000 203.875000 ;
      RECT 219.580000 205.035000 224.455000 205.205000 ;
      RECT 219.585000 204.255000 224.455000 204.425000 ;
      RECT 219.585000 205.815000 224.455000 205.985000 ;
      RECT 219.620000  69.905000 220.150000  70.075000 ;
      RECT 219.630000 236.215000 224.120000 236.315000 ;
      RECT 219.695000  83.405000 219.865000  83.660000 ;
      RECT 219.695000  83.660000 220.225000  83.830000 ;
      RECT 219.695000  83.830000 219.865000  84.415000 ;
      RECT 219.700000  37.870000 219.870000  40.870000 ;
      RECT 219.700000  57.300000 219.870000  60.300000 ;
      RECT 219.765000  31.635000 219.935000  35.825000 ;
      RECT 219.765000  46.165000 220.095000  47.015000 ;
      RECT 219.765000  51.155000 220.095000  52.005000 ;
      RECT 219.785000  42.840000 219.955000  44.010000 ;
      RECT 219.785000  54.160000 219.955000  55.330000 ;
      RECT 219.815000  61.800000 219.985000  67.420000 ;
      RECT 219.845000  47.015000 220.015000  47.625000 ;
      RECT 219.845000  50.545000 220.015000  51.155000 ;
      RECT 219.850000  79.240000 220.760000  79.310000 ;
      RECT 219.850000  79.310000 220.250000  83.060000 ;
      RECT 219.850000 228.370000 222.825000 228.865000 ;
      RECT 219.850000 229.815000 222.825000 230.425000 ;
      RECT 219.850000 231.375000 222.825000 231.985000 ;
      RECT 219.850000 232.935000 222.825000 233.545000 ;
      RECT 219.850000 234.495000 222.825000 234.990000 ;
      RECT 219.850000 235.275000 223.315000 235.770000 ;
      RECT 219.870000  79.140000 220.760000  79.240000 ;
      RECT 219.920000  45.280000 220.595000  45.450000 ;
      RECT 219.920000  52.720000 220.595000  52.890000 ;
      RECT 219.980000  68.885000 220.150000  69.905000 ;
      RECT 219.980000  70.075000 220.150000  73.635000 ;
      RECT 220.040000  42.470000 221.390000  42.640000 ;
      RECT 220.040000  42.640000 221.290000  42.670000 ;
      RECT 220.040000  55.500000 221.290000  55.530000 ;
      RECT 220.040000  55.530000 221.390000  55.700000 ;
      RECT 220.055000  84.030000 220.645000  84.200000 ;
      RECT 220.080000  84.555000 220.250000  85.565000 ;
      RECT 220.085000  61.175000 220.595000  61.505000 ;
      RECT 220.085000  67.585000 220.595000  67.915000 ;
      RECT 220.105000  32.135000 220.825000  33.645000 ;
      RECT 220.105000  33.815000 220.825000  34.145000 ;
      RECT 220.105000  34.315000 220.275000  35.325000 ;
      RECT 220.115000 229.035000 222.825000 229.645000 ;
      RECT 220.115000 230.595000 222.825000 231.205000 ;
      RECT 220.115000 232.155000 222.825000 232.765000 ;
      RECT 220.115000 233.715000 222.825000 234.325000 ;
      RECT 220.120000  76.165000 220.290000  78.340000 ;
      RECT 220.120000  78.340000 220.650000  78.510000 ;
      RECT 220.120000  78.510000 220.290000  78.875000 ;
      RECT 220.155000  61.505000 220.525000  67.585000 ;
      RECT 220.215000  42.840000 220.385000  44.180000 ;
      RECT 220.215000  44.180000 221.775000  44.350000 ;
      RECT 220.215000  53.820000 221.775000  53.990000 ;
      RECT 220.215000  53.990000 220.385000  55.330000 ;
      RECT 220.230000   7.195000 220.930000  14.325000 ;
      RECT 220.230000  17.965000 220.930000  25.095000 ;
      RECT 220.300000  85.850000 220.830000  86.020000 ;
      RECT 220.415000  75.775000 223.415000  75.945000 ;
      RECT 220.420000  84.615000 221.080000  85.575000 ;
      RECT 220.420000  85.575000 220.830000  85.850000 ;
      RECT 220.425000  44.580000 220.595000  45.280000 ;
      RECT 220.425000  45.450000 220.595000  45.590000 ;
      RECT 220.425000  46.100000 220.595000  48.550000 ;
      RECT 220.425000  49.620000 220.595000  52.070000 ;
      RECT 220.425000  52.580000 220.595000  52.720000 ;
      RECT 220.425000  52.890000 220.595000  53.590000 ;
      RECT 220.475000  81.395000 221.665000  81.565000 ;
      RECT 220.475000  81.565000 220.645000  84.030000 ;
      RECT 220.475000  84.200000 220.645000  84.415000 ;
      RECT 220.530000  68.205000 223.765000  68.375000 ;
      RECT 220.530000  68.375000 220.700000  71.015000 ;
      RECT 220.530000  71.015000 221.060000  71.185000 ;
      RECT 220.530000  71.185000 220.700000  73.635000 ;
      RECT 220.585000 206.610000 220.755000 217.810000 ;
      RECT 220.585000 217.810000 225.035000 217.980000 ;
      RECT 220.645000  42.840000 220.815000  44.010000 ;
      RECT 220.645000  54.160000 220.815000  55.330000 ;
      RECT 220.655000  32.125000 220.825000  32.135000 ;
      RECT 220.655000  34.145000 220.825000  35.165000 ;
      RECT 220.655000  35.165000 221.185000  35.335000 ;
      RECT 220.695000  61.675000 220.865000  62.740000 ;
      RECT 220.695000  62.910000 220.865000  63.285000 ;
      RECT 220.695000  63.905000 220.865000  64.235000 ;
      RECT 220.695000  64.405000 220.865000  67.115000 ;
      RECT 220.780000 173.755000 221.450000 173.925000 ;
      RECT 220.780000 174.115000 221.450000 174.285000 ;
      RECT 220.780000 175.785000 221.450000 175.955000 ;
      RECT 220.780000 176.325000 221.450000 176.495000 ;
      RECT 220.780000 177.995000 221.450000 178.165000 ;
      RECT 220.780000 178.535000 221.450000 178.705000 ;
      RECT 220.780000 180.205000 221.450000 180.375000 ;
      RECT 220.780000 180.745000 221.450000 180.915000 ;
      RECT 220.780000 182.415000 221.450000 188.785000 ;
      RECT 220.780000 189.915000 221.450000 192.565000 ;
      RECT 220.850000 173.705000 221.380000 173.755000 ;
      RECT 220.860000  82.050000 221.135000  83.060000 ;
      RECT 220.860000  83.060000 221.080000  84.615000 ;
      RECT 220.865000 192.875000 222.730000 193.405000 ;
      RECT 220.865000 193.605000 226.570000 194.135000 ;
      RECT 220.900000  75.945000 221.070000  78.875000 ;
      RECT 220.965000  79.540000 221.135000  80.985000 ;
      RECT 220.990000  61.385000 221.545000  61.505000 ;
      RECT 220.990000  61.505000 221.520000  61.555000 ;
      RECT 221.000000  85.870000 221.670000  86.040000 ;
      RECT 221.035000  61.175000 221.545000  61.385000 ;
      RECT 221.035000  67.585000 221.545000  67.915000 ;
      RECT 221.045000  37.765000 221.215000  40.845000 ;
      RECT 221.045000  57.325000 221.215000  60.405000 ;
      RECT 221.075000  42.840000 221.245000  44.180000 ;
      RECT 221.075000  53.990000 221.245000  55.330000 ;
      RECT 221.105000  61.555000 221.475000  67.585000 ;
      RECT 221.125000  69.905000 221.655000  70.075000 ;
      RECT 221.165000 207.380000 221.335000 217.230000 ;
      RECT 221.245000  46.335000 221.775000  46.505000 ;
      RECT 221.245000  51.665000 221.775000  51.835000 ;
      RECT 221.250000  84.485000 221.420000  85.870000 ;
      RECT 221.310000  68.885000 221.480000  69.905000 ;
      RECT 221.310000  70.075000 221.480000  74.525000 ;
      RECT 221.330000  83.310000 222.680000  83.480000 ;
      RECT 221.370000  41.265000 222.335000  41.435000 ;
      RECT 221.370000  41.435000 221.680000  42.130000 ;
      RECT 221.370000  42.130000 221.900000  42.300000 ;
      RECT 221.370000  55.870000 221.900000  56.040000 ;
      RECT 221.370000  56.040000 221.680000  56.735000 ;
      RECT 221.370000  56.735000 222.335000  56.905000 ;
      RECT 221.455000 206.800000 224.165000 206.980000 ;
      RECT 221.455000 217.440000 224.165000 217.620000 ;
      RECT 221.470000 113.195000 222.140000 113.525000 ;
      RECT 221.495000 245.655000 222.345000 250.435000 ;
      RECT 221.505000  42.840000 221.675000  44.010000 ;
      RECT 221.505000  54.160000 221.675000  55.330000 ;
      RECT 221.505000 206.980000 221.775000 217.440000 ;
      RECT 221.510000  38.155000 221.795000  40.865000 ;
      RECT 221.510000  40.865000 221.680000  41.095000 ;
      RECT 221.510000  57.075000 221.680000  57.305000 ;
      RECT 221.510000  57.305000 221.795000  60.015000 ;
      RECT 221.510000  78.340000 222.040000  78.510000 ;
      RECT 221.555000  83.735000 222.085000  84.070000 ;
      RECT 221.555000  84.070000 222.445000  84.240000 ;
      RECT 221.560000  31.595000 224.175000  31.765000 ;
      RECT 221.560000  32.710000 223.475000  32.785000 ;
      RECT 221.560000  32.785000 222.450000  33.600000 ;
      RECT 221.560000  35.565000 222.450000  35.945000 ;
      RECT 221.560000  35.945000 232.945000  36.455000 ;
      RECT 221.580000  28.555000 270.960000  29.190000 ;
      RECT 221.580000  29.190000 225.455000  30.145000 ;
      RECT 221.580000  30.145000 226.035000  31.485000 ;
      RECT 221.580000  31.485000 224.175000  31.595000 ;
      RECT 221.580000  31.765000 223.475000  32.710000 ;
      RECT 221.580000  33.600000 222.430000  35.565000 ;
      RECT 221.595000 113.910000 224.595000 164.900000 ;
      RECT 221.605000  44.350000 221.775000  45.760000 ;
      RECT 221.605000  46.100000 221.775000  46.335000 ;
      RECT 221.605000  46.505000 221.775000  48.380000 ;
      RECT 221.605000  49.790000 221.775000  51.665000 ;
      RECT 221.605000  51.835000 221.775000  52.070000 ;
      RECT 221.605000  52.410000 221.775000  53.820000 ;
      RECT 221.605000  74.745000 229.415000  74.915000 ;
      RECT 221.640000  84.555000 221.810000  84.595000 ;
      RECT 221.640000  84.595000 222.250000  84.765000 ;
      RECT 221.640000  84.765000 221.810000  85.565000 ;
      RECT 221.645000  61.675000 221.815000  66.145000 ;
      RECT 221.680000  76.165000 221.850000  78.340000 ;
      RECT 221.680000  78.510000 221.850000  78.875000 ;
      RECT 221.690000   5.735000 222.390000  15.795000 ;
      RECT 221.690000  16.495000 222.390000  26.555000 ;
      RECT 221.850000  37.335000 224.105000  37.505000 ;
      RECT 221.850000  41.085000 222.520000  41.255000 ;
      RECT 221.850000  41.255000 222.335000  41.265000 ;
      RECT 221.850000  41.760000 222.380000  41.930000 ;
      RECT 221.850000  56.240000 222.380000  56.410000 ;
      RECT 221.850000  56.905000 222.335000  56.915000 ;
      RECT 221.850000  56.915000 222.520000  57.085000 ;
      RECT 221.850000  60.665000 224.105000  60.835000 ;
      RECT 221.875000  81.480000 222.545000  81.650000 ;
      RECT 221.895000  67.115000 222.425000  67.285000 ;
      RECT 221.900000  71.015000 222.430000  71.185000 ;
      RECT 221.915000  61.175000 222.425000  61.505000 ;
      RECT 221.915000  67.585000 222.425000  67.915000 ;
      RECT 221.945000 207.380000 222.115000 217.230000 ;
      RECT 221.955000  81.395000 222.485000  81.480000 ;
      RECT 221.965000  37.505000 224.105000  37.595000 ;
      RECT 221.965000  37.595000 222.335000  41.085000 ;
      RECT 221.965000  43.110000 222.495000  43.280000 ;
      RECT 221.965000  54.890000 222.495000  55.060000 ;
      RECT 221.965000  57.085000 222.335000  60.575000 ;
      RECT 221.965000  60.575000 224.105000  60.665000 ;
      RECT 221.975000   0.710000 228.165000   0.880000 ;
      RECT 221.975000   0.880000 222.145000   5.035000 ;
      RECT 221.985000  61.505000 222.355000  67.115000 ;
      RECT 221.985000  67.285000 222.355000  67.585000 ;
      RECT 222.045000  81.820000 222.575000  81.990000 ;
      RECT 222.045000  81.990000 222.215000  83.060000 ;
      RECT 222.060000 192.395000 222.730000 192.875000 ;
      RECT 222.070000  41.930000 222.380000  43.110000 ;
      RECT 222.070000  55.060000 222.380000  56.240000 ;
      RECT 222.090000  68.375000 222.260000  71.015000 ;
      RECT 222.090000  71.185000 222.260000  73.635000 ;
      RECT 222.185000  43.280000 222.355000  48.390000 ;
      RECT 222.185000  49.780000 222.355000  54.890000 ;
      RECT 222.285000 206.980000 222.555000 217.440000 ;
      RECT 222.335000  98.675000 223.185000 106.775000 ;
      RECT 222.420000  84.555000 222.590000  86.210000 ;
      RECT 222.460000  75.945000 222.630000  78.875000 ;
      RECT 222.505000  37.765000 222.675000  40.865000 ;
      RECT 222.505000  57.305000 222.675000  60.405000 ;
      RECT 222.550000  41.445000 223.015000  41.615000 ;
      RECT 222.550000  41.615000 222.720000  42.520000 ;
      RECT 222.550000  42.520000 222.835000  42.690000 ;
      RECT 222.550000  55.480000 222.835000  55.650000 ;
      RECT 222.550000  55.650000 222.720000  56.555000 ;
      RECT 222.550000  56.555000 223.015000  56.725000 ;
      RECT 222.595000  61.675000 222.765000  62.725000 ;
      RECT 222.595000  62.955000 222.765000  63.285000 ;
      RECT 222.595000  63.905000 222.765000  64.235000 ;
      RECT 222.595000  64.405000 222.765000  67.420000 ;
      RECT 222.665000  42.690000 222.835000  43.615000 ;
      RECT 222.665000  54.555000 222.835000  55.480000 ;
      RECT 222.680000  69.905000 223.210000  70.075000 ;
      RECT 222.725000 207.380000 222.895000 217.230000 ;
      RECT 222.755000  81.395000 223.425000  81.565000 ;
      RECT 222.845000  40.395000 223.555000  40.865000 ;
      RECT 222.845000  40.865000 223.015000  41.445000 ;
      RECT 222.845000  56.725000 223.015000  57.305000 ;
      RECT 222.845000  57.305000 223.555000  57.775000 ;
      RECT 222.870000  68.885000 223.040000  69.905000 ;
      RECT 222.870000  70.075000 223.040000  73.635000 ;
      RECT 222.880000  78.340000 223.410000  78.510000 ;
      RECT 222.890000  41.785000 223.510000  42.115000 ;
      RECT 222.890000  56.055000 223.510000  56.385000 ;
      RECT 222.900000  84.745000 229.690000  84.915000 ;
      RECT 222.905000   1.640000 227.235000   1.810000 ;
      RECT 222.905000   1.810000 223.075000   4.080000 ;
      RECT 222.905000   4.080000 227.235000   4.250000 ;
      RECT 222.995000 228.700000 223.315000 235.275000 ;
      RECT 223.065000  82.050000 223.435000  83.895000 ;
      RECT 223.065000  83.895000 226.540000  84.405000 ;
      RECT 223.065000 206.980000 223.335000 217.440000 ;
      RECT 223.105000 244.045000 223.955000 252.535000 ;
      RECT 223.115000  48.350000 226.485000  48.520000 ;
      RECT 223.115000  49.650000 226.485000  49.820000 ;
      RECT 223.145000  61.675000 223.315000  63.495000 ;
      RECT 223.145000  64.405000 223.315000  67.115000 ;
      RECT 223.150000   6.495000 227.525000   7.195000 ;
      RECT 223.150000   7.195000 223.850000  14.325000 ;
      RECT 223.150000  14.325000 227.525000  15.035000 ;
      RECT 223.150000  17.255000 227.525000  17.965000 ;
      RECT 223.150000  17.965000 223.850000  25.095000 ;
      RECT 223.150000  25.095000 227.525000  25.795000 ;
      RECT 223.155000  45.290000 223.325000  48.000000 ;
      RECT 223.155000  50.170000 223.325000  52.880000 ;
      RECT 223.185000  41.360000 224.105000  41.530000 ;
      RECT 223.185000  41.530000 223.510000  41.785000 ;
      RECT 223.185000  56.385000 223.510000  56.640000 ;
      RECT 223.185000  56.640000 224.105000  56.810000 ;
      RECT 223.210000  35.165000 231.785000  35.335000 ;
      RECT 223.240000  76.165000 223.410000  78.340000 ;
      RECT 223.240000  78.510000 223.410000  78.875000 ;
      RECT 223.275000  48.215000 226.325000  48.350000 ;
      RECT 223.275000  49.820000 226.325000  49.955000 ;
      RECT 223.285000  79.635000 223.455000  80.790000 ;
      RECT 223.285000  80.790000 227.875000  80.960000 ;
      RECT 223.285000  80.960000 223.455000  80.985000 ;
      RECT 223.305000  33.860000 223.475000  34.915000 ;
      RECT 223.315000   2.435000 223.485000   3.445000 ;
      RECT 223.325000  63.695000 223.855000  63.865000 ;
      RECT 223.385000  38.155000 223.555000  40.395000 ;
      RECT 223.385000  57.775000 223.555000  60.015000 ;
      RECT 223.415000  61.175000 223.925000  61.505000 ;
      RECT 223.415000  67.585000 223.925000  67.915000 ;
      RECT 223.460000  71.015000 223.990000  71.185000 ;
      RECT 223.485000  61.505000 223.855000  63.695000 ;
      RECT 223.485000  63.865000 223.855000  67.585000 ;
      RECT 223.485000 228.585000 224.335000 231.315000 ;
      RECT 223.485000 231.315000 225.015000 235.420000 ;
      RECT 223.505000 207.380000 223.675000 217.230000 ;
      RECT 223.545000  42.605000 223.715000  44.400000 ;
      RECT 223.545000  53.770000 223.715000  55.565000 ;
      RECT 223.560000  45.030000 224.105000  45.200000 ;
      RECT 223.560000  52.970000 224.105000  53.140000 ;
      RECT 223.595000  68.375000 223.765000  68.885000 ;
      RECT 223.595000  68.885000 223.820000  71.015000 ;
      RECT 223.595000  71.185000 223.820000  73.345000 ;
      RECT 223.605000  83.310000 224.955000  83.480000 ;
      RECT 223.650000  44.570000 224.660000  44.740000 ;
      RECT 223.650000  44.740000 224.180000  44.800000 ;
      RECT 223.650000  53.370000 224.180000  53.430000 ;
      RECT 223.650000  53.430000 224.660000  53.600000 ;
      RECT 223.650000  73.345000 223.820000  73.635000 ;
      RECT 223.725000  37.595000 224.105000  38.615000 ;
      RECT 223.725000  59.555000 224.105000  60.575000 ;
      RECT 223.765000  42.000000 224.435000  42.170000 ;
      RECT 223.765000  56.000000 224.435000  56.170000 ;
      RECT 223.790000  76.165000 223.960000  78.875000 ;
      RECT 223.835000  42.170000 224.365000  42.300000 ;
      RECT 223.835000  55.870000 224.365000  56.000000 ;
      RECT 223.835000  79.140000 224.640000  79.310000 ;
      RECT 223.835000  79.310000 224.005000  80.475000 ;
      RECT 223.845000 206.980000 224.115000 217.440000 ;
      RECT 223.935000  40.195000 224.105000  41.360000 ;
      RECT 223.935000  45.000000 224.105000  45.030000 ;
      RECT 223.935000  45.200000 224.105000  48.000000 ;
      RECT 223.935000  50.170000 224.105000  52.970000 ;
      RECT 223.935000  53.140000 224.105000  53.170000 ;
      RECT 223.935000  56.810000 224.105000  57.975000 ;
      RECT 223.935000  68.205000 226.645000  68.375000 ;
      RECT 223.950000  97.045000 235.725000 102.920000 ;
      RECT 223.950000 102.920000 271.970000 103.770000 ;
      RECT 223.950000 103.770000 236.175000 108.380000 ;
      RECT 223.950000 108.380000 271.970000 108.735000 ;
      RECT 224.005000   2.220000 226.765000   2.390000 ;
      RECT 224.005000   3.500000 226.715000   3.670000 ;
      RECT 224.025000  61.800000 224.195000  67.420000 ;
      RECT 224.030000 113.195000 224.700000 113.525000 ;
      RECT 224.035000  38.970000 225.565000  39.720000 ;
      RECT 224.035000  58.450000 225.565000  59.200000 ;
      RECT 224.065000  42.505000 224.595000  42.675000 ;
      RECT 224.065000  55.495000 224.595000  55.665000 ;
      RECT 224.085000  75.775000 226.795000  75.945000 ;
      RECT 224.175000  32.165000 224.755000  32.335000 ;
      RECT 224.205000  81.395000 224.795000  81.940000 ;
      RECT 224.205000  81.940000 224.375000  83.060000 ;
      RECT 224.245000  70.335000 224.775000  70.505000 ;
      RECT 224.275000  37.765000 225.325000  38.970000 ;
      RECT 224.275000  39.720000 225.325000  40.865000 ;
      RECT 224.275000  57.305000 225.325000  58.450000 ;
      RECT 224.275000  59.200000 225.325000  60.405000 ;
      RECT 224.285000 207.380000 224.455000 217.230000 ;
      RECT 224.295000  61.175000 224.805000  61.505000 ;
      RECT 224.295000  67.585000 224.805000  67.915000 ;
      RECT 224.325000   8.065000 224.865000  13.460000 ;
      RECT 224.325000  18.830000 224.865000  24.225000 ;
      RECT 224.365000  61.505000 224.735000  63.455000 ;
      RECT 224.365000  63.455000 224.985000  63.625000 ;
      RECT 224.365000  63.625000 224.735000  67.585000 ;
      RECT 224.395000  78.340000 224.925000  78.510000 ;
      RECT 224.425000  42.675000 224.595000  43.615000 ;
      RECT 224.425000  54.555000 224.595000  55.495000 ;
      RECT 224.430000  68.375000 224.600000  70.335000 ;
      RECT 224.430000  70.505000 224.600000  73.635000 ;
      RECT 224.485000  80.695000 227.875000  80.790000 ;
      RECT 224.485000  80.960000 227.875000  81.205000 ;
      RECT 224.505000 221.910000 224.810000 230.710000 ;
      RECT 224.505000 230.710000 227.505000 230.990000 ;
      RECT 224.505000 236.270000 224.675000 236.485000 ;
      RECT 224.505000 236.655000 224.675000 239.660000 ;
      RECT 224.570000  75.945000 224.740000  78.340000 ;
      RECT 224.570000  78.510000 224.740000  78.875000 ;
      RECT 224.585000  31.775000 224.755000  32.165000 ;
      RECT 224.585000  32.335000 224.755000  34.915000 ;
      RECT 224.670000  13.630000 225.995000  14.040000 ;
      RECT 224.670000  18.250000 225.995000  18.660000 ;
      RECT 224.715000  45.290000 224.885000  48.000000 ;
      RECT 224.715000  50.170000 224.885000  52.880000 ;
      RECT 224.715000 242.435000 225.565000 244.355000 ;
      RECT 224.715000 244.355000 236.945000 247.105000 ;
      RECT 224.715000 247.105000 346.520000 251.735000 ;
      RECT 224.865000 198.235000 225.035000 206.440000 ;
      RECT 224.865000 206.610000 225.035000 213.855000 ;
      RECT 224.865000 213.855000 229.315000 214.025000 ;
      RECT 224.865000 214.025000 225.035000 217.810000 ;
      RECT 224.905000  61.675000 225.075000  62.740000 ;
      RECT 224.905000  62.910000 225.075000  63.285000 ;
      RECT 224.905000  63.905000 225.075000  64.235000 ;
      RECT 224.905000  64.405000 225.075000  67.115000 ;
      RECT 224.925000  31.485000 226.035000  31.735000 ;
      RECT 224.925000  33.255000 226.615000  33.425000 ;
      RECT 224.940000  44.570000 225.950000  44.740000 ;
      RECT 224.940000  53.430000 225.950000  53.600000 ;
      RECT 224.980000 221.215000 227.080000 230.235000 ;
      RECT 225.005000  42.505000 225.535000  42.675000 ;
      RECT 225.005000  42.675000 225.175000  43.615000 ;
      RECT 225.005000  54.555000 225.175000  55.495000 ;
      RECT 225.005000  55.495000 225.535000  55.665000 ;
      RECT 225.020000  71.015000 225.550000  71.185000 ;
      RECT 225.125000  82.050000 225.910000  83.895000 ;
      RECT 225.165000  42.000000 225.835000  42.170000 ;
      RECT 225.165000  56.000000 225.835000  56.170000 ;
      RECT 225.165000  81.430000 227.875000  81.600000 ;
      RECT 225.175000  61.175000 225.685000  61.505000 ;
      RECT 225.175000  67.585000 225.685000  67.915000 ;
      RECT 225.185000 230.990000 226.075000 238.295000 ;
      RECT 225.210000  68.885000 225.380000  71.015000 ;
      RECT 225.210000  71.185000 225.380000  73.635000 ;
      RECT 225.235000  42.170000 225.765000  42.300000 ;
      RECT 225.235000  55.870000 225.765000  56.000000 ;
      RECT 225.245000  61.505000 225.615000  67.585000 ;
      RECT 225.350000  76.165000 225.520000  78.875000 ;
      RECT 225.420000  44.740000 225.950000  44.800000 ;
      RECT 225.420000  53.370000 225.950000  53.430000 ;
      RECT 225.445000 198.815000 225.615000 205.605000 ;
      RECT 225.445000 206.465000 225.615000 213.315000 ;
      RECT 225.455000 238.575000 248.345000 239.105000 ;
      RECT 225.455000 239.105000 225.625000 240.355000 ;
      RECT 225.495000  37.335000 227.750000  37.505000 ;
      RECT 225.495000  37.505000 227.635000  37.595000 ;
      RECT 225.495000  37.595000 225.875000  38.615000 ;
      RECT 225.495000  40.195000 225.665000  41.360000 ;
      RECT 225.495000  41.360000 226.415000  41.530000 ;
      RECT 225.495000  45.000000 225.665000  45.030000 ;
      RECT 225.495000  45.030000 226.040000  45.200000 ;
      RECT 225.495000  45.200000 225.665000  48.000000 ;
      RECT 225.495000  50.170000 225.665000  52.970000 ;
      RECT 225.495000  52.970000 226.040000  53.140000 ;
      RECT 225.495000  53.140000 225.665000  53.170000 ;
      RECT 225.495000  56.640000 226.415000  56.810000 ;
      RECT 225.495000  56.810000 225.665000  57.975000 ;
      RECT 225.495000  59.555000 225.875000  60.575000 ;
      RECT 225.495000  60.575000 227.635000  60.665000 ;
      RECT 225.495000  60.665000 227.750000  60.835000 ;
      RECT 225.735000 198.425000 228.445000 198.595000 ;
      RECT 225.735000 205.815000 228.445000 206.245000 ;
      RECT 225.785000  61.800000 225.955000  67.420000 ;
      RECT 225.785000 198.595000 226.055000 205.815000 ;
      RECT 225.795000 214.785000 231.675000 218.740000 ;
      RECT 225.800000   8.065000 226.340000  13.460000 ;
      RECT 225.800000  18.830000 226.340000  24.225000 ;
      RECT 225.800000  70.335000 226.330000  70.505000 ;
      RECT 225.850000 251.735000 346.520000 251.760000 ;
      RECT 225.865000  31.735000 226.035000  32.855000 ;
      RECT 225.865000  33.860000 226.035000  34.915000 ;
      RECT 225.885000  42.605000 226.055000  44.400000 ;
      RECT 225.885000  53.770000 226.055000  55.565000 ;
      RECT 225.900000 192.285000 226.570000 193.605000 ;
      RECT 225.960000  78.340000 226.490000  78.510000 ;
      RECT 225.990000  68.375000 226.160000  70.335000 ;
      RECT 225.990000  70.505000 226.160000  73.635000 ;
      RECT 226.045000  38.155000 226.215000  40.395000 ;
      RECT 226.045000  40.395000 226.755000  40.865000 ;
      RECT 226.045000  57.305000 226.755000  57.775000 ;
      RECT 226.045000  57.775000 226.215000  60.015000 ;
      RECT 226.055000  61.175000 226.565000  61.505000 ;
      RECT 226.055000  67.585000 226.655000  67.685000 ;
      RECT 226.055000  67.685000 226.565000  67.915000 ;
      RECT 226.090000  41.530000 226.415000  41.785000 ;
      RECT 226.090000  41.785000 226.710000  42.115000 ;
      RECT 226.090000  56.055000 226.710000  56.385000 ;
      RECT 226.090000  56.385000 226.415000  56.640000 ;
      RECT 226.105000 113.910000 229.105000 164.900000 ;
      RECT 226.110000  83.310000 226.780000  83.480000 ;
      RECT 226.125000  61.505000 226.495000  67.515000 ;
      RECT 226.125000  67.515000 226.655000  67.585000 ;
      RECT 226.130000  75.945000 226.300000  78.340000 ;
      RECT 226.130000  78.510000 226.300000  78.875000 ;
      RECT 226.195000  81.770000 226.725000  81.940000 ;
      RECT 226.215000 239.550000 228.040000 241.160000 ;
      RECT 226.215000 241.160000 227.870000 241.240000 ;
      RECT 226.215000 242.030000 228.620000 243.720000 ;
      RECT 226.225000 198.815000 226.395000 205.605000 ;
      RECT 226.225000 206.465000 226.395000 213.255000 ;
      RECT 226.245000 231.160000 227.070000 231.605000 ;
      RECT 226.245000 231.605000 248.345000 232.050000 ;
      RECT 226.245000 232.050000 227.070000 238.575000 ;
      RECT 226.275000  45.290000 226.445000  48.000000 ;
      RECT 226.275000  50.170000 226.445000  52.880000 ;
      RECT 226.300000  29.425000 226.970000  29.595000 ;
      RECT 226.365000  81.940000 226.535000  83.060000 ;
      RECT 226.380000  29.595000 226.910000  29.745000 ;
      RECT 226.410000  71.015000 226.940000  71.185000 ;
      RECT 226.565000 198.595000 226.835000 205.815000 ;
      RECT 226.585000  40.865000 226.755000  41.445000 ;
      RECT 226.585000  41.445000 227.050000  41.615000 ;
      RECT 226.585000  56.555000 227.050000  56.725000 ;
      RECT 226.585000  56.725000 226.755000  57.305000 ;
      RECT 226.665000  61.675000 226.835000  63.495000 ;
      RECT 226.665000  64.405000 226.835000  67.115000 ;
      RECT 226.765000  42.520000 227.050000  42.690000 ;
      RECT 226.765000  42.690000 226.935000  43.615000 ;
      RECT 226.765000  52.095000 226.935000  55.480000 ;
      RECT 226.765000  55.480000 227.050000  55.650000 ;
      RECT 226.770000  68.885000 226.940000  71.015000 ;
      RECT 226.770000  71.185000 226.940000  73.635000 ;
      RECT 226.825000   7.195000 227.525000  14.325000 ;
      RECT 226.825000  17.965000 227.525000  25.095000 ;
      RECT 226.880000  41.615000 227.050000  42.520000 ;
      RECT 226.880000  55.650000 227.050000  56.555000 ;
      RECT 226.910000  76.165000 227.080000  78.875000 ;
      RECT 226.925000  37.765000 227.095000  40.865000 ;
      RECT 226.925000  57.305000 227.095000  60.405000 ;
      RECT 226.965000  33.255000 227.495000  33.425000 ;
      RECT 226.980000  83.290000 229.310000  83.460000 ;
      RECT 226.980000  83.460000 229.250000  84.745000 ;
      RECT 227.005000 198.815000 227.175000 205.605000 ;
      RECT 227.005000 206.465000 227.175000 213.255000 ;
      RECT 227.065000   1.810000 227.235000   4.080000 ;
      RECT 227.080000  41.085000 227.750000  41.255000 ;
      RECT 227.080000  56.915000 227.750000  57.085000 ;
      RECT 227.105000  43.110000 227.635000  48.390000 ;
      RECT 227.105000  54.890000 227.635000  55.060000 ;
      RECT 227.115000 173.235000 300.630000 176.145000 ;
      RECT 227.115000 176.145000 227.965000 194.305000 ;
      RECT 227.145000  30.145000 227.315000  33.255000 ;
      RECT 227.145000  33.425000 227.315000  34.915000 ;
      RECT 227.205000  79.250000 229.915000  79.595000 ;
      RECT 227.210000  79.140000 229.900000  79.250000 ;
      RECT 227.215000  61.675000 227.385000  63.695000 ;
      RECT 227.215000  63.695000 227.745000  63.865000 ;
      RECT 227.215000  63.865000 227.385000  67.115000 ;
      RECT 227.220000  41.760000 227.750000  41.930000 ;
      RECT 227.220000  41.930000 227.530000  43.110000 ;
      RECT 227.220000  55.060000 227.530000  56.240000 ;
      RECT 227.220000  56.240000 227.750000  56.410000 ;
      RECT 227.240000 232.550000 227.605000 238.030000 ;
      RECT 227.245000  49.780000 227.415000  54.890000 ;
      RECT 227.250000 221.910000 227.505000 230.710000 ;
      RECT 227.260000  68.635000 227.430000  71.415000 ;
      RECT 227.260000  71.415000 228.150000  72.305000 ;
      RECT 227.260000  72.305000 227.430000  73.575000 ;
      RECT 227.265000  37.595000 227.635000  41.085000 ;
      RECT 227.265000  41.255000 227.750000  41.265000 ;
      RECT 227.265000  41.265000 228.230000  41.435000 ;
      RECT 227.265000  56.735000 228.230000  56.905000 ;
      RECT 227.265000  56.905000 227.750000  56.915000 ;
      RECT 227.265000  57.085000 227.635000  60.575000 ;
      RECT 227.330000  78.340000 227.860000  78.510000 ;
      RECT 227.335000 238.030000 227.505000 238.050000 ;
      RECT 227.345000 198.595000 227.615000 205.815000 ;
      RECT 227.445000  82.050000 227.615000  83.060000 ;
      RECT 227.450000  67.885000 227.980000  68.055000 ;
      RECT 227.465000  61.255000 227.995000  61.425000 ;
      RECT 227.485000  32.885000 228.015000  33.055000 ;
      RECT 227.485000  61.175000 227.995000  61.255000 ;
      RECT 227.485000  61.425000 227.995000  61.505000 ;
      RECT 227.555000  61.505000 227.925000  61.885000 ;
      RECT 227.555000  66.015000 227.925000  67.885000 ;
      RECT 227.690000  76.165000 227.860000  78.340000 ;
      RECT 227.690000  78.510000 227.860000  78.875000 ;
      RECT 227.695000  30.145000 227.865000  32.885000 ;
      RECT 227.695000  33.055000 227.865000  34.915000 ;
      RECT 227.700000  42.130000 228.230000  42.300000 ;
      RECT 227.700000  55.870000 228.230000  56.040000 ;
      RECT 227.750000  68.885000 227.920000  71.415000 ;
      RECT 227.750000  72.305000 227.920000  73.635000 ;
      RECT 227.785000 198.815000 227.955000 205.605000 ;
      RECT 227.785000 206.465000 227.955000 213.255000 ;
      RECT 227.805000  38.155000 228.090000  40.865000 ;
      RECT 227.805000  57.305000 228.090000  60.015000 ;
      RECT 227.825000  44.180000 229.385000  44.350000 ;
      RECT 227.825000  44.350000 227.995000  45.760000 ;
      RECT 227.825000  45.760000 230.355000  45.930000 ;
      RECT 227.825000  46.100000 227.995000  46.335000 ;
      RECT 227.825000  46.335000 228.355000  46.505000 ;
      RECT 227.825000  46.505000 227.995000  48.380000 ;
      RECT 227.825000  49.790000 227.995000  51.665000 ;
      RECT 227.825000  51.665000 228.355000  51.835000 ;
      RECT 227.825000  51.835000 227.995000  52.070000 ;
      RECT 227.825000  52.240000 230.355000  52.410000 ;
      RECT 227.825000  52.410000 227.995000  53.820000 ;
      RECT 227.825000  53.820000 229.385000  53.990000 ;
      RECT 227.920000  40.865000 228.090000  41.095000 ;
      RECT 227.920000  41.435000 228.230000  42.130000 ;
      RECT 227.920000  56.040000 228.230000  56.735000 ;
      RECT 227.920000  57.075000 228.090000  57.305000 ;
      RECT 227.925000  42.840000 228.095000  44.010000 ;
      RECT 227.925000  54.160000 228.095000  55.330000 ;
      RECT 227.995000   0.880000 228.165000   5.035000 ;
      RECT 228.040000 232.885000 247.765000 233.495000 ;
      RECT 228.055000  33.255000 230.085000  33.425000 ;
      RECT 228.055000 221.465000 247.765000 222.075000 ;
      RECT 228.055000 222.245000 247.765000 222.855000 ;
      RECT 228.055000 223.025000 247.765000 223.635000 ;
      RECT 228.055000 223.805000 247.765000 224.415000 ;
      RECT 228.055000 224.585000 247.765000 225.195000 ;
      RECT 228.055000 225.365000 247.765000 225.975000 ;
      RECT 228.055000 226.145000 247.765000 226.755000 ;
      RECT 228.055000 226.925000 247.765000 227.535000 ;
      RECT 228.055000 227.705000 247.765000 228.315000 ;
      RECT 228.055000 228.485000 247.765000 229.095000 ;
      RECT 228.055000 229.265000 247.765000 229.875000 ;
      RECT 228.055000 230.045000 247.765000 230.655000 ;
      RECT 228.055000 230.825000 247.765000 231.435000 ;
      RECT 228.055000 232.220000 247.765000 232.715000 ;
      RECT 228.055000 233.665000 247.765000 234.160000 ;
      RECT 228.055000 234.330000 247.765000 234.825000 ;
      RECT 228.055000 234.995000 247.765000 235.605000 ;
      RECT 228.055000 235.775000 247.765000 236.270000 ;
      RECT 228.055000 236.465000 247.765000 236.960000 ;
      RECT 228.055000 237.130000 247.765000 237.740000 ;
      RECT 228.055000 237.910000 247.765000 238.405000 ;
      RECT 228.060000  29.420000 228.730000  29.590000 ;
      RECT 228.075000  68.205000 233.845000  68.525000 ;
      RECT 228.095000  61.675000 228.265000  62.685000 ;
      RECT 228.095000  62.955000 228.265000  63.285000 ;
      RECT 228.095000  63.905000 228.265000  64.235000 ;
      RECT 228.095000  64.405000 228.265000  67.115000 ;
      RECT 228.115000  79.900000 228.285000  80.475000 ;
      RECT 228.125000 198.595000 228.395000 205.815000 ;
      RECT 228.140000  29.590000 228.670000  30.115000 ;
      RECT 228.165000  81.770000 228.695000  81.940000 ;
      RECT 228.210000  42.470000 229.560000  42.640000 ;
      RECT 228.210000  55.530000 229.560000  55.700000 ;
      RECT 228.285000   5.735000 228.985000  15.795000 ;
      RECT 228.285000  16.495000 228.985000  26.555000 ;
      RECT 228.310000  42.640000 229.560000  42.670000 ;
      RECT 228.310000  55.500000 229.560000  55.530000 ;
      RECT 228.340000  71.015000 228.870000  71.185000 ;
      RECT 228.350000  67.585000 228.860000  67.915000 ;
      RECT 228.355000  42.840000 228.525000  44.180000 ;
      RECT 228.355000  53.990000 228.525000  55.330000 ;
      RECT 228.355000  61.255000 228.885000  61.425000 ;
      RECT 228.385000  37.765000 228.555000  40.845000 ;
      RECT 228.385000  57.325000 228.555000  60.405000 ;
      RECT 228.435000  61.175000 228.805000  61.255000 ;
      RECT 228.435000  61.425000 228.805000  67.585000 ;
      RECT 228.470000  76.165000 228.640000  78.875000 ;
      RECT 228.525000  81.940000 228.695000  83.060000 ;
      RECT 228.530000  68.885000 228.700000  71.015000 ;
      RECT 228.530000  71.185000 228.700000  73.635000 ;
      RECT 228.565000 198.815000 228.735000 205.605000 ;
      RECT 228.565000 206.465000 228.735000 213.255000 ;
      RECT 228.585000 239.550000 237.205000 241.240000 ;
      RECT 228.605000  80.695000 231.655000  80.865000 ;
      RECT 228.785000  42.840000 228.955000  44.010000 ;
      RECT 228.785000  54.160000 228.955000  55.330000 ;
      RECT 228.975000  30.145000 232.945000  31.535000 ;
      RECT 228.975000  31.535000 230.085000  31.735000 ;
      RECT 228.975000  31.735000 229.145000  32.855000 ;
      RECT 228.975000  33.860000 229.145000  34.915000 ;
      RECT 228.975000  64.405000 229.145000  67.115000 ;
      RECT 229.005000  44.580000 229.175000  45.280000 ;
      RECT 229.005000  45.280000 229.680000  45.450000 ;
      RECT 229.005000  45.450000 229.175000  45.590000 ;
      RECT 229.005000  46.100000 229.175000  48.550000 ;
      RECT 229.005000  48.550000 231.895000  48.720000 ;
      RECT 229.005000  49.450000 231.895000  49.620000 ;
      RECT 229.005000  49.620000 229.175000  52.070000 ;
      RECT 229.005000  52.580000 229.175000  52.720000 ;
      RECT 229.005000  52.720000 229.680000  52.890000 ;
      RECT 229.005000  52.890000 229.175000  53.590000 ;
      RECT 229.080000  78.340000 229.610000  78.510000 ;
      RECT 229.145000 198.235000 229.315000 198.485000 ;
      RECT 229.145000 198.485000 230.260000 198.655000 ;
      RECT 229.145000 198.655000 229.315000 213.855000 ;
      RECT 229.155000  63.415000 229.685000  63.585000 ;
      RECT 229.200000  71.415000 229.760000  72.305000 ;
      RECT 229.205000 176.905000 298.850000 178.210000 ;
      RECT 229.205000 178.210000 344.705000 178.905000 ;
      RECT 229.205000 178.905000 230.055000 196.425000 ;
      RECT 229.215000  42.840000 229.385000  44.180000 ;
      RECT 229.215000  53.990000 229.385000  55.330000 ;
      RECT 229.240000  67.585000 229.750000  67.915000 ;
      RECT 229.245000  80.865000 229.775000  83.070000 ;
      RECT 229.250000  76.165000 229.420000  78.340000 ;
      RECT 229.250000  78.510000 229.420000  78.875000 ;
      RECT 229.310000  68.885000 229.760000  71.415000 ;
      RECT 229.310000  72.305000 229.760000  74.515000 ;
      RECT 229.315000  63.585000 229.685000  67.585000 ;
      RECT 229.505000  46.165000 229.835000  47.015000 ;
      RECT 229.505000  51.155000 229.835000  52.005000 ;
      RECT 229.555000  29.190000 270.960000  29.405000 ;
      RECT 229.555000  29.405000 232.945000  30.145000 ;
      RECT 229.585000  47.015000 229.755000  47.625000 ;
      RECT 229.585000  50.545000 229.755000  51.155000 ;
      RECT 229.590000  74.515000 229.760000  74.525000 ;
      RECT 229.645000  42.840000 229.815000  44.010000 ;
      RECT 229.645000  54.160000 229.815000  55.330000 ;
      RECT 229.730000  37.870000 229.900000  40.870000 ;
      RECT 229.730000  57.300000 229.900000  60.300000 ;
      RECT 229.795000  84.010000 230.325000  84.180000 ;
      RECT 229.855000  61.675000 230.025000  65.585000 ;
      RECT 229.855000  65.585000 230.385000  65.755000 ;
      RECT 229.855000  65.755000 230.025000  67.420000 ;
      RECT 229.910000   3.840000 231.930000   4.590000 ;
      RECT 229.910000  14.420000 231.930000  15.170000 ;
      RECT 229.915000  42.470000 231.265000  42.475000 ;
      RECT 229.915000  42.475000 232.575000  42.645000 ;
      RECT 229.915000  55.525000 232.575000  55.695000 ;
      RECT 229.915000  55.695000 231.265000  55.700000 ;
      RECT 229.930000  71.015000 230.460000  71.185000 ;
      RECT 229.930000 197.515000 230.260000 198.485000 ;
      RECT 229.930000 208.205000 230.655000 208.735000 ;
      RECT 229.950000  41.360000 230.480000  41.530000 ;
      RECT 229.950000  56.640000 230.480000  56.810000 ;
      RECT 230.030000  76.165000 230.200000  78.875000 ;
      RECT 230.075000  42.840000 230.245000  44.180000 ;
      RECT 230.075000  44.180000 231.895000  44.350000 ;
      RECT 230.075000  53.820000 231.895000  53.990000 ;
      RECT 230.075000  53.990000 230.245000  55.330000 ;
      RECT 230.075000 209.275000 231.675000 214.785000 ;
      RECT 230.090000  68.885000 230.260000  71.015000 ;
      RECT 230.090000  71.185000 230.260000  73.635000 ;
      RECT 230.115000  61.255000 230.645000  61.425000 ;
      RECT 230.125000  61.175000 230.635000  61.255000 ;
      RECT 230.125000  61.425000 230.635000  61.505000 ;
      RECT 230.140000 112.085000 230.670000 112.255000 ;
      RECT 230.150000 112.000000 230.660000 112.085000 ;
      RECT 230.150000 112.255000 230.660000 112.330000 ;
      RECT 230.155000  81.285000 230.325000  84.010000 ;
      RECT 230.155000  84.180000 230.325000  84.465000 ;
      RECT 230.155000  84.465000 230.765000  84.795000 ;
      RECT 230.170000  74.255000 236.610000  74.505000 ;
      RECT 230.170000  75.700000 230.840000  75.785000 ;
      RECT 230.170000  75.785000 230.900000  75.870000 ;
      RECT 230.185000  44.580000 230.355000  45.760000 ;
      RECT 230.185000  45.930000 230.355000  47.080000 ;
      RECT 230.185000  47.370000 231.055000  48.380000 ;
      RECT 230.185000  49.790000 231.055000  50.800000 ;
      RECT 230.185000  51.090000 230.355000  52.240000 ;
      RECT 230.185000  52.410000 230.355000  53.590000 ;
      RECT 230.195000  61.505000 230.565000  61.880000 ;
      RECT 230.195000  63.455000 230.525000  63.695000 ;
      RECT 230.195000  63.695000 230.725000  63.865000 ;
      RECT 230.195000  63.865000 230.525000  63.965000 ;
      RECT 230.255000  31.775000 230.425000  34.915000 ;
      RECT 230.310000  37.840000 234.550000  38.010000 ;
      RECT 230.310000  38.010000 230.480000  41.360000 ;
      RECT 230.310000  56.810000 230.480000  60.160000 ;
      RECT 230.310000  60.160000 234.550000  60.330000 ;
      RECT 230.370000  75.870000 230.900000  75.955000 ;
      RECT 230.490000 113.195000 231.160000 113.525000 ;
      RECT 230.505000  42.840000 230.675000  44.010000 ;
      RECT 230.505000  54.160000 230.675000  55.330000 ;
      RECT 230.525000  46.335000 231.055000  47.370000 ;
      RECT 230.525000  50.800000 231.055000  51.835000 ;
      RECT 230.535000  37.335000 232.565000  37.505000 ;
      RECT 230.535000  60.665000 232.565000  60.835000 ;
      RECT 230.615000 113.910000 233.615000 164.900000 ;
      RECT 230.735000  64.405000 230.905000  67.115000 ;
      RECT 230.810000  76.165000 230.980000  78.265000 ;
      RECT 230.810000  78.265000 231.420000  78.435000 ;
      RECT 230.810000  78.435000 230.980000  78.875000 ;
      RECT 230.825000 197.275000 231.675000 209.275000 ;
      RECT 230.835000  31.535000 232.945000  31.735000 ;
      RECT 230.870000  68.885000 231.040000  74.255000 ;
      RECT 230.885000 239.105000 239.335000 239.275000 ;
      RECT 230.935000  42.840000 231.105000  44.180000 ;
      RECT 230.935000  53.990000 231.105000  55.330000 ;
      RECT 230.935000  81.285000 231.105000  84.380000 ;
      RECT 230.935000  84.380000 234.460000  84.545000 ;
      RECT 230.935000  84.545000 234.475000  84.560000 ;
      RECT 230.935000  84.780000 231.525000  84.950000 ;
      RECT 230.935000  84.950000 231.105000  85.465000 ;
      RECT 231.005000  45.280000 231.535000  45.450000 ;
      RECT 231.005000  52.720000 231.535000  52.890000 ;
      RECT 231.005000  61.175000 231.515000  61.285000 ;
      RECT 231.005000  61.285000 231.535000  61.455000 ;
      RECT 231.005000  61.455000 231.515000  61.505000 ;
      RECT 231.015000 242.030000 237.065000 242.090000 ;
      RECT 231.015000 242.090000 237.185000 243.700000 ;
      RECT 231.015000 243.700000 237.065000 243.720000 ;
      RECT 231.020000  67.585000 231.530000  67.915000 ;
      RECT 231.075000  61.505000 231.445000  67.585000 ;
      RECT 231.150000  75.775000 232.160000  75.945000 ;
      RECT 231.155000 179.155000 293.520000 180.175000 ;
      RECT 231.155000 180.175000 234.110000 183.525000 ;
      RECT 231.155000 183.525000 249.755000 184.375000 ;
      RECT 231.155000 184.375000 234.110000 188.010000 ;
      RECT 231.155000 188.010000 249.755000 188.860000 ;
      RECT 231.155000 188.860000 234.110000 192.620000 ;
      RECT 231.155000 192.620000 235.245000 192.950000 ;
      RECT 231.155000 192.950000 234.110000 193.515000 ;
      RECT 231.155000 193.515000 283.670000 194.595000 ;
      RECT 231.155000 194.595000 342.805000 195.440000 ;
      RECT 231.190000  38.180000 231.450000  41.160000 ;
      RECT 231.190000  57.010000 231.450000  59.990000 ;
      RECT 231.365000  42.840000 231.535000  44.010000 ;
      RECT 231.365000  44.580000 231.535000  45.280000 ;
      RECT 231.365000  45.450000 231.535000  47.080000 ;
      RECT 231.365000  47.370000 231.895000  48.550000 ;
      RECT 231.365000  49.620000 231.895000  50.800000 ;
      RECT 231.365000  51.090000 231.535000  52.720000 ;
      RECT 231.365000  52.890000 231.535000  53.590000 ;
      RECT 231.365000  54.160000 231.535000  55.330000 ;
      RECT 231.460000  71.015000 231.990000  71.185000 ;
      RECT 231.485000  80.865000 231.655000  83.995000 ;
      RECT 231.535000  31.735000 232.945000  32.785000 ;
      RECT 231.535000  33.860000 231.705000  34.915000 ;
      RECT 231.590000  76.165000 231.760000  78.875000 ;
      RECT 231.615000  61.675000 231.785000  62.725000 ;
      RECT 231.615000  62.955000 231.785000  63.285000 ;
      RECT 231.615000  63.905000 231.785000  64.235000 ;
      RECT 231.615000  64.405000 231.785000  67.115000 ;
      RECT 231.650000  38.180000 231.910000  41.160000 ;
      RECT 231.650000  57.010000 231.910000  59.990000 ;
      RECT 231.650000  68.885000 231.820000  71.015000 ;
      RECT 231.650000  71.185000 231.820000  73.635000 ;
      RECT 231.705000  43.095000 232.235000  43.265000 ;
      RECT 231.705000  44.350000 231.895000  47.370000 ;
      RECT 231.705000  50.800000 231.895000  53.820000 ;
      RECT 231.705000  54.905000 232.235000  55.075000 ;
      RECT 231.765000  84.560000 234.475000  84.715000 ;
      RECT 231.825000  41.360000 232.355000  41.530000 ;
      RECT 231.825000  56.640000 232.355000  56.810000 ;
      RECT 231.855000  85.025000 234.225000  86.210000 ;
      RECT 232.005000  41.530000 232.175000  42.305000 ;
      RECT 232.005000  55.865000 232.175000  56.640000 ;
      RECT 232.065000  43.265000 232.235000  48.390000 ;
      RECT 232.065000  49.780000 232.235000  54.905000 ;
      RECT 232.090000  80.770000 232.620000  80.940000 ;
      RECT 232.135000  63.415000 232.665000  63.585000 ;
      RECT 232.265000  80.940000 232.435000  83.995000 ;
      RECT 232.345000  15.225000 237.195000  15.395000 ;
      RECT 232.345000  16.505000 237.095000  16.675000 ;
      RECT 232.370000  76.165000 232.540000  79.140000 ;
      RECT 232.370000  79.140000 232.945000  79.310000 ;
      RECT 232.405000  42.645000 232.575000  43.405000 ;
      RECT 232.405000  43.405000 233.055000  44.415000 ;
      RECT 232.405000  53.755000 233.055000  54.765000 ;
      RECT 232.405000  54.765000 232.575000  55.525000 ;
      RECT 232.430000  68.885000 232.600000  74.255000 ;
      RECT 232.435000  32.785000 232.945000  35.945000 ;
      RECT 232.495000  61.675000 232.665000  63.415000 ;
      RECT 232.495000  63.585000 232.665000  67.115000 ;
      RECT 232.525000  41.290000 233.195000  41.460000 ;
      RECT 232.525000  46.335000 233.055000  46.505000 ;
      RECT 232.525000  51.665000 233.055000  51.835000 ;
      RECT 232.525000  56.710000 233.195000  56.880000 ;
      RECT 232.545000  47.855000 232.715000  48.465000 ;
      RECT 232.545000  48.465000 238.075000  48.635000 ;
      RECT 232.545000  49.535000 235.395000  49.705000 ;
      RECT 232.545000  49.705000 232.715000  50.315000 ;
      RECT 232.585000  42.030000 233.115000  42.200000 ;
      RECT 232.585000  55.970000 233.115000  56.140000 ;
      RECT 232.620000  38.180000 232.790000  41.290000 ;
      RECT 232.620000  41.460000 233.115000  42.030000 ;
      RECT 232.620000  56.140000 233.115000  56.710000 ;
      RECT 232.620000  56.880000 232.790000  59.990000 ;
      RECT 232.675000 198.275000 307.965000 199.125000 ;
      RECT 232.675000 199.125000 236.585000 217.365000 ;
      RECT 232.675000 217.365000 307.965000 218.215000 ;
      RECT 232.775000  37.335000 233.445000  37.505000 ;
      RECT 232.775000  60.665000 233.445000  60.835000 ;
      RECT 232.885000  44.415000 233.055000  46.335000 ;
      RECT 232.885000  46.505000 233.055000  48.085000 ;
      RECT 232.885000  50.085000 233.055000  51.665000 ;
      RECT 232.885000  51.835000 233.055000  53.755000 ;
      RECT 232.920000  76.165000 233.090000  78.350000 ;
      RECT 232.920000  78.350000 233.450000  78.520000 ;
      RECT 232.920000  78.520000 233.090000  78.875000 ;
      RECT 233.015000  71.015000 233.545000  71.185000 ;
      RECT 233.045000  61.675000 233.215000  63.415000 ;
      RECT 233.045000  63.415000 233.575000  63.585000 ;
      RECT 233.045000  63.585000 233.215000  67.115000 ;
      RECT 233.045000  81.285000 233.215000  83.995000 ;
      RECT 233.050000 113.195000 233.720000 113.525000 ;
      RECT 233.210000  68.885000 233.380000  71.015000 ;
      RECT 233.210000  71.185000 233.380000  73.635000 ;
      RECT 233.225000  45.000000 233.755000  45.170000 ;
      RECT 233.225000  53.000000 233.755000  53.170000 ;
      RECT 233.245000  75.775000 234.255000  75.945000 ;
      RECT 233.285000  41.635000 233.535000  42.305000 ;
      RECT 233.285000  55.865000 233.535000  56.535000 ;
      RECT 233.320000  41.580000 233.535000  41.635000 ;
      RECT 233.320000  42.305000 233.490000  43.405000 ;
      RECT 233.320000  43.405000 233.515000  44.415000 ;
      RECT 233.320000  53.755000 233.515000  54.765000 ;
      RECT 233.320000  54.765000 233.490000  55.865000 ;
      RECT 233.320000  56.535000 233.535000  56.590000 ;
      RECT 233.345000  45.170000 233.515000  48.085000 ;
      RECT 233.345000  50.085000 233.515000  53.000000 ;
      RECT 233.365000  38.180000 233.670000  40.890000 ;
      RECT 233.365000  40.890000 233.535000  41.580000 ;
      RECT 233.365000  56.590000 233.535000  57.280000 ;
      RECT 233.365000  57.280000 233.670000  59.990000 ;
      RECT 233.465000  80.770000 233.995000  80.940000 ;
      RECT 233.575000  19.055000 233.745000  26.470000 ;
      RECT 233.575000  26.470000 239.325000  26.640000 ;
      RECT 233.685000  42.400000 234.215000  42.570000 ;
      RECT 233.685000  42.570000 234.095000  44.585000 ;
      RECT 233.685000  44.585000 234.225000  44.740000 ;
      RECT 233.685000  45.375000 234.225000  45.665000 ;
      RECT 233.685000  45.665000 233.975000  48.085000 ;
      RECT 233.685000  50.085000 233.975000  52.505000 ;
      RECT 233.685000  52.505000 234.225000  52.795000 ;
      RECT 233.685000  53.430000 234.225000  53.585000 ;
      RECT 233.685000  53.585000 234.095000  55.600000 ;
      RECT 233.685000  55.600000 234.215000  55.770000 ;
      RECT 233.700000  75.945000 233.870000  79.620000 ;
      RECT 233.700000  79.620000 235.790000  79.790000 ;
      RECT 233.705000  42.030000 234.735000  42.200000 ;
      RECT 233.705000  55.970000 234.735000  56.140000 ;
      RECT 233.725000  37.335000 234.395000  37.505000 ;
      RECT 233.725000  60.665000 236.835000  60.835000 ;
      RECT 233.755000  71.415000 234.650000  72.305000 ;
      RECT 233.805000  41.290000 234.550000  41.460000 ;
      RECT 233.805000  56.710000 234.550000  56.880000 ;
      RECT 233.825000  80.940000 233.995000  83.995000 ;
      RECT 233.875000  41.460000 234.405000  41.530000 ;
      RECT 233.875000  56.640000 234.405000  56.710000 ;
      RECT 233.925000  44.740000 234.225000  45.375000 ;
      RECT 233.925000  52.795000 234.225000  53.430000 ;
      RECT 233.925000  61.675000 234.095000  62.725000 ;
      RECT 233.925000  62.955000 234.095000  63.285000 ;
      RECT 233.925000  63.905000 234.095000  64.235000 ;
      RECT 233.925000  64.405000 234.095000  67.115000 ;
      RECT 233.980000  31.565000 235.205000  31.735000 ;
      RECT 233.990000  68.635000 234.650000  71.415000 ;
      RECT 233.990000  72.305000 234.650000  74.255000 ;
      RECT 234.125000  22.010000 234.385000  22.655000 ;
      RECT 234.170000  19.080000 234.340000  22.010000 ;
      RECT 234.170000  22.655000 234.340000  25.870000 ;
      RECT 234.170000  61.285000 234.705000  61.455000 ;
      RECT 234.175000  48.105000 234.930000  48.275000 ;
      RECT 234.175000  49.895000 234.930000  50.065000 ;
      RECT 234.180000  67.585000 234.690000  67.915000 ;
      RECT 234.195000  61.175000 234.705000  61.285000 ;
      RECT 234.195000  61.455000 234.705000  61.505000 ;
      RECT 234.265000  43.405000 234.435000  44.415000 ;
      RECT 234.265000  53.755000 234.435000  54.765000 ;
      RECT 234.265000  61.505000 234.635000  67.585000 ;
      RECT 234.305000  78.350000 234.835000  78.520000 ;
      RECT 234.340000  30.285000 235.205000  31.565000 ;
      RECT 234.340000  31.735000 235.205000  31.795000 ;
      RECT 234.340000  32.515000 235.205000  35.725000 ;
      RECT 234.340000  35.725000 234.510000  36.025000 ;
      RECT 234.380000  38.010000 234.550000  41.290000 ;
      RECT 234.380000  56.880000 234.550000  60.160000 ;
      RECT 234.400000  46.335000 234.930000  46.505000 ;
      RECT 234.400000  51.665000 234.930000  51.835000 ;
      RECT 234.420000  44.630000 234.590000  45.300000 ;
      RECT 234.420000  52.870000 234.590000  53.540000 ;
      RECT 234.460000  42.510000 234.995000  43.085000 ;
      RECT 234.460000  55.085000 234.995000  55.660000 ;
      RECT 234.480000  76.165000 234.650000  78.350000 ;
      RECT 234.480000  78.520000 234.650000  78.875000 ;
      RECT 234.490000  18.650000 238.435000  18.820000 ;
      RECT 234.565000  41.635000 234.735000  42.030000 ;
      RECT 234.565000  42.200000 234.735000  42.305000 ;
      RECT 234.565000  55.865000 234.735000  55.970000 ;
      RECT 234.565000  56.140000 234.735000  56.535000 ;
      RECT 234.725000  43.405000 234.930000  44.415000 ;
      RECT 234.725000  53.755000 234.930000  54.765000 ;
      RECT 234.735000  14.655000 239.945000  14.825000 ;
      RECT 234.760000  44.415000 234.930000  46.335000 ;
      RECT 234.760000  46.505000 234.930000  48.105000 ;
      RECT 234.760000  50.065000 234.930000  51.665000 ;
      RECT 234.760000  51.835000 234.930000  53.755000 ;
      RECT 234.780000  80.895000 235.450000  81.065000 ;
      RECT 234.805000  64.405000 234.975000  67.115000 ;
      RECT 234.805000  75.775000 236.210000  75.945000 ;
      RECT 234.840000  80.800000 235.370000  80.895000 ;
      RECT 234.840000  81.285000 235.010000  86.270000 ;
      RECT 234.865000 180.765000 249.815000 180.935000 ;
      RECT 234.865000 181.545000 249.815000 181.715000 ;
      RECT 234.865000 182.325000 249.815000 182.495000 ;
      RECT 234.865000 185.395000 249.815000 185.565000 ;
      RECT 234.865000 186.175000 249.815000 186.345000 ;
      RECT 234.865000 186.955000 249.815000 187.125000 ;
      RECT 234.865000 189.805000 249.815000 189.975000 ;
      RECT 234.865000 190.585000 249.815000 190.755000 ;
      RECT 234.865000 191.365000 249.815000 191.535000 ;
      RECT 234.965000  71.015000 235.495000  71.185000 ;
      RECT 234.970000  68.885000 235.140000  71.015000 ;
      RECT 234.970000  71.185000 235.140000  73.635000 ;
      RECT 234.985000  63.695000 235.515000  63.865000 ;
      RECT 235.035000  31.795000 235.205000  31.895000 ;
      RECT 235.065000  61.255000 235.595000  61.425000 ;
      RECT 235.075000  61.175000 235.585000  61.255000 ;
      RECT 235.075000  61.425000 235.585000  61.505000 ;
      RECT 235.105000   4.515000 243.425000   4.685000 ;
      RECT 235.105000   4.685000 235.275000  10.055000 ;
      RECT 235.125000 113.910000 238.125000 164.900000 ;
      RECT 235.145000  61.505000 235.515000  61.880000 ;
      RECT 235.185000  63.455000 235.515000  63.695000 ;
      RECT 235.185000  63.865000 235.515000  63.965000 ;
      RECT 235.205000  23.495000 235.465000  25.000000 ;
      RECT 235.225000  37.870000 235.395000  44.425000 ;
      RECT 235.225000  45.065000 235.395000  48.465000 ;
      RECT 235.225000  49.705000 235.395000  52.000000 ;
      RECT 235.225000  52.610000 235.395000  58.725000 ;
      RECT 235.225000  58.725000 235.410000  59.255000 ;
      RECT 235.225000  59.255000 235.395000  60.320000 ;
      RECT 235.250000  19.080000 235.420000  23.495000 ;
      RECT 235.250000  25.000000 235.420000  25.870000 ;
      RECT 235.260000  76.165000 235.430000  79.140000 ;
      RECT 235.260000  79.140000 236.460000  79.370000 ;
      RECT 235.295000  68.205000 241.065000  68.555000 ;
      RECT 235.305000  29.785000 235.815000  30.115000 ;
      RECT 235.305000  36.195000 235.815000  36.525000 ;
      RECT 235.325000  65.585000 235.855000  65.755000 ;
      RECT 235.375000  30.115000 235.745000  36.195000 ;
      RECT 235.560000  72.535000 236.090000  72.705000 ;
      RECT 235.565000  10.860000 236.095000  11.030000 ;
      RECT 235.620000  79.790000 235.790000  86.035000 ;
      RECT 235.625000  42.510000 236.160000  43.085000 ;
      RECT 235.680000  78.350000 236.210000  78.520000 ;
      RECT 235.685000   5.035000 235.855000   8.850000 ;
      RECT 235.685000   8.850000 236.215000   9.020000 ;
      RECT 235.685000   9.020000 235.855000   9.785000 ;
      RECT 235.685000  10.855000 235.855000  10.860000 ;
      RECT 235.685000  11.030000 235.855000  14.185000 ;
      RECT 235.685000  14.185000 239.355000  14.355000 ;
      RECT 235.685000  61.675000 235.855000  65.585000 ;
      RECT 235.685000  65.755000 235.855000  67.420000 ;
      RECT 235.690000  43.405000 235.895000  44.415000 ;
      RECT 235.690000  44.415000 235.860000  46.335000 ;
      RECT 235.690000  46.335000 236.220000  46.505000 ;
      RECT 235.690000  46.505000 235.860000  48.105000 ;
      RECT 235.690000  48.105000 236.445000  48.275000 ;
      RECT 235.750000  68.555000 235.920000  72.535000 ;
      RECT 235.750000  72.705000 235.920000  73.635000 ;
      RECT 235.885000  41.635000 236.055000  42.030000 ;
      RECT 235.885000  42.030000 236.915000  42.200000 ;
      RECT 235.885000  42.200000 236.055000  42.305000 ;
      RECT 235.915000  30.285000 236.085000  36.025000 ;
      RECT 235.960000  67.585000 236.470000  67.915000 ;
      RECT 235.960000  80.895000 236.630000  81.065000 ;
      RECT 236.025000  63.415000 236.555000  63.585000 ;
      RECT 236.025000  63.585000 236.395000  67.585000 ;
      RECT 236.030000  44.630000 236.200000  45.300000 ;
      RECT 236.040000  75.945000 236.210000  78.350000 ;
      RECT 236.040000  78.520000 236.210000  78.875000 ;
      RECT 236.040000  80.800000 236.570000  80.895000 ;
      RECT 236.070000  37.840000 240.310000  38.010000 ;
      RECT 236.070000  38.010000 236.240000  41.290000 ;
      RECT 236.070000  41.290000 236.815000  41.460000 ;
      RECT 236.120000  50.330000 245.210000  59.670000 ;
      RECT 236.185000  29.785000 237.575000  30.085000 ;
      RECT 236.185000  30.085000 236.695000  30.115000 ;
      RECT 236.185000  36.195000 236.695000  36.225000 ;
      RECT 236.185000  36.225000 237.580000  36.525000 ;
      RECT 236.185000  43.405000 236.355000  44.415000 ;
      RECT 236.215000  41.460000 236.745000  41.530000 ;
      RECT 236.225000  37.335000 236.895000  37.505000 ;
      RECT 236.255000  30.115000 236.625000  36.195000 ;
      RECT 236.260000  79.370000 236.460000  80.145000 ;
      RECT 236.260000  80.145000 236.565000  80.475000 ;
      RECT 236.265000  10.795000 236.435000  14.185000 ;
      RECT 236.285000  19.565000 236.545000  20.600000 ;
      RECT 236.330000  19.080000 236.500000  19.565000 ;
      RECT 236.330000  20.600000 236.500000  25.870000 ;
      RECT 236.335000  71.015000 236.865000  71.185000 ;
      RECT 236.365000 180.935000 245.665000 181.375000 ;
      RECT 236.365000 181.885000 245.665000 182.325000 ;
      RECT 236.365000 185.565000 245.665000 186.005000 ;
      RECT 236.365000 186.515000 245.665000 186.955000 ;
      RECT 236.365000 189.975000 245.665000 190.415000 ;
      RECT 236.365000 190.925000 245.665000 191.365000 ;
      RECT 236.395000  44.585000 236.935000  44.740000 ;
      RECT 236.395000  44.740000 236.695000  45.375000 ;
      RECT 236.395000  45.375000 236.935000  45.665000 ;
      RECT 236.400000  81.285000 236.570000  86.270000 ;
      RECT 236.405000  42.400000 236.935000  42.570000 ;
      RECT 236.465000   5.035000 236.635000   9.220000 ;
      RECT 236.465000   9.220000 237.000000   9.390000 ;
      RECT 236.465000   9.390000 236.635000  10.015000 ;
      RECT 236.465000  10.015000 237.215000  10.185000 ;
      RECT 236.525000  42.570000 236.935000  44.585000 ;
      RECT 236.530000  68.885000 236.700000  71.015000 ;
      RECT 236.530000  71.185000 236.700000  73.635000 ;
      RECT 236.555000  95.265000 299.555000 102.115000 ;
      RECT 236.565000  64.405000 236.735000  67.115000 ;
      RECT 236.630000  75.525000 236.800000  79.145000 ;
      RECT 236.645000  45.665000 236.935000  48.085000 ;
      RECT 236.735000  18.820000 237.160000  26.185000 ;
      RECT 236.795000  30.285000 236.965000  31.895000 ;
      RECT 236.795000  32.515000 236.965000  35.725000 ;
      RECT 236.825000  61.255000 237.355000  61.425000 ;
      RECT 236.850000  67.585000 237.535000  67.685000 ;
      RECT 236.850000  67.685000 237.360000  67.915000 ;
      RECT 236.865000  45.000000 237.395000  45.170000 ;
      RECT 236.905000  61.175000 237.275000  61.255000 ;
      RECT 236.905000  61.425000 237.275000  67.515000 ;
      RECT 236.905000  67.515000 237.535000  67.585000 ;
      RECT 236.940000 104.530000 248.875000 104.700000 ;
      RECT 236.940000 104.700000 237.110000 107.450000 ;
      RECT 236.940000 107.450000 248.875000 107.620000 ;
      RECT 236.950000  38.180000 237.255000  40.890000 ;
      RECT 237.045000  10.185000 237.215000  11.360000 ;
      RECT 237.045000  11.360000 237.575000  11.530000 ;
      RECT 237.045000  11.530000 237.215000  13.505000 ;
      RECT 237.065000  30.085000 237.575000  30.115000 ;
      RECT 237.070000  36.195000 237.580000  36.225000 ;
      RECT 237.085000  40.890000 237.255000  41.580000 ;
      RECT 237.085000  41.580000 237.300000  41.635000 ;
      RECT 237.085000  41.635000 237.335000  42.305000 ;
      RECT 237.095000 200.495000 237.625000 215.995000 ;
      RECT 237.105000  43.405000 237.300000  44.415000 ;
      RECT 237.105000  45.170000 237.275000  48.085000 ;
      RECT 237.120000  72.535000 237.650000  72.705000 ;
      RECT 237.130000  42.305000 237.300000  43.405000 ;
      RECT 237.135000  30.115000 237.505000  36.195000 ;
      RECT 237.175000  37.335000 237.845000  37.505000 ;
      RECT 237.245000   5.035000 237.415000   8.850000 ;
      RECT 237.245000   8.850000 237.775000   9.020000 ;
      RECT 237.245000   9.020000 237.415000   9.785000 ;
      RECT 237.260000  60.665000 237.790000  60.835000 ;
      RECT 237.310000  68.555000 237.480000  72.535000 ;
      RECT 237.310000  72.705000 237.480000  73.635000 ;
      RECT 237.350000 105.375000 237.520000 106.360000 ;
      RECT 237.350000 106.360000 237.880000 106.530000 ;
      RECT 237.350000 106.530000 237.520000 106.725000 ;
      RECT 237.365000  23.495000 237.625000  25.000000 ;
      RECT 237.365000 243.890000 240.460000 244.175000 ;
      RECT 237.365000 244.175000 237.735000 244.345000 ;
      RECT 237.365000 244.345000 238.115000 246.365000 ;
      RECT 237.365000 246.365000 237.735000 246.535000 ;
      RECT 237.365000 246.535000 240.460000 246.935000 ;
      RECT 237.380000  74.400000 237.550000  81.020000 ;
      RECT 237.410000  19.080000 237.580000  23.495000 ;
      RECT 237.410000  25.000000 237.580000  25.870000 ;
      RECT 237.425000  41.290000 238.095000  41.460000 ;
      RECT 237.445000  61.675000 237.615000  62.685000 ;
      RECT 237.445000  62.955000 237.615000  63.285000 ;
      RECT 237.445000  63.905000 237.615000  64.235000 ;
      RECT 237.445000  64.405000 237.615000  67.115000 ;
      RECT 237.450000 105.035000 248.355000 105.205000 ;
      RECT 237.450000 106.940000 248.355000 107.110000 ;
      RECT 237.480000  81.950000 237.650000  87.070000 ;
      RECT 237.505000  10.295000 239.525000  10.465000 ;
      RECT 237.505000  41.460000 238.000000  42.030000 ;
      RECT 237.505000  42.030000 238.035000  42.200000 ;
      RECT 237.565000  43.405000 238.215000  44.415000 ;
      RECT 237.565000  44.415000 237.735000  46.335000 ;
      RECT 237.565000  46.335000 238.095000  46.505000 ;
      RECT 237.565000  46.505000 237.735000  48.085000 ;
      RECT 237.575000  15.350000 240.135000  18.455000 ;
      RECT 237.585000   9.590000 237.855000  10.295000 ;
      RECT 237.585000  36.975000 237.755000  37.335000 ;
      RECT 237.665000   9.220000 238.195000   9.390000 ;
      RECT 237.675000  30.285000 237.845000  36.025000 ;
      RECT 237.715000  61.175000 238.225000  61.255000 ;
      RECT 237.715000  61.255000 238.245000  61.425000 ;
      RECT 237.715000  61.425000 238.225000  61.505000 ;
      RECT 237.720000  77.400000 238.140000  78.240000 ;
      RECT 237.720000  78.240000 238.560000  78.410000 ;
      RECT 237.720000  78.410000 238.140000  78.750000 ;
      RECT 237.720000  78.750000 237.890000  79.730000 ;
      RECT 237.720000  79.730000 238.140000  81.080000 ;
      RECT 237.725000 239.550000 243.390000 241.240000 ;
      RECT 237.750000  22.940000 238.280000  23.110000 ;
      RECT 237.785000  61.505000 238.155000  61.885000 ;
      RECT 237.815000  18.820000 238.240000  22.940000 ;
      RECT 237.815000  23.110000 238.240000  26.185000 ;
      RECT 237.825000  10.795000 237.995000  14.185000 ;
      RECT 237.825000 242.030000 243.050000 243.720000 ;
      RECT 237.830000  38.180000 238.000000  41.290000 ;
      RECT 237.895000  71.015000 238.425000  71.185000 ;
      RECT 237.905000  47.855000 238.075000  48.465000 ;
      RECT 237.945000  29.785000 239.335000  30.085000 ;
      RECT 237.945000  30.085000 238.455000  30.115000 ;
      RECT 237.945000  36.195000 238.455000  36.225000 ;
      RECT 237.945000  36.225000 239.335000  36.525000 ;
      RECT 237.965000  63.695000 238.495000  63.865000 ;
      RECT 237.970000  74.420000 238.140000  76.020000 ;
      RECT 237.970000  81.890000 238.140000  83.290000 ;
      RECT 237.970000  83.290000 238.500000  83.460000 ;
      RECT 237.970000  83.460000 238.140000  86.640000 ;
      RECT 238.000000 105.205000 242.750000 105.280000 ;
      RECT 238.000000 105.990000 242.750000 106.160000 ;
      RECT 238.000000 106.870000 242.750000 106.940000 ;
      RECT 238.015000  30.115000 238.385000  36.195000 ;
      RECT 238.025000   5.035000 238.195000   9.220000 ;
      RECT 238.025000   9.390000 238.195000   9.785000 ;
      RECT 238.045000  42.475000 240.705000  42.645000 ;
      RECT 238.045000  42.645000 238.215000  43.405000 ;
      RECT 238.055000  37.335000 240.085000  37.505000 ;
      RECT 238.055000 199.685000 238.715000 200.085000 ;
      RECT 238.055000 200.085000 238.725000 200.255000 ;
      RECT 238.055000 216.235000 238.725000 216.405000 ;
      RECT 238.090000  68.885000 238.260000  71.015000 ;
      RECT 238.090000  71.185000 238.260000  73.635000 ;
      RECT 238.105000  79.075000 238.615000  79.120000 ;
      RECT 238.105000  79.120000 238.670000  79.290000 ;
      RECT 238.105000  79.290000 238.615000  79.405000 ;
      RECT 238.115000  60.665000 240.085000  60.835000 ;
      RECT 238.215000  76.370000 241.945000  76.540000 ;
      RECT 238.245000  11.360000 238.775000  11.530000 ;
      RECT 238.260000  87.150000 240.290000  87.320000 ;
      RECT 238.265000  41.360000 238.795000  41.530000 ;
      RECT 238.285000 244.175000 240.460000 246.535000 ;
      RECT 238.325000  61.675000 238.495000  63.695000 ;
      RECT 238.325000  63.865000 238.495000  67.115000 ;
      RECT 238.385000  43.095000 238.915000  43.265000 ;
      RECT 238.385000  43.265000 238.555000  48.390000 ;
      RECT 238.445000   8.850000 238.975000   9.020000 ;
      RECT 238.445000  19.565000 238.705000  20.600000 ;
      RECT 238.445000  41.530000 238.615000  42.305000 ;
      RECT 238.490000  19.080000 238.660000  19.565000 ;
      RECT 238.490000  20.600000 238.660000  25.870000 ;
      RECT 238.555000  30.285000 238.725000  31.895000 ;
      RECT 238.555000  32.515000 238.725000  35.725000 ;
      RECT 238.605000  10.795000 238.775000  11.360000 ;
      RECT 238.605000  11.530000 238.775000  13.505000 ;
      RECT 238.660000  75.100000 242.050000  75.270000 ;
      RECT 238.680000  72.535000 239.210000  72.705000 ;
      RECT 238.710000  38.180000 238.970000  41.160000 ;
      RECT 238.725000  44.180000 240.545000  44.350000 ;
      RECT 238.725000  44.350000 238.915000  47.370000 ;
      RECT 238.725000  47.370000 239.255000  48.550000 ;
      RECT 238.725000  48.550000 241.615000  48.720000 ;
      RECT 238.805000   5.035000 238.975000   8.850000 ;
      RECT 238.805000   9.020000 238.975000   9.785000 ;
      RECT 238.825000  30.085000 239.335000  30.115000 ;
      RECT 238.825000  36.195000 239.335000  36.225000 ;
      RECT 238.850000  81.890000 239.020000  86.640000 ;
      RECT 238.870000  68.555000 239.040000  72.535000 ;
      RECT 238.870000  72.705000 239.040000  73.635000 ;
      RECT 238.875000  61.675000 239.045000  62.725000 ;
      RECT 238.875000  62.955000 239.045000  63.285000 ;
      RECT 238.875000  63.905000 239.045000  64.235000 ;
      RECT 238.875000  64.405000 239.045000  67.420000 ;
      RECT 238.895000  30.115000 239.265000  36.195000 ;
      RECT 238.905000  77.010000 241.195000  77.180000 ;
      RECT 238.905000  81.300000 241.195000  81.470000 ;
      RECT 238.965000  77.180000 239.790000  79.150000 ;
      RECT 238.965000  79.150000 241.195000  79.320000 ;
      RECT 238.965000  79.320000 239.790000  81.250000 ;
      RECT 238.965000  81.250000 241.195000  81.300000 ;
      RECT 239.005000  10.860000 239.535000  11.030000 ;
      RECT 239.085000  42.840000 239.255000  44.010000 ;
      RECT 239.085000  44.580000 239.255000  45.280000 ;
      RECT 239.085000  45.280000 239.615000  45.450000 ;
      RECT 239.085000  45.450000 239.255000  47.080000 ;
      RECT 239.155000  24.800000 244.845000  24.970000 ;
      RECT 239.155000  24.970000 239.325000  26.470000 ;
      RECT 239.155000 200.495000 239.685000 215.995000 ;
      RECT 239.170000  38.180000 239.430000  41.160000 ;
      RECT 239.185000  10.855000 239.355000  10.860000 ;
      RECT 239.185000  11.030000 239.355000  14.185000 ;
      RECT 239.215000  61.175000 239.725000  61.505000 ;
      RECT 239.215000  67.115000 239.745000  67.285000 ;
      RECT 239.215000  67.585000 239.725000  67.915000 ;
      RECT 239.285000  61.505000 239.655000  67.115000 ;
      RECT 239.285000  67.285000 239.655000  67.585000 ;
      RECT 239.355000   5.035000 239.525000  10.295000 ;
      RECT 239.355000  42.470000 240.705000  42.475000 ;
      RECT 239.435000  30.285000 239.605000  36.025000 ;
      RECT 239.455000  71.015000 239.985000  71.185000 ;
      RECT 239.500000  22.015000 239.760000  22.655000 ;
      RECT 239.510000 113.195000 240.180000 113.525000 ;
      RECT 239.515000  42.840000 239.685000  44.180000 ;
      RECT 239.545000  19.530000 239.715000  22.015000 ;
      RECT 239.545000  22.655000 239.715000  24.280000 ;
      RECT 239.560000  83.290000 240.090000  83.460000 ;
      RECT 239.565000  46.335000 240.095000  47.370000 ;
      RECT 239.565000  47.370000 240.435000  48.380000 ;
      RECT 239.605000  25.475000 239.775000  27.495000 ;
      RECT 239.635000 113.910000 242.635000 164.900000 ;
      RECT 239.650000  68.885000 239.820000  71.015000 ;
      RECT 239.650000  71.185000 239.820000  73.635000 ;
      RECT 239.695000   9.960000 240.225000  10.130000 ;
      RECT 239.705000  10.130000 240.225000  10.965000 ;
      RECT 239.705000  29.785000 241.095000  30.085000 ;
      RECT 239.705000  30.085000 240.215000  30.115000 ;
      RECT 239.705000  36.195000 240.215000  36.225000 ;
      RECT 239.705000  36.225000 241.095000  36.525000 ;
      RECT 239.730000  81.890000 239.900000  83.290000 ;
      RECT 239.730000  83.460000 239.900000  86.640000 ;
      RECT 239.770000  18.850000 244.790000  19.020000 ;
      RECT 239.775000  30.115000 240.145000  36.195000 ;
      RECT 239.825000  61.675000 239.995000  66.135000 ;
      RECT 239.945000  42.840000 240.115000  44.010000 ;
      RECT 239.960000  77.400000 240.130000  78.750000 ;
      RECT 239.960000  79.540000 240.130000  81.080000 ;
      RECT 240.075000  61.285000 240.605000  61.455000 ;
      RECT 240.095000  61.175000 240.605000  61.285000 ;
      RECT 240.095000  61.455000 240.605000  61.505000 ;
      RECT 240.095000  67.585000 240.605000  67.915000 ;
      RECT 240.115000 200.085000 240.785000 200.255000 ;
      RECT 240.115000 216.235000 240.785000 216.405000 ;
      RECT 240.135000   4.685000 240.305000   9.785000 ;
      RECT 240.140000  38.010000 240.310000  41.360000 ;
      RECT 240.140000  41.360000 240.670000  41.530000 ;
      RECT 240.165000  61.505000 240.535000  67.585000 ;
      RECT 240.240000  72.535000 240.770000  72.705000 ;
      RECT 240.265000  44.580000 240.435000  45.760000 ;
      RECT 240.265000  45.760000 242.795000  45.930000 ;
      RECT 240.265000  45.930000 240.435000  47.080000 ;
      RECT 240.280000  20.875000 240.540000  21.515000 ;
      RECT 240.285000  25.390000 245.035000  25.560000 ;
      RECT 240.285000  26.470000 245.035000  26.640000 ;
      RECT 240.285000  27.550000 245.035000  27.720000 ;
      RECT 240.300000  77.180000 241.195000  79.150000 ;
      RECT 240.300000  79.320000 241.195000  81.250000 ;
      RECT 240.315000  30.285000 240.485000  31.895000 ;
      RECT 240.315000  32.515000 240.485000  35.725000 ;
      RECT 240.325000  19.530000 240.495000  20.875000 ;
      RECT 240.325000  21.515000 240.495000  24.280000 ;
      RECT 240.360000  17.235000 241.250000  17.615000 ;
      RECT 240.375000  42.840000 240.545000  44.180000 ;
      RECT 240.415000  10.295000 243.125000  10.465000 ;
      RECT 240.430000  68.555000 240.600000  72.535000 ;
      RECT 240.430000  72.705000 240.600000  73.635000 ;
      RECT 240.460000  15.140000 241.130000  15.310000 ;
      RECT 240.585000  30.085000 241.095000  30.115000 ;
      RECT 240.585000  36.195000 241.095000  36.225000 ;
      RECT 240.610000  81.890000 240.780000  86.640000 ;
      RECT 240.655000  30.115000 241.025000  36.195000 ;
      RECT 240.720000  37.870000 240.890000  40.870000 ;
      RECT 240.775000  61.675000 240.945000  62.725000 ;
      RECT 240.775000  62.955000 240.945000  63.285000 ;
      RECT 240.775000  63.905000 240.945000  64.235000 ;
      RECT 240.775000  64.405000 240.945000  67.115000 ;
      RECT 240.785000  46.165000 241.115000  47.015000 ;
      RECT 240.805000  42.840000 240.975000  44.010000 ;
      RECT 240.845000  71.015000 241.405000  71.185000 ;
      RECT 240.850000 112.085000 241.380000 112.255000 ;
      RECT 240.855000  87.150000 241.525000  87.320000 ;
      RECT 240.860000 112.000000 241.370000 112.085000 ;
      RECT 240.860000 112.255000 241.370000 112.330000 ;
      RECT 240.865000  47.015000 241.035000  47.625000 ;
      RECT 240.915000   5.035000 241.085000   8.850000 ;
      RECT 240.915000   8.850000 241.445000   9.020000 ;
      RECT 240.915000   9.020000 241.085000   9.785000 ;
      RECT 240.940000  45.280000 241.615000  45.450000 ;
      RECT 241.045000  61.175000 241.555000  61.505000 ;
      RECT 241.045000  67.585000 241.555000  67.915000 ;
      RECT 241.060000  22.015000 241.320000  22.655000 ;
      RECT 241.060000  42.470000 242.410000  42.640000 ;
      RECT 241.060000  42.640000 242.310000  42.670000 ;
      RECT 241.105000  19.530000 241.275000  22.015000 ;
      RECT 241.105000  22.655000 241.275000  24.280000 ;
      RECT 241.110000  83.290000 241.660000  83.460000 ;
      RECT 241.115000  61.505000 241.485000  67.585000 ;
      RECT 241.195000  30.285000 241.365000  36.025000 ;
      RECT 241.210000  68.885000 241.405000  71.015000 ;
      RECT 241.210000  71.185000 241.405000  73.345000 ;
      RECT 241.210000  73.345000 241.380000  73.635000 ;
      RECT 241.215000 200.495000 241.745000 215.995000 ;
      RECT 241.235000  42.840000 241.405000  44.180000 ;
      RECT 241.235000  44.180000 242.795000  44.350000 ;
      RECT 241.235000  68.205000 248.290000  68.385000 ;
      RECT 241.235000  68.385000 241.405000  68.885000 ;
      RECT 241.445000  44.580000 241.615000  45.280000 ;
      RECT 241.445000  45.450000 241.615000  45.590000 ;
      RECT 241.445000  46.100000 241.615000  48.550000 ;
      RECT 241.465000  29.785000 241.975000  30.115000 ;
      RECT 241.465000  36.195000 241.975000  36.525000 ;
      RECT 241.475000  75.270000 242.005000  75.330000 ;
      RECT 241.475000  79.110000 242.005000  79.280000 ;
      RECT 241.485000  79.075000 241.995000  79.110000 ;
      RECT 241.485000  79.280000 241.995000  79.405000 ;
      RECT 241.490000  81.890000 241.660000  83.290000 ;
      RECT 241.490000  83.460000 241.660000  86.640000 ;
      RECT 241.530000  78.240000 242.435000  78.410000 ;
      RECT 241.535000  30.115000 241.905000  36.195000 ;
      RECT 241.655000  61.675000 241.825000  67.415000 ;
      RECT 241.665000  42.840000 241.835000  44.010000 ;
      RECT 241.695000   4.685000 241.865000   9.785000 ;
      RECT 241.700000  68.635000 242.360000  71.040000 ;
      RECT 241.700000  71.040000 242.690000  71.240000 ;
      RECT 241.700000  71.240000 242.620000  72.305000 ;
      RECT 241.700000  72.305000 242.360000  73.635000 ;
      RECT 241.815000  11.600000 241.985000  13.410000 ;
      RECT 241.815000  13.830000 241.985000  18.040000 ;
      RECT 241.815000  18.040000 242.600000  18.440000 ;
      RECT 241.815000  18.440000 245.790000  18.660000 ;
      RECT 241.840000  20.875000 242.100000  21.515000 ;
      RECT 241.885000  19.530000 242.055000  20.875000 ;
      RECT 241.885000  21.515000 242.055000  24.280000 ;
      RECT 241.910000  61.260000 242.440000  61.430000 ;
      RECT 241.925000  61.175000 242.435000  61.260000 ;
      RECT 241.925000  61.430000 242.435000  61.505000 ;
      RECT 241.925000  67.585000 242.435000  67.915000 ;
      RECT 241.960000  77.400000 242.435000  78.240000 ;
      RECT 241.960000  78.410000 242.435000  78.750000 ;
      RECT 241.960000  79.730000 242.435000  81.080000 ;
      RECT 241.995000  61.505000 242.365000  67.585000 ;
      RECT 242.065000  37.765000 242.235000  40.845000 ;
      RECT 242.070000 113.195000 242.740000 113.525000 ;
      RECT 242.075000  30.285000 242.245000  31.895000 ;
      RECT 242.075000  32.515000 242.245000  35.725000 ;
      RECT 242.090000  83.290000 243.320000  83.460000 ;
      RECT 242.095000  42.840000 242.265000  44.180000 ;
      RECT 242.115000   8.850000 242.645000   9.020000 ;
      RECT 242.175000 200.085000 242.845000 200.255000 ;
      RECT 242.175000 216.235000 242.845000 216.405000 ;
      RECT 242.180000  81.920000 242.510000  83.290000 ;
      RECT 242.180000  86.430000 243.340000  86.940000 ;
      RECT 242.250000  74.400000 242.420000  74.930000 ;
      RECT 242.250000  75.430000 242.420000  76.020000 ;
      RECT 242.265000  46.335000 242.795000  46.505000 ;
      RECT 242.265000  78.750000 242.435000  79.730000 ;
      RECT 242.345000  29.785000 242.855000  30.115000 ;
      RECT 242.345000  36.195000 242.855000  36.525000 ;
      RECT 242.390000  41.265000 243.355000  41.435000 ;
      RECT 242.390000  41.435000 242.700000  42.130000 ;
      RECT 242.390000  42.130000 242.920000  42.300000 ;
      RECT 242.415000  30.115000 242.785000  36.195000 ;
      RECT 242.475000   5.035000 242.645000   8.850000 ;
      RECT 242.475000   9.020000 242.645000   9.785000 ;
      RECT 242.510000  11.600000 242.680000  17.345000 ;
      RECT 242.520000  68.385000 248.290000  68.555000 ;
      RECT 242.525000  42.840000 242.695000  44.010000 ;
      RECT 242.530000  38.155000 242.815000  40.865000 ;
      RECT 242.530000  40.865000 242.700000  41.095000 ;
      RECT 242.535000  61.675000 242.705000  62.740000 ;
      RECT 242.535000  62.910000 242.705000  63.285000 ;
      RECT 242.535000  63.905000 242.705000  64.235000 ;
      RECT 242.535000  64.405000 242.705000  67.115000 ;
      RECT 242.620000  22.015000 242.880000  22.655000 ;
      RECT 242.625000  44.350000 242.795000  45.760000 ;
      RECT 242.625000  46.100000 242.795000  46.335000 ;
      RECT 242.625000  46.505000 242.795000  48.380000 ;
      RECT 242.665000  19.530000 242.835000  22.015000 ;
      RECT 242.665000  22.655000 242.835000  24.280000 ;
      RECT 242.730000  78.240000 243.320000  78.410000 ;
      RECT 242.730000  78.950000 243.320000  79.120000 ;
      RECT 242.770000  17.510000 243.300000  18.270000 ;
      RECT 242.780000  11.100000 243.290000  11.430000 ;
      RECT 242.805000  61.175000 243.315000  61.505000 ;
      RECT 242.805000  67.585000 243.315000  67.590000 ;
      RECT 242.805000  67.590000 244.195000  67.915000 ;
      RECT 242.815000   8.830000 243.085000  10.295000 ;
      RECT 242.850000  11.430000 243.220000  17.510000 ;
      RECT 242.865000 106.360000 243.395000 106.530000 ;
      RECT 242.870000  37.335000 245.125000  37.505000 ;
      RECT 242.870000  41.085000 243.540000  41.255000 ;
      RECT 242.870000  41.255000 243.355000  41.265000 ;
      RECT 242.870000  41.760000 243.400000  41.930000 ;
      RECT 242.875000  61.505000 243.245000  67.585000 ;
      RECT 242.955000  30.285000 243.125000  36.025000 ;
      RECT 242.955000 105.400000 243.125000 106.360000 ;
      RECT 242.955000 106.530000 243.125000 106.750000 ;
      RECT 242.970000  68.555000 243.140000  73.635000 ;
      RECT 242.985000  37.505000 245.125000  37.595000 ;
      RECT 242.985000  37.595000 243.355000  41.085000 ;
      RECT 242.985000  43.110000 243.515000  48.390000 ;
      RECT 242.990000  74.920000 243.320000  78.240000 ;
      RECT 242.990000  78.410000 243.320000  78.440000 ;
      RECT 242.990000  79.120000 243.320000  83.290000 ;
      RECT 242.990000  83.460000 243.320000  83.830000 ;
      RECT 243.090000  41.930000 243.400000  43.110000 ;
      RECT 243.225000  29.785000 244.615000  30.085000 ;
      RECT 243.225000  30.085000 243.735000  30.115000 ;
      RECT 243.225000  36.195000 243.735000  36.225000 ;
      RECT 243.225000  36.225000 244.620000  36.525000 ;
      RECT 243.240000  19.565000 243.500000  24.340000 ;
      RECT 243.255000   4.685000 243.425000   9.785000 ;
      RECT 243.275000 200.495000 243.805000 215.995000 ;
      RECT 243.285000  19.530000 243.455000  19.565000 ;
      RECT 243.295000  30.115000 243.665000  36.195000 ;
      RECT 243.390000  11.600000 243.560000  13.210000 ;
      RECT 243.390000  13.830000 243.560000  14.160000 ;
      RECT 243.390000  14.330000 243.560000  17.040000 ;
      RECT 243.415000  61.800000 243.585000  67.420000 ;
      RECT 243.470000  18.040000 245.790000  18.440000 ;
      RECT 243.525000  37.765000 243.695000  40.865000 ;
      RECT 243.570000  41.445000 244.035000  41.615000 ;
      RECT 243.570000  41.615000 243.740000  42.520000 ;
      RECT 243.570000  42.520000 243.855000  42.690000 ;
      RECT 243.580000 242.025000 248.775000 243.720000 ;
      RECT 243.605000 105.205000 248.355000 105.280000 ;
      RECT 243.605000 105.990000 248.355000 106.160000 ;
      RECT 243.605000 106.870000 248.355000 106.940000 ;
      RECT 243.650000  11.260000 244.180000  11.430000 ;
      RECT 243.660000  11.100000 244.170000  11.260000 ;
      RECT 243.660000  17.510000 244.170000  17.840000 ;
      RECT 243.685000  42.690000 243.855000  43.615000 ;
      RECT 243.685000  61.175000 244.195000  61.505000 ;
      RECT 243.685000  67.585000 244.195000  67.590000 ;
      RECT 243.730000  11.430000 244.100000  17.510000 ;
      RECT 243.750000  68.885000 243.920000  73.635000 ;
      RECT 243.755000  61.505000 244.125000  63.695000 ;
      RECT 243.755000  63.695000 244.285000  63.865000 ;
      RECT 243.755000  63.865000 244.125000  67.585000 ;
      RECT 243.780000  86.430000 244.940000  86.940000 ;
      RECT 243.800000  74.920000 244.130000  78.240000 ;
      RECT 243.800000  78.240000 244.390000  78.410000 ;
      RECT 243.800000  78.410000 244.130000  78.440000 ;
      RECT 243.800000  78.950000 244.390000  79.120000 ;
      RECT 243.800000  79.120000 244.130000  83.290000 ;
      RECT 243.800000  83.290000 245.030000  83.460000 ;
      RECT 243.800000  83.460000 244.130000  83.830000 ;
      RECT 243.835000  30.285000 244.005000  31.895000 ;
      RECT 243.835000  32.515000 244.005000  35.725000 ;
      RECT 243.865000  40.395000 244.575000  40.865000 ;
      RECT 243.865000  40.865000 244.035000  41.445000 ;
      RECT 243.910000  41.785000 244.530000  42.115000 ;
      RECT 243.910000 239.550000 248.775000 241.240000 ;
      RECT 243.970000   4.515000 245.365000   8.840000 ;
      RECT 243.970000   8.840000 247.970000  10.760000 ;
      RECT 243.970000  10.760000 252.915000  10.930000 ;
      RECT 244.020000  22.700000 244.280000  23.340000 ;
      RECT 244.065000  19.530000 244.235000  22.700000 ;
      RECT 244.065000  23.340000 244.235000  24.280000 ;
      RECT 244.105000  30.085000 244.615000  30.115000 ;
      RECT 244.110000  36.195000 244.620000  36.225000 ;
      RECT 244.135000  48.350000 247.505000  48.520000 ;
      RECT 244.145000 113.910000 247.145000 164.900000 ;
      RECT 244.175000  30.115000 244.545000  36.195000 ;
      RECT 244.175000  45.290000 244.345000  48.000000 ;
      RECT 244.205000  41.360000 245.125000  41.530000 ;
      RECT 244.205000  41.530000 244.530000  41.785000 ;
      RECT 244.235000 200.085000 244.905000 200.255000 ;
      RECT 244.235000 216.235000 244.905000 216.405000 ;
      RECT 244.270000  11.725000 244.440000  17.345000 ;
      RECT 244.295000  48.215000 247.345000  48.350000 ;
      RECT 244.295000  61.645000 244.675000  61.815000 ;
      RECT 244.295000  61.815000 244.465000  63.495000 ;
      RECT 244.295000  64.405000 244.465000  67.115000 ;
      RECT 244.365000  61.260000 244.895000  61.430000 ;
      RECT 244.405000  38.155000 244.575000  40.395000 ;
      RECT 244.490000  87.885000 245.290000  90.920000 ;
      RECT 244.490000  90.920000 265.275000  91.465000 ;
      RECT 244.490000  91.465000 290.580000  91.720000 ;
      RECT 244.505000  61.430000 244.675000  61.645000 ;
      RECT 244.530000  68.555000 244.700000  73.635000 ;
      RECT 244.540000  11.100000 245.050000  11.430000 ;
      RECT 244.540000  17.510000 245.050000  17.840000 ;
      RECT 244.565000  42.605000 244.735000  44.400000 ;
      RECT 244.580000  45.030000 245.125000  45.200000 ;
      RECT 244.610000  11.430000 244.980000  17.295000 ;
      RECT 244.610000  17.295000 245.140000  17.465000 ;
      RECT 244.610000  17.465000 245.050000  17.510000 ;
      RECT 244.610000  81.920000 244.940000  83.290000 ;
      RECT 244.670000  44.570000 245.680000  44.740000 ;
      RECT 244.670000  44.740000 245.200000  44.800000 ;
      RECT 244.685000  77.400000 245.160000  78.240000 ;
      RECT 244.685000  78.240000 245.590000  78.410000 ;
      RECT 244.685000  78.410000 245.160000  78.750000 ;
      RECT 244.685000  78.750000 244.855000  79.730000 ;
      RECT 244.685000  79.730000 245.160000  81.080000 ;
      RECT 244.700000  74.400000 244.870000  74.930000 ;
      RECT 244.700000  75.430000 244.870000  76.020000 ;
      RECT 244.715000  30.285000 244.885000  36.025000 ;
      RECT 244.745000  37.595000 245.125000  38.615000 ;
      RECT 244.785000  42.000000 245.455000  42.170000 ;
      RECT 244.800000  19.565000 245.060000  24.340000 ;
      RECT 244.845000  19.530000 245.015000  19.565000 ;
      RECT 244.845000  61.675000 245.015000  63.495000 ;
      RECT 244.845000  64.405000 245.015000  67.115000 ;
      RECT 244.855000  42.170000 245.385000  42.300000 ;
      RECT 244.955000  40.195000 245.125000  41.360000 ;
      RECT 244.955000  45.000000 245.125000  45.030000 ;
      RECT 244.955000  45.200000 245.125000  48.000000 ;
      RECT 244.985000  29.785000 246.375000  30.085000 ;
      RECT 244.985000  30.085000 245.495000  30.115000 ;
      RECT 244.985000  36.195000 245.495000  36.225000 ;
      RECT 244.985000  36.225000 246.375000  36.525000 ;
      RECT 245.055000  30.115000 245.425000  36.195000 ;
      RECT 245.055000  38.970000 246.585000  39.720000 ;
      RECT 245.070000  75.100000 248.460000  75.270000 ;
      RECT 245.085000  42.505000 245.615000  42.675000 ;
      RECT 245.115000  61.175000 245.625000  61.505000 ;
      RECT 245.115000  67.585000 245.625000  67.915000 ;
      RECT 245.115000  75.270000 245.645000  75.330000 ;
      RECT 245.115000  79.110000 245.645000  79.280000 ;
      RECT 245.125000  79.075000 245.635000  79.110000 ;
      RECT 245.125000  79.280000 245.635000  79.405000 ;
      RECT 245.150000  11.600000 245.320000  13.420000 ;
      RECT 245.150000  14.330000 245.320000  17.040000 ;
      RECT 245.175000  76.370000 248.905000  76.540000 ;
      RECT 245.185000  61.075000 245.355000  61.175000 ;
      RECT 245.185000  61.505000 245.555000  67.585000 ;
      RECT 245.230000  18.660000 245.610000  18.855000 ;
      RECT 245.230000  18.855000 249.860000  18.880000 ;
      RECT 245.230000  18.880000 255.935000  18.920000 ;
      RECT 245.230000  18.920000 255.820000  19.030000 ;
      RECT 245.230000  19.030000 253.325000  19.135000 ;
      RECT 245.230000  19.135000 245.610000  21.150000 ;
      RECT 245.295000  37.765000 246.345000  38.970000 ;
      RECT 245.295000  39.720000 246.345000  40.865000 ;
      RECT 245.305000  22.190000 245.695000  22.840000 ;
      RECT 245.305000  22.840000 247.250000  23.235000 ;
      RECT 245.310000  68.885000 245.480000  73.635000 ;
      RECT 245.335000 200.495000 245.865000 215.995000 ;
      RECT 245.445000  42.675000 245.615000  43.615000 ;
      RECT 245.445000 192.620000 245.955000 192.700000 ;
      RECT 245.445000 192.700000 245.985000 192.870000 ;
      RECT 245.445000 192.870000 245.955000 192.950000 ;
      RECT 245.460000  81.890000 245.630000  83.290000 ;
      RECT 245.460000  83.290000 246.010000  83.460000 ;
      RECT 245.460000  83.460000 245.630000  86.640000 ;
      RECT 245.595000  30.285000 245.765000  31.895000 ;
      RECT 245.595000  32.515000 245.765000  35.725000 ;
      RECT 245.595000  87.150000 246.265000  87.320000 ;
      RECT 245.700000  11.600000 245.870000  13.420000 ;
      RECT 245.700000  14.330000 245.870000  17.040000 ;
      RECT 245.710000  25.675000 245.970000  26.655000 ;
      RECT 245.725000  61.800000 245.895000  67.420000 ;
      RECT 245.735000  45.290000 245.905000  48.000000 ;
      RECT 245.755000  23.885000 245.925000  25.675000 ;
      RECT 245.815000  26.945000 252.840000  27.115000 ;
      RECT 245.830000  61.175000 246.505000  61.345000 ;
      RECT 245.835000 181.885000 250.545000 182.155000 ;
      RECT 245.835000 185.735000 250.545000 186.005000 ;
      RECT 245.835000 190.925000 250.545000 191.195000 ;
      RECT 245.865000  30.085000 246.375000  30.115000 ;
      RECT 245.865000  36.195000 246.375000  36.225000 ;
      RECT 245.925000  77.010000 246.935000  77.180000 ;
      RECT 245.925000  81.300000 246.935000  81.470000 ;
      RECT 245.935000  30.115000 246.305000  36.195000 ;
      RECT 245.960000  17.510000 246.490000  18.670000 ;
      RECT 245.960000  44.570000 246.970000  44.740000 ;
      RECT 245.970000  11.100000 246.480000  11.430000 ;
      RECT 245.995000  61.345000 246.505000  61.505000 ;
      RECT 245.995000  67.585000 246.505000  67.915000 ;
      RECT 246.005000  76.895000 246.535000  77.010000 ;
      RECT 246.015000   4.600000 271.435000   4.770000 ;
      RECT 246.015000  19.325000 246.605000  20.815000 ;
      RECT 246.015000  20.815000 246.690000  21.145000 ;
      RECT 246.015000  21.145000 246.605000  22.080000 ;
      RECT 246.015000  22.080000 248.660000  22.670000 ;
      RECT 246.025000  42.505000 246.555000  42.675000 ;
      RECT 246.025000  42.675000 246.195000  43.615000 ;
      RECT 246.040000  11.430000 246.410000  17.510000 ;
      RECT 246.065000  61.505000 246.435000  67.585000 ;
      RECT 246.090000  68.555000 246.260000  73.635000 ;
      RECT 246.090000  88.610000 246.260000  88.895000 ;
      RECT 246.090000  88.895000 246.620000  89.065000 ;
      RECT 246.095000   5.020000 246.265000   6.280000 ;
      RECT 246.095000   7.150000 246.265000   8.840000 ;
      RECT 246.175000  80.875000 246.705000  81.300000 ;
      RECT 246.185000  42.000000 246.855000  42.170000 ;
      RECT 246.240000  89.870000 267.165000  90.110000 ;
      RECT 246.255000  42.170000 246.785000  42.300000 ;
      RECT 246.285000  56.670000 246.455000  60.405000 ;
      RECT 246.295000 200.085000 246.965000 200.255000 ;
      RECT 246.295000 216.235000 246.965000 216.405000 ;
      RECT 246.315000  89.285000 266.110000  89.455000 ;
      RECT 246.340000  81.890000 246.510000  86.640000 ;
      RECT 246.340000 243.890000 248.695000 244.175000 ;
      RECT 246.340000 244.175000 247.775000 246.535000 ;
      RECT 246.340000 246.535000 248.695000 246.935000 ;
      RECT 246.440000  44.740000 246.970000  44.800000 ;
      RECT 246.475000  30.285000 246.645000  36.025000 ;
      RECT 246.490000  23.405000 247.680000  23.710000 ;
      RECT 246.490000  23.710000 246.750000  26.595000 ;
      RECT 246.500000 191.905000 283.670000 193.515000 ;
      RECT 246.515000  37.335000 248.770000  37.505000 ;
      RECT 246.515000  37.505000 248.655000  37.595000 ;
      RECT 246.515000  37.595000 246.895000  38.615000 ;
      RECT 246.515000  40.195000 246.685000  41.360000 ;
      RECT 246.515000  41.360000 247.435000  41.530000 ;
      RECT 246.515000  45.000000 246.685000  45.030000 ;
      RECT 246.515000  45.030000 247.060000  45.200000 ;
      RECT 246.515000  45.200000 246.685000  48.000000 ;
      RECT 246.575000  54.555000 246.745000  55.495000 ;
      RECT 246.575000  55.495000 247.105000  55.665000 ;
      RECT 246.580000  11.725000 246.750000  17.345000 ;
      RECT 246.605000  61.675000 246.775000  62.740000 ;
      RECT 246.605000  62.910000 246.775000  63.285000 ;
      RECT 246.605000  63.905000 246.775000  64.235000 ;
      RECT 246.605000  64.405000 246.775000  67.115000 ;
      RECT 246.625000  55.835000 247.295000  55.895000 ;
      RECT 246.625000  55.895000 247.340000  56.065000 ;
      RECT 246.625000  56.065000 247.295000  56.345000 ;
      RECT 246.625000  56.345000 246.895000  58.805000 ;
      RECT 246.625000  58.805000 247.235000  60.665000 ;
      RECT 246.625000  60.665000 249.390000  60.835000 ;
      RECT 246.660000  18.040000 249.860000  18.855000 ;
      RECT 246.745000  29.785000 248.135000  30.085000 ;
      RECT 246.745000  30.085000 247.255000  30.115000 ;
      RECT 246.745000  36.195000 247.255000  36.225000 ;
      RECT 246.745000  36.225000 248.135000  36.525000 ;
      RECT 246.785000  63.455000 247.315000  63.625000 ;
      RECT 246.815000  30.115000 247.185000  36.195000 ;
      RECT 246.830000  87.150000 248.860000  87.320000 ;
      RECT 246.850000  11.100000 247.360000  11.430000 ;
      RECT 246.850000  17.510000 247.360000  17.840000 ;
      RECT 246.870000  68.885000 247.040000  73.635000 ;
      RECT 246.875000  61.175000 247.385000  61.505000 ;
      RECT 246.875000  67.585000 247.385000  67.915000 ;
      RECT 246.905000  42.605000 247.075000  44.400000 ;
      RECT 246.920000  11.430000 247.290000  17.510000 ;
      RECT 246.945000  61.505000 247.315000  63.455000 ;
      RECT 246.945000  63.625000 247.315000  67.585000 ;
      RECT 246.990000  77.400000 247.160000  78.750000 ;
      RECT 246.990000  79.540000 247.160000  81.080000 ;
      RECT 247.030000  83.290000 247.560000  83.460000 ;
      RECT 247.065000  38.155000 247.235000  40.395000 ;
      RECT 247.065000  40.395000 247.775000  40.865000 ;
      RECT 247.065000  56.515000 248.270000  56.700000 ;
      RECT 247.065000  56.700000 247.235000  57.680000 ;
      RECT 247.110000  20.240000 247.370000  21.310000 ;
      RECT 247.110000  41.530000 247.435000  41.785000 ;
      RECT 247.110000  41.785000 247.730000  42.115000 ;
      RECT 247.115000  19.775000 252.825000  19.945000 ;
      RECT 247.195000  19.135000 253.325000  19.500000 ;
      RECT 247.205000  77.010000 248.215000  77.180000 ;
      RECT 247.205000  81.300000 248.215000  81.470000 ;
      RECT 247.220000  81.890000 247.390000  83.290000 ;
      RECT 247.220000  83.460000 247.390000  86.640000 ;
      RECT 247.270000  25.675000 247.530000  26.655000 ;
      RECT 247.285000  76.895000 247.815000  77.010000 ;
      RECT 247.295000  45.290000 247.465000  48.000000 ;
      RECT 247.315000  23.885000 247.485000  25.675000 ;
      RECT 247.355000  30.285000 247.525000  31.895000 ;
      RECT 247.355000  32.515000 247.525000  35.725000 ;
      RECT 247.375000   4.970000 247.905000   5.140000 ;
      RECT 247.375000   5.140000 247.545000   8.160000 ;
      RECT 247.395000 200.495000 247.925000 215.995000 ;
      RECT 247.420000  22.670000 247.680000  23.405000 ;
      RECT 247.455000  53.770000 247.985000  53.935000 ;
      RECT 247.455000  53.935000 248.945000  54.055000 ;
      RECT 247.455000  54.055000 250.105000  54.385000 ;
      RECT 247.455000  54.385000 247.985000  54.660000 ;
      RECT 247.455000  54.660000 247.625000  55.565000 ;
      RECT 247.455000  80.875000 247.985000  81.300000 ;
      RECT 247.460000  11.600000 247.630000  13.210000 ;
      RECT 247.460000  13.830000 247.630000  14.160000 ;
      RECT 247.460000  14.330000 247.630000  17.040000 ;
      RECT 247.485000  61.675000 247.655000  63.695000 ;
      RECT 247.485000  63.695000 248.745000  63.865000 ;
      RECT 247.485000  63.865000 247.655000  67.420000 ;
      RECT 247.605000  40.865000 247.775000  41.445000 ;
      RECT 247.605000  41.445000 248.070000  41.615000 ;
      RECT 247.625000  30.085000 248.135000  30.115000 ;
      RECT 247.625000  36.195000 248.135000  36.225000 ;
      RECT 247.635000  50.865000 247.805000  53.770000 ;
      RECT 247.650000  68.555000 247.820000  73.635000 ;
      RECT 247.695000  30.115000 248.065000  36.195000 ;
      RECT 247.715000   6.510000 249.405000   6.680000 ;
      RECT 247.715000  56.870000 248.610000  57.040000 ;
      RECT 247.715000  57.040000 247.885000  60.015000 ;
      RECT 247.730000  11.100000 248.240000  11.430000 ;
      RECT 247.730000  17.510000 248.240000  17.840000 ;
      RECT 247.740000  56.265000 248.270000  56.515000 ;
      RECT 247.760000  55.735000 248.270000  56.265000 ;
      RECT 247.785000  42.520000 248.070000  42.690000 ;
      RECT 247.785000  42.690000 247.955000  43.615000 ;
      RECT 247.800000  11.430000 248.170000  17.510000 ;
      RECT 247.890000  21.125000 248.150000  21.765000 ;
      RECT 247.890000  23.495000 248.150000  26.595000 ;
      RECT 247.900000  41.615000 248.070000  42.520000 ;
      RECT 247.935000  20.300000 248.105000  21.125000 ;
      RECT 247.945000  37.765000 248.115000  40.865000 ;
      RECT 247.945000 244.345000 248.695000 246.365000 ;
      RECT 247.985000 181.105000 250.545000 181.375000 ;
      RECT 247.985000 186.515000 250.545000 186.785000 ;
      RECT 247.985000 190.145000 250.545000 190.415000 ;
      RECT 248.035000  61.675000 248.205000  63.495000 ;
      RECT 248.035000  64.405000 248.205000  67.115000 ;
      RECT 248.065000  52.355000 248.575000  52.685000 ;
      RECT 248.100000  41.085000 248.770000  41.255000 ;
      RECT 248.100000  81.890000 248.270000  86.640000 ;
      RECT 248.125000  43.110000 248.655000  48.390000 ;
      RECT 248.175000 221.215000 248.345000 231.605000 ;
      RECT 248.175000 232.050000 248.345000 238.575000 ;
      RECT 248.235000  30.285000 248.405000  36.025000 ;
      RECT 248.240000  41.760000 248.770000  41.930000 ;
      RECT 248.240000  41.930000 248.550000  43.110000 ;
      RECT 248.275000  50.535000 249.365000  50.705000 ;
      RECT 248.275000  50.705000 248.445000  52.355000 ;
      RECT 248.275000  52.685000 248.445000  52.840000 ;
      RECT 248.285000  37.595000 248.655000  41.085000 ;
      RECT 248.285000  41.255000 248.770000  41.265000 ;
      RECT 248.285000  41.265000 249.250000  41.435000 ;
      RECT 248.305000  61.175000 248.815000  61.505000 ;
      RECT 248.305000  67.585000 248.815000  67.590000 ;
      RECT 248.305000  67.590000 249.695000  67.915000 ;
      RECT 248.325000 244.175000 248.695000 244.345000 ;
      RECT 248.325000 246.365000 248.695000 246.535000 ;
      RECT 248.335000  54.555000 248.610000  54.920000 ;
      RECT 248.335000  54.920000 248.865000  55.090000 ;
      RECT 248.335000  55.090000 248.610000  55.565000 ;
      RECT 248.340000  11.600000 248.510000  17.345000 ;
      RECT 248.355000 200.085000 249.025000 200.255000 ;
      RECT 248.355000 216.235000 249.025000 216.405000 ;
      RECT 248.375000  61.505000 248.745000  63.695000 ;
      RECT 248.375000  63.865000 248.745000  67.585000 ;
      RECT 248.430000  68.885000 248.600000  73.635000 ;
      RECT 248.440000  55.565000 248.610000  56.870000 ;
      RECT 248.450000  79.120000 249.015000  79.290000 ;
      RECT 248.460000  11.260000 248.990000  11.430000 ;
      RECT 248.470000  49.415000 249.140000  50.365000 ;
      RECT 248.495000  57.305000 248.665000  60.405000 ;
      RECT 248.505000  29.785000 249.015000  30.115000 ;
      RECT 248.505000  36.195000 249.015000  36.525000 ;
      RECT 248.505000  79.075000 249.015000  79.120000 ;
      RECT 248.505000  79.290000 249.015000  79.405000 ;
      RECT 248.530000 113.195000 249.200000 113.525000 ;
      RECT 248.560000  78.240000 249.400000  78.410000 ;
      RECT 248.575000  30.115000 248.945000  36.195000 ;
      RECT 248.620000  83.290000 249.150000  83.460000 ;
      RECT 248.655000   5.020000 248.825000   6.280000 ;
      RECT 248.655000   7.080000 248.825000   9.790000 ;
      RECT 248.655000  68.205000 249.325000  68.555000 ;
      RECT 248.655000 113.910000 251.655000 164.900000 ;
      RECT 248.670000  20.240000 248.930000  21.310000 ;
      RECT 248.670000  25.675000 248.930000  26.655000 ;
      RECT 248.705000 104.700000 248.875000 107.450000 ;
      RECT 248.715000  23.885000 248.885000  25.675000 ;
      RECT 248.720000  42.130000 249.250000  42.300000 ;
      RECT 248.735000  50.875000 248.945000  51.885000 ;
      RECT 248.735000  52.875000 248.945000  53.935000 ;
      RECT 248.745000  51.885000 248.945000  52.875000 ;
      RECT 248.780000  54.385000 250.105000  54.660000 ;
      RECT 248.780000  55.525000 249.310000  57.005000 ;
      RECT 248.780000  57.005000 249.445000  57.175000 ;
      RECT 248.810000  57.175000 249.445000  57.205000 ;
      RECT 248.820000  11.430000 248.990000  11.600000 ;
      RECT 248.820000  11.600000 249.060000  17.345000 ;
      RECT 248.825000  38.155000 249.110000  40.865000 ;
      RECT 248.845000  44.180000 250.405000  44.350000 ;
      RECT 248.845000  44.350000 249.015000  45.760000 ;
      RECT 248.845000  45.760000 251.375000  45.930000 ;
      RECT 248.845000  46.100000 249.015000  46.335000 ;
      RECT 248.845000  46.335000 249.375000  46.505000 ;
      RECT 248.845000  46.505000 249.015000  48.380000 ;
      RECT 248.915000  61.800000 249.085000  67.420000 ;
      RECT 248.940000  22.080000 250.220000  22.670000 ;
      RECT 248.940000  40.865000 249.110000  41.095000 ;
      RECT 248.940000  41.435000 249.250000  42.130000 ;
      RECT 248.945000  42.840000 249.115000  44.010000 ;
      RECT 248.980000  74.420000 249.150000  76.020000 ;
      RECT 248.980000  77.400000 249.400000  78.240000 ;
      RECT 248.980000  78.410000 249.400000  78.750000 ;
      RECT 248.980000  79.730000 249.400000  81.080000 ;
      RECT 248.980000  81.890000 249.150000  83.290000 ;
      RECT 248.980000  83.460000 249.150000  86.640000 ;
      RECT 249.105000 220.065000 346.520000 220.085000 ;
      RECT 249.105000 220.085000 249.955000 247.105000 ;
      RECT 249.115000  30.285000 249.285000  31.895000 ;
      RECT 249.115000  32.515000 249.285000  35.725000 ;
      RECT 249.150000  10.390000 249.680000  10.560000 ;
      RECT 249.160000  11.100000 249.670000  11.430000 ;
      RECT 249.160000  17.510000 249.670000  17.840000 ;
      RECT 249.170000  10.260000 249.680000  10.390000 ;
      RECT 249.170000  10.560000 249.680000  10.590000 ;
      RECT 249.185000  61.175000 249.695000  61.505000 ;
      RECT 249.185000  67.585000 249.695000  67.590000 ;
      RECT 249.195000  50.705000 249.365000  51.885000 ;
      RECT 249.195000  52.875000 249.365000  53.885000 ;
      RECT 249.210000  68.885000 249.380000  73.635000 ;
      RECT 249.220000  52.230000 249.750000  52.400000 ;
      RECT 249.230000  11.430000 249.600000  17.510000 ;
      RECT 249.230000  42.470000 250.580000  42.640000 ;
      RECT 249.230000  78.750000 249.400000  79.730000 ;
      RECT 249.255000  61.505000 249.625000  67.585000 ;
      RECT 249.275000  57.205000 249.445000  60.015000 ;
      RECT 249.330000  42.640000 250.580000  42.670000 ;
      RECT 249.375000  42.840000 249.545000  44.180000 ;
      RECT 249.385000  29.785000 249.895000  30.115000 ;
      RECT 249.385000  36.195000 249.895000  36.525000 ;
      RECT 249.405000  37.765000 249.575000  40.845000 ;
      RECT 249.420000  52.095000 249.750000  52.230000 ;
      RECT 249.420000  52.400000 249.750000  52.605000 ;
      RECT 249.455000  30.115000 249.825000  36.195000 ;
      RECT 249.455000 200.495000 249.985000 215.995000 ;
      RECT 249.470000  81.950000 249.640000  85.820000 ;
      RECT 249.470000  85.820000 249.650000  86.350000 ;
      RECT 249.470000  86.350000 249.640000  86.765000 ;
      RECT 249.495000  20.300000 249.665000  21.655000 ;
      RECT 249.495000  23.670000 249.665000  26.595000 ;
      RECT 249.550000  70.860000 250.360000  71.415000 ;
      RECT 249.550000  71.415000 250.440000  72.305000 ;
      RECT 249.550000  72.305000 250.360000  72.365000 ;
      RECT 249.570000  74.400000 249.740000  81.020000 ;
      RECT 249.575000  51.740000 250.105000  51.910000 ;
      RECT 249.575000  53.770000 250.105000  54.055000 ;
      RECT 249.640000 103.770000 249.810000 108.380000 ;
      RECT 249.655000  50.875000 250.105000  51.740000 ;
      RECT 249.655000  52.775000 250.105000  53.770000 ;
      RECT 249.700000  68.635000 249.870000  68.925000 ;
      RECT 249.700000  68.925000 250.360000  70.860000 ;
      RECT 249.700000  72.365000 250.360000  73.610000 ;
      RECT 249.755000   6.510000 250.285000   6.680000 ;
      RECT 249.770000  11.600000 249.940000  13.210000 ;
      RECT 249.770000  13.830000 249.940000  14.160000 ;
      RECT 249.770000  14.330000 249.940000  17.040000 ;
      RECT 249.795000  61.675000 249.965000  62.740000 ;
      RECT 249.795000  62.910000 249.965000  63.285000 ;
      RECT 249.795000  63.905000 249.965000  64.235000 ;
      RECT 249.795000  64.405000 249.965000  67.115000 ;
      RECT 249.805000  42.840000 249.975000  44.010000 ;
      RECT 249.885000  63.455000 250.505000  63.625000 ;
      RECT 249.900000  81.450000 250.570000  81.940000 ;
      RECT 249.915000  56.265000 250.445000  56.435000 ;
      RECT 249.920000  51.910000 250.105000  52.775000 ;
      RECT 249.935000   5.020000 250.105000   6.510000 ;
      RECT 249.935000   6.680000 250.105000   9.790000 ;
      RECT 249.955000  57.325000 250.125000  60.405000 ;
      RECT 249.960000  82.180000 250.130000  86.930000 ;
      RECT 249.995000  30.285000 250.165000  36.045000 ;
      RECT 250.025000  44.580000 250.195000  45.280000 ;
      RECT 250.025000  45.280000 250.700000  45.450000 ;
      RECT 250.025000  45.450000 250.195000  45.590000 ;
      RECT 250.025000  46.100000 250.195000  48.550000 ;
      RECT 250.025000  48.550000 252.915000  48.720000 ;
      RECT 250.025000  74.000000 250.700000  74.170000 ;
      RECT 250.030000  17.510000 250.560000  18.670000 ;
      RECT 250.035000 181.075000 250.545000 181.105000 ;
      RECT 250.035000 181.375000 250.545000 181.405000 ;
      RECT 250.035000 181.855000 250.545000 181.885000 ;
      RECT 250.035000 182.155000 250.545000 182.185000 ;
      RECT 250.035000 185.705000 250.545000 185.735000 ;
      RECT 250.035000 186.005000 250.545000 186.035000 ;
      RECT 250.035000 186.485000 250.545000 186.515000 ;
      RECT 250.035000 186.785000 250.545000 186.815000 ;
      RECT 250.035000 190.115000 250.545000 190.145000 ;
      RECT 250.035000 190.415000 250.545000 190.445000 ;
      RECT 250.035000 190.895000 250.545000 190.925000 ;
      RECT 250.035000 191.195000 250.545000 191.225000 ;
      RECT 250.040000  11.100000 250.550000  11.430000 ;
      RECT 250.065000  61.175000 250.575000  61.505000 ;
      RECT 250.065000  67.585000 250.575000  67.915000 ;
      RECT 250.110000  11.430000 250.480000  17.510000 ;
      RECT 250.135000  61.505000 250.505000  63.455000 ;
      RECT 250.135000  63.625000 250.505000  67.585000 ;
      RECT 250.160000  68.205000 250.830000  68.375000 ;
      RECT 250.160000  68.375000 250.910000  68.545000 ;
      RECT 250.230000  20.240000 250.490000  21.310000 ;
      RECT 250.230000  25.675000 250.490000  26.655000 ;
      RECT 250.235000  42.840000 250.405000  44.180000 ;
      RECT 250.250000  87.150000 251.600000  87.320000 ;
      RECT 250.265000  29.785000 251.655000  30.115000 ;
      RECT 250.265000  36.195000 251.655000  36.525000 ;
      RECT 250.275000  23.885000 250.445000  25.675000 ;
      RECT 250.275000  50.845000 250.445000  53.370000 ;
      RECT 250.275000  53.370000 250.805000  53.540000 ;
      RECT 250.275000  53.540000 250.445000  56.265000 ;
      RECT 250.305000   6.880000 250.835000   7.050000 ;
      RECT 250.335000  30.115000 250.705000  36.195000 ;
      RECT 250.415000 200.085000 251.085000 200.255000 ;
      RECT 250.415000 216.235000 251.085000 216.405000 ;
      RECT 250.430000  49.090000 251.100000  50.625000 ;
      RECT 250.445000  73.930000 250.700000  74.000000 ;
      RECT 250.445000  74.170000 250.700000  74.200000 ;
      RECT 250.445000  74.200000 250.615000  74.760000 ;
      RECT 250.445000  74.760000 250.730000  75.770000 ;
      RECT 250.470000  77.080000 251.000000  77.250000 ;
      RECT 250.485000   5.020000 250.655000   6.880000 ;
      RECT 250.485000   7.050000 250.655000   9.790000 ;
      RECT 250.490000  76.575000 250.660000  77.080000 ;
      RECT 250.500000  22.080000 252.380000  22.670000 ;
      RECT 250.525000  46.165000 250.855000  47.015000 ;
      RECT 250.530000  73.490000 251.140000  73.660000 ;
      RECT 250.530000  73.660000 250.700000  73.930000 ;
      RECT 250.575000 104.530000 268.095000 104.700000 ;
      RECT 250.575000 104.700000 250.745000 107.065000 ;
      RECT 250.575000 107.065000 267.055000 107.090000 ;
      RECT 250.575000 107.090000 268.095000 107.620000 ;
      RECT 250.605000  47.015000 250.775000  47.625000 ;
      RECT 250.630000  53.995000 250.960000  54.325000 ;
      RECT 250.635000  55.785000 250.965000  55.895000 ;
      RECT 250.635000  55.895000 251.165000  56.065000 ;
      RECT 250.635000  56.065000 250.965000  56.295000 ;
      RECT 250.650000  11.725000 250.820000  17.345000 ;
      RECT 250.665000  42.840000 250.835000  44.010000 ;
      RECT 250.670000  83.690000 251.200000  83.860000 ;
      RECT 250.675000  61.675000 250.845000  67.415000 ;
      RECT 250.715000 181.235000 250.885000 181.560000 ;
      RECT 250.715000 181.560000 251.245000 182.730000 ;
      RECT 250.715000 182.730000 268.770000 185.070000 ;
      RECT 250.715000 185.070000 251.245000 187.295000 ;
      RECT 250.715000 187.295000 268.770000 189.635000 ;
      RECT 250.715000 189.635000 251.245000 190.805000 ;
      RECT 250.720000 221.230000 341.150000 222.080000 ;
      RECT 250.720000 222.080000 251.570000 245.255000 ;
      RECT 250.720000 245.255000 341.150000 246.105000 ;
      RECT 250.730000  18.040000 258.600000  18.210000 ;
      RECT 250.730000  18.210000 255.935000  18.880000 ;
      RECT 250.740000  78.075000 250.910000  81.430000 ;
      RECT 250.740000  81.430000 251.010000  81.600000 ;
      RECT 250.750000  37.870000 250.920000  40.870000 ;
      RECT 250.785000  74.370000 254.905000  74.540000 ;
      RECT 250.840000  81.600000 251.010000  83.690000 ;
      RECT 250.840000  83.860000 251.010000  86.930000 ;
      RECT 250.845000   6.510000 252.875000   6.680000 ;
      RECT 250.865000  77.700000 251.535000  77.870000 ;
      RECT 250.870000  73.830000 252.190000  74.370000 ;
      RECT 250.875000  30.285000 251.045000  31.895000 ;
      RECT 250.875000  32.515000 251.045000  35.725000 ;
      RECT 250.910000   9.990000 251.440000  10.590000 ;
      RECT 250.910000  11.260000 251.440000  11.430000 ;
      RECT 250.920000  11.100000 251.430000  11.260000 ;
      RECT 250.920000  17.510000 251.430000  17.840000 ;
      RECT 250.935000  42.470000 252.285000  42.475000 ;
      RECT 250.935000  42.475000 253.595000  42.645000 ;
      RECT 250.945000  61.175000 251.455000  61.505000 ;
      RECT 250.945000  67.585000 251.455000  67.915000 ;
      RECT 250.970000  41.360000 251.500000  41.530000 ;
      RECT 250.970000  72.600000 251.140000  72.935000 ;
      RECT 250.970000  72.935000 251.500000  73.105000 ;
      RECT 250.970000  73.105000 251.140000  73.490000 ;
      RECT 250.990000  11.430000 251.360000  17.510000 ;
      RECT 251.015000  61.505000 251.385000  67.585000 ;
      RECT 251.055000  20.300000 251.225000  21.570000 ;
      RECT 251.055000  23.670000 251.225000  26.595000 ;
      RECT 251.075000 181.235000 251.245000 181.560000 ;
      RECT 251.090000 113.195000 251.760000 113.525000 ;
      RECT 251.095000  42.840000 251.265000  44.180000 ;
      RECT 251.095000  44.180000 252.915000  44.350000 ;
      RECT 251.095000 105.040000 267.585000 105.210000 ;
      RECT 251.095000 105.210000 255.845000 105.280000 ;
      RECT 251.095000 105.990000 255.845000 106.160000 ;
      RECT 251.095000 106.870000 256.210000 106.920000 ;
      RECT 251.095000 106.920000 267.055000 107.065000 ;
      RECT 251.120000  70.655000 251.995000  71.185000 ;
      RECT 251.120000  71.185000 251.630000  72.250000 ;
      RECT 251.155000  50.845000 251.325000  55.525000 ;
      RECT 251.165000  58.725000 252.055000  59.255000 ;
      RECT 251.170000  76.420000 256.070000  76.590000 ;
      RECT 251.170000  77.300000 256.450000  77.480000 ;
      RECT 251.205000  44.580000 251.375000  45.760000 ;
      RECT 251.205000  45.930000 251.375000  47.080000 ;
      RECT 251.205000  47.370000 252.075000  48.380000 ;
      RECT 251.205000  56.755000 252.055000  58.725000 ;
      RECT 251.205000  59.255000 252.055000  60.485000 ;
      RECT 251.215000  30.115000 251.585000  36.195000 ;
      RECT 251.250000  74.790000 251.780000  74.960000 ;
      RECT 251.270000  76.065000 252.320000  76.190000 ;
      RECT 251.270000  76.190000 252.160000  76.235000 ;
      RECT 251.330000  37.840000 255.570000  38.010000 ;
      RECT 251.330000  38.010000 251.500000  41.360000 ;
      RECT 251.380000  49.005000 252.580000  49.175000 ;
      RECT 251.380000  49.175000 252.050000  50.625000 ;
      RECT 251.380000  55.785000 251.710000  56.265000 ;
      RECT 251.380000  56.265000 251.910000  56.435000 ;
      RECT 251.415000 181.075000 251.925000 181.105000 ;
      RECT 251.415000 181.105000 253.975000 181.375000 ;
      RECT 251.415000 181.375000 251.925000 181.405000 ;
      RECT 251.415000 181.855000 251.925000 181.885000 ;
      RECT 251.415000 181.885000 256.125000 182.155000 ;
      RECT 251.415000 182.155000 251.925000 182.185000 ;
      RECT 251.415000 185.705000 251.925000 185.735000 ;
      RECT 251.415000 185.735000 256.125000 186.005000 ;
      RECT 251.415000 186.005000 251.925000 186.035000 ;
      RECT 251.415000 186.485000 251.925000 186.515000 ;
      RECT 251.415000 186.515000 253.975000 186.785000 ;
      RECT 251.415000 186.785000 251.925000 186.815000 ;
      RECT 251.440000  74.760000 251.610000  74.790000 ;
      RECT 251.440000  74.960000 251.610000  75.770000 ;
      RECT 251.515000 200.495000 252.045000 215.995000 ;
      RECT 251.525000  42.840000 251.695000  44.010000 ;
      RECT 251.530000  11.600000 251.700000  13.420000 ;
      RECT 251.530000  14.330000 251.700000  17.040000 ;
      RECT 251.545000  46.335000 252.075000  47.370000 ;
      RECT 251.555000  37.335000 253.585000  37.505000 ;
      RECT 251.555000  61.675000 251.725000  62.725000 ;
      RECT 251.555000  62.955000 251.725000  63.285000 ;
      RECT 251.555000  63.905000 251.725000  64.235000 ;
      RECT 251.555000  64.405000 251.725000  67.115000 ;
      RECT 251.620000  78.075000 251.790000  80.785000 ;
      RECT 251.650000  76.020000 252.320000  76.065000 ;
      RECT 251.720000  82.180000 251.890000  86.930000 ;
      RECT 251.750000  72.600000 251.970000  73.610000 ;
      RECT 251.755000  30.285000 251.925000  36.030000 ;
      RECT 251.765000   5.020000 251.935000   6.280000 ;
      RECT 251.765000   7.080000 251.935000   9.790000 ;
      RECT 251.790000  20.240000 252.050000  21.310000 ;
      RECT 251.790000  25.675000 252.050000  26.655000 ;
      RECT 251.800000  71.380000 251.970000  72.600000 ;
      RECT 251.835000  23.885000 252.005000  25.675000 ;
      RECT 251.865000  77.700000 252.535000  77.870000 ;
      RECT 251.885000  55.895000 252.415000  56.065000 ;
      RECT 251.920000  68.205000 252.590000  68.545000 ;
      RECT 251.955000  42.840000 252.125000  44.180000 ;
      RECT 251.980000  81.400000 252.510000  81.430000 ;
      RECT 251.980000  81.430000 252.650000  81.600000 ;
      RECT 252.005000  29.945000 252.535000  30.115000 ;
      RECT 252.025000  29.785000 252.535000  29.945000 ;
      RECT 252.025000  36.195000 252.535000  36.525000 ;
      RECT 252.025000  45.280000 252.555000  45.450000 ;
      RECT 252.035000  50.845000 252.870000  54.705000 ;
      RECT 252.035000  54.705000 252.205000  55.895000 ;
      RECT 252.080000  11.600000 252.250000  13.420000 ;
      RECT 252.080000  14.330000 252.250000  17.040000 ;
      RECT 252.095000  30.115000 252.465000  36.195000 ;
      RECT 252.105000  61.675000 252.275000  63.495000 ;
      RECT 252.105000  64.405000 252.275000  67.115000 ;
      RECT 252.145000 180.765000 267.095000 180.935000 ;
      RECT 252.145000 181.545000 267.095000 181.715000 ;
      RECT 252.145000 182.325000 267.095000 182.495000 ;
      RECT 252.145000 185.395000 267.095000 185.565000 ;
      RECT 252.145000 186.175000 267.095000 186.345000 ;
      RECT 252.145000 186.955000 267.095000 187.125000 ;
      RECT 252.210000  38.180000 252.470000  41.160000 ;
      RECT 252.235000 189.805000 267.185000 189.975000 ;
      RECT 252.235000 190.585000 267.185000 190.755000 ;
      RECT 252.235000 191.365000 267.185000 191.535000 ;
      RECT 252.240000  83.690000 252.770000  83.860000 ;
      RECT 252.320000  74.760000 253.030000  75.770000 ;
      RECT 252.335000 222.845000 339.535000 223.695000 ;
      RECT 252.335000 223.695000 253.185000 243.640000 ;
      RECT 252.335000 243.640000 339.535000 244.490000 ;
      RECT 252.340000  17.700000 252.870000  17.870000 ;
      RECT 252.350000  11.100000 252.860000  11.430000 ;
      RECT 252.350000  17.510000 252.860000  17.700000 ;
      RECT 252.375000  61.175000 252.885000  61.505000 ;
      RECT 252.375000  67.585000 252.885000  67.915000 ;
      RECT 252.385000  42.840000 252.555000  44.010000 ;
      RECT 252.385000  44.580000 252.555000  45.280000 ;
      RECT 252.385000  45.450000 252.555000  47.080000 ;
      RECT 252.385000  47.370000 252.915000  48.550000 ;
      RECT 252.390000  68.925000 252.740000  74.000000 ;
      RECT 252.390000  74.000000 252.980000  74.170000 ;
      RECT 252.420000  11.430000 252.790000  17.510000 ;
      RECT 252.445000  61.505000 252.815000  67.585000 ;
      RECT 252.475000 200.085000 253.145000 200.255000 ;
      RECT 252.475000 216.235000 253.145000 216.405000 ;
      RECT 252.490000  75.770000 253.030000  76.420000 ;
      RECT 252.495000 244.490000 331.140000 244.520000 ;
      RECT 252.500000  78.075000 252.670000  80.785000 ;
      RECT 252.600000  82.180000 252.770000  83.690000 ;
      RECT 252.600000  83.860000 252.770000  86.930000 ;
      RECT 252.615000  20.300000 252.785000  21.570000 ;
      RECT 252.615000  23.670000 252.785000  26.595000 ;
      RECT 252.635000  30.285000 252.805000  31.895000 ;
      RECT 252.635000  32.515000 252.805000  35.725000 ;
      RECT 252.665000  55.085000 255.195000  55.285000 ;
      RECT 252.665000  55.285000 252.835000  60.365000 ;
      RECT 252.670000  38.180000 252.930000  41.160000 ;
      RECT 252.700000  49.955000 252.870000  50.845000 ;
      RECT 252.725000  43.095000 253.255000  43.265000 ;
      RECT 252.725000  44.350000 252.915000  47.370000 ;
      RECT 252.745000   8.840000 256.200000   9.010000 ;
      RECT 252.745000   9.010000 252.915000  10.760000 ;
      RECT 252.835000  77.480000 253.725000  77.620000 ;
      RECT 252.845000  41.360000 253.375000  41.530000 ;
      RECT 252.885000  29.575000 253.415000  30.115000 ;
      RECT 252.905000  36.195000 253.415000  36.525000 ;
      RECT 252.930000  60.535000 256.660000  60.855000 ;
      RECT 252.935000  49.595000 255.815000  49.765000 ;
      RECT 252.960000  11.725000 253.130000  17.345000 ;
      RECT 252.960000  69.125000 253.490000  71.415000 ;
      RECT 252.960000  71.415000 253.850000  72.305000 ;
      RECT 252.960000  72.305000 253.490000  72.365000 ;
      RECT 252.960000  73.405000 253.510000  73.575000 ;
      RECT 252.975000  30.115000 253.345000  36.195000 ;
      RECT 252.980000  73.120000 253.510000  73.405000 ;
      RECT 252.985000  61.800000 253.155000  67.420000 ;
      RECT 253.025000  41.530000 253.195000  42.305000 ;
      RECT 253.045000   5.020000 253.215000   8.160000 ;
      RECT 253.085000  43.265000 253.255000  48.390000 ;
      RECT 253.160000  78.130000 253.330000  81.050000 ;
      RECT 253.160000  81.950000 253.330000  84.850000 ;
      RECT 253.165000 113.910000 256.165000 164.900000 ;
      RECT 253.200000  74.760000 253.370000  74.790000 ;
      RECT 253.200000  74.790000 253.730000  74.960000 ;
      RECT 253.200000  74.960000 253.370000  75.770000 ;
      RECT 253.220000  17.700000 253.750000  17.870000 ;
      RECT 253.230000  11.100000 253.740000  11.430000 ;
      RECT 253.230000  17.510000 253.740000  17.700000 ;
      RECT 253.255000  61.175000 253.765000  61.505000 ;
      RECT 253.255000  67.585000 253.765000  67.915000 ;
      RECT 253.265000  20.410000 253.435000  25.940000 ;
      RECT 253.300000  11.430000 253.670000  17.510000 ;
      RECT 253.325000  61.505000 253.695000  67.585000 ;
      RECT 253.385000   4.970000 253.915000   6.680000 ;
      RECT 253.410000  76.020000 254.080000  76.190000 ;
      RECT 253.425000  42.645000 253.595000  43.405000 ;
      RECT 253.425000  43.405000 254.075000  44.415000 ;
      RECT 253.455000  85.555000 256.430000  85.785000 ;
      RECT 253.455000  85.785000 256.565000  86.315000 ;
      RECT 253.455000  86.315000 256.430000  87.700000 ;
      RECT 253.480000  49.955000 253.650000  55.085000 ;
      RECT 253.515000  30.260000 253.895000  36.030000 ;
      RECT 253.545000  41.290000 254.215000  41.460000 ;
      RECT 253.545000  46.335000 254.075000  46.505000 ;
      RECT 253.565000  47.855000 253.735000  48.465000 ;
      RECT 253.565000  48.465000 259.095000  48.635000 ;
      RECT 253.575000 200.495000 254.105000 215.995000 ;
      RECT 253.585000  29.945000 254.115000  30.115000 ;
      RECT 253.585000  30.115000 253.895000  30.260000 ;
      RECT 253.605000  42.030000 254.135000  42.200000 ;
      RECT 253.615000  21.340000 254.025000  22.850000 ;
      RECT 253.615000  22.850000 255.065000  23.360000 ;
      RECT 253.615000  23.360000 254.025000  23.375000 ;
      RECT 253.640000  38.180000 253.810000  41.290000 ;
      RECT 253.640000  41.460000 254.135000  42.030000 ;
      RECT 253.650000  81.810000 254.870000  81.980000 ;
      RECT 253.650000  81.980000 253.820000  84.280000 ;
      RECT 253.650000  84.280000 254.180000  84.450000 ;
      RECT 253.650000  84.450000 253.820000  84.930000 ;
      RECT 253.680000  68.635000 253.850000  71.415000 ;
      RECT 253.680000  72.305000 253.850000  73.575000 ;
      RECT 253.715000  81.325000 254.385000  81.570000 ;
      RECT 253.735000 189.975000 263.035000 190.415000 ;
      RECT 253.735000 190.925000 263.035000 191.365000 ;
      RECT 253.795000  37.335000 254.465000  37.505000 ;
      RECT 253.810000 223.695000 254.420000 225.350000 ;
      RECT 253.820000  78.070000 253.990000  80.780000 ;
      RECT 253.840000  11.600000 254.010000  13.210000 ;
      RECT 253.840000  13.830000 254.010000  14.160000 ;
      RECT 253.840000  14.330000 254.010000  17.040000 ;
      RECT 253.845000  55.455000 254.015000  60.365000 ;
      RECT 253.865000  61.675000 254.035000  62.740000 ;
      RECT 253.865000  62.910000 254.035000  63.285000 ;
      RECT 253.865000  63.905000 254.035000  64.235000 ;
      RECT 253.865000  64.405000 254.035000  67.115000 ;
      RECT 253.905000  44.415000 254.075000  46.335000 ;
      RECT 253.905000  46.505000 254.075000  48.085000 ;
      RECT 253.910000 225.650000 254.080000 226.630000 ;
      RECT 253.910000 226.630000 313.675000 227.730000 ;
      RECT 253.910000 227.730000 314.225000 228.050000 ;
      RECT 253.910000 228.220000 313.205000 229.255000 ;
      RECT 253.910000 232.355000 313.205000 233.390000 ;
      RECT 253.910000 233.560000 323.690000 234.410000 ;
      RECT 253.910000 234.410000 313.675000 234.980000 ;
      RECT 253.910000 234.980000 254.080000 235.960000 ;
      RECT 253.910000 237.100000 254.080000 238.080000 ;
      RECT 253.910000 238.080000 301.130000 239.500000 ;
      RECT 253.910000 239.670000 301.260000 240.705000 ;
      RECT 253.945000  77.700000 254.615000  77.870000 ;
      RECT 253.965000  53.370000 254.495000  53.540000 ;
      RECT 254.065000  30.285000 254.235000  32.105000 ;
      RECT 254.065000  33.015000 254.235000  35.725000 ;
      RECT 254.080000  74.760000 254.780000  75.770000 ;
      RECT 254.110000  11.100000 254.620000  11.430000 ;
      RECT 254.110000  17.510000 254.620000  17.840000 ;
      RECT 254.110000  19.550000 255.630000  21.085000 ;
      RECT 254.145000  23.610000 254.315000  26.080000 ;
      RECT 254.180000  11.430000 254.550000  17.510000 ;
      RECT 254.245000  45.000000 254.775000  45.170000 ;
      RECT 254.245000  49.955000 254.415000  53.370000 ;
      RECT 254.245000  53.540000 254.415000  54.705000 ;
      RECT 254.250000  75.770000 254.780000  76.250000 ;
      RECT 254.305000  41.635000 254.555000  42.305000 ;
      RECT 254.325000   5.020000 254.495000   6.280000 ;
      RECT 254.325000   7.150000 254.495000   8.840000 ;
      RECT 254.325000  36.195000 254.855000  36.845000 ;
      RECT 254.335000  29.785000 254.845000  30.115000 ;
      RECT 254.340000  41.580000 254.555000  41.635000 ;
      RECT 254.340000  42.305000 254.510000  43.405000 ;
      RECT 254.340000  43.405000 254.535000  44.415000 ;
      RECT 254.365000  45.170000 254.535000  48.085000 ;
      RECT 254.385000  38.180000 254.690000  40.890000 ;
      RECT 254.385000  40.890000 254.555000  41.580000 ;
      RECT 254.405000  30.115000 254.775000  36.195000 ;
      RECT 254.530000  82.220000 254.700000  83.300000 ;
      RECT 254.530000  83.300000 255.230000  83.470000 ;
      RECT 254.530000  83.470000 254.700000  84.930000 ;
      RECT 254.535000 200.085000 255.205000 200.255000 ;
      RECT 254.535000 216.235000 255.205000 216.405000 ;
      RECT 254.560000  73.405000 255.090000  73.575000 ;
      RECT 254.575000  23.360000 255.065000  24.795000 ;
      RECT 254.575000  24.795000 257.655000  25.310000 ;
      RECT 254.600000  69.125000 255.650000  69.295000 ;
      RECT 254.700000  78.070000 254.870000  81.810000 ;
      RECT 254.705000  42.400000 255.235000  42.570000 ;
      RECT 254.705000  42.570000 255.115000  44.585000 ;
      RECT 254.705000  44.585000 255.245000  44.740000 ;
      RECT 254.705000  45.375000 255.245000  45.665000 ;
      RECT 254.705000  45.665000 254.995000  48.085000 ;
      RECT 254.720000  11.600000 254.890000  13.590000 ;
      RECT 254.720000  13.590000 255.980000  13.850000 ;
      RECT 254.720000  13.850000 254.890000  17.345000 ;
      RECT 254.725000  42.030000 255.755000  42.200000 ;
      RECT 254.745000  37.335000 255.415000  37.505000 ;
      RECT 254.820000  85.150000 256.170000  85.320000 ;
      RECT 254.825000  41.290000 255.570000  41.460000 ;
      RECT 254.850000 224.125000 264.850000 226.460000 ;
      RECT 254.850000 229.425000 264.850000 232.185000 ;
      RECT 254.850000 235.150000 264.850000 237.910000 ;
      RECT 254.850000 240.875000 264.850000 243.210000 ;
      RECT 254.895000  41.460000 255.425000  41.530000 ;
      RECT 254.935000   3.200000 260.025000   3.370000 ;
      RECT 254.935000   3.660000 259.685000   3.830000 ;
      RECT 254.935000   4.120000 260.025000   4.290000 ;
      RECT 254.945000  30.410000 255.115000  36.045000 ;
      RECT 254.945000  44.740000 255.245000  45.375000 ;
      RECT 254.945000  77.700000 255.615000  77.870000 ;
      RECT 254.955000   2.680000 279.030000   2.850000 ;
      RECT 254.960000  74.760000 255.610000  74.930000 ;
      RECT 254.960000  74.930000 255.130000  75.770000 ;
      RECT 255.025000  49.955000 255.815000  54.705000 ;
      RECT 255.025000  55.285000 255.195000  60.365000 ;
      RECT 255.195000  48.105000 255.950000  48.275000 ;
      RECT 255.205000  81.030000 256.215000  81.545000 ;
      RECT 255.215000  29.785000 255.725000  30.115000 ;
      RECT 255.215000  36.195000 259.325000  36.525000 ;
      RECT 255.240000  26.165000 255.410000  26.835000 ;
      RECT 255.270000  11.600000 255.440000  13.420000 ;
      RECT 255.270000  14.330000 255.440000  17.040000 ;
      RECT 255.280000  73.405000 255.650000  73.575000 ;
      RECT 255.280000  73.575000 255.610000  74.760000 ;
      RECT 255.285000  30.115000 255.655000  36.195000 ;
      RECT 255.285000  43.405000 255.455000  44.415000 ;
      RECT 255.285000  49.045000 255.815000  49.595000 ;
      RECT 255.400000  38.010000 255.570000  41.290000 ;
      RECT 255.410000  82.140000 255.580000  84.930000 ;
      RECT 255.420000  46.335000 255.950000  46.505000 ;
      RECT 255.425000   4.990000 255.955000   5.160000 ;
      RECT 255.440000  44.630000 255.610000  45.300000 ;
      RECT 255.460000  21.085000 255.630000  24.200000 ;
      RECT 255.470000  27.175000 256.750000  28.305000 ;
      RECT 255.480000  42.510000 256.015000  43.085000 ;
      RECT 255.540000  11.100000 256.050000  11.430000 ;
      RECT 255.540000  17.510000 256.050000  17.840000 ;
      RECT 255.580000  78.070000 255.750000  80.780000 ;
      RECT 255.585000  41.635000 255.755000  42.030000 ;
      RECT 255.585000  42.200000 255.755000  42.305000 ;
      RECT 255.605000   5.160000 255.775000   8.160000 ;
      RECT 255.610000  11.430000 255.980000  13.590000 ;
      RECT 255.610000  13.850000 255.980000  17.510000 ;
      RECT 255.635000 200.495000 256.165000 215.995000 ;
      RECT 255.645000  54.705000 255.815000  60.365000 ;
      RECT 255.745000  43.405000 255.950000  44.415000 ;
      RECT 255.760000  83.300000 256.460000  83.470000 ;
      RECT 255.780000  44.415000 255.950000  46.335000 ;
      RECT 255.780000  46.505000 255.950000  48.105000 ;
      RECT 255.780000  74.000000 259.980000  74.540000 ;
      RECT 255.780000  74.540000 256.070000  76.420000 ;
      RECT 255.800000  19.960000 256.310000  24.415000 ;
      RECT 255.825000  30.285000 255.995000  31.350000 ;
      RECT 255.825000  31.520000 255.995000  31.895000 ;
      RECT 255.825000  32.515000 255.995000  35.725000 ;
      RECT 255.860000  25.730000 256.440000  26.865000 ;
      RECT 255.905000  70.200000 256.435000  70.370000 ;
      RECT 255.920000  77.480000 256.450000  78.010000 ;
      RECT 255.945000   6.510000 257.635000   6.680000 ;
      RECT 255.985000  49.595000 256.655000  60.535000 ;
      RECT 256.000000  69.485000 256.170000  70.200000 ;
      RECT 256.000000  70.370000 256.170000  73.215000 ;
      RECT 256.030000   9.010000 256.200000  10.760000 ;
      RECT 256.030000  10.760000 261.145000  10.930000 ;
      RECT 256.055000 106.360000 256.585000 106.530000 ;
      RECT 256.150000  11.725000 256.320000  17.345000 ;
      RECT 256.175000  61.675000 256.345000  62.725000 ;
      RECT 256.175000  62.955000 256.345000  63.285000 ;
      RECT 256.175000  63.905000 256.345000  64.235000 ;
      RECT 256.175000  64.405000 256.345000  67.115000 ;
      RECT 256.240000  74.760000 256.410000  75.160000 ;
      RECT 256.240000  75.160000 256.770000  75.330000 ;
      RECT 256.240000  75.330000 256.410000  75.770000 ;
      RECT 256.240000  76.070000 256.410000  77.300000 ;
      RECT 256.240000  78.010000 256.410000  80.820000 ;
      RECT 256.245000  37.870000 256.415000  44.425000 ;
      RECT 256.245000  45.065000 256.415000  48.465000 ;
      RECT 256.290000  82.220000 256.460000  83.300000 ;
      RECT 256.290000  83.470000 256.460000  84.930000 ;
      RECT 256.295000 180.935000 265.595000 181.375000 ;
      RECT 256.295000 181.885000 265.595000 182.325000 ;
      RECT 256.295000 185.565000 265.595000 186.005000 ;
      RECT 256.295000 186.515000 265.595000 186.955000 ;
      RECT 256.335000 105.400000 256.505000 106.360000 ;
      RECT 256.335000 106.530000 256.505000 106.750000 ;
      RECT 256.410000  17.700000 256.940000  17.870000 ;
      RECT 256.420000  11.100000 256.930000  11.430000 ;
      RECT 256.420000  17.510000 256.930000  17.700000 ;
      RECT 256.445000  61.175000 256.955000  61.505000 ;
      RECT 256.445000  67.585000 256.955000  67.915000 ;
      RECT 256.465000  81.330000 257.135000  81.500000 ;
      RECT 256.490000  11.430000 256.860000  17.510000 ;
      RECT 256.515000  61.505000 256.885000  67.585000 ;
      RECT 256.535000  21.225000 257.080000  21.395000 ;
      RECT 256.595000 200.085000 257.265000 200.255000 ;
      RECT 256.595000 216.235000 257.265000 216.405000 ;
      RECT 256.605000  68.810000 257.855000  69.700000 ;
      RECT 256.605000  69.700000 257.795000  73.365000 ;
      RECT 256.630000 106.870000 261.815000 106.920000 ;
      RECT 256.645000  42.510000 257.180000  43.085000 ;
      RECT 256.700000  89.690000 267.165000  89.870000 ;
      RECT 256.700000 105.210000 261.450000 105.280000 ;
      RECT 256.700000 105.990000 261.450000 106.160000 ;
      RECT 256.705000  33.015000 256.875000  35.725000 ;
      RECT 256.710000  43.405000 256.915000  44.415000 ;
      RECT 256.710000  44.415000 256.880000  46.335000 ;
      RECT 256.710000  46.335000 257.240000  46.505000 ;
      RECT 256.710000  46.505000 256.880000  48.105000 ;
      RECT 256.710000  48.105000 257.465000  48.275000 ;
      RECT 256.780000  81.950000 256.950000  84.850000 ;
      RECT 256.800000  26.165000 256.970000  26.835000 ;
      RECT 256.825000  49.985000 256.995000  60.365000 ;
      RECT 256.885000   5.020000 257.055000   6.280000 ;
      RECT 256.885000   7.080000 257.055000   9.790000 ;
      RECT 256.905000  41.635000 257.075000  42.030000 ;
      RECT 256.905000  42.030000 257.935000  42.200000 ;
      RECT 256.905000  42.200000 257.075000  42.305000 ;
      RECT 257.030000  11.600000 257.200000  13.210000 ;
      RECT 257.030000  13.830000 257.200000  14.160000 ;
      RECT 257.030000  14.330000 257.200000  17.040000 ;
      RECT 257.050000  44.630000 257.220000  45.300000 ;
      RECT 257.055000  61.675000 257.225000  67.420000 ;
      RECT 257.070000  85.760000 257.240000  85.770000 ;
      RECT 257.070000  85.770000 257.720000  86.780000 ;
      RECT 257.090000  37.840000 261.330000  38.010000 ;
      RECT 257.090000  38.010000 257.260000  41.290000 ;
      RECT 257.090000  41.290000 257.835000  41.460000 ;
      RECT 257.120000  18.210000 258.010000  18.300000 ;
      RECT 257.120000  75.990000 257.650000  76.160000 ;
      RECT 257.120000  76.160000 257.290000  80.820000 ;
      RECT 257.175000  49.985000 257.615000  60.365000 ;
      RECT 257.205000  43.405000 257.375000  44.415000 ;
      RECT 257.225000  25.310000 257.655000  25.360000 ;
      RECT 257.225000  25.360000 257.765000  28.030000 ;
      RECT 257.225000  28.030000 257.755000  28.200000 ;
      RECT 257.235000  41.460000 257.765000  41.530000 ;
      RECT 257.245000  37.335000 257.915000  37.505000 ;
      RECT 257.270000  82.220000 257.440000  83.290000 ;
      RECT 257.270000  83.290000 257.880000  83.460000 ;
      RECT 257.270000  83.460000 257.440000  84.930000 ;
      RECT 257.300000  11.100000 257.810000  11.430000 ;
      RECT 257.300000  17.510000 257.810000  17.840000 ;
      RECT 257.300000  21.330000 257.595000  22.705000 ;
      RECT 257.305000  18.940000 257.595000  21.330000 ;
      RECT 257.330000  74.790000 257.860000  74.960000 ;
      RECT 257.370000  11.430000 257.740000  17.510000 ;
      RECT 257.375000  22.705000 257.545000  24.320000 ;
      RECT 257.380000   9.215000 257.910000  10.590000 ;
      RECT 257.415000  44.585000 257.955000  44.740000 ;
      RECT 257.415000  44.740000 257.715000  45.375000 ;
      RECT 257.415000  45.375000 257.955000  45.665000 ;
      RECT 257.425000  42.400000 257.955000  42.570000 ;
      RECT 257.520000  74.760000 257.690000  74.790000 ;
      RECT 257.520000  74.960000 257.690000  75.770000 ;
      RECT 257.530000  81.190000 258.115000  81.335000 ;
      RECT 257.530000  81.335000 258.540000  81.505000 ;
      RECT 257.545000  42.570000 257.955000  44.585000 ;
      RECT 257.550000 113.195000 258.220000 113.525000 ;
      RECT 257.585000  30.285000 257.755000  31.335000 ;
      RECT 257.585000  33.015000 257.755000  35.725000 ;
      RECT 257.585000  81.020000 258.115000  81.190000 ;
      RECT 257.605000  61.675000 257.775000  63.495000 ;
      RECT 257.605000  64.405000 257.775000  67.115000 ;
      RECT 257.610000  76.420000 261.010000  76.590000 ;
      RECT 257.610000  77.200000 260.320000  77.370000 ;
      RECT 257.625000  49.045000 258.295000  49.765000 ;
      RECT 257.625000  60.555000 258.295000  60.615000 ;
      RECT 257.625000  60.615000 259.685000  60.785000 ;
      RECT 257.665000  45.665000 257.955000  48.085000 ;
      RECT 257.665000  85.150000 258.675000  85.320000 ;
      RECT 257.675000 113.910000 260.675000 164.900000 ;
      RECT 257.695000 200.495000 258.225000 215.995000 ;
      RECT 257.710000  29.785000 259.240000  30.115000 ;
      RECT 257.735000  78.070000 257.905000  80.780000 ;
      RECT 257.800000  19.625000 258.480000  19.795000 ;
      RECT 257.800000  19.795000 258.415000  21.225000 ;
      RECT 257.800000  21.225000 258.475000  21.395000 ;
      RECT 257.860000  77.680000 258.530000  77.850000 ;
      RECT 257.875000  24.955000 258.805000  25.215000 ;
      RECT 257.875000  49.985000 258.045000  54.895000 ;
      RECT 257.875000  55.455000 258.045000  60.365000 ;
      RECT 257.875000  61.175000 258.385000  61.505000 ;
      RECT 257.875000  67.585000 258.385000  67.915000 ;
      RECT 257.885000  45.000000 258.415000  45.170000 ;
      RECT 257.910000  11.725000 258.080000  17.345000 ;
      RECT 257.910000  76.370000 260.240000  76.420000 ;
      RECT 257.910000  77.080000 260.240000  77.200000 ;
      RECT 257.925000  30.115000 258.295000  36.195000 ;
      RECT 257.945000  61.505000 258.315000  67.585000 ;
      RECT 257.945000  87.005000 261.715000  87.175000 ;
      RECT 257.970000  38.180000 258.275000  40.890000 ;
      RECT 257.970000  87.000000 261.700000  87.005000 ;
      RECT 257.985000   6.510000 258.515000   6.680000 ;
      RECT 258.050000  82.140000 258.220000  84.930000 ;
      RECT 258.100000  26.090000 258.270000  26.780000 ;
      RECT 258.100000  26.780000 258.740000  27.040000 ;
      RECT 258.100000  27.040000 258.270000  27.100000 ;
      RECT 258.105000  40.890000 258.275000  41.580000 ;
      RECT 258.105000  41.580000 258.320000  41.635000 ;
      RECT 258.105000  41.635000 258.355000  42.305000 ;
      RECT 258.125000  43.405000 258.320000  44.415000 ;
      RECT 258.125000  45.170000 258.295000  48.085000 ;
      RECT 258.150000  42.305000 258.320000  43.405000 ;
      RECT 258.165000   5.020000 258.335000   6.510000 ;
      RECT 258.165000   6.680000 258.335000   9.790000 ;
      RECT 258.180000  11.100000 258.690000  11.430000 ;
      RECT 258.180000  17.510000 258.690000  17.515000 ;
      RECT 258.180000  17.515000 259.440000  17.840000 ;
      RECT 258.195000  37.335000 258.865000  37.505000 ;
      RECT 258.250000  11.430000 258.620000  17.510000 ;
      RECT 258.305000  49.985000 265.915000  50.345000 ;
      RECT 258.305000  50.345000 260.870000  50.995000 ;
      RECT 258.305000  50.995000 259.055000  60.365000 ;
      RECT 258.325000  27.350000 262.765000  27.520000 ;
      RECT 258.445000  41.290000 259.115000  41.460000 ;
      RECT 258.465000  30.285000 258.635000  35.725000 ;
      RECT 258.485000  61.800000 258.655000  67.420000 ;
      RECT 258.515000  71.440000 259.405000  72.330000 ;
      RECT 258.525000  41.460000 259.020000  42.030000 ;
      RECT 258.525000  42.030000 259.055000  42.200000 ;
      RECT 258.535000   6.880000 259.065000   7.050000 ;
      RECT 258.545000  25.215000 258.805000  26.145000 ;
      RECT 258.545000  26.145000 259.685000  26.405000 ;
      RECT 258.555000  68.460000 259.405000  71.440000 ;
      RECT 258.555000  72.330000 259.405000  72.450000 ;
      RECT 258.555000  72.450000 260.395000  73.365000 ;
      RECT 258.585000  43.405000 259.235000  44.415000 ;
      RECT 258.585000  44.415000 258.755000  46.335000 ;
      RECT 258.585000  46.335000 259.115000  46.505000 ;
      RECT 258.585000  46.505000 258.755000  48.085000 ;
      RECT 258.615000  78.070000 258.785000  80.950000 ;
      RECT 258.615000  80.950000 259.780000  81.120000 ;
      RECT 258.650000  19.745000 258.910000  20.385000 ;
      RECT 258.650000  83.290000 259.180000  83.460000 ;
      RECT 258.655000  21.610000 258.825000  24.645000 ;
      RECT 258.655000 200.085000 259.325000 200.255000 ;
      RECT 258.655000 216.235000 259.325000 216.405000 ;
      RECT 258.665000  18.945000 258.865000  19.745000 ;
      RECT 258.695000  20.385000 258.865000  21.025000 ;
      RECT 258.715000   5.020000 258.885000   6.880000 ;
      RECT 258.715000   7.050000 258.885000   9.790000 ;
      RECT 258.755000  61.175000 259.265000  61.505000 ;
      RECT 258.755000  67.585000 259.265000  67.915000 ;
      RECT 258.790000  11.600000 258.960000  13.420000 ;
      RECT 258.790000  14.330000 258.960000  17.040000 ;
      RECT 258.800000  74.760000 258.970000  75.180000 ;
      RECT 258.800000  75.180000 259.340000  75.350000 ;
      RECT 258.800000  75.350000 258.970000  75.770000 ;
      RECT 258.805000  30.115000 259.175000  36.195000 ;
      RECT 258.825000  61.505000 259.195000  67.585000 ;
      RECT 258.830000  82.220000 259.000000  83.290000 ;
      RECT 258.830000  83.460000 259.000000  84.930000 ;
      RECT 258.850000  38.180000 259.020000  41.290000 ;
      RECT 258.860000  77.680000 259.530000  77.850000 ;
      RECT 258.885000  49.805000 265.335000  49.985000 ;
      RECT 258.885000  60.365000 259.055000  60.445000 ;
      RECT 258.925000  47.855000 259.095000  48.465000 ;
      RECT 259.035000  17.840000 259.440000  18.875000 ;
      RECT 259.035000  18.875000 259.565000  19.045000 ;
      RECT 259.065000  42.475000 261.725000  42.645000 ;
      RECT 259.065000  42.645000 259.235000  43.405000 ;
      RECT 259.075000   6.510000 261.105000   6.680000 ;
      RECT 259.075000  37.335000 261.105000  37.505000 ;
      RECT 259.130000  85.150000 260.140000  85.320000 ;
      RECT 259.150000  10.390000 259.680000  10.560000 ;
      RECT 259.160000  10.260000 259.670000  10.390000 ;
      RECT 259.160000  10.560000 259.670000  10.590000 ;
      RECT 259.250000  25.130000 259.455000  25.570000 ;
      RECT 259.250000  25.570000 265.515000  25.740000 ;
      RECT 259.275000  52.630000 259.805000  52.800000 ;
      RECT 259.280000  26.090000 259.450000  26.145000 ;
      RECT 259.280000  26.405000 259.450000  27.100000 ;
      RECT 259.285000  19.350000 285.170000  19.520000 ;
      RECT 259.285000  19.520000 259.455000  20.525000 ;
      RECT 259.285000  24.090000 259.455000  25.130000 ;
      RECT 259.285000  25.740000 263.930000  25.815000 ;
      RECT 259.285000  41.360000 259.815000  41.530000 ;
      RECT 259.295000  51.955000 259.685000  52.630000 ;
      RECT 259.295000  52.800000 259.685000  54.985000 ;
      RECT 259.295000  54.985000 259.805000  55.315000 ;
      RECT 259.320000  51.235000 259.990000  51.785000 ;
      RECT 259.340000  11.600000 259.510000  17.345000 ;
      RECT 259.345000  30.285000 259.515000  31.335000 ;
      RECT 259.345000  33.015000 259.515000  35.725000 ;
      RECT 259.365000  61.675000 259.535000  62.740000 ;
      RECT 259.365000  62.910000 259.535000  63.285000 ;
      RECT 259.365000  63.905000 259.535000  64.235000 ;
      RECT 259.365000  64.405000 259.535000  67.115000 ;
      RECT 259.405000  43.095000 259.935000  43.265000 ;
      RECT 259.405000  43.265000 259.575000  48.390000 ;
      RECT 259.440000  84.280000 259.970000  84.450000 ;
      RECT 259.465000  41.530000 259.635000  42.305000 ;
      RECT 259.495000  78.070000 259.665000  80.780000 ;
      RECT 259.515000  55.785000 259.685000  60.615000 ;
      RECT 259.605000  32.140000 260.135000  32.310000 ;
      RECT 259.610000  11.100000 260.120000  11.430000 ;
      RECT 259.610000  17.510000 260.120000  17.840000 ;
      RECT 259.610000  81.120000 259.780000  84.280000 ;
      RECT 259.610000  84.450000 259.780000  84.930000 ;
      RECT 259.660000  74.790000 260.250000  74.960000 ;
      RECT 259.680000  11.430000 260.050000  17.510000 ;
      RECT 259.705000  61.175000 260.215000  61.505000 ;
      RECT 259.705000  67.585000 260.215000  67.915000 ;
      RECT 259.730000  18.040000 260.870000  18.210000 ;
      RECT 259.730000  38.180000 259.990000  41.160000 ;
      RECT 259.745000  44.180000 261.565000  44.350000 ;
      RECT 259.745000  44.350000 259.935000  47.370000 ;
      RECT 259.745000  47.370000 260.275000  48.550000 ;
      RECT 259.745000  48.550000 262.635000  48.720000 ;
      RECT 259.755000 200.495000 260.285000 215.995000 ;
      RECT 259.775000  61.505000 260.145000  67.585000 ;
      RECT 259.805000  18.210000 260.695000  18.270000 ;
      RECT 259.855000   3.370000 260.025000   4.120000 ;
      RECT 259.855000  59.125000 264.365000  60.315000 ;
      RECT 259.865000  19.870000 260.035000  24.620000 ;
      RECT 259.950000  81.335000 260.620000  81.570000 ;
      RECT 259.950000  83.290000 260.560000  83.460000 ;
      RECT 259.965000  30.285000 260.135000  32.140000 ;
      RECT 259.965000  32.310000 260.135000  36.030000 ;
      RECT 259.975000  51.955000 260.145000  58.495000 ;
      RECT 259.995000   5.020000 260.165000   6.280000 ;
      RECT 259.995000   7.080000 260.165000   9.790000 ;
      RECT 260.080000  74.760000 260.250000  74.790000 ;
      RECT 260.080000  74.960000 260.250000  75.770000 ;
      RECT 260.090000  25.130000 263.995000  25.300000 ;
      RECT 260.090000  59.115000 264.220000  59.125000 ;
      RECT 260.105000  42.840000 260.275000  44.010000 ;
      RECT 260.105000  44.580000 260.275000  45.280000 ;
      RECT 260.105000  45.280000 260.635000  45.450000 ;
      RECT 260.105000  45.450000 260.275000  47.080000 ;
      RECT 260.105000  68.620000 260.275000  71.130000 ;
      RECT 260.110000 113.195000 260.780000 113.525000 ;
      RECT 260.145000  78.090000 260.695000  81.090000 ;
      RECT 260.190000  38.180000 260.450000  41.160000 ;
      RECT 260.195000   3.430000 260.365000   4.430000 ;
      RECT 260.200000  51.235000 260.870000  51.405000 ;
      RECT 260.200000  58.715000 261.550000  58.885000 ;
      RECT 260.220000  11.600000 260.390000  13.210000 ;
      RECT 260.220000  13.830000 260.390000  14.160000 ;
      RECT 260.220000  14.330000 260.390000  17.040000 ;
      RECT 260.225000  26.780000 260.865000  27.040000 ;
      RECT 260.235000  29.785000 260.745000  30.115000 ;
      RECT 260.235000  36.195000 260.745000  36.525000 ;
      RECT 260.305000  30.115000 260.675000  36.195000 ;
      RECT 260.315000  51.405000 260.585000  58.715000 ;
      RECT 260.315000  61.675000 260.485000  66.145000 ;
      RECT 260.375000  42.470000 261.725000  42.475000 ;
      RECT 260.390000  82.220000 260.560000  83.290000 ;
      RECT 260.390000  83.460000 260.560000  84.930000 ;
      RECT 260.440000  71.350000 264.170000  71.520000 ;
      RECT 260.445000  68.385000 264.255000  68.400000 ;
      RECT 260.445000  68.400000 264.215000  68.555000 ;
      RECT 260.445000  70.985000 264.170000  71.350000 ;
      RECT 260.460000  26.090000 260.630000  26.780000 ;
      RECT 260.460000  27.040000 260.630000  27.100000 ;
      RECT 260.485000  68.230000 264.255000  68.385000 ;
      RECT 260.535000   3.200000 265.625000   3.370000 ;
      RECT 260.535000   3.370000 260.705000   4.120000 ;
      RECT 260.535000   4.120000 265.625000   4.290000 ;
      RECT 260.535000  42.840000 260.705000  44.180000 ;
      RECT 260.585000  46.335000 261.115000  47.370000 ;
      RECT 260.585000  47.370000 261.455000  48.380000 ;
      RECT 260.585000  61.175000 261.095000  61.505000 ;
      RECT 260.585000  67.585000 261.095000  67.915000 ;
      RECT 260.645000  19.870000 260.815000  24.620000 ;
      RECT 260.655000  61.505000 261.025000  67.585000 ;
      RECT 260.715000 200.085000 261.385000 200.255000 ;
      RECT 260.715000 216.235000 261.385000 216.405000 ;
      RECT 260.755000  51.765000 261.210000  51.935000 ;
      RECT 260.755000  51.935000 260.925000  58.495000 ;
      RECT 260.770000  11.600000 260.940000  13.420000 ;
      RECT 260.770000  14.330000 260.940000  17.040000 ;
      RECT 260.840000  76.590000 261.010000  77.155000 ;
      RECT 260.845000  30.285000 261.015000  31.335000 ;
      RECT 260.845000  31.565000 261.015000  31.895000 ;
      RECT 260.845000  32.515000 261.015000  32.845000 ;
      RECT 260.845000  33.015000 261.015000  35.725000 ;
      RECT 260.875000   3.660000 266.075000   3.830000 ;
      RECT 260.920000  32.140000 261.555000  32.310000 ;
      RECT 260.965000  42.840000 261.135000  44.010000 ;
      RECT 260.975000   8.840000 264.430000   9.010000 ;
      RECT 260.975000   9.010000 261.145000  10.760000 ;
      RECT 261.040000  11.100000 261.550000  11.430000 ;
      RECT 261.040000  17.510000 261.550000  18.465000 ;
      RECT 261.040000  18.465000 261.575000  18.635000 ;
      RECT 261.040000  50.515000 261.210000  51.765000 ;
      RECT 261.050000  71.775000 261.220000  74.940000 ;
      RECT 261.095000  52.210000 261.365000  58.715000 ;
      RECT 261.110000  11.430000 261.480000  17.510000 ;
      RECT 261.110000  26.145000 261.810000  26.405000 ;
      RECT 261.115000  29.785000 264.265000  30.115000 ;
      RECT 261.115000  36.195000 261.625000  36.220000 ;
      RECT 261.115000  36.220000 264.265000  36.525000 ;
      RECT 261.140000  81.950000 261.310000  84.850000 ;
      RECT 261.160000  38.010000 261.330000  41.360000 ;
      RECT 261.160000  41.360000 261.690000  41.530000 ;
      RECT 261.170000  78.070000 261.340000  79.055000 ;
      RECT 261.170000  79.055000 261.870000  79.225000 ;
      RECT 261.170000  79.225000 261.340000  80.780000 ;
      RECT 261.185000  30.115000 261.555000  32.140000 ;
      RECT 261.185000  32.310000 261.555000  36.195000 ;
      RECT 261.265000  61.675000 261.985000  62.725000 ;
      RECT 261.265000  62.955000 261.985000  63.285000 ;
      RECT 261.265000  63.905000 261.985000  64.235000 ;
      RECT 261.265000  64.405000 261.435000  67.420000 ;
      RECT 261.275000   5.020000 261.445000   8.160000 ;
      RECT 261.285000  44.580000 261.455000  45.760000 ;
      RECT 261.285000  45.760000 263.815000  45.930000 ;
      RECT 261.285000  45.930000 261.455000  47.080000 ;
      RECT 261.380000  50.345000 262.840000  50.995000 ;
      RECT 261.395000  42.840000 261.565000  44.180000 ;
      RECT 261.425000  19.870000 261.595000  24.620000 ;
      RECT 261.460000  77.680000 262.810000  77.850000 ;
      RECT 261.460000  81.335000 262.810000  81.805000 ;
      RECT 261.490000  81.805000 262.810000  81.940000 ;
      RECT 261.535000  51.955000 261.705000  58.495000 ;
      RECT 261.630000  72.250000 261.800000  74.000000 ;
      RECT 261.630000  74.000000 262.160000  74.170000 ;
      RECT 261.630000  74.170000 261.800000  75.880000 ;
      RECT 261.630000  75.880000 264.155000  76.050000 ;
      RECT 261.630000  76.220000 261.800000  77.360000 ;
      RECT 261.630000  82.220000 261.800000  84.070000 ;
      RECT 261.630000  84.070000 262.160000  84.240000 ;
      RECT 261.630000  84.240000 261.800000  84.930000 ;
      RECT 261.640000  26.090000 261.810000  26.145000 ;
      RECT 261.640000  26.405000 261.810000  27.100000 ;
      RECT 261.650000  11.725000 261.820000  17.345000 ;
      RECT 261.660000 106.360000 262.190000 106.530000 ;
      RECT 261.720000  18.040000 275.225000  18.210000 ;
      RECT 261.725000  30.285000 261.895000  36.030000 ;
      RECT 261.740000  37.870000 261.910000  40.870000 ;
      RECT 261.805000  46.165000 262.135000  47.015000 ;
      RECT 261.815000  64.405000 261.985000  67.420000 ;
      RECT 261.815000 200.495000 262.345000 215.995000 ;
      RECT 261.825000  42.840000 261.995000  44.010000 ;
      RECT 261.830000  85.770000 262.000000  86.780000 ;
      RECT 261.885000  47.015000 262.055000  47.625000 ;
      RECT 261.910000  17.700000 262.440000  17.870000 ;
      RECT 261.920000  11.100000 262.430000  11.430000 ;
      RECT 261.920000  17.510000 262.430000  17.700000 ;
      RECT 261.940000 105.400000 262.110000 106.360000 ;
      RECT 261.940000 106.530000 262.110000 106.750000 ;
      RECT 261.960000  45.280000 262.635000  45.450000 ;
      RECT 261.970000  75.160000 262.500000  75.330000 ;
      RECT 261.990000  11.430000 262.360000  17.510000 ;
      RECT 261.995000  36.195000 263.385000  36.220000 ;
      RECT 262.025000  51.665000 262.195000  58.425000 ;
      RECT 262.040000  26.315000 262.570000  27.350000 ;
      RECT 262.045000  85.150000 263.735000  85.320000 ;
      RECT 262.050000  78.070000 262.220000  80.950000 ;
      RECT 262.050000  80.950000 263.360000  81.165000 ;
      RECT 262.060000  75.330000 262.390000  75.690000 ;
      RECT 262.065000  30.115000 262.435000  36.195000 ;
      RECT 262.080000  42.470000 263.430000  42.640000 ;
      RECT 262.080000  42.640000 263.330000  42.670000 ;
      RECT 262.140000  67.885000 263.545000  67.915000 ;
      RECT 262.140000  67.915000 262.670000  68.055000 ;
      RECT 262.155000  61.175000 262.665000  61.505000 ;
      RECT 262.155000  67.585000 263.545000  67.885000 ;
      RECT 262.165000  87.000000 265.895000  87.005000 ;
      RECT 262.165000  87.005000 265.935000  87.175000 ;
      RECT 262.185000 113.910000 265.185000 164.900000 ;
      RECT 262.205000  19.870000 262.375000  24.620000 ;
      RECT 262.225000  61.505000 262.595000  67.585000 ;
      RECT 262.235000 106.870000 267.055000 106.920000 ;
      RECT 262.255000  42.840000 262.425000  44.180000 ;
      RECT 262.255000  44.180000 263.815000  44.350000 ;
      RECT 262.305000 105.210000 267.055000 105.280000 ;
      RECT 262.305000 105.990000 267.055000 106.160000 ;
      RECT 262.410000  82.200000 262.580000  84.930000 ;
      RECT 262.465000  44.580000 262.635000  45.280000 ;
      RECT 262.465000  45.450000 262.635000  45.590000 ;
      RECT 262.465000  46.100000 262.635000  48.550000 ;
      RECT 262.515000  51.955000 262.685000  58.495000 ;
      RECT 262.530000  11.600000 262.700000  13.210000 ;
      RECT 262.530000  13.830000 262.700000  14.160000 ;
      RECT 262.530000  14.330000 262.700000  17.040000 ;
      RECT 262.555000   5.020000 262.725000   6.280000 ;
      RECT 262.555000   7.150000 262.725000   8.840000 ;
      RECT 262.580000  76.050000 262.750000  77.230000 ;
      RECT 262.605000  30.285000 262.775000  31.335000 ;
      RECT 262.605000  31.565000 262.775000  31.895000 ;
      RECT 262.605000  32.515000 262.775000  32.845000 ;
      RECT 262.605000  33.015000 262.775000  35.725000 ;
      RECT 262.670000  58.715000 264.020000  58.885000 ;
      RECT 262.685000  42.840000 262.855000  44.010000 ;
      RECT 262.760000  79.055000 263.290000  79.225000 ;
      RECT 262.765000  61.675000 262.935000  66.145000 ;
      RECT 262.775000 200.085000 263.445000 200.255000 ;
      RECT 262.775000 216.235000 263.445000 216.405000 ;
      RECT 262.795000  18.210000 267.285000  18.265000 ;
      RECT 262.800000  11.100000 263.310000  11.430000 ;
      RECT 262.800000  17.510000 263.310000  17.840000 ;
      RECT 262.820000  26.090000 262.990000  26.780000 ;
      RECT 262.820000  26.780000 263.475000  27.040000 ;
      RECT 262.820000  27.040000 262.990000  27.100000 ;
      RECT 262.835000  75.160000 263.365000  75.330000 ;
      RECT 262.855000  52.210000 263.125000  58.715000 ;
      RECT 262.870000  11.430000 263.240000  17.510000 ;
      RECT 262.930000  78.070000 263.100000  79.055000 ;
      RECT 262.930000  79.225000 263.100000  80.780000 ;
      RECT 262.940000  75.330000 263.270000  75.690000 ;
      RECT 262.945000  30.115000 263.315000  36.195000 ;
      RECT 262.960000  84.070000 263.490000  84.240000 ;
      RECT 263.010000  50.515000 263.180000  51.765000 ;
      RECT 263.010000  51.765000 263.465000  51.935000 ;
      RECT 263.035000  61.175000 263.545000  61.505000 ;
      RECT 263.045000  27.350000 263.945000  27.520000 ;
      RECT 263.085000  37.765000 263.255000  40.845000 ;
      RECT 263.105000  61.505000 263.475000  67.585000 ;
      RECT 263.115000  42.840000 263.285000  44.180000 ;
      RECT 263.190000  81.165000 263.360000  84.070000 ;
      RECT 263.190000  84.240000 263.360000  84.930000 ;
      RECT 263.205000 190.925000 267.915000 191.195000 ;
      RECT 263.220000  77.680000 264.570000  77.850000 ;
      RECT 263.285000  46.335000 263.815000  46.505000 ;
      RECT 263.295000  51.935000 263.465000  58.495000 ;
      RECT 263.350000  50.345000 265.915000  50.995000 ;
      RECT 263.350000  51.235000 264.020000  51.405000 ;
      RECT 263.410000  11.600000 263.580000  13.590000 ;
      RECT 263.410000  13.590000 264.670000  13.850000 ;
      RECT 263.410000  13.850000 263.580000  17.345000 ;
      RECT 263.410000  41.265000 264.375000  41.435000 ;
      RECT 263.410000  41.435000 263.720000  42.130000 ;
      RECT 263.410000  42.130000 263.940000  42.300000 ;
      RECT 263.485000  19.870000 263.655000  24.620000 ;
      RECT 263.485000  30.285000 263.655000  36.030000 ;
      RECT 263.530000  11.260000 264.060000  11.430000 ;
      RECT 263.530000  71.775000 263.700000  74.960000 ;
      RECT 263.530000  76.220000 263.700000  77.360000 ;
      RECT 263.545000  42.840000 263.715000  44.010000 ;
      RECT 263.550000  38.155000 263.835000  40.865000 ;
      RECT 263.550000  40.865000 263.720000  41.095000 ;
      RECT 263.625000  68.725000 264.555000  69.905000 ;
      RECT 263.625000  69.905000 264.155000  70.075000 ;
      RECT 263.635000  51.405000 263.905000  58.715000 ;
      RECT 263.645000  44.350000 263.815000  45.760000 ;
      RECT 263.645000  46.100000 263.815000  46.335000 ;
      RECT 263.645000  46.505000 263.815000  48.380000 ;
      RECT 263.655000   7.365000 264.185000   7.535000 ;
      RECT 263.715000  61.675000 263.885000  62.725000 ;
      RECT 263.715000  62.955000 263.885000  63.285000 ;
      RECT 263.715000  63.905000 263.885000  64.235000 ;
      RECT 263.715000  64.405000 263.885000  67.115000 ;
      RECT 263.755000  36.195000 264.265000  36.220000 ;
      RECT 263.810000  78.070000 263.980000  80.780000 ;
      RECT 263.825000  30.115000 264.195000  36.195000 ;
      RECT 263.825000  75.180000 264.155000  75.880000 ;
      RECT 263.835000   5.020000 264.005000   7.365000 ;
      RECT 263.835000   7.535000 264.005000   8.160000 ;
      RECT 263.875000 200.495000 264.405000 215.995000 ;
      RECT 263.890000  11.430000 264.060000  11.600000 ;
      RECT 263.890000  11.600000 264.130000  13.420000 ;
      RECT 263.890000  37.335000 266.145000  37.505000 ;
      RECT 263.890000  41.085000 264.560000  41.255000 ;
      RECT 263.890000  41.255000 264.375000  41.265000 ;
      RECT 263.890000  41.760000 264.420000  41.930000 ;
      RECT 263.960000  14.330000 264.130000  17.040000 ;
      RECT 263.970000  82.200000 264.140000  84.930000 ;
      RECT 263.985000  21.120000 264.515000  21.220000 ;
      RECT 263.985000  21.220000 264.530000  23.410000 ;
      RECT 263.985000  61.175000 264.495000  61.505000 ;
      RECT 263.985000  67.585000 264.495000  67.915000 ;
      RECT 264.000000  26.060000 264.530000  27.100000 ;
      RECT 264.005000  37.505000 266.145000  37.595000 ;
      RECT 264.005000  37.595000 264.375000  41.085000 ;
      RECT 264.005000  43.110000 264.535000  48.390000 ;
      RECT 264.055000  61.505000 264.425000  67.585000 ;
      RECT 264.075000  51.955000 264.245000  58.495000 ;
      RECT 264.110000  41.930000 264.420000  43.110000 ;
      RECT 264.160000  79.055000 264.860000  79.225000 ;
      RECT 264.175000   6.510000 265.865000   6.680000 ;
      RECT 264.215000  81.320000 264.885000  81.340000 ;
      RECT 264.215000  81.340000 265.165000  81.490000 ;
      RECT 264.230000  11.100000 264.740000  11.430000 ;
      RECT 264.230000  17.510000 264.740000  17.840000 ;
      RECT 264.230000  51.235000 264.900000  51.785000 ;
      RECT 264.260000   9.010000 264.430000  10.760000 ;
      RECT 264.260000  10.760000 275.555000  10.930000 ;
      RECT 264.275000  81.490000 265.165000  81.510000 ;
      RECT 264.300000  11.430000 264.670000  13.590000 ;
      RECT 264.300000  13.850000 264.670000  17.510000 ;
      RECT 264.365000  30.285000 264.535000  31.335000 ;
      RECT 264.365000  31.565000 264.535000  31.895000 ;
      RECT 264.365000  32.515000 264.535000  32.845000 ;
      RECT 264.365000  33.015000 264.535000  35.725000 ;
      RECT 264.385000  68.620000 264.555000  68.725000 ;
      RECT 264.385000  70.120000 264.555000  71.945000 ;
      RECT 264.390000  84.070000 264.920000  84.240000 ;
      RECT 264.405000  75.570000 264.935000  75.740000 ;
      RECT 264.415000  52.630000 264.945000  52.800000 ;
      RECT 264.415000  54.985000 264.925000  55.315000 ;
      RECT 264.475000  91.720000 290.580000  92.265000 ;
      RECT 264.480000  72.250000 264.650000  75.570000 ;
      RECT 264.480000  75.740000 264.650000  77.230000 ;
      RECT 264.535000  51.955000 264.925000  52.630000 ;
      RECT 264.535000  52.800000 264.925000  54.985000 ;
      RECT 264.535000  55.785000 264.705000  60.615000 ;
      RECT 264.535000  60.615000 266.595000  60.785000 ;
      RECT 264.545000  37.765000 264.715000  40.865000 ;
      RECT 264.590000  41.445000 265.055000  41.615000 ;
      RECT 264.590000  41.615000 264.760000  42.520000 ;
      RECT 264.590000  42.520000 264.875000  42.690000 ;
      RECT 264.595000  61.675000 264.765000  67.415000 ;
      RECT 264.615000  32.140000 265.145000  32.310000 ;
      RECT 264.690000  78.070000 264.860000  79.055000 ;
      RECT 264.690000  79.225000 264.860000  80.780000 ;
      RECT 264.705000  29.785000 265.215000  30.115000 ;
      RECT 264.705000  36.195000 265.215000  36.525000 ;
      RECT 264.705000  42.690000 264.875000  43.615000 ;
      RECT 264.750000  82.220000 264.920000  84.070000 ;
      RECT 264.750000  84.240000 264.920000  84.930000 ;
      RECT 264.760000  25.740000 265.140000  25.815000 ;
      RECT 264.765000  19.870000 264.935000  24.620000 ;
      RECT 264.775000  30.115000 265.145000  32.140000 ;
      RECT 264.775000  32.310000 265.145000  36.195000 ;
      RECT 264.835000 200.085000 265.505000 200.255000 ;
      RECT 264.835000 216.235000 265.505000 216.405000 ;
      RECT 264.840000  11.725000 265.010000  17.345000 ;
      RECT 264.865000  61.175000 265.375000  61.505000 ;
      RECT 264.865000  67.585000 265.375000  67.915000 ;
      RECT 264.885000  40.395000 265.595000  40.865000 ;
      RECT 264.885000  40.865000 265.055000  41.445000 ;
      RECT 264.930000  41.785000 265.550000  42.115000 ;
      RECT 264.935000  61.505000 265.305000  67.585000 ;
      RECT 264.935000  68.620000 265.105000  70.305000 ;
      RECT 264.935000  70.305000 265.465000  70.475000 ;
      RECT 264.935000  70.475000 265.105000  71.330000 ;
      RECT 265.100000  11.260000 265.630000  11.430000 ;
      RECT 265.110000  11.100000 265.620000  11.260000 ;
      RECT 265.110000  17.510000 265.620000  17.840000 ;
      RECT 265.115000   5.020000 265.285000   6.280000 ;
      RECT 265.115000   7.080000 265.285000   9.790000 ;
      RECT 265.150000  68.230000 267.450000  68.400000 ;
      RECT 265.155000  48.350000 268.525000  48.520000 ;
      RECT 265.165000  50.995000 265.915000  60.365000 ;
      RECT 265.165000  60.365000 265.335000  60.445000 ;
      RECT 265.180000  11.430000 265.550000  17.510000 ;
      RECT 265.195000  45.290000 265.365000  48.000000 ;
      RECT 265.205000  88.075000 268.600000  88.360000 ;
      RECT 265.205000  88.360000 265.870000  89.285000 ;
      RECT 265.210000  72.490000 267.105000  74.940000 ;
      RECT 265.225000  41.360000 266.145000  41.530000 ;
      RECT 265.225000  41.530000 265.550000  41.785000 ;
      RECT 265.265000  71.415000 267.105000  72.490000 ;
      RECT 265.280000  78.130000 265.450000  81.050000 ;
      RECT 265.280000  81.950000 265.450000  84.850000 ;
      RECT 265.280000 223.695000 266.130000 225.350000 ;
      RECT 265.280000 229.255000 266.130000 232.355000 ;
      RECT 265.280000 240.705000 266.130000 243.640000 ;
      RECT 265.315000  30.285000 265.485000  34.755000 ;
      RECT 265.315000  48.215000 268.365000  48.350000 ;
      RECT 265.330000  25.740000 265.515000  26.920000 ;
      RECT 265.330000  26.920000 284.775000  27.090000 ;
      RECT 265.345000  23.560000 265.515000  25.570000 ;
      RECT 265.355000 190.145000 267.915000 190.415000 ;
      RECT 265.425000  38.155000 265.595000  40.395000 ;
      RECT 265.455000  70.675000 266.045000  70.845000 ;
      RECT 265.475000  61.675000 265.645000  62.725000 ;
      RECT 265.475000  62.955000 265.645000  63.285000 ;
      RECT 265.475000  63.905000 265.645000  64.235000 ;
      RECT 265.475000  64.405000 265.645000  67.115000 ;
      RECT 265.500000  35.110000 266.030000  35.280000 ;
      RECT 265.585000  29.785000 266.095000  30.115000 ;
      RECT 265.585000  36.195000 266.095000  36.525000 ;
      RECT 265.585000  42.605000 265.755000  44.400000 ;
      RECT 265.600000  45.030000 266.145000  45.200000 ;
      RECT 265.610000  10.390000 266.140000  10.560000 ;
      RECT 265.620000 225.650000 265.790000 226.630000 ;
      RECT 265.620000 234.980000 265.790000 235.960000 ;
      RECT 265.620000 237.100000 265.790000 238.080000 ;
      RECT 265.630000  10.260000 266.140000  10.390000 ;
      RECT 265.630000  10.560000 266.140000  10.590000 ;
      RECT 265.635000  68.400000 266.045000  70.675000 ;
      RECT 265.655000  30.115000 266.025000  35.110000 ;
      RECT 265.655000  35.280000 266.025000  36.195000 ;
      RECT 265.690000  44.570000 266.700000  44.740000 ;
      RECT 265.690000  44.740000 266.220000  44.800000 ;
      RECT 265.720000  11.600000 265.890000  13.210000 ;
      RECT 265.720000  13.830000 265.890000  14.160000 ;
      RECT 265.720000  14.330000 265.890000  17.040000 ;
      RECT 265.745000  61.175000 266.255000  61.505000 ;
      RECT 265.745000  67.585000 266.255000  67.915000 ;
      RECT 265.765000  37.595000 266.145000  38.615000 ;
      RECT 265.805000  42.000000 266.475000  42.170000 ;
      RECT 265.815000  61.505000 266.185000  67.585000 ;
      RECT 265.875000  42.170000 266.405000  42.300000 ;
      RECT 265.905000   3.200000 271.095000   3.370000 ;
      RECT 265.905000   3.370000 266.075000   3.660000 ;
      RECT 265.905000   3.830000 266.075000   4.120000 ;
      RECT 265.905000   4.120000 271.095000   4.290000 ;
      RECT 265.925000  19.870000 266.095000  22.580000 ;
      RECT 265.925000  23.850000 266.095000  26.560000 ;
      RECT 265.925000  49.045000 266.595000  49.765000 ;
      RECT 265.925000  60.555000 266.595000  60.615000 ;
      RECT 265.935000 200.495000 266.465000 215.995000 ;
      RECT 265.960000  86.580000 266.490000  86.750000 ;
      RECT 265.975000  40.195000 266.145000  41.360000 ;
      RECT 265.975000  45.000000 266.145000  45.030000 ;
      RECT 265.975000  45.200000 266.145000  48.000000 ;
      RECT 265.990000  11.100000 266.500000  11.430000 ;
      RECT 265.990000  17.510000 266.500000  17.840000 ;
      RECT 266.025000  22.750000 278.670000  23.680000 ;
      RECT 266.060000  11.430000 266.430000  17.510000 ;
      RECT 266.075000  38.970000 267.605000  39.720000 ;
      RECT 266.105000  42.505000 266.635000  42.675000 ;
      RECT 266.110000  85.770000 266.280000  86.580000 ;
      RECT 266.110000  86.750000 266.280000  86.780000 ;
      RECT 266.120000  90.110000 267.165000  90.460000 ;
      RECT 266.120000  90.460000 288.200000  90.700000 ;
      RECT 266.175000  49.985000 266.345000  54.895000 ;
      RECT 266.175000  55.455000 266.345000  60.365000 ;
      RECT 266.215000   6.510000 266.745000   6.680000 ;
      RECT 266.215000  68.620000 266.385000  71.415000 ;
      RECT 266.245000   3.660000 271.095000   3.830000 ;
      RECT 266.265000  30.285000 266.435000  31.335000 ;
      RECT 266.265000  31.565000 266.435000  31.895000 ;
      RECT 266.265000  32.515000 266.435000  32.845000 ;
      RECT 266.265000  33.015000 266.435000  36.030000 ;
      RECT 266.315000  37.765000 267.365000  38.970000 ;
      RECT 266.315000  39.720000 267.365000  40.865000 ;
      RECT 266.355000  61.675000 266.525000  67.415000 ;
      RECT 266.370000  88.610000 267.165000  89.690000 ;
      RECT 266.395000   5.020000 266.565000   6.510000 ;
      RECT 266.395000   6.680000 266.565000   9.790000 ;
      RECT 266.465000  42.675000 266.635000  43.615000 ;
      RECT 266.560000 224.125000 276.560000 226.460000 ;
      RECT 266.560000 229.425000 276.560000 232.185000 ;
      RECT 266.560000 235.150000 276.560000 237.910000 ;
      RECT 266.560000 240.875000 276.560000 243.210000 ;
      RECT 266.570000 113.195000 267.240000 113.525000 ;
      RECT 266.600000  11.600000 266.770000  17.345000 ;
      RECT 266.605000  49.985000 267.045000  60.365000 ;
      RECT 266.625000  61.175000 267.135000  61.505000 ;
      RECT 266.625000  67.585000 267.135000  67.915000 ;
      RECT 266.660000  84.070000 266.830000  84.970000 ;
      RECT 266.660000  84.970000 267.190000  85.140000 ;
      RECT 266.660000  85.140000 266.830000  86.780000 ;
      RECT 266.695000  61.505000 267.065000  67.585000 ;
      RECT 266.695000 113.910000 269.695000 164.900000 ;
      RECT 266.720000  11.260000 267.250000  11.430000 ;
      RECT 266.755000  45.290000 266.925000  48.000000 ;
      RECT 266.765000   6.880000 267.295000   7.050000 ;
      RECT 266.875000  87.000000 267.885000  87.170000 ;
      RECT 266.885000  30.285000 267.055000  31.335000 ;
      RECT 266.885000  31.565000 267.055000  31.895000 ;
      RECT 266.885000  32.515000 267.055000  32.845000 ;
      RECT 266.885000  33.015000 267.055000  35.725000 ;
      RECT 266.895000 200.085000 267.565000 200.255000 ;
      RECT 266.895000 216.235000 267.565000 216.405000 ;
      RECT 266.945000   5.020000 267.115000   6.880000 ;
      RECT 266.945000   7.050000 267.115000   9.790000 ;
      RECT 266.980000  44.570000 267.990000  44.740000 ;
      RECT 267.045000  42.505000 267.575000  42.675000 ;
      RECT 267.045000  42.675000 267.215000  43.615000 ;
      RECT 267.050000  85.340000 267.700000  87.000000 ;
      RECT 267.075000  32.075000 267.665000  32.245000 ;
      RECT 267.080000  11.430000 267.250000  11.600000 ;
      RECT 267.080000  11.600000 267.320000  12.610000 ;
      RECT 267.150000  12.610000 267.320000  17.345000 ;
      RECT 267.155000 106.360000 267.685000 106.530000 ;
      RECT 267.205000  19.870000 267.375000  22.580000 ;
      RECT 267.205000  23.850000 267.375000  26.560000 ;
      RECT 267.205000  29.575000 267.735000  29.745000 ;
      RECT 267.205000  42.000000 267.875000  42.170000 ;
      RECT 267.210000  75.510000 267.875000  82.880000 ;
      RECT 267.225000  29.745000 267.735000  30.115000 ;
      RECT 267.225000  36.195000 267.735000  36.525000 ;
      RECT 267.225000  49.985000 267.395000  60.365000 ;
      RECT 267.235000  61.675000 267.405000  62.725000 ;
      RECT 267.235000  62.955000 267.405000  63.285000 ;
      RECT 267.235000  63.905000 267.405000  64.235000 ;
      RECT 267.235000  64.405000 267.405000  67.115000 ;
      RECT 267.275000  42.170000 267.805000  42.300000 ;
      RECT 267.295000  30.115000 267.665000  32.075000 ;
      RECT 267.295000  32.245000 267.665000  36.195000 ;
      RECT 267.305000   6.510000 269.335000   6.680000 ;
      RECT 267.310000  72.550000 267.875000  75.510000 ;
      RECT 267.345000  70.675000 267.875000  70.845000 ;
      RECT 267.390000  10.260000 267.900000  10.390000 ;
      RECT 267.390000  10.390000 268.000000  10.560000 ;
      RECT 267.390000  10.560000 267.900000  10.590000 ;
      RECT 267.405000  89.285000 287.220000  89.455000 ;
      RECT 267.405000 190.115000 267.915000 190.145000 ;
      RECT 267.405000 190.415000 267.915000 190.445000 ;
      RECT 267.405000 190.895000 267.915000 190.925000 ;
      RECT 267.405000 191.195000 267.915000 191.225000 ;
      RECT 267.420000  11.100000 267.930000  11.430000 ;
      RECT 267.420000  17.510000 267.930000  17.840000 ;
      RECT 267.460000  44.740000 267.990000  44.800000 ;
      RECT 267.480000 185.070000 268.770000 187.295000 ;
      RECT 267.490000  11.430000 267.860000  17.510000 ;
      RECT 267.495000  68.620000 267.665000  70.675000 ;
      RECT 267.495000  70.845000 267.665000  71.330000 ;
      RECT 267.515000 105.400000 267.685000 106.360000 ;
      RECT 267.515000 106.530000 267.685000 106.750000 ;
      RECT 267.535000  37.335000 269.790000  37.505000 ;
      RECT 267.535000  37.505000 269.675000  37.595000 ;
      RECT 267.535000  37.595000 267.915000  38.615000 ;
      RECT 267.535000  40.195000 267.705000  41.360000 ;
      RECT 267.535000  41.360000 268.455000  41.530000 ;
      RECT 267.535000  45.000000 267.705000  45.030000 ;
      RECT 267.535000  45.030000 268.080000  45.200000 ;
      RECT 267.535000  45.200000 267.705000  48.000000 ;
      RECT 267.560000  60.535000 271.290000  60.855000 ;
      RECT 267.565000  49.595000 268.235000  60.535000 ;
      RECT 267.575000  61.175000 268.085000  61.505000 ;
      RECT 267.575000  67.585000 268.965000  67.915000 ;
      RECT 267.645000  61.505000 268.015000  67.585000 ;
      RECT 267.665000 180.175000 293.520000 180.515000 ;
      RECT 267.835000  30.285000 268.005000  34.755000 ;
      RECT 267.895000  88.360000 268.600000  89.285000 ;
      RECT 267.925000  42.605000 268.095000  44.400000 ;
      RECT 267.925000 104.700000 268.095000 107.090000 ;
      RECT 267.940000  84.070000 268.110000  86.780000 ;
      RECT 267.995000 200.495000 268.525000 215.995000 ;
      RECT 268.030000  11.600000 268.200000  13.210000 ;
      RECT 268.030000  13.830000 268.200000  14.160000 ;
      RECT 268.030000  14.330000 268.200000  17.040000 ;
      RECT 268.035000  69.905000 268.565000  70.075000 ;
      RECT 268.045000  68.950000 268.215000  69.905000 ;
      RECT 268.045000  70.075000 268.215000  71.660000 ;
      RECT 268.080000  72.820000 268.250000  73.325000 ;
      RECT 268.080000  73.325000 268.610000  73.495000 ;
      RECT 268.080000  73.495000 268.250000  77.570000 ;
      RECT 268.080000  78.120000 268.250000  81.770000 ;
      RECT 268.080000  81.770000 268.610000  81.940000 ;
      RECT 268.080000  81.940000 268.250000  82.870000 ;
      RECT 268.085000  38.155000 268.255000  40.395000 ;
      RECT 268.085000  40.395000 268.795000  40.865000 ;
      RECT 268.085000 189.635000 268.770000 190.805000 ;
      RECT 268.090000  36.265000 268.620000  36.435000 ;
      RECT 268.105000  29.785000 268.615000  30.115000 ;
      RECT 268.105000  36.195000 268.615000  36.265000 ;
      RECT 268.105000  36.435000 268.615000  36.525000 ;
      RECT 268.130000  41.530000 268.455000  41.785000 ;
      RECT 268.130000  41.785000 268.750000  42.115000 ;
      RECT 268.165000  87.000000 269.175000  87.170000 ;
      RECT 268.175000  30.115000 268.545000  36.195000 ;
      RECT 268.185000  61.675000 268.355000  66.145000 ;
      RECT 268.225000   5.020000 268.395000   6.280000 ;
      RECT 268.225000   7.080000 268.395000   9.790000 ;
      RECT 268.235000  72.140000 268.905000  72.310000 ;
      RECT 268.235000  83.090000 268.905000  83.490000 ;
      RECT 268.290000  17.700000 268.820000  17.870000 ;
      RECT 268.300000  11.100000 268.810000  11.430000 ;
      RECT 268.300000  17.510000 268.810000  17.700000 ;
      RECT 268.315000  45.290000 268.485000  48.000000 ;
      RECT 268.325000  68.230000 271.040000  68.555000 ;
      RECT 268.335000  84.570000 268.865000  84.740000 ;
      RECT 268.335000  84.740000 268.690000  86.580000 ;
      RECT 268.335000  86.580000 268.985000  87.000000 ;
      RECT 268.365000  66.745000 268.895000  66.915000 ;
      RECT 268.370000  11.430000 268.740000  17.510000 ;
      RECT 268.405000  49.955000 269.195000  54.705000 ;
      RECT 268.405000  54.705000 268.575000  60.365000 ;
      RECT 268.420000  72.310000 268.790000  73.155000 ;
      RECT 268.455000  61.175000 268.965000  61.505000 ;
      RECT 268.485000  19.870000 268.655000  22.580000 ;
      RECT 268.485000  23.850000 268.655000  26.560000 ;
      RECT 268.525000  61.505000 268.895000  66.745000 ;
      RECT 268.525000  66.915000 268.895000  67.585000 ;
      RECT 268.625000  40.865000 268.795000  41.445000 ;
      RECT 268.625000  41.445000 269.090000  41.615000 ;
      RECT 268.635000  70.675000 269.165000  70.845000 ;
      RECT 268.785000  30.285000 268.955000  31.335000 ;
      RECT 268.785000  31.565000 268.955000  31.895000 ;
      RECT 268.785000  32.515000 268.955000  32.845000 ;
      RECT 268.785000  33.015000 268.955000  36.030000 ;
      RECT 268.805000  42.520000 269.090000  42.690000 ;
      RECT 268.805000  42.690000 268.975000  43.615000 ;
      RECT 268.825000  68.950000 268.995000  70.675000 ;
      RECT 268.825000  70.845000 268.995000  71.660000 ;
      RECT 268.860000  85.340000 269.390000  85.510000 ;
      RECT 268.860000 103.770000 271.970000 108.380000 ;
      RECT 268.910000  11.725000 269.080000  17.345000 ;
      RECT 268.920000  41.615000 269.090000  42.520000 ;
      RECT 268.940000 180.515000 293.520000 183.710000 ;
      RECT 268.940000 183.710000 342.805000 185.670000 ;
      RECT 268.940000 185.670000 309.875000 186.220000 ;
      RECT 268.940000 186.220000 283.670000 188.775000 ;
      RECT 268.940000 188.775000 283.675000 189.945000 ;
      RECT 268.940000 189.945000 283.670000 191.905000 ;
      RECT 268.955000 200.085000 269.625000 200.255000 ;
      RECT 268.955000 216.235000 269.625000 216.405000 ;
      RECT 268.960000  72.820000 269.130000  77.570000 ;
      RECT 268.960000  78.120000 269.130000  82.870000 ;
      RECT 268.965000  37.765000 269.135000  40.865000 ;
      RECT 269.025000  55.085000 271.555000  55.285000 ;
      RECT 269.025000  55.285000 269.195000  60.365000 ;
      RECT 269.120000  41.085000 269.790000  41.255000 ;
      RECT 269.130000 113.195000 269.800000 113.525000 ;
      RECT 269.135000  61.675000 269.305000  62.725000 ;
      RECT 269.135000  62.955000 270.700000  63.285000 ;
      RECT 269.135000  63.905000 270.700000  64.235000 ;
      RECT 269.135000  64.405000 269.305000  67.420000 ;
      RECT 269.145000  43.110000 269.675000  48.390000 ;
      RECT 269.170000  17.700000 269.700000  17.870000 ;
      RECT 269.180000  11.100000 269.690000  11.430000 ;
      RECT 269.180000  17.510000 269.690000  17.700000 ;
      RECT 269.195000  72.140000 270.885000  72.310000 ;
      RECT 269.205000   8.840000 273.255000   9.270000 ;
      RECT 269.205000   9.270000 273.795000   9.645000 ;
      RECT 269.205000   9.645000 275.555000  10.760000 ;
      RECT 269.220000  84.070000 269.390000  85.340000 ;
      RECT 269.220000  85.510000 269.390000  86.780000 ;
      RECT 269.250000  11.430000 269.620000  17.510000 ;
      RECT 269.255000  49.595000 271.285000  49.765000 ;
      RECT 269.260000  41.760000 269.790000  41.930000 ;
      RECT 269.260000  41.930000 269.570000  43.110000 ;
      RECT 269.300000  72.310000 269.670000  73.155000 ;
      RECT 269.305000  37.595000 269.675000  41.085000 ;
      RECT 269.305000  41.255000 269.790000  41.265000 ;
      RECT 269.305000  41.265000 270.270000  41.435000 ;
      RECT 269.325000   7.380000 269.855000   7.550000 ;
      RECT 269.380000  83.090000 272.770000  83.510000 ;
      RECT 269.420000  69.905000 269.950000  70.075000 ;
      RECT 269.480000  30.285000 269.650000  31.795000 ;
      RECT 269.480000  32.515000 269.650000  36.025000 ;
      RECT 269.505000   5.020000 269.675000   7.380000 ;
      RECT 269.505000   7.550000 269.675000   8.160000 ;
      RECT 269.605000  68.950000 269.775000  69.905000 ;
      RECT 269.605000  70.075000 269.775000  71.660000 ;
      RECT 269.670000  73.325000 270.200000  73.495000 ;
      RECT 269.670000  81.770000 270.200000  81.940000 ;
      RECT 269.695000  48.990000 270.225000  49.595000 ;
      RECT 269.720000  61.675000 269.890000  62.955000 ;
      RECT 269.720000  64.235000 270.700000  67.115000 ;
      RECT 269.720000  67.115000 269.890000  67.415000 ;
      RECT 269.725000  53.370000 270.255000  53.540000 ;
      RECT 269.740000  42.130000 270.270000  42.300000 ;
      RECT 269.765000  19.870000 269.935000  22.580000 ;
      RECT 269.765000  23.850000 269.935000  26.560000 ;
      RECT 269.770000  83.730000 273.060000  83.900000 ;
      RECT 269.770000  83.900000 269.940000  86.780000 ;
      RECT 269.790000  11.600000 269.960000  13.420000 ;
      RECT 269.790000  14.330000 269.960000  17.040000 ;
      RECT 269.805000  49.955000 269.975000  53.370000 ;
      RECT 269.805000  53.540000 269.975000  54.705000 ;
      RECT 269.840000  72.820000 270.010000  73.325000 ;
      RECT 269.840000  73.495000 270.010000  77.570000 ;
      RECT 269.840000  78.120000 270.010000  81.770000 ;
      RECT 269.840000  81.940000 270.010000  82.870000 ;
      RECT 269.845000  38.155000 270.130000  40.865000 ;
      RECT 269.865000  44.180000 271.425000  44.350000 ;
      RECT 269.865000  44.350000 270.035000  45.760000 ;
      RECT 269.865000  45.760000 272.395000  45.930000 ;
      RECT 269.865000  46.100000 270.035000  46.335000 ;
      RECT 269.865000  46.335000 270.395000  46.505000 ;
      RECT 269.865000  46.505000 270.035000  48.380000 ;
      RECT 269.960000  40.865000 270.130000  41.095000 ;
      RECT 269.960000  41.435000 270.270000  42.130000 ;
      RECT 269.965000  42.840000 270.135000  44.010000 ;
      RECT 270.010000  83.690000 273.060000  83.730000 ;
      RECT 270.050000  87.000000 272.760000  87.005000 ;
      RECT 270.050000  87.005000 272.765000  87.170000 ;
      RECT 270.055000 200.495000 270.585000 215.995000 ;
      RECT 270.075000  87.170000 272.765000  87.175000 ;
      RECT 270.180000  72.310000 270.550000  73.155000 ;
      RECT 270.195000  70.305000 270.725000  70.475000 ;
      RECT 270.205000  55.455000 270.375000  60.365000 ;
      RECT 270.250000  42.470000 271.600000  42.640000 ;
      RECT 270.350000  42.640000 271.600000  42.670000 ;
      RECT 270.360000  85.340000 270.890000  85.510000 ;
      RECT 270.385000  68.950000 270.555000  70.305000 ;
      RECT 270.385000  70.475000 270.555000  71.660000 ;
      RECT 270.395000  42.840000 270.565000  44.180000 ;
      RECT 270.425000  37.765000 270.595000  40.845000 ;
      RECT 270.530000  61.675000 270.700000  62.725000 ;
      RECT 270.550000  84.070000 270.720000  85.340000 ;
      RECT 270.550000  85.510000 270.720000  86.780000 ;
      RECT 270.570000  49.955000 270.740000  55.085000 ;
      RECT 270.720000  72.820000 270.890000  77.570000 ;
      RECT 270.720000  78.120000 270.890000  82.870000 ;
      RECT 270.785000   5.020000 270.955000   6.280000 ;
      RECT 270.785000   7.150000 270.955000   8.840000 ;
      RECT 270.800000  61.175000 271.310000  61.505000 ;
      RECT 270.800000  67.585000 271.310000  67.915000 ;
      RECT 270.805000  69.905000 271.375000  70.075000 ;
      RECT 270.825000  42.840000 270.995000  44.010000 ;
      RECT 270.870000  61.505000 271.240000  67.585000 ;
      RECT 270.915000  10.930000 275.555000  11.370000 ;
      RECT 270.955000  11.720000 271.125000  12.900000 ;
      RECT 270.955000  12.900000 272.885000  13.180000 ;
      RECT 271.015000 200.085000 271.685000 200.255000 ;
      RECT 271.015000 216.235000 271.685000 216.405000 ;
      RECT 271.045000  19.870000 271.215000  22.580000 ;
      RECT 271.045000  23.850000 271.215000  26.560000 ;
      RECT 271.045000  44.580000 271.215000  45.280000 ;
      RECT 271.045000  45.280000 271.720000  45.450000 ;
      RECT 271.045000  45.450000 271.215000  45.590000 ;
      RECT 271.045000  46.100000 271.215000  48.550000 ;
      RECT 271.045000  48.550000 273.935000  48.720000 ;
      RECT 271.050000   6.470000 272.590000   6.640000 ;
      RECT 271.085000  68.950000 271.375000  69.905000 ;
      RECT 271.085000  70.075000 271.375000  71.960000 ;
      RECT 271.085000  71.960000 271.690000  72.250000 ;
      RECT 271.085000 199.300000 271.615000 200.085000 ;
      RECT 271.205000 113.910000 274.205000 164.900000 ;
      RECT 271.240000  73.325000 271.770000  73.495000 ;
      RECT 271.240000  81.770000 271.770000  81.940000 ;
      RECT 271.245000   6.810000 273.255000   6.980000 ;
      RECT 271.245000   6.980000 271.415000   8.160000 ;
      RECT 271.255000  13.900000 271.425000  17.270000 ;
      RECT 271.255000  17.270000 275.225000  18.040000 ;
      RECT 271.255000  42.840000 271.425000  44.180000 ;
      RECT 271.265000   4.770000 271.435000   6.040000 ;
      RECT 271.315000   3.410000 272.590000   4.080000 ;
      RECT 271.330000  83.900000 271.500000  86.780000 ;
      RECT 271.350000  49.955000 271.520000  50.845000 ;
      RECT 271.350000  50.845000 272.185000  54.705000 ;
      RECT 271.385000  55.285000 271.555000  60.365000 ;
      RECT 271.410000  61.675000 271.580000  67.415000 ;
      RECT 271.480000  72.250000 271.690000  72.820000 ;
      RECT 271.480000  72.820000 271.770000  73.325000 ;
      RECT 271.480000  73.495000 271.770000  77.570000 ;
      RECT 271.545000  46.165000 271.875000  47.015000 ;
      RECT 271.600000  78.120000 271.770000  81.770000 ;
      RECT 271.600000  81.940000 271.770000  82.870000 ;
      RECT 271.625000  47.015000 271.795000  47.625000 ;
      RECT 271.680000  61.175000 272.190000  61.505000 ;
      RECT 271.680000  67.585000 272.190000  67.915000 ;
      RECT 271.685000  42.840000 271.855000  44.010000 ;
      RECT 271.705000   7.150000 271.875000   8.840000 ;
      RECT 271.750000  61.505000 272.120000  67.585000 ;
      RECT 271.770000  37.870000 271.940000  40.870000 ;
      RECT 271.805000  55.895000 272.335000  56.065000 ;
      RECT 271.835000  11.720000 272.005000  12.730000 ;
      RECT 271.835000  14.210000 272.005000  16.920000 ;
      RECT 271.860000  68.490000 272.030000  72.305000 ;
      RECT 271.920000  84.970000 272.450000  85.140000 ;
      RECT 271.955000  42.470000 273.305000  42.475000 ;
      RECT 271.955000  42.475000 274.615000  42.645000 ;
      RECT 271.990000  41.360000 272.520000  41.530000 ;
      RECT 272.010000   4.080000 272.590000   6.470000 ;
      RECT 272.015000  54.705000 272.185000  55.895000 ;
      RECT 272.080000  13.180000 272.360000  13.760000 ;
      RECT 272.080000  13.760000 272.885000  14.040000 ;
      RECT 272.110000  84.070000 272.280000  84.970000 ;
      RECT 272.110000  85.140000 272.280000  86.780000 ;
      RECT 272.115000  42.840000 272.285000  44.180000 ;
      RECT 272.115000  44.180000 273.935000  44.350000 ;
      RECT 272.115000 200.495000 272.645000 215.995000 ;
      RECT 272.165000   6.980000 272.335000   8.160000 ;
      RECT 272.165000  56.755000 273.015000  58.725000 ;
      RECT 272.165000  58.725000 273.055000  59.255000 ;
      RECT 272.165000  59.255000 273.015000  60.485000 ;
      RECT 272.170000  49.085000 272.840000  50.625000 ;
      RECT 272.170000  72.545000 272.885000  78.155000 ;
      RECT 272.170000  78.155000 287.460000  78.570000 ;
      RECT 272.170000  78.570000 272.885000  82.850000 ;
      RECT 272.225000  44.580000 272.395000  45.760000 ;
      RECT 272.225000  45.930000 272.395000  47.080000 ;
      RECT 272.225000  47.370000 273.095000  48.380000 ;
      RECT 272.290000  61.675000 272.460000  62.740000 ;
      RECT 272.290000  62.910000 272.460000  63.285000 ;
      RECT 272.290000  63.905000 272.460000  64.235000 ;
      RECT 272.290000  64.405000 272.460000  67.115000 ;
      RECT 272.295000 199.685000 272.825000 200.255000 ;
      RECT 272.310000  56.265000 272.840000  56.435000 ;
      RECT 272.325000  19.870000 272.495000  22.580000 ;
      RECT 272.325000  23.850000 272.495000  26.560000 ;
      RECT 272.350000  37.840000 276.590000  38.010000 ;
      RECT 272.350000  38.010000 272.520000  41.360000 ;
      RECT 272.355000  14.040000 272.885000  14.160000 ;
      RECT 272.355000  50.625000 272.725000  55.420000 ;
      RECT 272.510000  55.785000 272.840000  56.265000 ;
      RECT 272.530000  13.350000 273.540000  13.520000 ;
      RECT 272.545000  42.840000 272.715000  44.010000 ;
      RECT 272.560000  61.175000 273.070000  61.505000 ;
      RECT 272.560000  67.585000 273.070000  67.590000 ;
      RECT 272.560000  67.590000 273.950000  67.920000 ;
      RECT 272.565000  46.335000 273.095000  47.370000 ;
      RECT 272.575000  37.045000 274.605000  37.505000 ;
      RECT 272.625000   7.150000 272.795000   8.840000 ;
      RECT 272.630000  61.505000 273.000000  67.585000 ;
      RECT 272.645000   3.040000 273.315000   3.210000 ;
      RECT 272.715000  11.720000 272.885000  12.900000 ;
      RECT 272.715000  14.160000 272.885000  16.920000 ;
      RECT 272.760000   3.210000 273.030000   5.115000 ;
      RECT 272.890000  83.900000 273.060000  86.780000 ;
      RECT 272.895000  50.845000 273.065000  55.525000 ;
      RECT 272.975000  42.840000 273.145000  44.180000 ;
      RECT 273.045000  45.280000 273.575000  45.450000 ;
      RECT 273.055000  55.895000 273.585000  56.065000 ;
      RECT 273.075000 200.085000 273.745000 200.255000 ;
      RECT 273.075000 216.235000 273.745000 216.405000 ;
      RECT 273.085000   6.980000 273.255000   8.160000 ;
      RECT 273.120000  49.090000 273.790000  50.625000 ;
      RECT 273.125000 102.115000 299.555000 107.805000 ;
      RECT 273.170000  61.800000 273.340000  67.420000 ;
      RECT 273.200000   3.760000 273.370000   6.470000 ;
      RECT 273.200000  79.090000 277.950000  79.260000 ;
      RECT 273.200000  79.970000 278.090000  80.135000 ;
      RECT 273.200000  80.135000 277.950000  80.140000 ;
      RECT 273.200000  80.850000 277.950000  81.020000 ;
      RECT 273.200000  81.730000 278.090000  81.895000 ;
      RECT 273.200000  81.895000 277.950000  81.900000 ;
      RECT 273.200000  82.610000 277.950000  82.780000 ;
      RECT 273.230000  38.180000 273.490000  41.160000 ;
      RECT 273.245000  53.995000 273.575000  54.325000 ;
      RECT 273.255000  55.785000 273.585000  55.895000 ;
      RECT 273.255000  56.065000 273.585000  56.295000 ;
      RECT 273.260000  13.520000 273.540000  13.720000 ;
      RECT 273.260000  13.720000 274.940000  13.770000 ;
      RECT 273.260000  13.770000 274.885000  14.000000 ;
      RECT 273.290000  74.765000 273.460000  77.080000 ;
      RECT 273.290000  77.080000 273.820000  77.250000 ;
      RECT 273.290000  77.250000 273.460000  77.475000 ;
      RECT 273.370000  83.610000 273.540000  86.760000 ;
      RECT 273.405000  42.840000 273.575000  44.010000 ;
      RECT 273.405000  44.580000 273.575000  45.280000 ;
      RECT 273.405000  45.450000 273.575000  47.080000 ;
      RECT 273.405000  47.370000 273.935000  48.550000 ;
      RECT 273.415000  53.370000 273.945000  53.540000 ;
      RECT 273.440000  61.175000 273.950000  61.505000 ;
      RECT 273.440000  67.585000 273.950000  67.590000 ;
      RECT 273.510000  61.505000 273.880000  64.025000 ;
      RECT 273.510000  64.025000 274.770000  64.235000 ;
      RECT 273.510000  64.235000 273.880000  67.585000 ;
      RECT 273.595000  11.370000 273.765000  12.730000 ;
      RECT 273.595000  14.210000 273.765000  16.920000 ;
      RECT 273.605000   6.840000 274.350000   7.010000 ;
      RECT 273.605000   7.010000 273.775000   8.760000 ;
      RECT 273.605000  19.870000 273.775000  22.580000 ;
      RECT 273.605000  23.850000 273.775000  26.560000 ;
      RECT 273.625000   4.440000 273.795000   4.505000 ;
      RECT 273.625000   4.505000 273.830000   4.970000 ;
      RECT 273.660000   4.970000 273.830000   5.175000 ;
      RECT 273.690000  38.180000 273.950000  41.160000 ;
      RECT 273.720000   5.660000 273.890000   6.670000 ;
      RECT 273.745000  43.095000 274.275000  43.265000 ;
      RECT 273.745000  44.350000 273.935000  47.370000 ;
      RECT 273.775000  50.845000 273.945000  53.370000 ;
      RECT 273.775000  53.540000 273.945000  56.265000 ;
      RECT 273.775000  56.265000 274.305000  56.435000 ;
      RECT 273.820000  13.350000 274.490000  13.520000 ;
      RECT 273.850000  84.275000 274.020000  87.055000 ;
      RECT 273.865000  41.360000 274.395000  41.530000 ;
      RECT 273.945000   7.180000 274.615000   7.260000 ;
      RECT 273.945000   7.260000 277.375000   7.380000 ;
      RECT 273.945000   7.380000 277.385000   7.430000 ;
      RECT 274.000000   3.275000 274.530000   3.295000 ;
      RECT 274.000000   3.295000 279.140000   3.445000 ;
      RECT 274.000000   4.740000 279.140000   4.910000 ;
      RECT 274.045000  41.530000 274.215000  42.305000 ;
      RECT 274.050000   3.445000 279.140000   3.465000 ;
      RECT 274.050000   3.755000 278.800000   3.925000 ;
      RECT 274.050000   4.280000 278.800000   4.450000 ;
      RECT 274.050000   5.200000 278.975000   5.390000 ;
      RECT 274.050000  49.015000 274.580000  49.785000 ;
      RECT 274.050000  49.785000 274.905000  49.955000 ;
      RECT 274.050000  61.675000 274.220000  63.855000 ;
      RECT 274.050000  64.405000 274.220000  67.115000 ;
      RECT 274.065000   7.750000 274.235000   8.760000 ;
      RECT 274.095000  57.325000 274.265000  60.405000 ;
      RECT 274.105000  43.265000 274.275000  49.015000 ;
      RECT 274.115000   4.450000 278.605000   4.455000 ;
      RECT 274.115000  50.875000 274.565000  51.740000 ;
      RECT 274.115000  51.740000 274.645000  51.910000 ;
      RECT 274.115000  51.910000 274.300000  52.775000 ;
      RECT 274.115000  52.775000 274.565000  53.770000 ;
      RECT 274.115000  53.770000 274.645000  54.055000 ;
      RECT 274.115000  54.055000 278.240000  54.385000 ;
      RECT 274.115000  54.385000 275.440000  54.660000 ;
      RECT 274.140000  68.085000 287.190000  68.255000 ;
      RECT 274.140000  68.255000 274.310000  73.625000 ;
      RECT 274.170000  74.340000 276.650000  74.595000 ;
      RECT 274.170000  74.595000 274.340000  77.475000 ;
      RECT 274.175000   6.670000 274.350000   6.840000 ;
      RECT 274.175000 199.300000 274.705000 200.255000 ;
      RECT 274.175000 200.495000 274.705000 215.995000 ;
      RECT 274.180000   5.660000 274.350000   6.670000 ;
      RECT 274.235000  87.275000 276.805000  87.475000 ;
      RECT 274.290000   9.010000 275.005000   9.180000 ;
      RECT 274.310000   3.675000 278.800000   3.755000 ;
      RECT 274.320000  79.965000 278.090000  79.970000 ;
      RECT 274.445000  42.645000 274.615000  43.405000 ;
      RECT 274.445000  43.405000 275.095000  44.415000 ;
      RECT 274.450000  85.230000 274.980000  85.400000 ;
      RECT 274.455000  81.725000 278.090000  81.730000 ;
      RECT 274.470000  52.095000 274.800000  52.230000 ;
      RECT 274.470000  52.230000 275.000000  52.400000 ;
      RECT 274.470000  52.400000 274.800000  52.605000 ;
      RECT 274.475000   9.180000 275.005000   9.475000 ;
      RECT 274.475000  11.720000 274.645000  12.725000 ;
      RECT 274.475000  12.725000 274.940000  13.005000 ;
      RECT 274.475000  14.000000 274.885000  14.210000 ;
      RECT 274.475000  14.210000 274.645000  16.920000 ;
      RECT 274.565000  41.290000 275.235000  41.460000 ;
      RECT 274.565000  46.335000 275.095000  46.505000 ;
      RECT 274.585000  47.855000 274.755000  48.465000 ;
      RECT 274.585000  48.465000 280.115000  48.635000 ;
      RECT 274.600000  61.675000 274.770000  64.025000 ;
      RECT 274.600000  64.235000 274.770000  67.420000 ;
      RECT 274.625000  42.030000 275.155000  42.200000 ;
      RECT 274.630000  84.345000 274.800000  85.230000 ;
      RECT 274.630000  85.400000 274.800000  87.055000 ;
      RECT 274.640000   5.390000 274.810000   6.670000 ;
      RECT 274.660000  13.005000 274.940000  13.720000 ;
      RECT 274.660000  38.180000 274.830000  41.290000 ;
      RECT 274.660000  41.460000 275.155000  42.030000 ;
      RECT 274.720000  68.605000 274.890000  69.905000 ;
      RECT 274.720000  69.905000 275.250000  70.075000 ;
      RECT 274.720000  70.075000 274.890000  74.340000 ;
      RECT 274.775000  57.005000 275.440000  57.175000 ;
      RECT 274.775000  57.175000 274.945000  60.015000 ;
      RECT 274.815000  37.335000 275.485000  37.505000 ;
      RECT 274.830000  60.665000 277.595000  60.835000 ;
      RECT 274.855000  50.535000 275.945000  50.705000 ;
      RECT 274.855000  50.705000 275.025000  51.885000 ;
      RECT 274.855000  52.875000 275.025000  53.885000 ;
      RECT 274.870000  61.175000 275.380000  61.505000 ;
      RECT 274.870000  67.585000 275.380000  67.915000 ;
      RECT 274.870000  77.080000 275.400000  77.250000 ;
      RECT 274.885000  19.870000 275.055000  22.580000 ;
      RECT 274.885000  23.850000 275.055000  26.560000 ;
      RECT 274.910000  55.525000 275.440000  57.005000 ;
      RECT 274.925000  44.415000 275.095000  46.335000 ;
      RECT 274.925000  46.505000 275.095000  48.085000 ;
      RECT 274.940000  61.505000 275.310000  67.585000 ;
      RECT 275.015000   6.920000 275.685000   7.090000 ;
      RECT 275.050000  74.765000 275.220000  77.080000 ;
      RECT 275.050000  77.250000 275.220000  77.475000 ;
      RECT 275.055000  13.900000 275.225000  17.270000 ;
      RECT 275.080000  49.415000 275.750000  50.365000 ;
      RECT 275.135000 200.085000 275.805000 200.255000 ;
      RECT 275.135000 216.235000 275.805000 216.405000 ;
      RECT 275.180000  39.675000 275.710000  39.845000 ;
      RECT 275.180000  73.865000 276.190000  74.035000 ;
      RECT 275.240000  73.600000 276.130000  73.865000 ;
      RECT 275.255000   7.720000 275.785000   9.070000 ;
      RECT 275.265000  45.000000 275.795000  45.170000 ;
      RECT 275.275000  50.875000 275.485000  51.885000 ;
      RECT 275.275000  51.885000 275.475000  52.875000 ;
      RECT 275.275000  52.875000 275.485000  53.935000 ;
      RECT 275.275000  53.935000 278.240000  54.055000 ;
      RECT 275.325000  41.635000 275.575000  42.305000 ;
      RECT 275.355000  11.720000 275.525000  12.730000 ;
      RECT 275.355000  54.905000 275.885000  55.075000 ;
      RECT 275.360000  41.580000 275.575000  41.635000 ;
      RECT 275.360000  42.305000 275.530000  43.405000 ;
      RECT 275.360000  43.405000 275.555000  44.415000 ;
      RECT 275.385000   9.380000 275.555000   9.645000 ;
      RECT 275.385000  45.170000 275.555000  48.085000 ;
      RECT 275.405000  38.180000 275.710000  39.675000 ;
      RECT 275.405000  39.845000 275.710000  40.890000 ;
      RECT 275.405000  40.890000 275.575000  41.580000 ;
      RECT 275.410000  84.275000 275.580000  87.055000 ;
      RECT 275.480000  61.675000 275.650000  62.740000 ;
      RECT 275.480000  62.910000 275.650000  63.285000 ;
      RECT 275.480000  63.905000 275.650000  64.235000 ;
      RECT 275.480000  64.405000 275.650000  67.115000 ;
      RECT 275.555000  57.305000 275.725000  60.405000 ;
      RECT 275.590000 113.195000 276.260000 113.525000 ;
      RECT 275.600000  68.255000 275.770000  73.355000 ;
      RECT 275.610000  54.555000 275.885000  54.905000 ;
      RECT 275.610000  55.075000 275.885000  55.565000 ;
      RECT 275.610000  55.565000 275.780000  56.870000 ;
      RECT 275.610000  56.870000 276.505000  57.040000 ;
      RECT 275.635000  14.170000 275.805000  18.920000 ;
      RECT 275.645000  52.355000 276.155000  52.685000 ;
      RECT 275.715000 113.910000 278.715000 164.900000 ;
      RECT 275.725000  42.400000 276.255000  42.570000 ;
      RECT 275.725000  42.570000 276.135000  44.585000 ;
      RECT 275.725000  44.585000 276.265000  44.740000 ;
      RECT 275.725000  45.375000 276.265000  45.665000 ;
      RECT 275.725000  45.665000 276.015000  48.085000 ;
      RECT 275.745000  42.030000 276.775000  42.200000 ;
      RECT 275.750000  61.175000 276.260000  61.435000 ;
      RECT 275.750000  61.435000 276.350000  61.505000 ;
      RECT 275.750000  67.585000 276.260000  67.915000 ;
      RECT 275.765000  37.335000 276.435000  37.505000 ;
      RECT 275.775000  50.705000 275.945000  52.355000 ;
      RECT 275.775000  52.685000 275.945000  52.840000 ;
      RECT 275.820000  61.505000 276.350000  61.605000 ;
      RECT 275.820000  61.605000 276.190000  67.585000 ;
      RECT 275.845000  41.290000 276.590000  41.460000 ;
      RECT 275.845000 195.440000 342.805000 195.445000 ;
      RECT 275.865000  36.980000 276.035000  37.335000 ;
      RECT 275.865000  37.505000 276.035000  37.510000 ;
      RECT 275.915000  41.460000 276.445000  41.530000 ;
      RECT 275.920000   5.660000 276.090000   7.070000 ;
      RECT 275.920000   7.070000 277.375000   7.260000 ;
      RECT 275.930000  74.595000 276.100000  77.475000 ;
      RECT 275.950000  55.735000 276.460000  56.265000 ;
      RECT 275.950000  56.265000 276.480000  56.515000 ;
      RECT 275.950000  56.515000 277.155000  56.700000 ;
      RECT 275.965000   7.720000 276.135000  12.470000 ;
      RECT 275.965000  44.740000 276.265000  45.375000 ;
      RECT 275.985000  13.490000 280.735000  13.570000 ;
      RECT 275.985000  13.570000 280.865000  13.660000 ;
      RECT 275.990000  86.680000 276.520000  86.850000 ;
      RECT 276.095000  49.735000 278.505000  49.760000 ;
      RECT 276.095000  49.760000 281.950000  49.790000 ;
      RECT 276.095000  49.790000 290.205000  49.975000 ;
      RECT 276.095000  49.975000 293.435000  50.405000 ;
      RECT 276.120000  12.950000 276.790000  13.120000 ;
      RECT 276.165000  19.870000 276.335000  22.580000 ;
      RECT 276.165000  23.850000 276.335000  26.560000 ;
      RECT 276.190000  84.345000 276.360000  86.680000 ;
      RECT 276.190000  86.850000 276.360000  87.055000 ;
      RECT 276.215000  48.105000 276.970000  48.275000 ;
      RECT 276.235000  53.770000 278.240000  53.935000 ;
      RECT 276.235000  54.385000 276.765000  54.660000 ;
      RECT 276.235000 199.685000 276.765000 200.255000 ;
      RECT 276.235000 200.495000 276.765000 215.995000 ;
      RECT 276.260000  12.910000 276.790000  12.950000 ;
      RECT 276.300000  69.905000 276.830000  70.075000 ;
      RECT 276.305000  43.405000 276.475000  44.415000 ;
      RECT 276.325000  49.280000 278.505000  49.735000 ;
      RECT 276.335000  57.040000 276.505000  60.015000 ;
      RECT 276.360000  61.800000 276.530000  67.420000 ;
      RECT 276.410000  50.405000 293.435000  50.600000 ;
      RECT 276.410000  50.600000 295.115000  51.555000 ;
      RECT 276.415000  51.555000 295.115000  53.600000 ;
      RECT 276.415000  53.600000 278.240000  53.770000 ;
      RECT 276.420000  38.010000 276.590000  41.290000 ;
      RECT 276.440000  46.335000 276.970000  46.505000 ;
      RECT 276.450000  77.080000 276.980000  77.250000 ;
      RECT 276.460000  44.630000 276.630000  45.300000 ;
      RECT 276.480000  68.605000 276.650000  69.905000 ;
      RECT 276.480000  70.075000 276.650000  73.815000 ;
      RECT 276.480000  73.815000 280.170000  73.985000 ;
      RECT 276.480000  73.985000 276.650000  74.340000 ;
      RECT 276.495000   6.510000 277.025000   6.680000 ;
      RECT 276.500000  42.510000 277.035000  43.085000 ;
      RECT 276.515000  14.170000 276.685000  18.920000 ;
      RECT 276.565000  61.065000 277.095000  61.175000 ;
      RECT 276.565000  61.175000 277.140000  61.235000 ;
      RECT 276.595000  54.660000 276.765000  55.565000 ;
      RECT 276.605000  41.635000 276.775000  42.030000 ;
      RECT 276.605000  42.200000 276.775000  42.305000 ;
      RECT 276.630000  61.235000 277.140000  61.505000 ;
      RECT 276.630000  67.585000 277.140000  67.915000 ;
      RECT 276.665000  11.320000 277.195000  11.490000 ;
      RECT 276.700000  61.505000 277.070000  67.585000 ;
      RECT 276.715000   5.680000 276.885000   6.510000 ;
      RECT 276.765000  43.405000 276.970000  44.415000 ;
      RECT 276.800000  44.415000 276.970000  46.335000 ;
      RECT 276.800000  46.505000 276.970000  48.105000 ;
      RECT 276.810000  74.765000 276.980000  77.080000 ;
      RECT 276.810000  77.250000 276.980000  77.475000 ;
      RECT 276.845000   7.720000 277.015000  11.320000 ;
      RECT 276.845000  11.490000 277.015000  12.470000 ;
      RECT 276.855000   7.430000 277.385000   7.550000 ;
      RECT 276.880000  55.895000 277.595000  56.065000 ;
      RECT 276.925000  55.835000 277.595000  55.895000 ;
      RECT 276.925000  56.065000 277.595000  56.345000 ;
      RECT 276.970000  84.275000 277.140000  87.055000 ;
      RECT 276.985000  56.700000 277.155000  57.680000 ;
      RECT 276.985000  58.805000 277.595000  60.665000 ;
      RECT 276.990000 223.695000 277.840000 225.350000 ;
      RECT 276.990000 229.255000 277.840000 232.355000 ;
      RECT 276.990000 240.705000 277.840000 243.640000 ;
      RECT 277.000000  37.870000 277.435000  40.870000 ;
      RECT 277.070000  12.950000 277.740000  13.120000 ;
      RECT 277.115000  55.495000 277.645000  55.665000 ;
      RECT 277.195000   5.390000 277.365000   6.700000 ;
      RECT 277.195000 200.085000 277.865000 200.255000 ;
      RECT 277.195000 216.235000 277.865000 216.405000 ;
      RECT 277.240000  61.675000 277.410000  63.495000 ;
      RECT 277.240000  64.405000 277.410000  67.115000 ;
      RECT 277.260000  13.120000 277.790000  13.320000 ;
      RECT 277.265000  40.870000 277.435000  44.425000 ;
      RECT 277.265000  47.855000 277.435000  48.465000 ;
      RECT 277.325000  56.345000 277.595000  58.805000 ;
      RECT 277.330000 225.650000 277.500000 226.630000 ;
      RECT 277.330000 234.980000 277.500000 235.960000 ;
      RECT 277.330000 237.100000 277.500000 238.080000 ;
      RECT 277.360000  68.255000 277.530000  73.355000 ;
      RECT 277.360000  74.400000 277.530000  78.155000 ;
      RECT 277.395000  14.170000 277.565000  18.920000 ;
      RECT 277.445000  19.870000 277.615000  22.580000 ;
      RECT 277.445000  23.850000 277.615000  26.560000 ;
      RECT 277.475000  54.555000 277.645000  55.495000 ;
      RECT 277.520000  84.215000 277.690000  86.925000 ;
      RECT 277.545000   7.010000 278.075000   7.180000 ;
      RECT 277.545000   8.900000 278.075000   9.070000 ;
      RECT 277.620000  37.335000 279.885000  37.505000 ;
      RECT 277.620000  37.505000 277.790000  39.510000 ;
      RECT 277.665000  42.510000 278.200000  43.085000 ;
      RECT 277.725000   5.690000 277.895000   7.010000 ;
      RECT 277.725000   7.180000 277.895000   8.900000 ;
      RECT 277.725000   9.070000 277.895000  12.470000 ;
      RECT 277.730000  43.405000 277.935000  44.415000 ;
      RECT 277.730000  44.415000 277.900000  46.335000 ;
      RECT 277.730000  46.335000 278.260000  46.505000 ;
      RECT 277.730000  46.505000 277.900000  48.105000 ;
      RECT 277.730000  48.105000 278.485000  48.275000 ;
      RECT 277.765000  56.670000 277.935000  60.405000 ;
      RECT 277.820000  74.405000 278.950000  74.575000 ;
      RECT 277.825000  61.675000 277.995000  62.955000 ;
      RECT 277.825000  62.955000 278.805000  63.285000 ;
      RECT 277.825000  63.905000 278.805000  67.115000 ;
      RECT 277.825000  67.115000 277.995000  67.415000 ;
      RECT 277.885000  87.275000 279.915000  87.445000 ;
      RECT 277.900000  74.575000 278.070000  75.690000 ;
      RECT 277.925000  41.635000 278.095000  42.030000 ;
      RECT 277.925000  42.030000 278.955000  42.200000 ;
      RECT 277.925000  42.200000 278.095000  42.305000 ;
      RECT 277.945000  87.445000 279.855000  87.455000 ;
      RECT 278.060000  69.905000 278.590000  70.075000 ;
      RECT 278.060000  77.080000 278.590000  77.250000 ;
      RECT 278.070000  12.950000 279.100000  13.150000 ;
      RECT 278.070000  13.150000 278.600000  13.320000 ;
      RECT 278.070000  44.520000 278.275000  45.300000 ;
      RECT 278.070000  54.385000 278.240000  55.575000 ;
      RECT 278.095000   7.380000 278.625000   7.550000 ;
      RECT 278.105000  43.405000 278.395000  44.415000 ;
      RECT 278.105000  44.415000 278.275000  44.520000 ;
      RECT 278.110000  37.840000 282.350000  38.010000 ;
      RECT 278.110000  38.010000 278.280000  41.290000 ;
      RECT 278.110000  41.290000 278.855000  41.460000 ;
      RECT 278.150000 113.195000 278.820000 113.525000 ;
      RECT 278.175000  29.500000 278.350000  30.030000 ;
      RECT 278.180000  30.030000 278.350000  30.500000 ;
      RECT 278.205000  32.095000 278.375000  33.375000 ;
      RECT 278.240000  68.605000 278.410000  69.905000 ;
      RECT 278.240000  70.075000 278.410000  73.815000 ;
      RECT 278.240000  74.765000 278.410000  77.080000 ;
      RECT 278.240000  77.250000 278.410000  77.475000 ;
      RECT 278.255000  41.460000 278.785000  41.530000 ;
      RECT 278.270000 224.125000 288.270000 226.460000 ;
      RECT 278.270000 229.425000 288.270000 232.185000 ;
      RECT 278.270000 235.150000 288.270000 237.910000 ;
      RECT 278.270000 240.875000 288.270000 243.210000 ;
      RECT 278.275000   5.690000 278.445000   7.380000 ;
      RECT 278.275000   7.550000 278.445000  12.470000 ;
      RECT 278.275000  14.170000 278.445000  18.920000 ;
      RECT 278.275000  81.955000 278.600000  83.800000 ;
      RECT 278.275000  83.800000 278.865000  83.970000 ;
      RECT 278.295000 199.300000 278.825000 200.255000 ;
      RECT 278.295000 200.495000 278.825000 215.995000 ;
      RECT 278.345000  56.690000 278.515000  60.405000 ;
      RECT 278.430000  79.315000 278.995000  81.675000 ;
      RECT 278.445000  42.400000 278.975000  42.570000 ;
      RECT 278.485000  44.585000 278.975000  44.740000 ;
      RECT 278.485000  44.740000 278.735000  45.375000 ;
      RECT 278.485000  45.375000 278.975000  45.665000 ;
      RECT 278.535000  13.660000 280.865000  13.740000 ;
      RECT 278.565000  42.570000 278.975000  44.585000 ;
      RECT 278.595000  31.870000 281.305000  32.040000 ;
      RECT 278.595000  32.650000 281.305000  32.820000 ;
      RECT 278.595000  33.430000 281.305000  33.600000 ;
      RECT 278.600000  85.230000 279.130000  85.400000 ;
      RECT 278.615000   7.010000 279.145000   7.040000 ;
      RECT 278.615000   7.040000 279.285000   7.210000 ;
      RECT 278.615000  34.015000 281.615000  34.325000 ;
      RECT 278.635000  61.675000 278.805000  62.725000 ;
      RECT 278.685000  32.605000 279.325000  32.650000 ;
      RECT 278.685000  32.820000 279.325000  32.865000 ;
      RECT 278.685000  45.665000 278.975000  48.085000 ;
      RECT 278.700000  30.555000 281.610000  30.725000 ;
      RECT 278.725000  19.870000 278.895000  22.580000 ;
      RECT 278.725000  23.850000 278.895000  26.560000 ;
      RECT 278.770000  81.675000 278.995000  83.310000 ;
      RECT 278.770000  83.310000 279.300000  83.480000 ;
      RECT 278.780000  74.575000 278.950000  75.690000 ;
      RECT 278.800000  84.215000 278.970000  85.230000 ;
      RECT 278.800000  85.400000 278.970000  86.925000 ;
      RECT 278.805000   5.390000 278.975000   6.700000 ;
      RECT 278.900000  29.275000 281.610000  29.445000 ;
      RECT 278.905000  45.000000 279.435000  45.170000 ;
      RECT 278.905000  61.175000 279.415000  61.505000 ;
      RECT 278.905000  67.585000 279.415000  67.915000 ;
      RECT 278.950000  22.750000 284.010000  23.680000 ;
      RECT 278.970000   3.465000 279.140000   4.740000 ;
      RECT 278.975000  11.320000 279.505000  11.490000 ;
      RECT 278.975000  61.505000 279.345000  67.585000 ;
      RECT 278.990000  38.180000 279.295000  40.890000 ;
      RECT 279.020000  87.870000 287.225000  87.885000 ;
      RECT 279.120000  68.255000 279.290000  73.355000 ;
      RECT 279.120000  74.400000 279.290000  78.155000 ;
      RECT 279.125000  40.890000 279.295000  41.580000 ;
      RECT 279.125000  41.580000 279.340000  41.635000 ;
      RECT 279.125000  41.635000 279.375000  42.305000 ;
      RECT 279.145000  43.405000 279.340000  44.415000 ;
      RECT 279.145000  45.170000 279.315000  48.085000 ;
      RECT 279.155000   7.720000 279.325000  11.320000 ;
      RECT 279.155000  11.490000 279.325000  12.470000 ;
      RECT 279.155000  14.170000 279.325000  18.920000 ;
      RECT 279.170000  42.305000 279.340000  43.405000 ;
      RECT 279.245000  79.265000 282.145000  79.435000 ;
      RECT 279.245000  80.045000 281.955000  80.215000 ;
      RECT 279.245000  80.925000 281.955000  80.930000 ;
      RECT 279.245000  80.930000 282.145000  81.095000 ;
      RECT 279.245000  81.805000 281.955000  81.975000 ;
      RECT 279.255000 200.085000 279.925000 200.255000 ;
      RECT 279.255000 216.235000 279.925000 216.405000 ;
      RECT 279.260000   6.510000 279.790000   6.680000 ;
      RECT 279.285000   5.680000 279.455000   6.510000 ;
      RECT 279.285000  53.600000 295.115000  54.780000 ;
      RECT 279.285000  54.780000 325.845000  55.295000 ;
      RECT 279.285000  55.295000 294.515000  56.185000 ;
      RECT 279.285000  56.185000 294.590000  56.715000 ;
      RECT 279.285000  56.715000 294.515000  58.725000 ;
      RECT 279.285000  58.725000 294.625000  59.255000 ;
      RECT 279.285000  59.255000 294.515000  60.605000 ;
      RECT 279.310000   2.995000 279.480000   4.160000 ;
      RECT 279.310000   4.500000 279.480000   5.170000 ;
      RECT 279.360000  81.775000 280.620000  81.805000 ;
      RECT 279.370000  12.900000 279.900000  12.950000 ;
      RECT 279.370000  12.950000 281.675000  13.070000 ;
      RECT 279.380000  13.070000 281.675000  13.120000 ;
      RECT 279.465000  41.290000 280.135000  41.460000 ;
      RECT 279.475000  82.625000 282.125000  83.565000 ;
      RECT 279.515000  61.675000 279.685000  67.415000 ;
      RECT 279.545000  41.460000 280.040000  42.030000 ;
      RECT 279.545000  42.030000 280.075000  42.200000 ;
      RECT 279.545000  74.405000 280.555000  74.575000 ;
      RECT 279.605000  19.870000 279.775000  22.580000 ;
      RECT 279.605000  23.850000 279.775000  26.560000 ;
      RECT 279.605000  43.405000 280.255000  44.415000 ;
      RECT 279.605000  44.415000 279.775000  46.335000 ;
      RECT 279.605000  46.335000 280.135000  46.505000 ;
      RECT 279.605000  46.505000 279.775000  48.085000 ;
      RECT 279.640000  69.905000 280.170000  70.075000 ;
      RECT 279.660000  74.575000 279.830000  75.690000 ;
      RECT 279.680000   3.295000 280.690000   3.465000 ;
      RECT 279.680000   3.755000 280.690000   3.925000 ;
      RECT 279.680000   4.215000 280.690000   4.385000 ;
      RECT 279.785000  61.175000 280.295000  61.505000 ;
      RECT 279.785000  67.585000 280.385000  67.685000 ;
      RECT 279.785000  67.685000 280.295000  67.915000 ;
      RECT 279.810000  31.820000 280.450000  31.870000 ;
      RECT 279.810000  32.040000 280.450000  32.080000 ;
      RECT 279.810000  33.385000 280.450000  33.430000 ;
      RECT 279.810000  33.600000 280.450000  33.645000 ;
      RECT 279.820000  77.080000 280.350000  77.250000 ;
      RECT 279.855000  61.505000 280.225000  67.515000 ;
      RECT 279.855000  67.515000 280.385000  67.585000 ;
      RECT 279.870000  38.180000 280.040000  41.290000 ;
      RECT 279.945000  47.855000 280.115000  48.465000 ;
      RECT 280.000000  68.605000 280.170000  69.905000 ;
      RECT 280.000000  70.075000 280.170000  73.815000 ;
      RECT 280.000000  74.765000 280.170000  77.080000 ;
      RECT 280.000000  77.250000 280.170000  77.475000 ;
      RECT 280.035000   7.200000 283.975000   7.370000 ;
      RECT 280.035000   7.370000 280.205000  12.650000 ;
      RECT 280.035000  14.170000 280.205000  18.920000 ;
      RECT 280.080000  84.215000 280.250000  86.925000 ;
      RECT 280.085000  42.475000 282.745000  42.645000 ;
      RECT 280.085000  42.645000 280.255000  43.405000 ;
      RECT 280.095000  37.335000 282.125000  37.505000 ;
      RECT 280.225000 113.910000 283.225000 164.900000 ;
      RECT 280.305000  41.360000 280.835000  41.530000 ;
      RECT 280.340000  74.575000 280.510000  75.690000 ;
      RECT 280.355000 199.685000 280.885000 200.255000 ;
      RECT 280.355000 200.495000 280.885000 215.995000 ;
      RECT 280.395000  61.675000 281.115000  62.725000 ;
      RECT 280.395000  62.955000 281.115000  63.285000 ;
      RECT 280.395000  63.905000 281.115000  64.235000 ;
      RECT 280.395000  64.235000 280.565000  67.115000 ;
      RECT 280.425000  43.095000 280.955000  43.265000 ;
      RECT 280.425000  43.265000 280.595000  48.390000 ;
      RECT 280.445000  87.275000 282.475000  87.445000 ;
      RECT 280.485000  19.870000 280.655000  22.580000 ;
      RECT 280.485000  23.850000 280.655000  26.560000 ;
      RECT 280.485000  41.530000 280.655000  42.305000 ;
      RECT 280.505000  87.445000 282.415000  87.455000 ;
      RECT 280.580000  68.255000 280.750000  73.625000 ;
      RECT 280.750000  38.180000 281.010000  41.160000 ;
      RECT 280.765000  44.180000 282.585000  44.350000 ;
      RECT 280.765000  44.350000 280.955000  47.370000 ;
      RECT 280.765000  47.370000 281.295000  48.550000 ;
      RECT 280.765000  48.550000 283.655000  48.720000 ;
      RECT 280.880000  74.400000 281.050000  78.155000 ;
      RECT 280.915000   7.720000 281.085000  11.320000 ;
      RECT 280.915000  11.320000 281.445000  11.490000 ;
      RECT 280.915000  11.490000 281.085000  12.470000 ;
      RECT 280.915000  14.170000 281.085000  18.920000 ;
      RECT 280.935000  81.095000 282.145000  81.100000 ;
      RECT 280.945000  64.405000 281.115000  67.420000 ;
      RECT 281.090000   3.515000 281.260000   5.885000 ;
      RECT 281.125000  42.840000 281.295000  44.010000 ;
      RECT 281.125000  44.580000 281.295000  45.280000 ;
      RECT 281.125000  45.280000 281.655000  45.450000 ;
      RECT 281.125000  45.450000 281.295000  47.080000 ;
      RECT 281.160000  68.255000 281.330000  73.355000 ;
      RECT 281.185000  86.680000 281.715000  86.850000 ;
      RECT 281.210000  38.180000 281.470000  41.160000 ;
      RECT 281.285000  61.175000 281.795000  61.505000 ;
      RECT 281.285000  67.585000 281.795000  67.915000 ;
      RECT 281.315000 200.085000 281.985000 200.255000 ;
      RECT 281.315000 216.235000 281.985000 216.405000 ;
      RECT 281.355000  61.505000 281.725000  67.585000 ;
      RECT 281.360000  84.215000 281.530000  86.680000 ;
      RECT 281.360000  86.850000 281.530000  86.925000 ;
      RECT 281.365000  19.870000 281.535000  22.580000 ;
      RECT 281.365000  23.850000 281.535000  26.560000 ;
      RECT 281.395000  42.470000 282.745000  42.475000 ;
      RECT 281.405000  74.405000 282.415000  74.575000 ;
      RECT 281.450000   3.295000 284.500000   3.465000 ;
      RECT 281.450000   4.175000 284.160000   4.345000 ;
      RECT 281.450000   5.055000 284.500000   5.225000 ;
      RECT 281.450000   5.935000 284.160000   6.105000 ;
      RECT 281.465000  14.170000 281.635000  18.920000 ;
      RECT 281.465000  74.000000 282.355000  74.405000 ;
      RECT 281.470000   2.715000 289.335000   2.885000 ;
      RECT 281.505000  13.490000 282.175000  13.660000 ;
      RECT 281.555000  42.840000 281.725000  44.180000 ;
      RECT 281.605000  46.335000 282.135000  47.370000 ;
      RECT 281.605000  47.370000 282.475000  48.380000 ;
      RECT 281.700000  77.080000 282.230000  77.250000 ;
      RECT 281.760000  74.765000 281.930000  77.080000 ;
      RECT 281.760000  77.250000 281.930000  77.475000 ;
      RECT 281.795000   7.370000 281.965000  12.650000 ;
      RECT 281.895000  61.675000 282.065000  66.145000 ;
      RECT 281.985000  42.840000 282.155000  44.010000 ;
      RECT 282.040000  68.605000 282.210000  69.905000 ;
      RECT 282.040000  69.905000 282.570000  70.075000 ;
      RECT 282.040000  70.075000 282.210000  73.355000 ;
      RECT 282.145000  61.175000 282.675000  61.345000 ;
      RECT 282.165000  61.345000 282.675000  61.505000 ;
      RECT 282.165000  67.585000 282.675000  67.915000 ;
      RECT 282.180000  38.010000 282.350000  41.360000 ;
      RECT 282.180000  41.360000 282.710000  41.530000 ;
      RECT 282.235000  61.505000 282.605000  67.585000 ;
      RECT 282.245000  19.870000 282.415000  22.580000 ;
      RECT 282.245000  23.850000 282.415000  26.560000 ;
      RECT 282.305000  44.580000 282.475000  45.760000 ;
      RECT 282.305000  45.760000 284.835000  45.930000 ;
      RECT 282.305000  45.930000 282.475000  47.080000 ;
      RECT 282.345000   7.720000 282.515000   9.730000 ;
      RECT 282.345000   9.730000 282.990000   9.900000 ;
      RECT 282.345000   9.900000 282.515000  18.920000 ;
      RECT 282.415000  42.840000 282.585000  44.180000 ;
      RECT 282.415000 199.300000 282.945000 200.255000 ;
      RECT 282.415000 200.495000 282.945000 215.995000 ;
      RECT 282.510000  80.270000 282.710000  82.645000 ;
      RECT 282.510000  82.645000 286.870000  82.845000 ;
      RECT 282.525000  79.260000 282.695000  79.990000 ;
      RECT 282.640000  74.400000 282.810000  78.155000 ;
      RECT 282.640000  84.215000 282.810000  86.925000 ;
      RECT 282.760000  37.870000 282.930000  40.870000 ;
      RECT 282.825000  46.165000 283.155000  47.015000 ;
      RECT 282.825000  83.800000 283.415000  83.970000 ;
      RECT 282.845000  42.840000 283.015000  44.010000 ;
      RECT 282.845000  61.675000 283.015000  62.725000 ;
      RECT 282.845000  62.955000 283.015000  63.285000 ;
      RECT 282.845000  63.905000 283.015000  64.235000 ;
      RECT 282.845000  64.405000 283.015000  67.115000 ;
      RECT 282.865000  11.320000 283.395000  11.490000 ;
      RECT 282.905000  47.015000 283.075000  47.625000 ;
      RECT 282.920000  68.255000 283.090000  73.355000 ;
      RECT 282.980000  45.280000 283.655000  45.450000 ;
      RECT 283.080000  83.970000 283.415000  87.015000 ;
      RECT 283.080000  87.015000 285.000000  87.210000 ;
      RECT 283.100000  42.470000 284.450000  42.640000 ;
      RECT 283.100000  42.640000 284.350000  42.670000 ;
      RECT 283.125000  19.870000 283.295000  22.580000 ;
      RECT 283.125000  23.850000 283.295000  26.560000 ;
      RECT 283.185000  61.175000 283.695000  61.505000 ;
      RECT 283.185000  67.585000 283.695000  67.915000 ;
      RECT 283.190000  74.765000 283.360000  77.645000 ;
      RECT 283.190000  77.645000 286.880000  77.815000 ;
      RECT 283.225000   7.720000 283.395000  11.320000 ;
      RECT 283.225000  11.490000 283.395000  12.470000 ;
      RECT 283.225000  14.170000 283.395000  18.920000 ;
      RECT 283.255000  61.505000 283.625000  67.585000 ;
      RECT 283.275000  42.840000 283.445000  44.180000 ;
      RECT 283.275000  44.180000 284.835000  44.350000 ;
      RECT 283.375000 200.085000 284.045000 200.255000 ;
      RECT 283.375000 216.235000 284.045000 216.405000 ;
      RECT 283.405000  79.755000 283.575000  82.465000 ;
      RECT 283.485000  44.580000 283.655000  45.280000 ;
      RECT 283.485000  45.450000 283.655000  45.590000 ;
      RECT 283.485000  46.100000 283.655000  48.550000 ;
      RECT 283.620000  69.905000 284.150000  70.075000 ;
      RECT 283.630000  82.845000 286.870000  82.855000 ;
      RECT 283.645000  83.815000 284.045000  86.825000 ;
      RECT 283.705000  42.840000 283.875000  44.010000 ;
      RECT 283.705000  83.755000 283.875000  83.815000 ;
      RECT 283.775000   7.720000 284.005000   8.950000 ;
      RECT 283.775000  11.700000 284.005000  12.710000 ;
      RECT 283.795000  61.675000 283.965000  66.145000 ;
      RECT 283.800000  68.605000 283.970000  69.905000 ;
      RECT 283.800000  70.075000 283.970000  74.765000 ;
      RECT 283.800000  74.765000 284.240000  74.935000 ;
      RECT 283.805000   7.370000 283.975000   7.720000 ;
      RECT 283.805000   8.950000 283.975000  11.700000 ;
      RECT 283.805000  12.710000 283.975000  12.740000 ;
      RECT 283.805000  13.900000 283.975000  18.900000 ;
      RECT 283.930000  83.365000 284.930000  83.535000 ;
      RECT 283.975000  66.375000 284.505000  66.545000 ;
      RECT 283.990000  83.535000 284.870000  83.625000 ;
      RECT 284.000000  87.210000 285.000000  87.215000 ;
      RECT 284.005000  19.870000 284.175000  22.580000 ;
      RECT 284.005000  23.850000 284.175000  26.560000 ;
      RECT 284.065000  61.175000 284.575000  61.505000 ;
      RECT 284.065000  67.585000 284.575000  67.915000 ;
      RECT 284.070000  74.935000 284.240000  77.475000 ;
      RECT 284.105000  37.765000 284.275000  40.845000 ;
      RECT 284.135000  42.840000 284.305000  44.180000 ;
      RECT 284.135000  61.505000 284.505000  66.375000 ;
      RECT 284.135000  66.545000 284.505000  67.585000 ;
      RECT 284.145000 186.390000 288.165000 187.365000 ;
      RECT 284.145000 192.960000 288.165000 193.710000 ;
      RECT 284.155000  73.865000 285.505000  74.035000 ;
      RECT 284.205000  73.600000 285.455000  73.865000 ;
      RECT 284.285000  79.755000 284.460000  80.540000 ;
      RECT 284.285000  80.540000 284.455000  82.465000 ;
      RECT 284.290000  79.525000 284.460000  79.755000 ;
      RECT 284.305000  46.335000 284.835000  46.505000 ;
      RECT 284.330000   3.465000 284.500000   5.055000 ;
      RECT 284.430000  41.265000 285.395000  41.435000 ;
      RECT 284.430000  41.435000 284.740000  42.130000 ;
      RECT 284.430000  42.130000 284.960000  42.300000 ;
      RECT 284.475000 199.685000 285.005000 200.255000 ;
      RECT 284.475000 200.495000 285.005000 215.995000 ;
      RECT 284.565000  42.840000 284.735000  44.010000 ;
      RECT 284.570000  38.155000 284.855000  40.865000 ;
      RECT 284.570000  40.865000 284.740000  41.095000 ;
      RECT 284.590000  19.520000 285.170000  24.735000 ;
      RECT 284.590000  24.735000 287.175000  24.905000 ;
      RECT 284.590000  24.905000 285.170000  25.750000 ;
      RECT 284.590000  25.750000 284.775000  26.920000 ;
      RECT 284.610000 113.195000 285.280000 113.525000 ;
      RECT 284.665000  44.350000 284.835000  45.760000 ;
      RECT 284.665000  46.100000 284.835000  46.335000 ;
      RECT 284.665000  46.505000 284.835000  48.380000 ;
      RECT 284.680000  68.255000 284.850000  73.355000 ;
      RECT 284.735000 113.910000 287.735000 164.900000 ;
      RECT 284.745000  61.675000 284.915000  62.725000 ;
      RECT 284.745000  62.955000 284.915000  63.285000 ;
      RECT 284.745000  63.905000 284.915000  64.235000 ;
      RECT 284.745000  64.405000 284.915000  67.420000 ;
      RECT 284.760000   2.885000 285.170000  19.350000 ;
      RECT 284.910000  37.335000 287.165000  37.505000 ;
      RECT 284.910000  41.085000 285.580000  41.255000 ;
      RECT 284.910000  41.255000 285.395000  41.265000 ;
      RECT 284.910000  41.760000 285.440000  41.930000 ;
      RECT 284.950000  74.765000 285.120000  77.645000 ;
      RECT 284.985000  83.755000 285.155000  85.105000 ;
      RECT 285.025000  37.505000 287.165000  37.595000 ;
      RECT 285.025000  37.595000 285.395000  41.085000 ;
      RECT 285.025000  43.110000 285.555000  43.280000 ;
      RECT 285.055000  85.740000 285.225000  86.825000 ;
      RECT 285.130000  41.930000 285.440000  43.110000 ;
      RECT 285.165000  79.755000 285.335000  82.465000 ;
      RECT 285.195000  69.905000 285.730000  70.075000 ;
      RECT 285.245000  43.280000 285.415000  48.390000 ;
      RECT 285.295000  61.675000 285.465000  67.420000 ;
      RECT 285.305000  74.405000 286.655000  74.575000 ;
      RECT 285.435000 200.085000 286.105000 200.255000 ;
      RECT 285.435000 216.235000 286.105000 216.405000 ;
      RECT 285.470000  77.080000 286.000000  77.250000 ;
      RECT 285.490000  74.575000 285.660000  75.690000 ;
      RECT 285.520000   3.395000 286.990000   3.655000 ;
      RECT 285.520000  23.765000 285.940000  24.295000 ;
      RECT 285.560000  68.605000 285.730000  69.905000 ;
      RECT 285.560000  70.075000 285.730000  73.355000 ;
      RECT 285.565000  37.765000 285.735000  40.865000 ;
      RECT 285.565000  61.175000 286.075000  61.505000 ;
      RECT 285.565000  67.585000 286.075000  67.915000 ;
      RECT 285.610000  41.445000 286.075000  41.615000 ;
      RECT 285.610000  41.615000 285.780000  42.520000 ;
      RECT 285.610000  42.520000 285.895000  42.690000 ;
      RECT 285.635000  61.505000 286.005000  67.585000 ;
      RECT 285.655000  83.765000 285.825000  86.475000 ;
      RECT 285.725000  42.690000 285.895000  43.615000 ;
      RECT 285.830000  74.765000 286.000000  77.080000 ;
      RECT 285.830000  77.250000 286.000000  77.475000 ;
      RECT 285.880000  83.375000 287.160000  83.545000 ;
      RECT 285.905000  40.395000 286.615000  40.865000 ;
      RECT 285.905000  40.865000 286.075000  41.445000 ;
      RECT 285.950000  41.785000 286.570000  42.115000 ;
      RECT 286.045000  79.755000 286.220000  80.540000 ;
      RECT 286.045000  80.540000 286.215000  82.465000 ;
      RECT 286.050000  79.525000 286.220000  79.755000 ;
      RECT 286.170000   3.825000 286.340000  23.710000 ;
      RECT 286.170000  74.575000 286.340000  75.690000 ;
      RECT 286.175000  48.350000 287.945000  48.385000 ;
      RECT 286.175000  48.385000 287.860000  48.520000 ;
      RECT 286.175000  61.675000 286.345000  62.725000 ;
      RECT 286.175000  62.955000 286.345000  63.285000 ;
      RECT 286.175000  63.905000 286.345000  64.235000 ;
      RECT 286.175000  64.405000 286.345000  67.115000 ;
      RECT 286.215000  45.290000 286.385000  48.000000 ;
      RECT 286.245000  41.360000 287.165000  41.530000 ;
      RECT 286.245000  41.530000 286.570000  41.785000 ;
      RECT 286.335000  48.215000 287.945000  48.350000 ;
      RECT 286.435000  83.765000 286.605000  86.475000 ;
      RECT 286.440000  68.255000 286.610000  73.355000 ;
      RECT 286.445000  38.155000 286.615000  40.395000 ;
      RECT 286.445000  61.175000 286.955000  61.505000 ;
      RECT 286.445000  67.585000 286.955000  67.915000 ;
      RECT 286.515000  61.505000 286.885000  67.585000 ;
      RECT 286.535000 199.300000 287.065000 200.255000 ;
      RECT 286.535000 200.495000 287.065000 215.995000 ;
      RECT 286.605000  42.605000 286.775000  44.570000 ;
      RECT 286.605000  44.570000 287.720000  44.740000 ;
      RECT 286.605000  44.740000 287.240000  44.800000 ;
      RECT 286.610000  23.765000 286.990000  24.275000 ;
      RECT 286.610000  24.275000 286.780000  24.295000 ;
      RECT 286.620000  45.030000 287.165000  45.200000 ;
      RECT 286.710000  74.765000 286.880000  77.645000 ;
      RECT 286.785000  37.595000 287.165000  38.615000 ;
      RECT 286.825000  42.000000 287.495000  42.170000 ;
      RECT 286.890000  88.725000 287.445000  88.895000 ;
      RECT 286.890000  89.715000 287.445000  89.885000 ;
      RECT 286.895000  42.170000 287.425000  42.300000 ;
      RECT 286.925000  79.755000 287.095000  82.465000 ;
      RECT 286.995000  40.195000 287.165000  41.360000 ;
      RECT 286.995000  45.000000 287.165000  45.030000 ;
      RECT 286.995000  45.200000 287.165000  48.000000 ;
      RECT 287.005000  24.905000 287.175000  36.235000 ;
      RECT 287.005000  36.235000 289.335000  36.405000 ;
      RECT 287.020000  68.255000 287.190000  73.625000 ;
      RECT 287.055000  61.675000 287.225000  67.415000 ;
      RECT 287.095000  38.970000 287.945000  39.720000 ;
      RECT 287.125000  42.505000 287.655000  42.675000 ;
      RECT 287.170000 113.195000 287.840000 113.525000 ;
      RECT 287.215000  83.765000 287.385000  86.475000 ;
      RECT 287.275000  88.610000 287.445000  88.725000 ;
      RECT 287.275000  88.895000 287.445000  88.940000 ;
      RECT 287.275000  89.650000 287.445000  89.715000 ;
      RECT 287.275000  89.885000 287.445000  89.980000 ;
      RECT 287.290000  74.400000 287.460000  78.155000 ;
      RECT 287.325000  61.175000 287.835000  61.505000 ;
      RECT 287.325000  67.585000 287.835000  67.915000 ;
      RECT 287.335000  37.765000 287.945000  38.970000 ;
      RECT 287.335000  39.720000 287.945000  40.865000 ;
      RECT 287.345000  88.205000 289.565000  88.425000 ;
      RECT 287.395000  61.505000 287.765000  67.585000 ;
      RECT 287.485000  42.675000 287.655000  43.615000 ;
      RECT 287.495000 200.085000 288.165000 200.255000 ;
      RECT 287.495000 216.235000 288.165000 216.405000 ;
      RECT 287.525000   3.295000 288.535000   3.465000 ;
      RECT 287.525000   3.755000 288.535000   3.925000 ;
      RECT 287.525000   4.215000 288.535000   4.385000 ;
      RECT 287.525000   4.675000 288.535000   4.845000 ;
      RECT 287.525000   5.135000 288.535000   5.305000 ;
      RECT 287.525000   5.595000 288.535000   5.765000 ;
      RECT 287.525000   6.055000 288.535000   6.225000 ;
      RECT 287.525000   6.515000 288.535000   6.685000 ;
      RECT 287.525000   6.975000 288.535000   7.145000 ;
      RECT 287.525000   7.345000 288.535000   7.605000 ;
      RECT 287.525000   7.985000 288.535000   8.155000 ;
      RECT 287.525000   8.485000 288.535000   8.685000 ;
      RECT 287.525000   9.065000 288.535000   9.235000 ;
      RECT 287.525000   9.595000 288.535000   9.765000 ;
      RECT 287.525000  10.125000 288.535000  10.295000 ;
      RECT 287.525000  13.745000 288.535000  13.915000 ;
      RECT 287.525000  15.025000 288.535000  15.195000 ;
      RECT 287.525000  16.305000 288.535000  16.475000 ;
      RECT 287.525000  16.855000 288.925000  17.025000 ;
      RECT 287.525000  18.135000 288.535000  18.305000 ;
      RECT 287.525000  19.415000 288.535000  19.585000 ;
      RECT 287.525000  19.965000 288.925000  20.135000 ;
      RECT 287.525000  21.245000 288.535000  21.415000 ;
      RECT 287.525000  22.525000 288.535000  22.695000 ;
      RECT 287.525000  23.075000 288.535000  23.245000 ;
      RECT 287.525000  23.245000 288.115000  24.055000 ;
      RECT 287.525000  24.355000 288.535000  24.560000 ;
      RECT 287.525000  24.560000 288.185000  24.755000 ;
      RECT 287.525000  25.435000 288.535000  25.605000 ;
      RECT 287.525000  26.515000 288.535000  26.685000 ;
      RECT 287.525000  27.595000 288.535000  27.765000 ;
      RECT 287.525000  28.675000 288.535000  28.845000 ;
      RECT 287.525000  29.755000 288.535000  29.925000 ;
      RECT 287.525000  30.835000 288.535000  31.005000 ;
      RECT 287.525000  31.385000 288.535000  31.555000 ;
      RECT 287.525000  32.465000 288.535000  32.635000 ;
      RECT 287.525000  33.545000 288.535000  33.715000 ;
      RECT 287.525000  34.095000 288.535000  34.265000 ;
      RECT 287.525000  34.875000 288.535000  35.045000 ;
      RECT 287.525000  35.655000 288.535000  35.825000 ;
      RECT 287.545000  10.875000 289.335000  12.745000 ;
      RECT 287.545000  13.165000 289.335000  13.335000 ;
      RECT 287.550000  10.830000 289.335000  10.875000 ;
      RECT 287.565000  82.140000 288.530000  82.810000 ;
      RECT 287.565000  82.810000 287.765000  86.995000 ;
      RECT 287.580000  86.995000 287.750000  87.340000 ;
      RECT 287.625000  78.890000 288.485000  79.420000 ;
      RECT 287.625000  79.420000 288.155000  79.960000 ;
      RECT 287.775000  45.290000 287.945000  48.000000 ;
      RECT 287.935000  61.675000 288.105000  62.725000 ;
      RECT 287.935000  62.955000 288.800000  63.285000 ;
      RECT 287.935000  63.905000 288.800000  63.975000 ;
      RECT 287.935000  63.975000 289.375000  67.115000 ;
      RECT 287.945000  80.595000 288.115000  81.180000 ;
      RECT 287.945000  81.435000 288.115000  81.965000 ;
      RECT 287.945000  83.000000 288.115000  84.335000 ;
      RECT 287.970000   9.765000 288.500000   9.770000 ;
      RECT 288.170000  80.160000 290.320000  80.405000 ;
      RECT 288.285000  32.080000 288.925000  32.250000 ;
      RECT 288.340000  23.630000 288.925000  24.160000 ;
      RECT 288.355000  86.930000 290.320000  87.285000 ;
      RECT 288.395000  25.065000 288.925000  25.235000 ;
      RECT 288.395000  27.225000 288.925000  27.395000 ;
      RECT 288.405000  79.610000 290.400000  79.945000 ;
      RECT 288.410000  84.925000 288.580000  85.935000 ;
      RECT 288.415000 199.685000 288.945000 200.255000 ;
      RECT 288.525000  68.505000 289.375000  76.025000 ;
      RECT 288.525000  76.025000 290.955000  76.195000 ;
      RECT 288.525000  76.195000 289.320000  76.345000 ;
      RECT 288.560000  84.535000 289.230000  84.705000 ;
      RECT 288.560000  84.705000 289.090000  84.735000 ;
      RECT 288.595000 200.495000 289.125000 215.995000 ;
      RECT 288.630000  61.675000 288.800000  62.955000 ;
      RECT 288.630000  67.115000 289.375000  68.505000 ;
      RECT 288.630000  76.345000 289.320000  77.785000 ;
      RECT 288.635000 186.220000 309.875000 187.450000 ;
      RECT 288.635000 187.450000 342.805000 187.620000 ;
      RECT 288.635000 187.620000 309.875000 189.190000 ;
      RECT 288.635000 189.190000 342.805000 189.360000 ;
      RECT 288.635000 189.360000 309.875000 190.930000 ;
      RECT 288.635000 190.930000 342.805000 191.100000 ;
      RECT 288.635000 191.100000 309.875000 191.955000 ;
      RECT 288.635000 191.955000 303.890000 194.500000 ;
      RECT 288.635000 194.500000 342.805000 194.595000 ;
      RECT 288.700000 223.695000 289.550000 225.350000 ;
      RECT 288.700000 229.255000 289.550000 232.355000 ;
      RECT 288.700000 240.705000 289.550000 243.640000 ;
      RECT 288.750000  80.615000 289.070000  81.925000 ;
      RECT 288.755000   3.520000 288.925000   6.000000 ;
      RECT 288.755000   6.280000 288.925000   6.915000 ;
      RECT 288.755000   6.915000 290.825000   7.085000 ;
      RECT 288.755000   7.085000 288.925000   7.380000 ;
      RECT 288.755000   7.910000 290.825000   8.080000 ;
      RECT 288.755000   8.080000 288.925000   8.660000 ;
      RECT 288.755000   8.870000 288.925000   9.225000 ;
      RECT 288.755000   9.225000 290.905000   9.450000 ;
      RECT 288.755000   9.450000 288.925000   9.540000 ;
      RECT 288.755000   9.820000 288.925000  10.570000 ;
      RECT 288.755000  13.970000 288.925000  14.970000 ;
      RECT 288.755000  15.250000 288.925000  16.855000 ;
      RECT 288.755000  17.195000 288.925000  18.080000 ;
      RECT 288.755000  18.360000 288.925000  19.965000 ;
      RECT 288.755000  20.305000 288.925000  21.190000 ;
      RECT 288.755000  21.755000 288.925000  23.460000 ;
      RECT 288.755000  24.160000 288.925000  24.300000 ;
      RECT 288.755000  24.580000 288.925000  25.065000 ;
      RECT 288.755000  25.235000 288.925000  26.460000 ;
      RECT 288.755000  26.740000 288.925000  27.225000 ;
      RECT 288.755000  27.395000 288.925000  28.620000 ;
      RECT 288.755000  28.900000 288.925000  30.780000 ;
      RECT 288.755000  31.610000 288.925000  32.080000 ;
      RECT 288.755000  32.250000 288.925000  32.410000 ;
      RECT 288.755000  32.690000 288.925000  33.490000 ;
      RECT 288.755000  34.320000 288.925000  35.600000 ;
      RECT 288.825000  80.595000 288.995000  80.615000 ;
      RECT 288.825000  83.000000 288.995000  84.010000 ;
      RECT 289.035000 216.180000 290.225000 216.405000 ;
      RECT 289.040000 225.650000 289.210000 226.630000 ;
      RECT 289.040000 234.980000 289.210000 235.960000 ;
      RECT 289.040000 237.100000 289.210000 238.080000 ;
      RECT 289.070000  87.870000 290.955000  87.885000 ;
      RECT 289.095000  78.830000 289.265000  79.420000 ;
      RECT 289.165000   2.885000 289.335000   6.745000 ;
      RECT 289.165000   7.255000 289.335000   7.740000 ;
      RECT 289.165000   8.250000 289.335000   8.815000 ;
      RECT 289.165000   8.815000 289.710000   8.985000 ;
      RECT 289.165000   8.985000 289.335000   8.995000 ;
      RECT 289.165000   9.700000 289.335000  10.830000 ;
      RECT 289.165000  13.335000 289.335000  36.235000 ;
      RECT 289.190000  84.925000 289.360000  85.030000 ;
      RECT 289.190000  85.030000 289.775000  85.200000 ;
      RECT 289.190000  85.200000 289.360000  85.935000 ;
      RECT 289.205000  37.870000 289.375000  42.475000 ;
      RECT 289.205000  43.510000 289.375000  44.400000 ;
      RECT 289.245000 113.910000 292.245000 164.900000 ;
      RECT 289.290000  82.140000 290.320000  82.810000 ;
      RECT 289.355000 200.085000 290.225000 200.255000 ;
      RECT 289.555000 200.255000 290.225000 216.180000 ;
      RECT 289.700000  83.090000 289.875000  83.945000 ;
      RECT 289.705000  83.000000 289.875000  83.090000 ;
      RECT 289.705000  83.945000 289.875000  84.010000 ;
      RECT 289.780000  87.885000 290.580000  91.465000 ;
      RECT 289.810000   9.640000 290.415000  10.050000 ;
      RECT 289.810000  10.050000 290.120000  10.585000 ;
      RECT 289.810000  10.585000 292.765000  10.895000 ;
      RECT 289.905000  80.405000 290.320000  82.140000 ;
      RECT 289.980000 224.125000 299.980000 226.460000 ;
      RECT 289.980000 229.425000 299.980000 232.185000 ;
      RECT 289.980000 235.150000 299.980000 237.910000 ;
      RECT 289.980000 240.875000 299.980000 243.210000 ;
      RECT 290.035000  46.500000 294.285000  46.990000 ;
      RECT 290.055000  82.810000 290.320000  86.930000 ;
      RECT 290.070000  78.225000 290.400000  79.610000 ;
      RECT 290.115000  46.990000 294.245000  47.125000 ;
      RECT 290.140000  60.605000 294.515000  62.780000 ;
      RECT 290.140000  62.780000 294.500000  63.070000 ;
      RECT 290.140000  74.525000 297.140000  75.535000 ;
      RECT 290.245000   2.815000 292.765000   2.985000 ;
      RECT 290.245000   2.985000 290.415000   6.745000 ;
      RECT 290.245000   7.255000 290.415000   7.740000 ;
      RECT 290.245000   8.250000 290.415000   8.885000 ;
      RECT 290.245000   8.885000 290.430000   8.995000 ;
      RECT 290.245000  13.265000 292.505000  13.435000 ;
      RECT 290.245000  13.435000 290.415000  25.915000 ;
      RECT 290.245000  25.915000 292.505000  26.085000 ;
      RECT 290.260000   8.995000 290.430000   9.055000 ;
      RECT 290.290000  10.245000 290.825000  10.415000 ;
      RECT 290.445000  34.640000 294.775000  34.845000 ;
      RECT 290.445000  34.845000 290.615000  41.465000 ;
      RECT 290.445000  41.465000 301.075000  41.635000 ;
      RECT 290.545000  28.410000 293.885000  28.765000 ;
      RECT 290.545000  28.765000 290.715000  31.785000 ;
      RECT 290.545000  31.785000 290.800000  31.995000 ;
      RECT 290.545000  31.995000 293.885000  32.165000 ;
      RECT 290.655000   3.520000 290.825000   6.000000 ;
      RECT 290.655000   6.280000 290.825000   6.915000 ;
      RECT 290.655000   7.085000 290.825000   7.380000 ;
      RECT 290.655000   8.080000 290.825000   8.990000 ;
      RECT 290.655000   9.745000 290.825000  10.245000 ;
      RECT 290.655000  13.970000 290.825000  14.445000 ;
      RECT 290.655000  14.445000 291.395000  14.615000 ;
      RECT 290.655000  14.615000 290.825000  14.970000 ;
      RECT 290.655000  15.250000 290.825000  16.855000 ;
      RECT 290.655000  16.855000 292.085000  17.025000 ;
      RECT 290.655000  17.195000 290.825000  18.080000 ;
      RECT 290.655000  18.360000 290.825000  19.965000 ;
      RECT 290.655000  19.965000 292.085000  20.135000 ;
      RECT 290.655000  20.305000 290.825000  21.190000 ;
      RECT 290.655000  21.470000 290.825000  23.460000 ;
      RECT 290.655000  23.630000 290.825000  23.970000 ;
      RECT 290.655000  23.970000 291.415000  24.140000 ;
      RECT 290.655000  24.140000 290.825000  24.300000 ;
      RECT 290.655000  24.580000 290.825000  25.065000 ;
      RECT 290.655000  25.065000 291.185000  25.235000 ;
      RECT 290.655000  25.235000 290.825000  25.380000 ;
      RECT 290.655000 200.495000 291.185000 215.995000 ;
      RECT 290.785000  76.195000 290.955000  87.700000 ;
      RECT 290.895000  35.155000 292.245000  35.325000 ;
      RECT 290.895000  36.235000 291.905000  36.405000 ;
      RECT 290.895000  37.315000 291.905000  37.485000 ;
      RECT 290.895000  37.865000 292.585000  38.035000 ;
      RECT 290.895000  38.645000 292.245000  38.815000 ;
      RECT 290.895000  39.425000 292.585000  39.595000 ;
      RECT 290.895000  40.205000 292.245000  40.375000 ;
      RECT 290.895000  40.985000 292.585000  41.155000 ;
      RECT 290.955000  29.380000 291.125000  29.755000 ;
      RECT 290.955000  29.755000 291.540000  29.925000 ;
      RECT 290.955000  29.925000 291.125000  31.380000 ;
      RECT 291.055000  13.665000 292.085000  13.915000 ;
      RECT 291.055000  16.305000 292.085000  16.475000 ;
      RECT 291.075000   3.295000 292.085000   3.465000 ;
      RECT 291.075000   3.755000 292.085000   3.925000 ;
      RECT 291.075000   4.215000 292.085000   4.385000 ;
      RECT 291.075000   4.675000 292.085000   4.845000 ;
      RECT 291.075000   5.135000 292.085000   5.305000 ;
      RECT 291.075000   5.595000 292.085000   5.765000 ;
      RECT 291.075000   6.055000 292.085000   6.225000 ;
      RECT 291.075000   6.515000 292.085000   6.685000 ;
      RECT 291.075000   6.975000 292.085000   7.145000 ;
      RECT 291.075000   7.435000 292.085000   7.605000 ;
      RECT 291.075000   7.985000 292.085000   8.180000 ;
      RECT 291.075000   8.485000 292.085000   8.685000 ;
      RECT 291.075000   9.045000 292.085000   9.215000 ;
      RECT 291.075000   9.575000 292.085000   9.745000 ;
      RECT 291.075000  10.105000 292.085000  10.275000 ;
      RECT 291.075000  15.025000 292.150000  15.195000 ;
      RECT 291.075000  18.135000 292.085000  18.305000 ;
      RECT 291.075000  19.415000 292.085000  19.585000 ;
      RECT 291.075000  21.245000 292.085000  21.415000 ;
      RECT 291.075000  22.525000 292.085000  22.695000 ;
      RECT 291.075000  23.075000 292.085000  23.245000 ;
      RECT 291.075000  24.355000 292.085000  24.525000 ;
      RECT 291.075000  25.435000 292.085000  25.605000 ;
      RECT 291.125000   7.345000 292.085000   7.435000 ;
      RECT 291.180000  88.625000 299.555000  92.010000 ;
      RECT 291.180000  92.010000 299.570000  93.070000 ;
      RECT 291.185000  75.535000 297.140000  85.300000 ;
      RECT 291.185000  85.300000 299.555000  88.625000 ;
      RECT 291.345000  29.095000 292.035000  29.405000 ;
      RECT 291.345000  31.435000 292.035000  31.665000 ;
      RECT 291.615000 200.085000 292.285000 200.255000 ;
      RECT 292.035000  63.070000 293.175000  69.040000 ;
      RECT 292.035000  69.040000 307.420000  70.420000 ;
      RECT 292.035000  70.420000 363.050000  71.040000 ;
      RECT 292.035000  71.040000 297.140000  74.525000 ;
      RECT 292.075000  35.325000 292.245000  36.460000 ;
      RECT 292.075000  36.460000 292.325000  37.260000 ;
      RECT 292.335000   2.985000 292.765000   7.485000 ;
      RECT 292.335000   7.485000 292.505000   8.025000 ;
      RECT 292.335000   8.025000 292.765000  10.585000 ;
      RECT 292.335000  13.435000 292.505000  25.915000 ;
      RECT 292.365000  29.095000 293.055000  29.955000 ;
      RECT 292.365000  31.435000 293.055000  31.665000 ;
      RECT 292.415000  38.035000 292.585000  39.425000 ;
      RECT 292.415000  39.595000 292.585000  40.985000 ;
      RECT 292.480000  35.380000 292.650000  36.370000 ;
      RECT 292.715000 200.495000 293.245000 215.995000 ;
      RECT 292.755000  38.090000 292.925000  38.730000 ;
      RECT 292.755000  38.730000 293.290000  38.900000 ;
      RECT 292.755000  38.900000 292.925000  39.370000 ;
      RECT 292.755000  39.650000 292.925000  40.575000 ;
      RECT 292.755000  40.575000 293.290000  40.745000 ;
      RECT 292.755000  40.745000 292.925000  40.930000 ;
      RECT 293.285000  29.040000 293.475000  31.380000 ;
      RECT 293.585000  35.705000 296.295000  35.875000 ;
      RECT 293.585000  36.585000 296.295000  36.755000 ;
      RECT 293.585000  37.465000 296.295000  37.635000 ;
      RECT 293.585000  38.345000 296.295000  38.515000 ;
      RECT 293.585000  39.225000 296.295000  39.395000 ;
      RECT 293.585000  40.105000 296.295000  40.275000 ;
      RECT 293.585000  40.985000 296.295000  41.155000 ;
      RECT 293.630000 113.195000 294.300000 113.525000 ;
      RECT 293.675000 200.085000 294.345000 200.255000 ;
      RECT 293.700000 113.165000 294.230000 113.195000 ;
      RECT 293.715000  28.765000 293.885000  31.995000 ;
      RECT 293.755000 113.910000 296.755000 164.900000 ;
      RECT 294.365000 178.905000 344.705000 182.950000 ;
      RECT 294.605000  34.845000 294.775000  35.040000 ;
      RECT 294.605000  35.040000 301.075000  35.395000 ;
      RECT 294.775000 200.495000 295.305000 215.995000 ;
      RECT 295.045000  44.300000 325.445000  44.470000 ;
      RECT 295.045000  44.470000 295.215000  49.840000 ;
      RECT 295.225000  21.015000 297.080000  21.285000 ;
      RECT 295.225000  21.285000 295.395000  21.605000 ;
      RECT 295.525000  44.820000 295.795000  50.840000 ;
      RECT 295.525000  50.840000 296.955000  51.140000 ;
      RECT 295.525000  51.140000 295.795000  54.430000 ;
      RECT 295.735000 200.085000 296.405000 200.255000 ;
      RECT 295.965000  45.575000 296.235000  50.000000 ;
      RECT 295.965000  50.000000 296.255000  50.670000 ;
      RECT 296.025000  64.435000 297.590000  64.605000 ;
      RECT 296.025000  64.605000 296.535000  67.865000 ;
      RECT 296.090000  56.625000 296.260000  63.475000 ;
      RECT 296.090000  63.475000 300.945000  63.645000 ;
      RECT 296.320000  13.520000 299.220000  13.640000 ;
      RECT 296.320000  13.640000 296.580000  14.585000 ;
      RECT 296.320000  16.000000 296.580000  16.900000 ;
      RECT 296.400000   4.635000 299.220000   4.815000 ;
      RECT 296.400000   4.815000 296.580000  12.515000 ;
      RECT 296.400000  12.515000 299.220000  12.695000 ;
      RECT 296.400000  13.460000 299.220000  13.520000 ;
      RECT 296.400000  14.585000 296.580000  16.000000 ;
      RECT 296.400000  16.900000 296.580000  17.085000 ;
      RECT 296.400000  17.300000 297.000000  17.485000 ;
      RECT 296.400000  17.485000 296.570000  17.830000 ;
      RECT 296.400000  18.055000 296.580000  19.485000 ;
      RECT 296.400000  19.485000 299.220000  19.770000 ;
      RECT 296.400000  20.535000 299.220000  20.715000 ;
      RECT 296.400000  20.715000 296.580000  20.845000 ;
      RECT 296.400000  21.455000 296.580000  24.345000 ;
      RECT 296.400000  24.345000 299.220000  24.525000 ;
      RECT 296.400000  25.500000 299.220000  25.680000 ;
      RECT 296.400000  25.680000 296.580000  34.060000 ;
      RECT 296.400000  34.060000 299.220000  34.240000 ;
      RECT 296.405000  44.470000 296.575000  49.570000 ;
      RECT 296.405000  51.720000 296.575000  54.780000 ;
      RECT 296.485000  50.035000 297.015000  50.205000 ;
      RECT 296.785000  50.015000 296.955000  50.035000 ;
      RECT 296.785000  50.205000 296.955000  50.840000 ;
      RECT 296.805000  57.440000 296.975000  62.290000 ;
      RECT 296.815000  55.765000 296.985000  55.965000 ;
      RECT 296.815000  55.965000 304.360000  56.295000 ;
      RECT 296.830000  16.385000 297.000000  17.300000 ;
      RECT 296.830000  26.145000 297.000000  26.815000 ;
      RECT 296.830000  27.970000 297.000000  29.905000 ;
      RECT 296.835000 200.495000 297.365000 215.995000 ;
      RECT 296.845000  35.930000 297.015000  36.955000 ;
      RECT 296.845000  36.955000 297.380000  37.125000 ;
      RECT 296.845000  37.125000 297.015000  37.410000 ;
      RECT 296.845000  37.690000 297.015000  40.575000 ;
      RECT 296.845000  40.575000 297.380000  40.745000 ;
      RECT 296.845000  40.745000 297.015000  40.930000 ;
      RECT 296.900000   5.450000 297.070000   8.690000 ;
      RECT 296.900000   9.520000 297.070000  11.985000 ;
      RECT 296.900000  18.000000 298.370000  18.170000 ;
      RECT 296.900000  18.170000 297.070000  18.955000 ;
      RECT 296.910000  21.285000 297.080000  23.710000 ;
      RECT 296.925000  49.665000 297.455000  49.835000 ;
      RECT 296.970000  14.105000 297.140000  15.520000 ;
      RECT 296.970000  15.520000 298.370000  15.690000 ;
      RECT 297.185000  44.820000 297.455000  49.665000 ;
      RECT 297.185000  49.835000 297.455000  54.430000 ;
      RECT 297.195000  56.635000 299.145000  56.805000 ;
      RECT 297.235000  35.705000 299.945000  35.875000 ;
      RECT 297.235000  36.585000 299.945000  36.755000 ;
      RECT 297.235000  37.465000 299.945000  37.635000 ;
      RECT 297.235000  38.345000 299.945000  38.515000 ;
      RECT 297.235000  39.225000 299.945000  39.395000 ;
      RECT 297.235000  40.105000 299.945000  40.275000 ;
      RECT 297.235000  40.985000 299.945000  41.155000 ;
      RECT 297.300000   5.225000 298.310000   5.395000 ;
      RECT 297.300000   6.105000 298.310000   6.275000 ;
      RECT 297.300000   6.985000 298.310000   7.155000 ;
      RECT 297.300000   7.865000 298.310000   8.035000 ;
      RECT 297.300000   8.745000 298.310000   8.915000 ;
      RECT 297.300000   9.295000 298.310000   9.465000 ;
      RECT 297.300000  10.175000 298.310000  10.345000 ;
      RECT 297.300000  11.055000 298.310000  11.225000 ;
      RECT 297.300000  11.935000 298.310000  12.105000 ;
      RECT 297.300000  21.125000 298.310000  21.295000 ;
      RECT 297.300000  22.005000 298.310000  22.175000 ;
      RECT 297.300000  22.885000 298.310000  23.055000 ;
      RECT 297.300000  23.765000 298.310000  23.935000 ;
      RECT 297.300000  28.200000 298.310000  28.370000 ;
      RECT 297.300000  29.080000 298.310000  29.250000 ;
      RECT 297.300000  29.960000 298.310000  30.130000 ;
      RECT 297.300000  30.840000 298.310000  31.010000 ;
      RECT 297.300000  31.720000 298.310000  31.890000 ;
      RECT 297.300000  32.600000 298.310000  32.770000 ;
      RECT 297.300000  33.480000 298.310000  33.650000 ;
      RECT 297.360000  14.050000 298.370000  14.140000 ;
      RECT 297.360000  14.140000 298.790000  14.310000 ;
      RECT 297.360000  14.830000 298.370000  15.000000 ;
      RECT 297.360000  15.690000 298.370000  15.780000 ;
      RECT 297.360000  16.160000 298.370000  16.330000 ;
      RECT 297.360000  16.620000 298.370000  16.790000 ;
      RECT 297.360000  17.080000 298.370000  17.250000 ;
      RECT 297.360000  17.540000 298.370000  17.710000 ;
      RECT 297.360000  18.550000 298.370000  18.720000 ;
      RECT 297.360000  19.010000 298.370000  19.180000 ;
      RECT 297.360000 111.435000 298.210000 166.535000 ;
      RECT 297.420000  26.090000 298.090000  26.260000 ;
      RECT 297.420000  26.870000 298.090000  27.040000 ;
      RECT 297.420000  27.650000 298.090000  27.820000 ;
      RECT 297.645000  65.155000 297.815000  67.865000 ;
      RECT 297.715000  44.820000 298.005000  49.740000 ;
      RECT 297.715000  49.740000 299.955000  49.910000 ;
      RECT 297.715000  49.910000 298.005000  51.240000 ;
      RECT 297.715000  51.240000 298.245000  51.410000 ;
      RECT 297.715000  51.410000 298.005000  54.430000 ;
      RECT 297.720000  55.295000 325.845000  55.645000 ;
      RECT 297.795000 200.085000 298.465000 200.255000 ;
      RECT 297.870000  64.435000 307.830000  64.605000 ;
      RECT 298.085000  57.440000 298.255000  62.290000 ;
      RECT 298.175000  50.405000 298.705000  50.575000 ;
      RECT 298.205000  50.080000 298.375000  50.405000 ;
      RECT 298.205000  50.575000 298.375000  50.750000 ;
      RECT 298.615000  44.470000 298.785000  49.570000 ;
      RECT 298.620000  14.310000 298.790000  15.725000 ;
      RECT 298.620000  16.420000 298.790000  18.435000 ;
      RECT 298.620000  26.870000 298.790000  27.595000 ;
      RECT 298.620000  30.185000 298.790000  33.425000 ;
      RECT 298.630000  64.425000 305.885000  64.435000 ;
      RECT 298.715000  51.720000 298.885000  54.780000 ;
      RECT 298.895000 200.495000 299.425000 215.995000 ;
      RECT 298.925000  65.155000 299.095000  67.865000 ;
      RECT 299.025000  50.960000 302.075000  51.130000 ;
      RECT 299.040000   4.815000 299.220000   7.175000 ;
      RECT 299.040000   7.175000 299.630000   7.345000 ;
      RECT 299.040000   7.345000 299.220000  12.515000 ;
      RECT 299.040000  13.640000 299.220000  19.485000 ;
      RECT 299.040000  20.715000 299.220000  24.345000 ;
      RECT 299.040000  25.680000 299.220000  34.060000 ;
      RECT 299.055000  50.080000 299.225000  50.960000 ;
      RECT 299.225000  48.845000 299.755000  49.015000 ;
      RECT 299.365000  57.440000 299.535000  62.290000 ;
      RECT 299.395000  44.820000 299.565000  48.845000 ;
      RECT 299.395000  49.015000 299.565000  49.570000 ;
      RECT 299.595000  51.720000 299.765000  53.000000 ;
      RECT 299.595000  53.000000 300.125000  53.170000 ;
      RECT 299.595000  53.170000 299.765000  54.430000 ;
      RECT 299.780000 109.585000 300.970000 127.885000 ;
      RECT 299.780000 127.885000 358.600000 128.205000 ;
      RECT 299.780000 128.205000 300.970000 143.735000 ;
      RECT 299.780000 143.735000 340.665000 143.905000 ;
      RECT 299.780000 143.905000 302.715000 159.150000 ;
      RECT 299.780000 159.150000 351.405000 160.000000 ;
      RECT 299.780000 160.000000 300.630000 168.145000 ;
      RECT 299.780000 176.145000 300.630000 176.600000 ;
      RECT 299.780000 176.600000 346.320000 177.450000 ;
      RECT 299.785000  49.910000 299.955000  50.670000 ;
      RECT 299.795000  71.685000 301.815000  72.435000 ;
      RECT 299.795000  82.265000 301.815000  83.015000 ;
      RECT 299.855000 200.085000 300.525000 200.255000 ;
      RECT 299.955000  57.440000 300.125000  62.290000 ;
      RECT 299.985000   4.635000 302.730000   4.815000 ;
      RECT 299.985000   4.815000 300.165000  18.835000 ;
      RECT 299.985000  19.705000 300.165000  34.060000 ;
      RECT 299.985000  34.060000 302.730000  34.240000 ;
      RECT 300.045000  19.005000 300.585000  19.535000 ;
      RECT 300.085000  56.635000 300.755000  56.805000 ;
      RECT 300.095000  40.575000 300.665000  40.745000 ;
      RECT 300.150000 234.980000 301.755000 235.745000 ;
      RECT 300.150000 235.745000 301.130000 238.080000 ;
      RECT 300.175000  44.470000 300.345000  49.570000 ;
      RECT 300.205000  65.155000 300.375000  67.865000 ;
      RECT 300.410000 223.695000 301.020000 225.350000 ;
      RECT 300.410000 229.255000 301.260000 232.355000 ;
      RECT 300.410000 240.705000 301.260000 242.540000 ;
      RECT 300.410000 242.540000 327.275000 243.460000 ;
      RECT 300.410000 243.460000 327.245000 243.640000 ;
      RECT 300.415000   5.450000 300.585000   9.890000 ;
      RECT 300.415000  10.840000 300.585000  12.280000 ;
      RECT 300.415000  13.325000 300.585000  15.785000 ;
      RECT 300.415000  16.420000 300.585000  18.255000 ;
      RECT 300.415000  19.535000 300.585000  19.725000 ;
      RECT 300.415000  20.295000 300.585000  21.735000 ;
      RECT 300.415000  22.570000 300.585000  27.125000 ;
      RECT 300.415000  27.955000 300.615000  28.955000 ;
      RECT 300.415000  30.405000 301.855000  30.575000 ;
      RECT 300.415000  30.575000 300.585000  31.665000 ;
      RECT 300.415000  31.840000 300.585000  33.425000 ;
      RECT 300.475000  51.720000 300.645000  54.780000 ;
      RECT 300.480000  50.000000 300.650000  50.670000 ;
      RECT 300.495000  35.930000 300.665000  37.520000 ;
      RECT 300.495000  37.690000 300.665000  40.575000 ;
      RECT 300.495000  40.745000 300.665000  40.930000 ;
      RECT 300.595000  48.845000 301.125000  49.015000 ;
      RECT 300.600000  29.235000 300.955000  30.235000 ;
      RECT 300.735000  57.440000 300.905000  62.290000 ;
      RECT 300.750000 225.650000 300.920000 226.630000 ;
      RECT 300.785000  28.885000 300.955000  29.235000 ;
      RECT 300.800000  83.975000 358.600000  84.825000 ;
      RECT 300.800000  84.825000 300.970000 108.735000 ;
      RECT 300.845000   5.225000 301.855000   5.395000 ;
      RECT 300.845000   6.405000 301.855000   6.575000 ;
      RECT 300.845000   7.585000 301.920000   7.755000 ;
      RECT 300.845000   8.765000 301.855000   8.935000 ;
      RECT 300.845000   9.945000 301.855000  10.115000 ;
      RECT 300.845000  10.615000 301.855000  10.785000 ;
      RECT 300.845000  11.045000 301.855000  11.215000 ;
      RECT 300.845000  11.475000 301.855000  11.645000 ;
      RECT 300.845000  11.905000 301.855000  12.105000 ;
      RECT 300.845000  12.335000 301.855000  12.505000 ;
      RECT 300.845000  13.590000 301.855000  13.760000 ;
      RECT 300.845000  14.050000 301.855000  14.220000 ;
      RECT 300.845000  14.510000 301.855000  14.680000 ;
      RECT 300.845000  14.970000 301.855000  15.140000 ;
      RECT 300.845000  15.430000 301.855000  15.600000 ;
      RECT 300.845000  15.890000 301.855000  16.060000 ;
      RECT 300.845000  16.350000 301.855000  16.520000 ;
      RECT 300.845000  16.810000 301.855000  16.980000 ;
      RECT 300.845000  17.360000 301.855000  17.530000 ;
      RECT 300.845000  17.820000 302.255000  17.990000 ;
      RECT 300.845000  18.370000 301.855000  18.540000 ;
      RECT 300.845000  18.830000 301.855000  19.000000 ;
      RECT 300.845000  19.290000 301.855000  19.460000 ;
      RECT 300.845000  20.070000 301.855000  20.240000 ;
      RECT 300.845000  20.500000 301.855000  20.670000 ;
      RECT 300.845000  20.930000 301.855000  21.100000 ;
      RECT 300.845000  21.360000 301.855000  21.530000 ;
      RECT 300.845000  21.790000 301.855000  21.960000 ;
      RECT 300.845000  22.460000 301.855000  22.630000 ;
      RECT 300.845000  23.640000 301.855000  23.810000 ;
      RECT 300.845000  24.820000 301.855000  24.990000 ;
      RECT 300.845000  26.000000 301.855000  26.170000 ;
      RECT 300.845000  27.180000 301.855000  27.350000 ;
      RECT 300.845000  30.840000 301.855000  31.010000 ;
      RECT 300.845000  31.720000 301.855000  31.890000 ;
      RECT 300.845000  32.600000 301.855000  32.770000 ;
      RECT 300.845000  33.480000 301.855000  33.650000 ;
      RECT 300.905000  35.395000 301.075000  41.465000 ;
      RECT 300.955000  44.820000 301.125000  48.845000 ;
      RECT 300.955000  49.015000 301.125000  50.080000 ;
      RECT 300.955000  50.080000 306.010000  50.265000 ;
      RECT 300.955000 200.495000 301.485000 215.995000 ;
      RECT 300.965000  20.470000 301.855000  20.500000 ;
      RECT 300.995000  53.000000 301.525000  53.170000 ;
      RECT 301.005000  50.440000 308.990000  50.610000 ;
      RECT 301.050000  50.610000 308.780000  50.665000 ;
      RECT 301.185000  27.730000 301.855000  27.900000 ;
      RECT 301.185000  29.010000 301.855000  29.180000 ;
      RECT 301.185000  30.100000 301.855000  30.405000 ;
      RECT 301.355000  51.720000 301.525000  53.000000 ;
      RECT 301.355000  53.170000 301.525000  54.430000 ;
      RECT 301.445000  39.185000 302.005000  39.355000 ;
      RECT 301.485000  65.155000 301.655000  67.865000 ;
      RECT 301.505000  44.470000 301.675000  49.570000 ;
      RECT 301.560000 161.460000 326.650000 162.310000 ;
      RECT 301.560000 162.310000 302.410000 174.990000 ;
      RECT 301.560000 174.990000 326.650000 175.840000 ;
      RECT 301.650000 200.085000 302.585000 200.255000 ;
      RECT 301.835000  35.125000 306.195000  35.295000 ;
      RECT 301.835000  35.295000 302.005000  39.185000 ;
      RECT 301.835000  39.355000 302.005000  41.565000 ;
      RECT 301.835000  41.565000 306.195000  41.735000 ;
      RECT 301.865000 160.000000 351.405000 160.220000 ;
      RECT 301.920000  35.040000 306.110000  35.125000 ;
      RECT 301.925000 224.125000 311.925000 226.460000 ;
      RECT 301.925000 229.425000 311.925000 232.185000 ;
      RECT 301.925000 235.150000 311.925000 237.910000 ;
      RECT 301.925000 240.875000 311.925000 242.110000 ;
      RECT 302.085000  14.275000 302.255000  15.375000 ;
      RECT 302.085000  15.655000 302.255000  16.755000 ;
      RECT 302.085000  17.990000 302.255000  18.775000 ;
      RECT 302.095000  48.355000 302.625000  48.525000 ;
      RECT 302.215000  86.040000 302.385000  87.360000 ;
      RECT 302.215000  87.360000 303.745000  87.530000 ;
      RECT 302.215000  87.530000 302.385000  87.910000 ;
      RECT 302.215000  87.910000 303.985000  88.080000 ;
      RECT 302.215000  88.080000 302.385000  89.970000 ;
      RECT 302.215000  89.970000 303.525000  90.140000 ;
      RECT 302.215000  90.140000 302.385000  96.450000 ;
      RECT 302.215000  96.450000 309.585000  97.225000 ;
      RECT 302.215000  97.225000 310.285000  97.815000 ;
      RECT 302.215000  97.815000 309.585000  98.390000 ;
      RECT 302.215000  98.390000 316.875000  98.560000 ;
      RECT 302.215000 113.960000 316.875000 114.130000 ;
      RECT 302.215000 114.130000 309.585000 114.715000 ;
      RECT 302.215000 114.715000 310.285000 115.305000 ;
      RECT 302.215000 115.305000 309.585000 116.070000 ;
      RECT 302.215000 116.070000 302.385000 122.380000 ;
      RECT 302.215000 122.380000 303.525000 122.550000 ;
      RECT 302.215000 122.550000 302.385000 124.440000 ;
      RECT 302.215000 124.440000 303.985000 124.610000 ;
      RECT 302.215000 124.610000 302.385000 126.480000 ;
      RECT 302.215000 129.450000 338.510000 129.620000 ;
      RECT 302.215000 129.620000 302.385000 142.385000 ;
      RECT 302.225000 104.770000 316.875000 104.940000 ;
      RECT 302.225000 104.940000 312.705000 107.580000 ;
      RECT 302.225000 107.580000 316.875000 107.750000 ;
      RECT 302.235000  51.720000 302.405000  54.780000 ;
      RECT 302.245000  35.930000 302.415000  36.955000 ;
      RECT 302.245000  36.955000 302.780000  37.125000 ;
      RECT 302.245000  37.125000 302.415000  37.410000 ;
      RECT 302.245000  37.690000 302.415000  39.610000 ;
      RECT 302.245000  39.610000 302.830000  39.780000 ;
      RECT 302.245000  39.780000 302.415000  40.930000 ;
      RECT 302.255000  99.140000 302.425000 103.890000 ;
      RECT 302.255000 108.340000 302.425000 113.205000 ;
      RECT 302.275000 129.415000 338.480000 129.450000 ;
      RECT 302.285000  44.820000 302.455000  48.355000 ;
      RECT 302.285000  48.525000 302.455000  49.570000 ;
      RECT 302.285000  74.465000 348.750000  75.120000 ;
      RECT 302.285000  75.120000 303.575000  82.955000 ;
      RECT 302.285000  82.955000 348.750000  83.975000 ;
      RECT 302.550000   4.815000 302.730000  34.060000 ;
      RECT 302.550000 113.550000 303.625000 113.720000 ;
      RECT 302.580000  94.730000 302.750000  95.090000 ;
      RECT 302.580000  95.090000 303.525000  95.260000 ;
      RECT 302.615000 104.350000 303.625000 104.520000 ;
      RECT 302.635000  35.705000 305.345000  35.875000 ;
      RECT 302.635000  36.585000 305.345000  36.755000 ;
      RECT 302.635000  37.465000 305.345000  37.635000 ;
      RECT 302.635000  38.345000 305.345000  38.515000 ;
      RECT 302.635000  39.225000 305.345000  39.395000 ;
      RECT 302.635000  40.105000 305.345000  40.275000 ;
      RECT 302.635000  40.985000 305.345000  41.155000 ;
      RECT 302.635000  92.530000 303.525000  92.700000 ;
      RECT 302.635000 119.820000 303.525000 119.990000 ;
      RECT 302.650000 166.450000 302.820000 170.850000 ;
      RECT 302.705000 117.260000 303.525000 117.430000 ;
      RECT 302.705000 117.430000 302.875000 117.790000 ;
      RECT 302.725000  86.080000 303.745000  86.250000 ;
      RECT 302.745000  91.250000 303.635000  91.420000 ;
      RECT 302.745000  93.810000 303.635000  93.980000 ;
      RECT 302.745000 118.540000 303.635000 118.710000 ;
      RECT 302.745000 121.100000 303.635000 121.270000 ;
      RECT 302.765000  65.155000 302.935000  67.865000 ;
      RECT 302.785000  51.720000 302.955000  53.370000 ;
      RECT 302.785000  53.370000 303.315000  53.540000 ;
      RECT 302.785000  53.540000 302.955000  54.430000 ;
      RECT 302.825000 130.030000 303.155000 130.540000 ;
      RECT 302.825000 135.540000 303.785000 136.050000 ;
      RECT 302.825000 136.430000 303.155000 136.940000 ;
      RECT 302.825000 141.940000 303.785000 142.450000 ;
      RECT 302.855000  88.690000 303.985000  88.860000 ;
      RECT 302.855000  95.870000 303.525000  96.040000 ;
      RECT 302.855000 116.480000 303.525000 116.650000 ;
      RECT 302.855000 123.660000 303.985000 123.830000 ;
      RECT 302.905000 130.540000 303.075000 130.600000 ;
      RECT 302.905000 136.940000 303.075000 137.000000 ;
      RECT 302.980000  96.040000 303.510000  96.090000 ;
      RECT 303.015000 200.495000 303.545000 215.995000 ;
      RECT 303.035000  99.140000 303.205000 103.890000 ;
      RECT 303.035000 108.340000 303.205000 113.090000 ;
      RECT 303.065000  44.470000 303.235000  49.570000 ;
      RECT 303.110000  50.865000 304.460000  51.170000 ;
      RECT 303.150000 160.565000 303.680000 160.895000 ;
      RECT 303.285000 162.480000 313.285000 165.195000 ;
      RECT 303.285000 172.105000 313.285000 174.820000 ;
      RECT 303.455000 130.030000 304.415000 130.540000 ;
      RECT 303.455000 136.430000 304.415000 136.940000 ;
      RECT 303.480000  53.000000 304.010000  53.170000 ;
      RECT 303.480000 145.155000 339.050000 145.325000 ;
      RECT 303.480000 145.325000 303.650000 158.215000 ;
      RECT 303.480000 158.215000 339.050000 158.385000 ;
      RECT 303.495000   4.635000 310.725000   4.815000 ;
      RECT 303.495000   4.815000 303.675000  28.605000 ;
      RECT 303.495000  28.605000 310.725000  28.785000 ;
      RECT 303.580000  56.465000 303.750000  57.515000 ;
      RECT 303.580000  57.745000 303.750000  58.075000 ;
      RECT 303.580000  58.695000 303.750000  59.025000 ;
      RECT 303.580000  59.195000 303.750000  61.905000 ;
      RECT 303.665000  51.720000 303.835000  53.000000 ;
      RECT 303.665000  53.170000 303.835000  54.430000 ;
      RECT 303.675000  48.355000 304.205000  48.525000 ;
      RECT 303.755000 116.325000 304.285000 116.495000 ;
      RECT 303.770000  95.920000 304.300000  96.090000 ;
      RECT 303.815000  87.850000 303.985000  87.910000 ;
      RECT 303.815000  88.080000 303.985000  88.520000 ;
      RECT 303.815000  88.860000 303.985000  94.870000 ;
      RECT 303.815000  95.430000 303.985000  95.920000 ;
      RECT 303.815000  96.090000 303.985000  96.100000 ;
      RECT 303.815000  99.140000 303.985000 103.890000 ;
      RECT 303.815000 108.340000 303.985000 113.205000 ;
      RECT 303.815000 116.495000 303.985000 117.090000 ;
      RECT 303.815000 117.650000 303.985000 123.660000 ;
      RECT 303.815000 124.000000 303.985000 124.440000 ;
      RECT 303.815000 124.610000 303.985000 124.670000 ;
      RECT 303.845000  44.820000 304.015000  48.355000 ;
      RECT 303.845000  48.525000 304.015000  49.570000 ;
      RECT 303.850000  62.375000 304.360000  62.705000 ;
      RECT 303.915000   5.370000 304.095000  28.050000 ;
      RECT 303.920000  56.295000 304.290000  62.375000 ;
      RECT 303.945000  86.305000 304.115000  87.305000 ;
      RECT 304.045000  65.155000 304.215000  67.865000 ;
      RECT 304.055000 199.125000 307.965000 217.365000 ;
      RECT 304.060000 146.750000 304.230000 156.600000 ;
      RECT 304.085000 135.540000 305.045000 136.050000 ;
      RECT 304.085000 141.940000 305.045000 142.450000 ;
      RECT 304.185000  75.880000 347.135000  76.050000 ;
      RECT 304.185000  76.050000 304.355000  82.020000 ;
      RECT 304.185000  82.020000 347.135000  82.190000 ;
      RECT 304.285000 157.010000 312.435000 157.180000 ;
      RECT 304.315000   5.225000 307.025000   5.395000 ;
      RECT 304.315000   7.505000 307.025000   7.675000 ;
      RECT 304.315000   9.785000 307.025000   9.955000 ;
      RECT 304.315000  12.065000 307.025000  12.235000 ;
      RECT 304.315000  14.345000 307.025000  14.515000 ;
      RECT 304.315000  16.625000 307.025000  16.795000 ;
      RECT 304.315000  18.905000 307.025000  19.075000 ;
      RECT 304.315000  21.185000 307.025000  21.355000 ;
      RECT 304.315000  23.465000 307.025000  23.635000 ;
      RECT 304.315000  25.745000 307.025000  25.915000 ;
      RECT 304.315000  28.025000 307.025000  28.195000 ;
      RECT 304.365000  99.140000 304.535000 104.360000 ;
      RECT 304.365000 104.360000 305.090000 104.530000 ;
      RECT 304.365000 108.340000 304.535000 113.550000 ;
      RECT 304.365000 113.550000 305.090000 113.720000 ;
      RECT 304.375000  53.370000 304.905000  53.540000 ;
      RECT 304.400000 146.360000 308.170000 146.530000 ;
      RECT 304.460000  56.465000 304.630000  58.250000 ;
      RECT 304.460000  58.250000 305.760000  58.495000 ;
      RECT 304.460000  58.495000 304.630000  62.210000 ;
      RECT 304.545000  51.720000 304.715000  53.370000 ;
      RECT 304.545000  53.540000 304.715000  54.430000 ;
      RECT 304.555000  85.710000 304.725000  95.560000 ;
      RECT 304.555000 116.770000 304.725000 126.620000 ;
      RECT 304.625000  44.470000 304.795000  49.570000 ;
      RECT 304.715000 130.030000 305.675000 130.540000 ;
      RECT 304.715000 136.430000 305.675000 136.940000 ;
      RECT 304.765000  76.400000 304.935000  81.150000 ;
      RECT 304.780000  85.370000 308.780000  85.540000 ;
      RECT 304.780000  95.920000 308.780000  96.090000 ;
      RECT 304.780000 116.430000 308.780000 116.600000 ;
      RECT 304.780000 126.980000 308.780000 127.150000 ;
      RECT 304.845000  51.000000 306.195000  51.410000 ;
      RECT 304.850000 192.925000 305.180000 192.970000 ;
      RECT 304.850000 192.970000 308.750000 193.740000 ;
      RECT 304.850000 193.740000 305.180000 193.775000 ;
      RECT 304.895000  85.540000 308.665000  95.920000 ;
      RECT 304.895000 116.600000 308.665000 126.980000 ;
      RECT 305.050000  56.465000 305.220000  57.515000 ;
      RECT 305.050000  57.745000 305.220000  58.075000 ;
      RECT 305.050000  58.695000 305.220000  59.025000 ;
      RECT 305.050000  59.195000 305.220000  61.905000 ;
      RECT 305.110000  81.610000 305.920000  81.780000 ;
      RECT 305.145000  99.140000 305.315000 104.005000 ;
      RECT 305.145000 108.340000 305.315000 113.205000 ;
      RECT 305.235000  48.370000 305.765000  48.540000 ;
      RECT 305.250000  82.615000 305.780000  82.785000 ;
      RECT 305.265000  51.640000 305.795000  51.810000 ;
      RECT 305.320000  55.965000 305.830000  56.295000 ;
      RECT 305.320000  62.375000 305.830000  62.705000 ;
      RECT 305.320000 192.630000 308.105000 192.800000 ;
      RECT 305.320000 193.910000 308.105000 194.080000 ;
      RECT 305.320000 194.080000 308.030000 194.500000 ;
      RECT 305.325000  65.155000 305.495000  67.865000 ;
      RECT 305.345000 135.540000 306.305000 136.050000 ;
      RECT 305.345000 141.940000 306.305000 142.450000 ;
      RECT 305.390000  56.295000 305.760000  58.250000 ;
      RECT 305.390000  58.495000 305.760000  62.375000 ;
      RECT 305.405000  44.820000 305.575000  48.370000 ;
      RECT 305.405000  48.540000 305.575000  49.570000 ;
      RECT 305.420000  71.040000 363.050000  71.560000 ;
      RECT 305.420000  71.560000 372.120000  71.830000 ;
      RECT 305.420000  71.830000 372.185000  72.420000 ;
      RECT 305.425000  51.810000 305.595000  54.430000 ;
      RECT 305.535000 104.360000 315.165000 104.530000 ;
      RECT 305.535000 113.550000 315.165000 113.720000 ;
      RECT 305.930000  56.465000 306.100000  62.205000 ;
      RECT 305.945000  53.370000 306.475000  53.540000 ;
      RECT 305.975000 130.030000 306.935000 130.540000 ;
      RECT 305.975000 136.430000 306.935000 136.940000 ;
      RECT 306.025000  35.295000 306.195000  41.565000 ;
      RECT 306.045000  76.400000 306.215000  81.150000 ;
      RECT 306.185000  44.470000 306.355000  49.570000 ;
      RECT 306.200000  55.965000 306.710000  56.295000 ;
      RECT 306.200000  62.375000 306.710000  62.705000 ;
      RECT 306.270000  56.295000 306.640000  62.375000 ;
      RECT 306.305000  51.720000 306.475000  53.370000 ;
      RECT 306.305000  53.540000 306.475000  54.430000 ;
      RECT 306.390000  81.610000 307.200000  81.780000 ;
      RECT 306.425000  99.140000 306.595000 103.890000 ;
      RECT 306.425000 108.340000 306.595000 113.090000 ;
      RECT 306.510000  81.180000 307.040000  81.610000 ;
      RECT 306.540000  50.095000 310.730000  50.265000 ;
      RECT 306.605000  65.155000 306.775000  67.865000 ;
      RECT 306.605000 135.540000 307.565000 136.050000 ;
      RECT 306.605000 141.940000 307.565000 142.450000 ;
      RECT 306.620000  50.080000 310.730000  50.095000 ;
      RECT 306.665000  30.775000 308.685000  31.525000 ;
      RECT 306.665000  41.355000 308.685000  42.105000 ;
      RECT 306.785000  47.570000 307.315000  47.740000 ;
      RECT 306.810000  56.465000 306.980000  57.515000 ;
      RECT 306.810000  57.745000 306.980000  58.075000 ;
      RECT 306.810000  58.695000 306.980000  59.025000 ;
      RECT 306.810000  59.195000 306.980000  61.905000 ;
      RECT 306.855000  51.720000 307.025000  54.780000 ;
      RECT 306.965000  44.820000 307.135000  47.570000 ;
      RECT 306.965000  47.740000 307.135000  49.570000 ;
      RECT 307.235000 130.030000 308.195000 130.540000 ;
      RECT 307.235000 136.430000 308.195000 136.940000 ;
      RECT 307.250000  51.310000 308.095000  51.170000 ;
      RECT 307.325000  76.400000 307.495000  81.150000 ;
      RECT 307.565000  53.370000 308.095000  53.540000 ;
      RECT 307.575000   5.430000 307.745000  15.680000 ;
      RECT 307.575000  16.265000 307.745000  27.990000 ;
      RECT 307.635000  58.310000 308.640000  58.480000 ;
      RECT 307.670000  81.610000 308.480000  81.780000 ;
      RECT 307.705000  99.140000 307.875000 104.005000 ;
      RECT 307.705000 108.340000 307.875000 113.205000 ;
      RECT 307.735000  51.720000 307.905000  53.370000 ;
      RECT 307.735000  53.540000 307.905000  54.430000 ;
      RECT 307.745000  44.470000 307.915000  49.570000 ;
      RECT 307.790000  81.180000 308.320000  81.610000 ;
      RECT 307.865000 135.540000 308.825000 136.050000 ;
      RECT 307.865000 141.940000 308.825000 142.450000 ;
      RECT 307.885000  65.155000 308.055000  67.865000 ;
      RECT 307.930000  56.465000 308.100000  57.515000 ;
      RECT 307.930000  57.745000 308.100000  58.075000 ;
      RECT 307.930000  58.695000 308.100000  59.025000 ;
      RECT 307.930000  59.195000 308.100000  61.905000 ;
      RECT 308.110000  64.435000 309.675000  64.605000 ;
      RECT 308.155000   5.375000 309.505000   5.545000 ;
      RECT 308.155000   7.655000 310.725000   7.825000 ;
      RECT 308.155000   8.435000 309.505000   8.605000 ;
      RECT 308.155000   9.215000 309.505000   9.385000 ;
      RECT 308.155000   9.995000 309.505000  10.165000 ;
      RECT 308.155000  10.775000 309.505000  10.945000 ;
      RECT 308.155000  11.555000 309.505000  11.725000 ;
      RECT 308.155000  12.335000 309.505000  12.505000 ;
      RECT 308.155000  13.115000 309.505000  13.285000 ;
      RECT 308.155000  13.895000 309.505000  14.065000 ;
      RECT 308.155000  14.675000 309.505000  14.845000 ;
      RECT 308.155000  15.145000 310.725000  15.315000 ;
      RECT 308.155000  15.315000 309.505000  15.625000 ;
      RECT 308.155000  16.235000 309.505000  16.405000 ;
      RECT 308.155000  17.015000 309.505000  17.185000 ;
      RECT 308.155000  17.795000 309.505000  17.965000 ;
      RECT 308.155000  18.575000 309.505000  18.745000 ;
      RECT 308.155000  19.355000 309.505000  19.525000 ;
      RECT 308.155000  20.135000 309.505000  20.305000 ;
      RECT 308.155000  20.855000 309.505000  21.085000 ;
      RECT 308.155000  21.695000 309.505000  21.865000 ;
      RECT 308.155000  22.475000 309.505000  22.645000 ;
      RECT 308.155000  23.255000 309.505000  23.425000 ;
      RECT 308.155000  24.035000 309.505000  24.205000 ;
      RECT 308.155000  24.815000 309.505000  24.985000 ;
      RECT 308.155000  25.595000 310.725000  25.765000 ;
      RECT 308.155000  27.875000 309.505000  28.045000 ;
      RECT 308.200000  55.965000 308.710000  56.295000 ;
      RECT 308.200000  62.375000 308.710000  62.705000 ;
      RECT 308.270000  56.295000 308.640000  58.310000 ;
      RECT 308.270000  58.480000 308.640000  62.375000 ;
      RECT 308.340000 146.750000 308.510000 156.600000 ;
      RECT 308.345000  47.570000 308.875000  47.740000 ;
      RECT 308.495000 130.030000 309.455000 130.540000 ;
      RECT 308.495000 136.430000 309.455000 136.940000 ;
      RECT 308.525000  44.820000 308.695000  47.570000 ;
      RECT 308.525000  47.740000 308.695000  49.570000 ;
      RECT 308.580000 192.845000 308.750000 192.970000 ;
      RECT 308.580000 193.740000 308.750000 193.855000 ;
      RECT 308.605000  76.400000 308.775000  81.150000 ;
      RECT 308.615000  51.720000 308.785000  54.780000 ;
      RECT 308.685000 146.360000 312.450000 146.530000 ;
      RECT 308.810000  56.465000 308.980000  62.210000 ;
      RECT 308.835000  85.710000 309.005000  95.560000 ;
      RECT 308.835000 116.770000 309.005000 126.620000 ;
      RECT 308.950000  81.610000 309.760000  81.780000 ;
      RECT 308.965000 197.275000 309.815000 219.215000 ;
      RECT 308.985000  99.140000 309.155000 103.890000 ;
      RECT 308.985000 108.340000 309.155000 113.090000 ;
      RECT 309.070000  81.180000 309.600000  81.610000 ;
      RECT 309.080000  55.965000 310.470000  56.295000 ;
      RECT 309.080000  62.375000 310.470000  62.705000 ;
      RECT 309.125000 135.540000 310.085000 136.050000 ;
      RECT 309.125000 141.940000 310.085000 142.450000 ;
      RECT 309.150000  56.295000 309.520000  62.375000 ;
      RECT 309.165000  64.605000 309.675000  67.865000 ;
      RECT 309.200000  50.265000 310.730000  51.000000 ;
      RECT 309.295000  36.440000 336.945000  36.610000 ;
      RECT 309.295000  36.610000 309.465000  43.350000 ;
      RECT 309.295000  43.350000 327.370000  43.520000 ;
      RECT 309.305000  44.470000 309.475000  49.570000 ;
      RECT 309.320000  53.370000 309.850000  53.540000 ;
      RECT 309.415000  85.730000 309.585000  96.450000 ;
      RECT 309.415000 116.070000 309.585000 126.790000 ;
      RECT 309.495000  51.720000 309.665000  53.370000 ;
      RECT 309.495000  53.540000 309.665000  54.430000 ;
      RECT 309.690000  56.465000 309.860000  57.515000 ;
      RECT 309.690000  57.745000 309.860000  58.075000 ;
      RECT 309.690000  58.695000 309.860000  59.025000 ;
      RECT 309.690000  59.195000 309.860000  61.905000 ;
      RECT 309.725000   7.825000 310.725000   8.295000 ;
      RECT 309.725000  14.985000 310.725000  15.145000 ;
      RECT 309.725000  15.520000 310.375000  16.125000 ;
      RECT 309.725000  18.105000 310.725000  18.435000 ;
      RECT 309.725000  25.125000 310.725000  25.595000 ;
      RECT 309.725000  47.570000 310.255000  47.740000 ;
      RECT 309.755000 130.030000 310.715000 130.540000 ;
      RECT 309.755000 136.430000 310.715000 136.940000 ;
      RECT 309.815000  36.980000 327.760000  37.310000 ;
      RECT 309.815000  37.610000 331.930000  37.940000 ;
      RECT 309.815000  37.940000 310.485000  38.240000 ;
      RECT 309.815000  38.240000 331.930000  38.570000 ;
      RECT 309.815000  38.870000 331.930000  39.200000 ;
      RECT 309.815000  39.200000 310.485000  39.500000 ;
      RECT 309.815000  39.500000 331.930000  39.830000 ;
      RECT 309.815000  40.130000 331.930000  40.460000 ;
      RECT 309.815000  40.460000 310.485000  40.760000 ;
      RECT 309.815000  40.760000 331.930000  41.090000 ;
      RECT 309.815000  41.390000 331.930000  41.720000 ;
      RECT 309.815000  41.720000 310.485000  42.020000 ;
      RECT 309.815000  42.020000 331.930000  42.350000 ;
      RECT 309.815000  42.650000 327.825000  42.980000 ;
      RECT 309.875000 192.815000 342.805000 192.985000 ;
      RECT 309.875000 192.985000 310.045000 194.500000 ;
      RECT 309.885000  76.400000 310.055000  81.150000 ;
      RECT 310.030000  56.295000 310.400000  62.375000 ;
      RECT 310.085000  44.820000 310.255000  47.570000 ;
      RECT 310.085000  47.740000 310.255000  49.570000 ;
      RECT 310.230000  81.610000 311.040000  81.780000 ;
      RECT 310.230000 186.330000 310.400000 187.000000 ;
      RECT 310.230000 188.070000 310.400000 188.740000 ;
      RECT 310.230000 189.805000 310.400000 190.475000 ;
      RECT 310.230000 191.550000 310.400000 192.220000 ;
      RECT 310.265000  99.140000 310.435000 104.005000 ;
      RECT 310.265000 108.340000 310.435000 113.205000 ;
      RECT 310.350000  81.180000 310.880000  81.610000 ;
      RECT 310.375000  51.720000 310.545000  54.780000 ;
      RECT 310.385000 135.540000 311.345000 136.050000 ;
      RECT 310.385000 141.940000 311.345000 142.450000 ;
      RECT 310.545000   4.815000 310.725000   7.655000 ;
      RECT 310.545000   8.295000 310.725000  14.985000 ;
      RECT 310.545000  15.315000 310.725000  18.105000 ;
      RECT 310.545000  18.435000 310.725000  25.125000 ;
      RECT 310.545000  25.765000 310.725000  28.605000 ;
      RECT 310.570000  56.465000 310.740000  62.210000 ;
      RECT 310.590000 193.680000 311.125000 193.850000 ;
      RECT 310.595000 193.605000 311.125000 193.680000 ;
      RECT 310.595000 193.850000 311.125000 193.965000 ;
      RECT 310.630000 186.190000 325.660000 186.360000 ;
      RECT 310.630000 186.970000 325.660000 187.140000 ;
      RECT 310.630000 188.710000 325.660000 188.880000 ;
      RECT 310.630000 190.450000 325.660000 190.620000 ;
      RECT 310.630000 192.190000 325.660000 192.360000 ;
      RECT 310.710000 187.930000 325.660000 188.100000 ;
      RECT 310.710000 189.670000 325.660000 189.840000 ;
      RECT 310.710000 191.410000 325.660000 191.580000 ;
      RECT 310.815000 198.455000 337.525000 199.305000 ;
      RECT 310.815000 199.305000 312.125000 199.985000 ;
      RECT 310.815000 199.985000 312.345000 214.935000 ;
      RECT 310.815000 214.935000 312.125000 215.605000 ;
      RECT 310.815000 215.605000 337.525000 218.285000 ;
      RECT 310.830000  84.825000 311.000000  96.855000 ;
      RECT 310.830000  96.855000 358.600000  97.145000 ;
      RECT 310.830000 115.375000 358.600000 115.675000 ;
      RECT 310.830000 115.675000 311.000000 127.885000 ;
      RECT 310.840000  55.965000 311.350000  56.295000 ;
      RECT 310.840000  62.375000 311.350000  62.705000 ;
      RECT 310.865000  44.470000 311.035000  49.570000 ;
      RECT 310.910000  56.295000 311.280000  62.375000 ;
      RECT 310.955000  50.440000 317.525000  50.610000 ;
      RECT 311.015000 130.030000 311.975000 130.540000 ;
      RECT 311.015000 136.430000 311.975000 136.940000 ;
      RECT 311.085000  53.370000 311.615000  53.540000 ;
      RECT 311.095000  50.610000 317.385000  50.665000 ;
      RECT 311.165000  76.400000 311.335000  81.150000 ;
      RECT 311.200000  50.080000 318.330000  50.095000 ;
      RECT 311.200000  50.095000 318.365000  50.250000 ;
      RECT 311.255000  51.720000 311.425000  53.370000 ;
      RECT 311.255000  53.540000 311.425000  54.430000 ;
      RECT 311.355000  50.250000 318.400000  50.265000 ;
      RECT 311.425000 130.540000 311.595000 130.600000 ;
      RECT 311.425000 136.940000 311.595000 137.000000 ;
      RECT 311.450000  56.465000 311.620000  57.515000 ;
      RECT 311.450000  57.745000 311.620000  58.075000 ;
      RECT 311.450000  58.695000 311.620000  59.025000 ;
      RECT 311.450000  59.195000 311.620000  61.905000 ;
      RECT 311.495000   4.670000 316.655000   4.885000 ;
      RECT 311.495000   4.885000 313.805000  12.670000 ;
      RECT 311.495000  12.670000 312.345000  20.495000 ;
      RECT 311.495000  20.495000 313.805000  28.535000 ;
      RECT 311.495000  28.535000 316.655000  28.705000 ;
      RECT 311.495000  28.705000 316.155000  29.870000 ;
      RECT 311.510000  81.610000 312.320000  81.780000 ;
      RECT 311.545000  99.140000 311.715000 103.890000 ;
      RECT 311.545000 108.340000 311.715000 113.090000 ;
      RECT 311.555000  47.555000 312.085000  47.725000 ;
      RECT 311.630000  81.180000 312.160000  81.610000 ;
      RECT 311.645000 135.540000 312.605000 136.050000 ;
      RECT 311.645000 141.940000 312.605000 142.450000 ;
      RECT 311.675000  63.645000 314.475000  69.665000 ;
      RECT 311.675000  69.665000 324.515000  69.835000 ;
      RECT 311.745000  44.820000 311.915000  47.555000 ;
      RECT 311.745000  47.725000 311.915000  49.570000 ;
      RECT 312.135000  51.720000 312.305000  54.780000 ;
      RECT 312.275000 130.030000 313.235000 130.540000 ;
      RECT 312.275000 136.430000 313.235000 136.940000 ;
      RECT 312.300000  88.500000 313.190000  93.375000 ;
      RECT 312.300000 119.145000 313.190000 124.020000 ;
      RECT 312.340000  85.710000 313.190000  88.500000 ;
      RECT 312.340000  93.375000 313.190000  95.620000 ;
      RECT 312.340000  95.620000 312.510000  95.730000 ;
      RECT 312.340000 116.790000 312.510000 116.900000 ;
      RECT 312.340000 116.900000 313.190000 119.145000 ;
      RECT 312.340000 124.020000 313.190000 126.810000 ;
      RECT 312.355000 229.255000 313.205000 232.355000 ;
      RECT 312.400000 199.505000 315.240000 199.675000 ;
      RECT 312.400000 215.155000 315.240000 215.385000 ;
      RECT 312.445000  76.400000 312.615000  81.150000 ;
      RECT 312.500000  51.000000 317.250000  51.170000 ;
      RECT 312.620000 146.750000 312.790000 156.600000 ;
      RECT 312.625000  44.470000 312.795000  49.570000 ;
      RECT 312.695000 225.650000 313.675000 226.630000 ;
      RECT 312.695000 234.980000 312.865000 235.960000 ;
      RECT 312.695000 237.100000 313.675000 239.845000 ;
      RECT 312.695000 239.845000 323.780000 240.135000 ;
      RECT 312.695000 240.135000 324.480000 240.705000 ;
      RECT 312.725000  55.645000 325.845000  56.075000 ;
      RECT 312.725000  56.075000 314.475000  63.645000 ;
      RECT 312.790000  81.610000 313.600000  81.780000 ;
      RECT 312.825000  13.230000 313.155000  14.250000 ;
      RECT 312.825000  19.170000 313.155000  19.935000 ;
      RECT 312.825000  99.140000 312.995000 104.005000 ;
      RECT 312.825000 108.340000 312.995000 113.205000 ;
      RECT 312.845000  51.810000 313.375000  51.980000 ;
      RECT 312.845000 157.010000 316.845000 157.180000 ;
      RECT 312.905000 135.540000 313.865000 136.050000 ;
      RECT 312.905000 141.940000 313.865000 142.450000 ;
      RECT 312.910000  81.180000 313.440000  81.610000 ;
      RECT 312.955000 199.965000 313.125000 214.935000 ;
      RECT 312.960000 146.360000 316.690000 146.530000 ;
      RECT 313.015000  51.720000 313.185000  51.810000 ;
      RECT 313.015000  51.980000 313.185000  54.430000 ;
      RECT 313.115000 105.760000 313.290000 106.425000 ;
      RECT 313.115000 106.425000 313.285000 106.770000 ;
      RECT 313.120000 105.455000 313.290000 105.760000 ;
      RECT 313.245000  85.370000 317.245000  85.540000 ;
      RECT 313.245000  95.920000 317.245000  96.090000 ;
      RECT 313.245000 116.430000 317.245000 116.600000 ;
      RECT 313.245000 126.980000 317.245000 127.150000 ;
      RECT 313.315000  47.555000 313.845000  47.725000 ;
      RECT 313.360000  85.540000 317.130000  95.920000 ;
      RECT 313.360000 116.600000 317.130000 126.980000 ;
      RECT 313.375000 228.050000 314.225000 228.830000 ;
      RECT 313.375000 228.830000 324.545000 229.680000 ;
      RECT 313.375000 232.355000 324.545000 232.985000 ;
      RECT 313.375000 232.985000 323.690000 233.560000 ;
      RECT 313.505000  44.820000 313.675000  47.555000 ;
      RECT 313.505000  47.725000 313.675000  49.570000 ;
      RECT 313.535000 130.030000 314.495000 130.540000 ;
      RECT 313.535000 136.430000 314.495000 136.940000 ;
      RECT 313.635000  12.670000 313.805000  20.495000 ;
      RECT 313.725000  76.400000 313.895000  81.150000 ;
      RECT 313.735000 199.985000 313.905000 214.985000 ;
      RECT 313.845000 225.160000 323.845000 227.480000 ;
      RECT 313.845000 230.445000 323.845000 232.185000 ;
      RECT 313.845000 235.150000 323.845000 237.910000 ;
      RECT 313.845000 240.875000 323.845000 242.110000 ;
      RECT 313.860000 160.565000 314.390000 160.895000 ;
      RECT 313.860000 167.825000 314.390000 168.355000 ;
      RECT 313.860000 168.880000 314.390000 169.410000 ;
      RECT 313.895000  51.720000 314.065000  54.780000 ;
      RECT 314.020000 224.260000 323.750000 224.590000 ;
      RECT 314.055000  14.950000 314.225000  18.470000 ;
      RECT 314.070000  81.610000 314.880000  81.780000 ;
      RECT 314.105000  99.140000 314.275000 103.890000 ;
      RECT 314.105000 108.340000 314.275000 113.090000 ;
      RECT 314.165000 135.540000 315.125000 136.050000 ;
      RECT 314.165000 141.940000 315.125000 142.450000 ;
      RECT 314.190000  81.180000 314.720000  81.610000 ;
      RECT 314.295000 105.760000 314.465000 107.065000 ;
      RECT 314.385000  44.470000 314.555000  49.570000 ;
      RECT 314.415000  12.625000 315.545000  12.795000 ;
      RECT 314.415000  12.795000 314.585000  13.650000 ;
      RECT 314.415000  26.925000 314.585000  27.780000 ;
      RECT 314.415000  27.780000 315.545000  27.950000 ;
      RECT 314.515000 199.965000 314.685000 214.935000 ;
      RECT 314.600000  51.810000 315.130000  51.980000 ;
      RECT 314.625000   5.385000 315.635000   5.555000 ;
      RECT 314.625000   6.165000 315.635000   6.335000 ;
      RECT 314.625000   6.945000 315.635000   7.115000 ;
      RECT 314.625000   7.725000 315.635000   7.895000 ;
      RECT 314.625000   8.505000 315.635000   8.675000 ;
      RECT 314.625000   9.285000 315.635000   9.455000 ;
      RECT 314.625000  10.065000 315.635000  10.235000 ;
      RECT 314.625000  14.725000 315.635000  14.895000 ;
      RECT 314.625000  15.185000 315.635000  15.355000 ;
      RECT 314.625000  15.705000 315.635000  15.875000 ;
      RECT 314.625000  16.165000 315.635000  16.335000 ;
      RECT 314.625000  17.085000 315.635000  17.255000 ;
      RECT 314.625000  17.545000 315.635000  17.715000 ;
      RECT 314.625000  18.065000 315.635000  18.235000 ;
      RECT 314.625000  18.525000 315.635000  18.695000 ;
      RECT 314.625000  20.790000 315.635000  20.960000 ;
      RECT 314.625000  21.570000 315.635000  21.740000 ;
      RECT 314.625000  22.350000 315.635000  22.520000 ;
      RECT 314.625000  23.130000 315.635000  23.300000 ;
      RECT 314.625000  23.910000 315.635000  24.080000 ;
      RECT 314.625000  24.690000 315.635000  24.860000 ;
      RECT 314.625000  25.470000 316.025000  25.640000 ;
      RECT 314.635000 106.950000 315.305000 107.120000 ;
      RECT 314.775000  51.720000 314.945000  51.810000 ;
      RECT 314.775000  51.980000 314.945000  54.430000 ;
      RECT 314.795000 130.030000 315.755000 130.540000 ;
      RECT 314.795000 136.430000 315.755000 136.940000 ;
      RECT 314.875000  13.705000 315.545000  13.875000 ;
      RECT 314.875000  26.700000 315.545000  26.870000 ;
      RECT 314.925000 162.480000 324.925000 165.195000 ;
      RECT 314.925000 172.105000 324.925000 174.820000 ;
      RECT 315.005000  76.400000 315.175000  81.150000 ;
      RECT 315.010000  58.795000 315.180000  68.685000 ;
      RECT 315.015000  29.870000 316.155000  30.380000 ;
      RECT 315.075000  47.555000 315.605000  47.725000 ;
      RECT 315.265000  44.820000 315.435000  47.555000 ;
      RECT 315.265000  47.725000 315.435000  49.570000 ;
      RECT 315.295000 199.985000 316.485000 214.935000 ;
      RECT 315.340000  58.375000 316.010000  58.545000 ;
      RECT 315.340000  69.085000 316.010000  69.255000 ;
      RECT 315.350000  81.610000 316.160000  81.780000 ;
      RECT 315.385000  99.140000 315.555000 100.235000 ;
      RECT 315.385000 100.235000 315.560000 103.890000 ;
      RECT 315.385000 108.340000 315.555000 113.205000 ;
      RECT 315.390000 103.890000 315.560000 104.005000 ;
      RECT 315.410000 199.305000 316.370000 199.985000 ;
      RECT 315.410000 214.935000 316.370000 215.605000 ;
      RECT 315.425000 135.540000 316.385000 136.050000 ;
      RECT 315.425000 141.940000 316.385000 142.450000 ;
      RECT 315.470000  81.180000 316.000000  81.610000 ;
      RECT 315.475000 105.455000 315.645000 106.770000 ;
      RECT 315.610000 104.360000 316.835000 104.530000 ;
      RECT 315.610000 113.550000 316.835000 113.720000 ;
      RECT 315.655000  51.720000 315.825000  54.780000 ;
      RECT 315.855000   5.610000 316.025000  10.010000 ;
      RECT 315.855000  21.015000 316.025000  25.470000 ;
      RECT 316.055000 104.940000 316.225000 107.580000 ;
      RECT 316.055000 130.030000 317.015000 130.540000 ;
      RECT 316.055000 136.430000 317.015000 136.940000 ;
      RECT 316.145000  44.470000 316.315000  49.570000 ;
      RECT 316.190000  58.795000 316.360000  68.685000 ;
      RECT 316.285000  76.400000 316.455000  81.150000 ;
      RECT 316.365000  51.810000 316.895000  51.980000 ;
      RECT 316.485000   4.885000 316.655000  28.535000 ;
      RECT 316.520000  58.375000 317.190000  58.545000 ;
      RECT 316.520000  69.085000 317.190000  69.255000 ;
      RECT 316.535000  51.720000 316.705000  51.810000 ;
      RECT 316.535000  51.980000 316.705000  54.430000 ;
      RECT 316.540000 199.505000 319.380000 199.675000 ;
      RECT 316.540000 215.155000 319.380000 215.385000 ;
      RECT 316.630000  81.610000 317.440000  81.780000 ;
      RECT 316.665000  99.140000 316.835000 104.360000 ;
      RECT 316.665000 108.340000 316.835000 113.550000 ;
      RECT 316.685000 135.540000 317.645000 136.050000 ;
      RECT 316.685000 141.940000 317.645000 142.450000 ;
      RECT 316.750000  81.180000 317.280000  81.610000 ;
      RECT 316.835000  47.555000 317.365000  47.725000 ;
      RECT 316.900000 146.750000 317.070000 156.600000 ;
      RECT 317.025000  44.820000 317.195000  47.555000 ;
      RECT 317.025000  47.725000 317.195000  49.570000 ;
      RECT 317.095000 199.965000 317.265000 214.935000 ;
      RECT 317.125000 157.010000 325.405000 157.180000 ;
      RECT 317.240000 146.360000 321.010000 146.530000 ;
      RECT 317.300000  85.710000 318.620000  95.620000 ;
      RECT 317.300000 116.900000 318.620000 126.810000 ;
      RECT 317.315000 130.030000 318.275000 130.540000 ;
      RECT 317.315000 136.430000 318.275000 136.940000 ;
      RECT 317.370000  58.795000 317.540000  68.685000 ;
      RECT 317.415000  51.720000 317.585000  54.780000 ;
      RECT 317.565000  76.400000 317.735000  81.150000 ;
      RECT 317.695000  50.265000 318.400000  50.660000 ;
      RECT 317.695000  50.660000 319.045000  51.170000 ;
      RECT 317.700000  58.375000 318.370000  58.545000 ;
      RECT 317.700000  69.085000 318.370000  69.255000 ;
      RECT 317.875000 199.985000 318.045000 214.985000 ;
      RECT 317.905000  44.470000 318.075000  49.570000 ;
      RECT 317.910000  81.610000 318.720000  81.780000 ;
      RECT 317.945000 135.540000 318.905000 136.050000 ;
      RECT 317.945000 141.940000 318.905000 142.450000 ;
      RECT 317.980000  25.605000 318.560000  26.000000 ;
      RECT 318.030000  81.180000 318.560000  81.610000 ;
      RECT 318.125000  52.180000 318.655000  52.350000 ;
      RECT 318.250000  97.145000 318.420000 106.160000 ;
      RECT 318.250000 106.160000 358.600000 106.360000 ;
      RECT 318.250000 106.360000 318.420000 115.375000 ;
      RECT 318.295000  51.720000 318.465000  52.180000 ;
      RECT 318.295000  52.350000 318.465000  54.430000 ;
      RECT 318.380000   0.750000 360.060000   0.930000 ;
      RECT 318.380000   0.930000 318.560000  25.605000 ;
      RECT 318.380000  26.000000 318.560000  29.320000 ;
      RECT 318.380000  29.320000 359.140000  29.490000 ;
      RECT 318.380000  29.490000 318.560000  34.290000 ;
      RECT 318.380000  34.290000 338.205000  34.470000 ;
      RECT 318.455000  44.820000 318.625000  48.355000 ;
      RECT 318.455000  48.355000 318.985000  48.525000 ;
      RECT 318.455000  48.525000 318.625000  49.570000 ;
      RECT 318.550000  58.795000 318.720000  68.685000 ;
      RECT 318.575000 130.030000 319.535000 130.540000 ;
      RECT 318.575000 136.430000 319.535000 136.940000 ;
      RECT 318.655000 199.965000 318.825000 214.935000 ;
      RECT 318.675000  85.370000 322.675000  85.540000 ;
      RECT 318.675000  95.920000 322.675000  96.090000 ;
      RECT 318.675000 116.430000 322.675000 116.600000 ;
      RECT 318.675000 126.980000 322.675000 127.150000 ;
      RECT 318.700000  50.080000 321.410000  50.095000 ;
      RECT 318.700000  50.095000 321.450000  50.250000 ;
      RECT 318.760000  50.250000 321.450000  50.265000 ;
      RECT 318.790000  85.540000 322.560000  95.920000 ;
      RECT 318.790000 116.600000 322.560000 126.980000 ;
      RECT 318.845000  76.400000 319.015000  81.150000 ;
      RECT 318.880000  58.375000 319.550000  58.545000 ;
      RECT 318.880000  69.085000 319.550000  69.255000 ;
      RECT 319.045000  47.555000 319.575000  47.725000 ;
      RECT 319.175000  51.720000 319.345000  54.780000 ;
      RECT 319.190000  81.610000 320.000000  81.780000 ;
      RECT 319.205000 135.540000 320.165000 136.050000 ;
      RECT 319.205000 141.940000 320.165000 142.450000 ;
      RECT 319.235000  44.820000 319.405000  47.555000 ;
      RECT 319.235000  47.725000 319.405000  49.570000 ;
      RECT 319.310000  81.180000 319.840000  81.610000 ;
      RECT 319.325000   4.010000 342.670000   4.190000 ;
      RECT 319.325000   4.190000 319.505000  10.480000 ;
      RECT 319.325000  10.480000 342.670000  10.990000 ;
      RECT 319.325000  10.990000 319.505000  11.865000 ;
      RECT 319.325000  11.865000 320.055000  12.535000 ;
      RECT 319.325000  12.535000 319.505000  19.635000 ;
      RECT 319.325000  19.635000 320.055000  20.305000 ;
      RECT 319.325000  20.305000 319.505000  21.175000 ;
      RECT 319.325000  21.175000 342.670000  21.685000 ;
      RECT 319.325000  21.685000 319.505000  28.375000 ;
      RECT 319.325000  28.375000 358.705000  28.555000 ;
      RECT 319.360000  28.555000 342.390000  28.565000 ;
      RECT 319.435000 199.985000 320.625000 214.935000 ;
      RECT 319.450000  30.880000 322.020000  31.050000 ;
      RECT 319.450000  31.050000 319.620000  33.355000 ;
      RECT 319.450000  33.355000 322.020000  33.525000 ;
      RECT 319.455000  50.265000 320.805000  51.170000 ;
      RECT 319.550000 199.305000 320.510000 199.985000 ;
      RECT 319.550000 214.935000 320.510000 215.605000 ;
      RECT 319.665000  98.390000 356.795000  98.560000 ;
      RECT 319.665000  98.560000 319.835000 104.760000 ;
      RECT 319.665000 104.760000 356.795000 104.930000 ;
      RECT 319.665000 107.590000 356.795000 107.760000 ;
      RECT 319.665000 107.760000 319.835000 113.960000 ;
      RECT 319.665000 113.960000 356.795000 114.130000 ;
      RECT 319.730000  58.795000 319.900000  68.685000 ;
      RECT 319.825000  48.355000 320.355000  48.525000 ;
      RECT 319.835000 130.030000 320.165000 130.540000 ;
      RECT 319.835000 136.430000 320.165000 136.940000 ;
      RECT 319.885000  13.665000 321.020000  14.335000 ;
      RECT 319.885000  14.845000 320.055000  15.020000 ;
      RECT 319.885000  15.020000 320.475000  15.190000 ;
      RECT 319.885000  15.190000 320.055000  15.515000 ;
      RECT 319.885000  16.680000 320.055000  16.710000 ;
      RECT 319.885000  16.710000 320.475000  16.880000 ;
      RECT 319.885000  16.880000 320.055000  17.350000 ;
      RECT 319.885000  17.860000 320.055000  18.085000 ;
      RECT 319.885000  18.085000 320.475000  18.255000 ;
      RECT 319.885000  18.255000 320.055000  18.530000 ;
      RECT 319.885000  52.180000 320.415000  52.350000 ;
      RECT 319.915000 130.540000 320.085000 130.600000 ;
      RECT 319.915000 136.940000 320.085000 137.000000 ;
      RECT 320.015000  44.820000 320.185000  48.355000 ;
      RECT 320.015000  48.525000 320.185000  49.570000 ;
      RECT 320.025000   4.620000 320.705000   4.950000 ;
      RECT 320.025000   5.250000 320.675000   5.580000 ;
      RECT 320.025000   5.880000 320.675000   6.210000 ;
      RECT 320.025000   6.510000 320.675000   6.840000 ;
      RECT 320.025000  25.785000 320.675000  26.115000 ;
      RECT 320.025000  26.415000 320.675000  26.745000 ;
      RECT 320.025000  27.045000 320.675000  27.375000 ;
      RECT 320.025000  27.675000 320.705000  28.005000 ;
      RECT 320.055000  51.720000 320.225000  52.180000 ;
      RECT 320.055000  52.350000 320.225000  54.430000 ;
      RECT 320.060000  31.575000 321.070000  31.745000 ;
      RECT 320.060000  32.755000 321.070000  32.925000 ;
      RECT 320.085000   8.400000 320.735000   8.480000 ;
      RECT 320.085000   8.480000 320.815000   8.650000 ;
      RECT 320.085000   8.650000 320.735000   8.730000 ;
      RECT 320.085000  23.895000 320.735000  23.975000 ;
      RECT 320.085000  23.975000 320.815000  24.145000 ;
      RECT 320.085000  24.145000 320.735000  24.225000 ;
      RECT 320.125000  76.400000 320.295000  81.150000 ;
      RECT 320.225000   7.770000 320.875000   8.100000 ;
      RECT 320.225000   9.030000 320.875000   9.360000 ;
      RECT 320.225000  23.265000 320.875000  23.595000 ;
      RECT 320.225000  24.525000 320.875000  24.855000 ;
      RECT 320.235000 101.080000 320.415000 101.970000 ;
      RECT 320.235000 110.280000 320.415000 111.170000 ;
      RECT 320.245000  98.800000 320.895000  98.970000 ;
      RECT 320.245000  98.970000 320.415000 101.080000 ;
      RECT 320.245000 101.970000 320.415000 104.350000 ;
      RECT 320.245000 104.350000 320.895000 104.520000 ;
      RECT 320.245000 108.000000 320.895000 108.170000 ;
      RECT 320.245000 108.170000 320.415000 110.280000 ;
      RECT 320.245000 111.170000 320.415000 113.550000 ;
      RECT 320.245000 113.550000 320.895000 113.720000 ;
      RECT 320.275000  11.525000 330.165000  11.695000 ;
      RECT 320.275000  12.705000 330.165000  12.875000 ;
      RECT 320.275000  13.325000 330.165000  13.495000 ;
      RECT 320.275000  14.505000 330.165000  14.675000 ;
      RECT 320.275000  15.685000 330.165000  15.855000 ;
      RECT 320.275000  16.315000 330.165000  16.485000 ;
      RECT 320.275000  17.495000 330.165000  17.665000 ;
      RECT 320.275000  18.675000 330.165000  18.845000 ;
      RECT 320.275000  19.295000 330.165000  19.465000 ;
      RECT 320.275000  20.475000 330.165000  20.645000 ;
      RECT 320.400000  21.165000 342.200000  21.175000 ;
      RECT 320.400000  21.685000 342.200000  21.695000 ;
      RECT 320.470000  81.610000 321.280000  81.780000 ;
      RECT 320.590000  81.180000 321.120000  81.610000 ;
      RECT 320.595000 130.030000 320.925000 130.540000 ;
      RECT 320.595000 135.540000 321.555000 136.050000 ;
      RECT 320.595000 136.430000 320.925000 136.940000 ;
      RECT 320.595000 141.940000 321.555000 142.450000 ;
      RECT 320.605000  47.555000 321.135000  47.725000 ;
      RECT 320.645000  98.970000 320.815000 104.350000 ;
      RECT 320.645000 108.170000 320.815000 113.550000 ;
      RECT 320.675000 130.540000 320.845000 130.600000 ;
      RECT 320.675000 136.940000 320.845000 137.000000 ;
      RECT 320.680000 199.505000 323.520000 199.675000 ;
      RECT 320.680000 215.155000 323.520000 215.385000 ;
      RECT 320.790000  57.285000 320.960000  59.995000 ;
      RECT 320.795000  44.820000 320.965000  47.555000 ;
      RECT 320.795000  47.725000 320.965000  49.570000 ;
      RECT 320.825000   9.660000 321.475000   9.990000 ;
      RECT 320.825000  22.635000 321.475000  22.965000 ;
      RECT 320.935000  51.720000 321.105000  54.780000 ;
      RECT 320.955000  61.640000 321.125000  64.350000 ;
      RECT 321.025000  99.140000 321.195000 103.890000 ;
      RECT 321.025000 108.340000 321.195000 113.090000 ;
      RECT 321.150000  56.500000 321.820000  56.670000 ;
      RECT 321.180000 146.750000 321.350000 156.600000 ;
      RECT 321.215000  51.000000 322.730000  51.170000 ;
      RECT 321.225000 130.030000 322.185000 130.540000 ;
      RECT 321.225000 136.430000 322.185000 136.940000 ;
      RECT 321.235000 199.965000 321.405000 214.935000 ;
      RECT 321.250000  98.800000 325.250000  98.970000 ;
      RECT 321.250000 104.350000 325.250000 104.520000 ;
      RECT 321.250000 108.000000 325.250000 108.170000 ;
      RECT 321.250000 113.550000 325.250000 113.720000 ;
      RECT 321.315000 193.605000 321.825000 193.685000 ;
      RECT 321.315000 193.685000 321.875000 193.855000 ;
      RECT 321.315000 193.855000 321.825000 193.935000 ;
      RECT 321.320000  31.890000 321.490000  32.560000 ;
      RECT 321.345000  61.250000 322.015000  61.420000 ;
      RECT 321.385000  48.355000 321.915000  48.525000 ;
      RECT 321.405000  76.400000 321.575000  81.150000 ;
      RECT 321.415000  61.235000 321.945000  61.250000 ;
      RECT 321.520000 146.360000 325.290000 146.530000 ;
      RECT 321.575000  44.820000 321.745000  48.355000 ;
      RECT 321.575000  48.525000 321.745000  49.570000 ;
      RECT 321.645000  52.180000 322.175000  52.350000 ;
      RECT 321.750000  81.610000 322.560000  81.780000 ;
      RECT 321.815000  51.720000 321.985000  52.180000 ;
      RECT 321.815000  52.350000 321.985000  54.430000 ;
      RECT 321.850000  31.050000 322.020000  33.355000 ;
      RECT 321.855000 135.540000 322.815000 136.050000 ;
      RECT 321.855000 141.940000 322.815000 142.450000 ;
      RECT 321.870000  81.180000 322.400000  81.610000 ;
      RECT 321.880000  50.080000 324.590000  50.250000 ;
      RECT 321.880000  50.250000 322.730000  51.000000 ;
      RECT 322.015000 199.985000 322.185000 214.985000 ;
      RECT 322.070000  57.285000 322.240000  59.995000 ;
      RECT 322.185000  47.970000 322.715000  48.140000 ;
      RECT 322.235000  61.640000 322.405000  64.350000 ;
      RECT 322.355000  44.820000 322.525000  47.970000 ;
      RECT 322.355000  48.140000 322.525000  49.570000 ;
      RECT 322.385000 192.985000 342.805000 194.500000 ;
      RECT 322.430000  56.500000 323.100000  56.670000 ;
      RECT 322.485000 130.030000 323.445000 130.540000 ;
      RECT 322.485000 136.430000 323.445000 136.940000 ;
      RECT 322.605000  98.970000 323.900000 104.350000 ;
      RECT 322.605000 108.170000 323.900000 113.550000 ;
      RECT 322.625000  61.250000 323.295000  61.420000 ;
      RECT 322.685000  76.400000 322.855000  81.150000 ;
      RECT 322.695000  51.720000 322.865000  54.780000 ;
      RECT 322.695000  61.235000 323.225000  61.250000 ;
      RECT 322.730000  85.710000 322.900000  95.560000 ;
      RECT 322.730000 116.960000 322.900000 126.810000 ;
      RECT 322.795000 199.965000 322.965000 214.935000 ;
      RECT 322.890000  29.490000 323.060000  34.290000 ;
      RECT 322.920000  50.440000 325.445000  50.610000 ;
      RECT 322.920000  50.610000 324.530000  50.665000 ;
      RECT 322.950000  48.355000 323.480000  48.525000 ;
      RECT 322.955000  85.370000 326.955000  85.540000 ;
      RECT 322.955000  95.920000 326.955000  96.090000 ;
      RECT 322.955000 116.430000 326.955000 116.600000 ;
      RECT 322.955000 126.980000 326.955000 127.150000 ;
      RECT 323.030000  81.610000 323.840000  81.780000 ;
      RECT 323.070000  85.540000 326.840000  95.920000 ;
      RECT 323.070000 116.600000 326.840000 126.980000 ;
      RECT 323.115000 135.540000 324.075000 136.050000 ;
      RECT 323.115000 141.940000 324.075000 142.450000 ;
      RECT 323.135000  44.820000 323.305000  48.355000 ;
      RECT 323.135000  48.525000 323.305000  49.570000 ;
      RECT 323.135000 199.675000 323.405000 215.155000 ;
      RECT 323.150000  81.180000 323.680000  81.610000 ;
      RECT 323.275000  51.410000 325.845000  54.780000 ;
      RECT 323.350000  57.285000 323.520000  59.995000 ;
      RECT 323.515000  61.640000 323.685000  64.350000 ;
      RECT 323.575000 199.985000 324.765000 214.935000 ;
      RECT 323.595000   7.770000 324.245000   8.100000 ;
      RECT 323.595000   8.400000 324.245000   8.730000 ;
      RECT 323.595000   9.030000 324.245000   9.360000 ;
      RECT 323.595000  23.265000 324.245000  23.595000 ;
      RECT 323.595000  23.895000 324.245000  24.225000 ;
      RECT 323.595000  24.525000 324.245000  24.855000 ;
      RECT 323.690000 199.305000 324.650000 199.985000 ;
      RECT 323.690000 214.935000 324.650000 215.605000 ;
      RECT 323.745000  47.970000 324.275000  48.140000 ;
      RECT 323.745000 130.030000 324.705000 130.540000 ;
      RECT 323.745000 136.430000 324.705000 136.940000 ;
      RECT 323.850000  30.880000 326.420000  31.050000 ;
      RECT 323.850000  31.050000 324.020000  33.355000 ;
      RECT 323.850000  33.355000 326.420000  33.525000 ;
      RECT 323.915000  44.820000 324.085000  47.970000 ;
      RECT 323.915000  48.140000 324.085000  49.570000 ;
      RECT 323.950000 224.340000 324.480000 224.510000 ;
      RECT 323.950000 239.795000 324.480000 239.965000 ;
      RECT 323.965000  76.400000 324.135000  81.150000 ;
      RECT 324.015000 224.510000 324.480000 226.750000 ;
      RECT 324.015000 226.750000 324.645000 228.050000 ;
      RECT 324.015000 229.680000 324.545000 232.355000 ;
      RECT 324.015000 233.170000 324.545000 234.660000 ;
      RECT 324.015000 234.660000 324.645000 235.960000 ;
      RECT 324.310000  81.610000 325.120000  81.780000 ;
      RECT 324.310000 237.100000 324.645000 238.400000 ;
      RECT 324.310000 238.400000 324.480000 239.795000 ;
      RECT 324.335000  48.355000 324.865000  48.525000 ;
      RECT 324.345000  56.075000 325.845000  58.085000 ;
      RECT 324.345000  58.085000 324.515000  69.665000 ;
      RECT 324.375000 135.540000 325.335000 136.050000 ;
      RECT 324.375000 141.940000 325.335000 142.450000 ;
      RECT 324.430000  81.180000 324.960000  81.610000 ;
      RECT 324.475000  31.575000 325.485000  31.745000 ;
      RECT 324.475000  32.755000 325.485000  32.925000 ;
      RECT 324.625000   7.770000 325.275000   8.100000 ;
      RECT 324.625000   8.400000 325.275000   8.730000 ;
      RECT 324.625000   9.030000 325.275000   9.360000 ;
      RECT 324.625000  23.265000 325.275000  23.595000 ;
      RECT 324.625000  23.895000 325.275000  24.225000 ;
      RECT 324.625000  24.525000 325.275000  24.855000 ;
      RECT 324.695000  44.820000 324.865000  48.355000 ;
      RECT 324.695000  48.525000 324.865000  49.570000 ;
      RECT 324.720000 224.260000 325.250000 224.590000 ;
      RECT 324.815000 224.590000 325.145000 240.725000 ;
      RECT 324.820000 199.505000 327.660000 199.675000 ;
      RECT 324.820000 215.155000 327.660000 215.385000 ;
      RECT 324.935000 199.675000 325.205000 215.155000 ;
      RECT 325.005000 130.030000 325.965000 130.540000 ;
      RECT 325.005000 136.430000 325.965000 136.940000 ;
      RECT 325.245000  76.400000 325.415000  81.150000 ;
      RECT 325.275000  44.470000 325.445000  50.440000 ;
      RECT 325.305000  99.140000 325.475000 103.890000 ;
      RECT 325.305000 108.340000 325.475000 113.090000 ;
      RECT 325.310000 223.865000 325.845000 224.035000 ;
      RECT 325.315000 224.760000 325.845000 230.315000 ;
      RECT 325.375000 199.965000 325.545000 214.935000 ;
      RECT 325.390000 166.450000 325.560000 170.850000 ;
      RECT 325.405000 230.570000 326.255000 239.805000 ;
      RECT 325.405000 239.805000 327.275000 242.540000 ;
      RECT 325.420000 224.035000 325.845000 224.760000 ;
      RECT 325.460000 146.750000 325.630000 156.600000 ;
      RECT 325.530000  98.800000 329.530000  98.970000 ;
      RECT 325.530000 104.350000 329.530000 104.520000 ;
      RECT 325.530000 108.000000 329.530000 108.170000 ;
      RECT 325.530000 113.550000 329.530000 113.720000 ;
      RECT 325.590000  81.610000 326.400000  81.780000 ;
      RECT 325.635000 135.540000 326.595000 136.050000 ;
      RECT 325.635000 141.940000 326.595000 142.450000 ;
      RECT 325.710000  81.180000 326.240000  81.610000 ;
      RECT 325.735000  31.890000 325.905000  32.560000 ;
      RECT 325.800000 162.310000 326.650000 174.990000 ;
      RECT 325.930000  58.760000 336.675000  58.790000 ;
      RECT 325.930000  58.790000 355.455000  58.960000 ;
      RECT 325.930000  58.960000 336.675000  58.990000 ;
      RECT 325.930000  58.990000 326.160000  68.100000 ;
      RECT 325.930000  68.100000 363.050000  68.330000 ;
      RECT 325.960000  68.330000 363.050000  70.420000 ;
      RECT 326.020000 145.325000 326.610000 158.215000 ;
      RECT 326.040000 223.865000 326.600000 224.205000 ;
      RECT 326.040000 224.205000 327.030000 224.735000 ;
      RECT 326.085000 224.905000 326.255000 230.570000 ;
      RECT 326.155000 199.985000 326.325000 214.985000 ;
      RECT 326.250000  31.050000 326.420000  33.355000 ;
      RECT 326.265000 130.030000 327.225000 130.540000 ;
      RECT 326.265000 136.430000 327.225000 136.940000 ;
      RECT 326.425000 186.190000 341.375000 186.360000 ;
      RECT 326.425000 186.970000 341.375000 187.140000 ;
      RECT 326.425000 187.930000 341.375000 188.100000 ;
      RECT 326.425000 188.710000 341.375000 188.880000 ;
      RECT 326.425000 189.670000 341.375000 189.840000 ;
      RECT 326.425000 190.450000 341.375000 190.620000 ;
      RECT 326.425000 191.410000 341.375000 191.580000 ;
      RECT 326.425000 192.190000 341.375000 192.360000 ;
      RECT 326.500000 224.735000 327.030000 237.925000 ;
      RECT 326.500000 237.925000 327.465000 239.225000 ;
      RECT 326.525000  76.400000 326.695000  81.150000 ;
      RECT 326.745000  46.610000 327.370000  46.705000 ;
      RECT 326.745000  46.705000 355.510000  46.875000 ;
      RECT 326.745000  46.875000 326.955000  54.460000 ;
      RECT 326.745000  54.460000 353.860000  54.670000 ;
      RECT 326.745000  54.670000 326.955000  58.760000 ;
      RECT 326.770000 223.865000 327.565000 224.035000 ;
      RECT 326.780000 146.390000 327.310000 146.560000 ;
      RECT 326.870000  81.610000 327.680000  81.780000 ;
      RECT 326.885000  98.970000 328.180000 104.350000 ;
      RECT 326.885000 108.170000 328.180000 113.550000 ;
      RECT 326.895000 135.540000 327.855000 136.050000 ;
      RECT 326.895000 141.940000 327.855000 142.450000 ;
      RECT 326.935000 199.965000 327.105000 214.935000 ;
      RECT 326.980000 146.560000 327.310000 147.065000 ;
      RECT 326.980000 151.465000 327.310000 152.865000 ;
      RECT 326.980000 157.265000 327.940000 157.775000 ;
      RECT 326.990000  81.180000 327.520000  81.610000 ;
      RECT 327.010000  85.710000 328.330000  95.620000 ;
      RECT 327.010000 116.900000 328.330000 126.810000 ;
      RECT 327.065000  43.520000 327.370000  45.835000 ;
      RECT 327.065000  45.835000 348.060000  46.165000 ;
      RECT 327.065000  46.165000 327.370000  46.610000 ;
      RECT 327.190000  29.490000 327.360000  34.290000 ;
      RECT 327.200000 224.035000 327.565000 233.745000 ;
      RECT 327.365000  47.305000 344.700000  50.015000 ;
      RECT 327.365000  50.955000 344.700000  53.665000 ;
      RECT 327.365000  55.340000 353.220000  58.050000 ;
      RECT 327.395000   6.510000 328.045000   6.840000 ;
      RECT 327.395000  25.785000 328.045000  26.115000 ;
      RECT 327.410000 160.220000 328.260000 176.600000 ;
      RECT 327.480000   1.885000 328.290000   2.985000 ;
      RECT 327.525000 130.030000 328.485000 130.540000 ;
      RECT 327.525000 136.430000 328.485000 136.940000 ;
      RECT 327.595000  50.560000 344.415000  50.730000 ;
      RECT 327.595000  54.980000 352.995000  55.150000 ;
      RECT 327.610000  65.805000 328.320000  66.055000 ;
      RECT 327.610000 146.555000 328.570000 147.065000 ;
      RECT 327.610000 151.465000 327.940000 152.865000 ;
      RECT 327.650000  50.530000 344.375000  50.560000 ;
      RECT 327.715000 199.985000 328.905000 214.935000 ;
      RECT 327.805000  76.400000 327.975000  81.150000 ;
      RECT 327.830000 199.305000 328.790000 199.985000 ;
      RECT 327.830000 214.935000 328.785000 215.605000 ;
      RECT 327.915000 224.125000 337.915000 226.445000 ;
      RECT 327.915000 228.735000 337.915000 230.645000 ;
      RECT 327.915000 232.935000 337.915000 235.255000 ;
      RECT 327.915000 236.415000 337.915000 238.735000 ;
      RECT 327.915000 241.700000 337.915000 242.935000 ;
      RECT 327.995000   9.030000 328.645000   9.360000 ;
      RECT 327.995000  23.265000 328.645000  23.595000 ;
      RECT 328.055000   8.480000 328.645000   8.650000 ;
      RECT 328.055000  23.975000 328.645000  24.145000 ;
      RECT 328.065000  65.765000 328.240000  65.805000 ;
      RECT 328.065000  66.055000 328.240000  66.095000 ;
      RECT 328.095000  43.945000 333.410000  44.275000 ;
      RECT 328.095000  44.275000 328.765000  44.575000 ;
      RECT 328.095000  44.575000 333.410000  44.905000 ;
      RECT 328.095000  45.245000 328.885000  45.495000 ;
      RECT 328.135000   8.400000 328.305000   8.480000 ;
      RECT 328.135000   8.650000 328.305000   8.730000 ;
      RECT 328.135000  23.895000 328.305000  23.975000 ;
      RECT 328.135000  24.145000 328.305000  24.225000 ;
      RECT 328.150000  81.610000 328.960000  81.780000 ;
      RECT 328.155000 135.540000 329.115000 136.050000 ;
      RECT 328.155000 141.940000 329.115000 142.450000 ;
      RECT 328.160000  30.880000 330.780000  31.050000 ;
      RECT 328.160000  31.050000 328.330000  33.355000 ;
      RECT 328.160000  33.355000 330.730000  33.525000 ;
      RECT 328.240000 151.465000 328.570000 152.865000 ;
      RECT 328.240000 157.265000 329.200000 157.775000 ;
      RECT 328.255000 116.430000 332.385000 116.600000 ;
      RECT 328.255000 126.980000 332.385000 127.150000 ;
      RECT 328.270000  81.180000 328.800000  81.610000 ;
      RECT 328.385000  85.370000 332.385000  85.540000 ;
      RECT 328.385000  95.920000 332.385000  96.090000 ;
      RECT 328.425000   6.510000 329.075000   6.840000 ;
      RECT 328.425000  25.785000 329.075000  26.115000 ;
      RECT 328.475000   8.400000 328.645000   8.480000 ;
      RECT 328.475000   8.650000 328.645000   8.730000 ;
      RECT 328.475000  23.895000 328.645000  23.975000 ;
      RECT 328.475000  24.145000 328.645000  24.225000 ;
      RECT 328.495000  45.205000 328.885000  45.245000 ;
      RECT 328.495000  45.495000 328.885000  45.535000 ;
      RECT 328.500000  85.540000 332.270000  95.920000 ;
      RECT 328.500000 116.600000 332.270000 126.980000 ;
      RECT 328.740000 146.390000 329.270000 146.555000 ;
      RECT 328.740000 146.555000 329.830000 146.560000 ;
      RECT 328.765000  31.575000 329.775000  31.745000 ;
      RECT 328.765000  32.755000 329.775000  32.925000 ;
      RECT 328.785000 130.030000 329.745000 130.540000 ;
      RECT 328.785000 136.430000 329.745000 136.940000 ;
      RECT 328.870000 146.560000 329.830000 147.065000 ;
      RECT 328.870000 151.465000 329.200000 152.865000 ;
      RECT 328.920000 168.645000 340.380000 169.345000 ;
      RECT 328.920000 169.345000 329.620000 175.240000 ;
      RECT 328.920000 175.240000 340.380000 175.940000 ;
      RECT 328.955000 215.155000 331.800000 215.385000 ;
      RECT 328.960000 199.505000 331.800000 199.675000 ;
      RECT 329.025000   8.400000 329.535000   8.480000 ;
      RECT 329.025000   8.480000 329.615000   8.650000 ;
      RECT 329.025000   8.650000 329.535000   8.730000 ;
      RECT 329.025000  23.895000 329.535000  23.975000 ;
      RECT 329.025000  23.975000 329.615000  24.145000 ;
      RECT 329.025000  24.145000 329.535000  24.225000 ;
      RECT 329.055000   7.850000 329.785000   8.020000 ;
      RECT 329.055000  24.605000 329.785000  24.775000 ;
      RECT 329.065000 161.195000 372.360000 162.215000 ;
      RECT 329.065000 162.215000 351.455000 162.385000 ;
      RECT 329.065000 162.385000 329.235000 163.295000 ;
      RECT 329.065000 163.295000 334.220000 163.625000 ;
      RECT 329.065000 163.625000 329.235000 165.455000 ;
      RECT 329.065000 165.455000 334.220000 165.785000 ;
      RECT 329.065000 165.785000 329.235000 167.705000 ;
      RECT 329.065000 167.705000 344.015000 167.875000 ;
      RECT 329.085000  76.400000 329.255000  81.150000 ;
      RECT 329.135000   7.770000 329.785000   7.850000 ;
      RECT 329.135000   8.020000 329.785000   8.100000 ;
      RECT 329.135000  24.525000 329.785000  24.605000 ;
      RECT 329.135000  24.775000 329.785000  24.855000 ;
      RECT 329.195000 130.540000 329.365000 130.600000 ;
      RECT 329.195000 136.940000 329.365000 137.000000 ;
      RECT 329.415000 135.540000 330.375000 136.050000 ;
      RECT 329.415000 141.940000 330.375000 142.450000 ;
      RECT 329.430000  81.610000 330.240000  81.780000 ;
      RECT 329.500000 151.465000 329.830000 152.865000 ;
      RECT 329.500000 157.265000 330.460000 157.775000 ;
      RECT 329.515000 199.965000 329.685000 214.935000 ;
      RECT 329.550000  81.180000 330.080000  81.610000 ;
      RECT 329.585000  99.140000 329.755000 103.890000 ;
      RECT 329.585000 108.340000 329.755000 113.090000 ;
      RECT 329.765000 164.015000 334.220000 164.345000 ;
      RECT 329.765000 164.345000 330.345000 164.735000 ;
      RECT 329.765000 164.735000 334.220000 165.065000 ;
      RECT 329.765000 166.175000 334.220000 166.505000 ;
      RECT 329.765000 166.505000 330.345000 166.895000 ;
      RECT 329.765000 166.895000 334.220000 167.225000 ;
      RECT 329.810000  98.800000 333.810000  98.970000 ;
      RECT 329.810000 104.350000 333.810000 104.520000 ;
      RECT 329.810000 108.000000 333.810000 108.170000 ;
      RECT 329.810000 113.550000 333.810000 113.720000 ;
      RECT 330.005000  13.725000 330.705000  13.895000 ;
      RECT 330.005000  14.915000 330.705000  15.085000 ;
      RECT 330.005000  16.710000 330.705000  16.880000 ;
      RECT 330.005000  18.275000 330.705000  18.445000 ;
      RECT 330.025000  31.890000 330.195000  32.560000 ;
      RECT 330.045000 130.030000 331.005000 130.540000 ;
      RECT 330.045000 136.430000 331.005000 136.940000 ;
      RECT 330.130000 146.555000 331.090000 147.065000 ;
      RECT 330.130000 151.465000 330.460000 152.865000 ;
      RECT 330.295000 199.985000 330.465000 214.985000 ;
      RECT 330.365000  76.400000 330.535000  81.150000 ;
      RECT 330.380000 170.105000 338.920000 170.805000 ;
      RECT 330.380000 170.805000 331.090000 173.780000 ;
      RECT 330.380000 173.780000 338.920000 174.480000 ;
      RECT 330.425000   7.140000 331.075000   7.470000 ;
      RECT 330.425000  25.155000 331.075000  25.485000 ;
      RECT 330.510000 162.755000 346.820000 163.075000 ;
      RECT 330.535000  13.665000 330.705000  13.725000 ;
      RECT 330.535000  13.895000 330.705000  14.915000 ;
      RECT 330.535000  15.085000 330.705000  15.515000 ;
      RECT 330.535000  16.655000 330.705000  16.710000 ;
      RECT 330.535000  16.880000 330.705000  18.275000 ;
      RECT 330.535000  18.445000 330.705000  18.505000 ;
      RECT 330.560000  31.050000 330.730000  33.355000 ;
      RECT 330.675000 135.540000 331.635000 136.050000 ;
      RECT 330.675000 141.940000 331.635000 142.450000 ;
      RECT 330.695000  37.055000 331.225000  37.225000 ;
      RECT 330.695000  42.755000 331.225000  42.925000 ;
      RECT 330.710000  81.610000 331.520000  81.780000 ;
      RECT 330.760000 151.465000 331.090000 152.865000 ;
      RECT 330.760000 157.265000 331.720000 157.775000 ;
      RECT 330.830000  81.180000 331.360000  81.610000 ;
      RECT 331.075000  13.665000 331.245000  13.705000 ;
      RECT 331.075000  13.705000 331.775000  13.875000 ;
      RECT 331.075000  13.875000 331.245000  15.285000 ;
      RECT 331.075000  15.285000 331.775000  15.455000 ;
      RECT 331.075000  15.455000 331.245000  15.515000 ;
      RECT 331.075000  16.655000 331.245000  16.720000 ;
      RECT 331.075000  16.720000 331.775000  16.890000 ;
      RECT 331.075000  16.890000 331.245000  18.120000 ;
      RECT 331.075000  18.120000 331.775000  18.290000 ;
      RECT 331.075000  18.290000 331.245000  18.505000 ;
      RECT 331.075000 199.965000 331.245000 214.935000 ;
      RECT 331.165000  98.970000 332.460000 104.350000 ;
      RECT 331.165000 108.170000 332.460000 113.550000 ;
      RECT 331.260000 146.390000 331.790000 146.555000 ;
      RECT 331.260000 146.555000 332.350000 146.560000 ;
      RECT 331.305000 130.030000 332.265000 130.540000 ;
      RECT 331.305000 136.430000 332.265000 136.940000 ;
      RECT 331.375000 171.625000 331.785000 172.950000 ;
      RECT 331.390000 146.560000 332.350000 147.065000 ;
      RECT 331.390000 151.465000 331.720000 152.865000 ;
      RECT 331.615000  11.525000 341.505000  11.695000 ;
      RECT 331.615000  12.705000 341.505000  12.875000 ;
      RECT 331.615000  13.325000 341.505000  13.495000 ;
      RECT 331.615000  14.505000 341.505000  14.675000 ;
      RECT 331.615000  15.685000 341.505000  15.855000 ;
      RECT 331.615000  16.315000 341.505000  16.485000 ;
      RECT 331.615000  17.495000 341.505000  17.665000 ;
      RECT 331.615000  18.675000 341.505000  18.845000 ;
      RECT 331.615000  19.295000 341.505000  19.465000 ;
      RECT 331.615000  20.475000 341.505000  20.645000 ;
      RECT 331.645000  76.400000 331.815000  81.150000 ;
      RECT 331.710000 163.075000 333.320000 163.125000 ;
      RECT 331.855000 199.985000 333.045000 214.935000 ;
      RECT 331.935000 135.540000 332.895000 136.050000 ;
      RECT 331.935000 141.940000 332.895000 142.450000 ;
      RECT 331.955000 171.280000 337.350000 171.820000 ;
      RECT 331.955000 172.755000 337.350000 173.295000 ;
      RECT 331.970000 199.305000 332.930000 199.985000 ;
      RECT 331.970000 214.935000 332.930000 215.605000 ;
      RECT 331.990000  81.610000 332.800000  81.780000 ;
      RECT 332.020000 151.465000 332.350000 152.865000 ;
      RECT 332.020000 157.265000 332.980000 157.775000 ;
      RECT 332.110000  81.180000 332.640000  81.610000 ;
      RECT 332.240000  29.490000 332.410000  34.290000 ;
      RECT 332.380000  45.270000 332.910000  45.440000 ;
      RECT 332.390000  45.205000 332.900000  45.270000 ;
      RECT 332.390000  45.440000 332.900000  45.535000 ;
      RECT 332.395000   8.400000 333.045000   8.730000 ;
      RECT 332.395000  23.895000 333.045000  24.225000 ;
      RECT 332.425000   9.030000 333.075000   9.360000 ;
      RECT 332.425000  23.265000 333.075000  23.595000 ;
      RECT 332.440000  85.710000 333.290000  88.500000 ;
      RECT 332.440000  88.500000 333.330000  93.375000 ;
      RECT 332.440000  93.375000 333.290000  95.620000 ;
      RECT 332.440000 116.900000 333.290000 119.145000 ;
      RECT 332.440000 119.145000 333.330000 124.020000 ;
      RECT 332.440000 124.020000 333.290000 126.810000 ;
      RECT 332.565000 130.030000 333.525000 130.540000 ;
      RECT 332.565000 136.430000 333.525000 136.940000 ;
      RECT 332.650000 146.555000 333.610000 147.065000 ;
      RECT 332.650000 151.465000 332.980000 152.865000 ;
      RECT 332.825000   7.770000 333.475000   8.100000 ;
      RECT 332.825000  24.525000 333.475000  24.855000 ;
      RECT 332.925000  76.400000 333.095000  81.150000 ;
      RECT 333.100000 199.505000 335.940000 199.675000 ;
      RECT 333.100000 215.155000 335.940000 215.385000 ;
      RECT 333.120000  95.620000 333.290000  95.730000 ;
      RECT 333.120000 116.790000 333.290000 116.900000 ;
      RECT 333.195000 135.540000 334.155000 136.050000 ;
      RECT 333.195000 141.940000 334.155000 142.450000 ;
      RECT 333.270000  81.610000 334.080000  81.780000 ;
      RECT 333.280000 151.465000 333.610000 152.865000 ;
      RECT 333.280000 157.265000 334.240000 157.775000 ;
      RECT 333.390000  81.180000 333.920000  81.610000 ;
      RECT 333.655000 199.965000 333.825000 214.935000 ;
      RECT 333.810000  30.880000 336.380000  31.050000 ;
      RECT 333.810000  31.050000 333.980000  33.355000 ;
      RECT 333.810000  33.355000 336.380000  33.525000 ;
      RECT 333.825000   8.400000 334.475000   8.730000 ;
      RECT 333.825000  23.895000 334.475000  24.225000 ;
      RECT 333.825000 130.030000 334.785000 130.540000 ;
      RECT 333.825000 136.430000 334.785000 136.940000 ;
      RECT 333.865000  99.140000 334.035000 103.890000 ;
      RECT 333.865000 108.340000 334.035000 113.090000 ;
      RECT 333.910000 146.390000 334.440000 146.560000 ;
      RECT 333.910000 146.560000 334.240000 147.065000 ;
      RECT 333.910000 151.465000 334.240000 152.865000 ;
      RECT 334.090000  98.800000 338.090000  98.970000 ;
      RECT 334.090000 104.350000 338.090000 104.520000 ;
      RECT 334.090000 108.000000 338.090000 108.170000 ;
      RECT 334.090000 113.550000 338.090000 113.720000 ;
      RECT 334.205000  76.400000 334.375000  81.150000 ;
      RECT 334.435000 199.985000 334.605000 214.985000 ;
      RECT 334.445000  31.575000 335.455000  31.745000 ;
      RECT 334.445000  32.755000 335.455000  32.925000 ;
      RECT 334.455000 135.540000 335.415000 136.050000 ;
      RECT 334.455000 141.940000 335.415000 142.450000 ;
      RECT 334.470000 163.295000 342.840000 163.625000 ;
      RECT 334.470000 164.015000 342.840000 164.345000 ;
      RECT 334.470000 164.735000 342.840000 165.065000 ;
      RECT 334.470000 165.455000 342.840000 165.785000 ;
      RECT 334.470000 166.175000 342.840000 166.505000 ;
      RECT 334.470000 166.895000 342.840000 167.225000 ;
      RECT 334.550000  81.610000 335.655000  81.780000 ;
      RECT 334.630000  84.825000 334.800000  96.855000 ;
      RECT 334.630000 115.675000 334.800000 127.885000 ;
      RECT 334.670000 145.325000 334.840000 158.215000 ;
      RECT 335.085000 130.030000 336.045000 130.540000 ;
      RECT 335.085000 136.430000 336.045000 136.940000 ;
      RECT 335.105000  44.020000 335.635000  44.190000 ;
      RECT 335.105000  44.640000 335.635000  44.810000 ;
      RECT 335.115000  43.945000 335.625000  44.020000 ;
      RECT 335.115000  44.190000 335.625000  44.275000 ;
      RECT 335.115000  44.575000 335.625000  44.640000 ;
      RECT 335.115000  44.810000 335.625000  44.905000 ;
      RECT 335.215000 199.965000 335.385000 214.935000 ;
      RECT 335.390000 147.505000 335.560000 157.355000 ;
      RECT 335.445000  98.970000 336.740000 104.350000 ;
      RECT 335.445000 108.170000 336.740000 113.550000 ;
      RECT 335.485000  76.400000 335.655000  81.610000 ;
      RECT 335.500000  36.980000 336.310000  37.310000 ;
      RECT 335.515000  42.650000 336.310000  42.980000 ;
      RECT 335.520000  37.610000 336.310000  37.940000 ;
      RECT 335.520000  38.240000 336.310000  39.200000 ;
      RECT 335.520000  39.500000 336.310000  40.460000 ;
      RECT 335.520000  40.760000 337.545000  41.090000 ;
      RECT 335.520000  41.390000 337.545000  41.720000 ;
      RECT 335.520000  42.020000 337.545000  42.350000 ;
      RECT 335.705000  31.890000 335.875000  32.560000 ;
      RECT 335.715000 135.540000 336.675000 136.050000 ;
      RECT 335.715000 141.940000 336.675000 142.450000 ;
      RECT 335.745000 146.815000 338.115000 146.985000 ;
      RECT 335.995000 199.985000 337.525000 214.935000 ;
      RECT 336.025000  77.050000 336.205000  80.460000 ;
      RECT 336.035000  76.400000 336.205000  77.050000 ;
      RECT 336.035000  80.460000 336.205000  81.150000 ;
      RECT 336.100000  89.620000 336.990000  94.495000 ;
      RECT 336.100000 118.025000 336.990000 122.900000 ;
      RECT 336.140000  85.710000 336.990000  89.620000 ;
      RECT 336.140000  94.495000 336.990000  95.620000 ;
      RECT 336.140000  95.620000 336.310000  95.730000 ;
      RECT 336.140000 116.790000 336.310000 116.900000 ;
      RECT 336.140000 116.900000 336.990000 118.025000 ;
      RECT 336.140000 122.900000 336.990000 126.810000 ;
      RECT 336.210000  31.050000 336.380000  33.355000 ;
      RECT 336.215000 199.305000 337.525000 199.985000 ;
      RECT 336.215000 214.935000 337.525000 215.605000 ;
      RECT 336.260000  81.320000 339.100000  81.780000 ;
      RECT 336.345000 130.030000 337.305000 130.540000 ;
      RECT 336.345000 136.430000 337.305000 136.940000 ;
      RECT 336.375000  80.750000 336.645000  81.320000 ;
      RECT 336.570000 147.505000 336.740000 157.355000 ;
      RECT 336.660000  36.610000 336.945000  39.575000 ;
      RECT 336.660000  39.575000 364.060000  39.745000 ;
      RECT 336.690000   2.235000 337.200000   2.755000 ;
      RECT 336.690000   2.755000 337.220000   2.925000 ;
      RECT 336.815000  76.400000 336.985000  81.150000 ;
      RECT 336.875000  40.130000 363.370000  40.460000 ;
      RECT 336.875000  42.650000 337.545000  43.610000 ;
      RECT 336.890000  45.270000 337.420000  45.440000 ;
      RECT 336.900000  45.205000 337.410000  45.270000 ;
      RECT 336.900000  45.440000 337.410000  45.535000 ;
      RECT 336.975000 135.540000 337.935000 136.050000 ;
      RECT 336.975000 141.940000 337.935000 142.450000 ;
      RECT 337.045000  85.370000 341.245000  85.540000 ;
      RECT 337.045000  95.920000 341.245000  96.090000 ;
      RECT 337.045000 116.430000 341.045000 116.600000 ;
      RECT 337.045000 126.980000 341.045000 127.150000 ;
      RECT 337.120000 147.505000 337.290000 157.355000 ;
      RECT 337.155000  80.750000 337.425000  81.320000 ;
      RECT 337.160000  85.540000 340.930000  95.920000 ;
      RECT 337.160000 116.600000 340.930000 126.980000 ;
      RECT 337.255000  29.490000 337.425000  34.290000 ;
      RECT 337.595000  76.400000 337.765000  81.150000 ;
      RECT 337.605000 130.030000 337.935000 130.540000 ;
      RECT 337.605000 136.430000 337.935000 136.940000 ;
      RECT 337.685000 130.540000 337.855000 130.600000 ;
      RECT 337.685000 136.940000 337.855000 137.000000 ;
      RECT 337.935000  80.750000 338.205000  81.320000 ;
      RECT 338.025000  34.470000 338.205000  37.515000 ;
      RECT 338.025000  37.515000 363.565000  37.695000 ;
      RECT 338.145000  99.140000 338.315000 103.890000 ;
      RECT 338.145000 108.340000 338.315000 113.090000 ;
      RECT 338.220000 170.805000 338.920000 173.780000 ;
      RECT 338.300000 147.505000 338.470000 157.355000 ;
      RECT 338.340000 129.620000 338.510000 142.385000 ;
      RECT 338.370000  98.800000 342.370000  98.970000 ;
      RECT 338.370000 104.350000 342.370000 104.520000 ;
      RECT 338.370000 108.000000 342.370000 108.170000 ;
      RECT 338.370000 113.550000 342.370000 113.720000 ;
      RECT 338.375000  76.400000 338.545000  81.150000 ;
      RECT 338.535000  30.255000 362.530000  30.425000 ;
      RECT 338.535000  30.425000 338.705000  36.590000 ;
      RECT 338.535000  36.590000 362.530000  36.750000 ;
      RECT 338.535000  36.750000 340.015000  36.760000 ;
      RECT 338.570000  82.390000 339.100000  82.560000 ;
      RECT 338.685000 223.695000 339.535000 243.640000 ;
      RECT 338.705000 197.275000 344.705000 199.885000 ;
      RECT 338.705000 199.885000 343.725000 216.295000 ;
      RECT 338.705000 216.295000 346.520000 219.215000 ;
      RECT 338.715000  80.750000 338.985000  81.315000 ;
      RECT 338.715000  81.315000 339.100000  81.320000 ;
      RECT 338.880000 145.325000 339.050000 158.215000 ;
      RECT 339.155000  76.400000 339.325000  81.150000 ;
      RECT 339.435000  31.485000 339.605000  32.155000 ;
      RECT 339.435000  32.665000 339.605000  33.335000 ;
      RECT 339.435000  33.845000 339.605000  34.515000 ;
      RECT 339.435000  35.025000 339.605000  35.695000 ;
      RECT 339.680000 169.345000 340.380000 175.240000 ;
      RECT 339.690000  77.050000 339.890000  80.860000 ;
      RECT 339.705000  76.400000 339.875000  77.050000 ;
      RECT 339.705000  80.860000 339.875000  81.610000 ;
      RECT 339.705000  81.610000 340.430000  81.780000 ;
      RECT 339.725000  98.970000 341.020000 104.350000 ;
      RECT 339.725000 108.170000 341.020000 113.550000 ;
      RECT 339.810000 146.790000 340.700000 147.135000 ;
      RECT 339.810000 148.365000 340.700000 151.055000 ;
      RECT 339.810000 152.475000 340.700000 157.925000 ;
      RECT 339.815000 143.905000 340.665000 146.790000 ;
      RECT 339.815000 147.135000 340.665000 148.365000 ;
      RECT 339.815000 151.055000 340.665000 152.475000 ;
      RECT 339.815000 157.925000 340.665000 159.150000 ;
      RECT 339.905000  36.580000 362.530000  36.590000 ;
      RECT 340.005000  31.155000 349.895000  31.325000 ;
      RECT 340.005000  32.335000 349.895000  32.505000 ;
      RECT 340.005000  33.515000 349.895000  33.685000 ;
      RECT 340.005000  34.695000 349.895000  34.865000 ;
      RECT 340.005000  35.875000 349.895000  36.045000 ;
      RECT 340.015000 128.205000 340.665000 143.735000 ;
      RECT 340.300000 222.080000 341.150000 245.255000 ;
      RECT 340.470000  77.050000 340.670000  80.860000 ;
      RECT 340.485000  76.400000 340.655000  77.050000 ;
      RECT 340.485000  80.860000 340.655000  81.150000 ;
      RECT 340.710000  81.555000 345.550000  81.835000 ;
      RECT 340.890000  16.720000 341.895000  16.890000 ;
      RECT 341.100000  85.710000 342.420000  95.620000 ;
      RECT 341.100000 116.900000 342.420000 126.810000 ;
      RECT 341.140000 167.875000 343.470000 168.225000 ;
      RECT 341.140000 168.225000 347.185000 168.395000 ;
      RECT 341.140000 168.395000 343.470000 169.785000 ;
      RECT 341.140000 169.785000 347.185000 169.955000 ;
      RECT 341.140000 169.955000 343.470000 171.345000 ;
      RECT 341.140000 171.345000 347.185000 171.515000 ;
      RECT 341.140000 171.515000 343.470000 172.905000 ;
      RECT 341.140000 172.905000 347.185000 173.485000 ;
      RECT 341.140000 173.485000 344.275000 174.055000 ;
      RECT 341.140000 174.055000 347.185000 174.835000 ;
      RECT 341.140000 174.835000 371.945000 176.430000 ;
      RECT 341.195000   4.620000 341.845000   4.950000 ;
      RECT 341.195000   5.250000 341.845000   5.580000 ;
      RECT 341.195000   5.880000 341.845000   6.210000 ;
      RECT 341.195000   6.510000 341.845000   6.840000 ;
      RECT 341.195000   7.140000 341.845000   7.470000 ;
      RECT 341.195000   7.770000 341.845000   8.100000 ;
      RECT 341.195000   8.400000 341.845000   8.730000 ;
      RECT 341.195000   9.030000 341.845000   9.360000 ;
      RECT 341.195000   9.660000 341.845000   9.990000 ;
      RECT 341.195000  15.095000 341.895000  15.265000 ;
      RECT 341.195000  18.120000 341.895000  18.290000 ;
      RECT 341.195000  22.635000 341.845000  22.965000 ;
      RECT 341.195000  23.265000 341.845000  23.595000 ;
      RECT 341.195000  23.895000 341.845000  24.225000 ;
      RECT 341.195000  24.525000 341.845000  24.855000 ;
      RECT 341.195000  25.155000 341.845000  25.485000 ;
      RECT 341.195000  25.785000 341.845000  26.115000 ;
      RECT 341.195000  26.415000 341.845000  26.745000 ;
      RECT 341.195000  27.045000 341.845000  27.375000 ;
      RECT 341.195000  27.675000 341.845000  28.005000 ;
      RECT 341.305000  13.705000 341.895000  13.875000 ;
      RECT 341.400000  44.025000 341.930000  44.195000 ;
      RECT 341.400000  44.640000 341.930000  44.810000 ;
      RECT 341.400000  45.270000 341.930000  45.440000 ;
      RECT 341.410000  43.945000 341.920000  44.025000 ;
      RECT 341.410000  44.195000 341.920000  44.275000 ;
      RECT 341.410000  44.575000 341.920000  44.640000 ;
      RECT 341.410000  44.810000 341.920000  44.905000 ;
      RECT 341.410000  45.205000 341.920000  45.270000 ;
      RECT 341.410000  45.440000 341.920000  45.535000 ;
      RECT 341.420000  16.655000 341.895000  16.720000 ;
      RECT 341.420000  16.890000 341.895000  17.325000 ;
      RECT 341.430000 129.450000 356.680000 129.620000 ;
      RECT 341.430000 129.620000 341.600000 131.490000 ;
      RECT 341.430000 131.490000 356.680000 131.660000 ;
      RECT 341.430000 131.660000 341.600000 147.335000 ;
      RECT 341.430000 147.335000 344.935000 147.505000 ;
      RECT 341.430000 147.505000 341.600000 150.925000 ;
      RECT 341.430000 150.925000 344.660000 151.095000 ;
      RECT 341.430000 151.095000 341.600000 152.685000 ;
      RECT 341.430000 152.685000 344.660000 152.855000 ;
      RECT 341.430000 152.855000 341.600000 158.215000 ;
      RECT 341.430000 158.215000 349.790000 158.590000 ;
      RECT 341.580000 186.475000 341.765000 187.000000 ;
      RECT 341.580000 187.000000 341.750000 187.005000 ;
      RECT 341.580000 188.140000 341.765000 188.670000 ;
      RECT 341.580000 189.880000 341.765000 190.410000 ;
      RECT 341.580000 191.620000 341.765000 192.150000 ;
      RECT 341.595000 186.330000 341.765000 186.475000 ;
      RECT 341.595000 188.070000 341.765000 188.140000 ;
      RECT 341.595000 188.670000 341.765000 188.740000 ;
      RECT 341.595000 189.810000 341.765000 189.880000 ;
      RECT 341.595000 190.410000 341.765000 190.480000 ;
      RECT 341.595000 191.550000 341.765000 191.620000 ;
      RECT 341.595000 192.150000 341.765000 192.220000 ;
      RECT 341.725000  11.865000 342.670000  12.535000 ;
      RECT 341.725000  13.665000 341.895000  13.705000 ;
      RECT 341.725000  13.875000 341.895000  14.335000 ;
      RECT 341.725000  14.845000 341.895000  15.095000 ;
      RECT 341.725000  15.265000 341.895000  15.515000 ;
      RECT 341.725000  17.835000 341.895000  18.120000 ;
      RECT 341.725000  18.290000 341.895000  18.505000 ;
      RECT 341.725000  19.635000 342.670000  20.305000 ;
      RECT 341.750000  77.110000 341.950000  80.920000 ;
      RECT 341.765000  76.400000 341.935000  77.110000 ;
      RECT 341.765000  80.920000 341.935000  81.555000 ;
      RECT 341.940000 154.515000 344.990000 154.685000 ;
      RECT 341.940000 154.685000 342.110000 156.075000 ;
      RECT 341.940000 156.075000 344.990000 156.245000 ;
      RECT 341.940000 156.245000 342.110000 157.635000 ;
      RECT 341.940000 157.635000 344.990000 157.805000 ;
      RECT 341.950000 143.300000 342.960000 143.795000 ;
      RECT 341.950000 145.905000 342.960000 146.075000 ;
      RECT 341.950000 146.455000 344.785000 146.625000 ;
      RECT 341.950000 148.215000 344.660000 148.385000 ;
      RECT 341.950000 149.095000 344.785000 149.265000 ;
      RECT 341.950000 149.645000 344.785000 149.815000 ;
      RECT 341.950000 151.805000 344.660000 151.975000 ;
      RECT 341.950000 153.965000 344.660000 154.135000 ;
      RECT 341.955000 185.670000 342.805000 187.450000 ;
      RECT 341.955000 187.620000 342.805000 189.190000 ;
      RECT 341.955000 189.360000 342.805000 190.930000 ;
      RECT 341.955000 191.100000 342.805000 192.815000 ;
      RECT 342.130000 132.010000 342.300000 141.970000 ;
      RECT 342.150000 220.085000 346.520000 247.105000 ;
      RECT 342.165000 142.270000 355.755000 142.440000 ;
      RECT 342.280000 155.295000 344.990000 155.465000 ;
      RECT 342.280000 156.855000 344.990000 157.025000 ;
      RECT 342.375000  67.005000 343.085000  67.255000 ;
      RECT 342.425000  99.140000 342.595000 103.890000 ;
      RECT 342.425000 108.340000 342.595000 113.090000 ;
      RECT 342.455000  66.965000 342.625000  67.005000 ;
      RECT 342.455000  67.255000 342.625000  67.295000 ;
      RECT 342.475000  85.370000 346.475000  85.540000 ;
      RECT 342.475000  95.920000 346.475000  96.090000 ;
      RECT 342.475000 116.430000 346.475000 116.600000 ;
      RECT 342.475000 126.980000 346.475000 127.150000 ;
      RECT 342.490000   4.190000 342.670000   5.235000 ;
      RECT 342.490000   5.235000 358.705000   5.415000 ;
      RECT 342.490000   5.415000 342.670000  10.480000 ;
      RECT 342.490000  10.990000 342.670000  11.865000 ;
      RECT 342.490000  12.535000 342.670000  19.635000 ;
      RECT 342.490000  20.305000 342.670000  21.175000 ;
      RECT 342.490000  21.685000 342.670000  28.375000 ;
      RECT 342.590000  85.540000 346.360000  95.920000 ;
      RECT 342.650000  98.800000 346.650000  98.970000 ;
      RECT 342.650000 104.350000 346.650000 104.520000 ;
      RECT 342.650000 108.000000 346.650000 108.170000 ;
      RECT 342.650000 113.550000 346.650000 113.720000 ;
      RECT 342.720000 116.600000 346.360000 126.980000 ;
      RECT 342.850000 142.930000 343.380000 143.100000 ;
      RECT 343.030000  77.050000 343.230000  80.860000 ;
      RECT 343.045000  76.400000 343.215000  77.050000 ;
      RECT 343.045000  80.860000 343.215000  81.150000 ;
      RECT 343.090000 163.295000 347.545000 163.625000 ;
      RECT 343.090000 164.015000 347.545000 164.345000 ;
      RECT 343.090000 164.735000 347.545000 164.815000 ;
      RECT 343.090000 164.815000 350.065000 164.985000 ;
      RECT 343.090000 164.985000 347.545000 165.065000 ;
      RECT 343.090000 165.455000 347.545000 165.785000 ;
      RECT 343.090000 166.175000 347.545000 166.505000 ;
      RECT 343.090000 166.895000 347.545000 166.955000 ;
      RECT 343.090000 166.955000 350.345000 167.125000 ;
      RECT 343.090000 167.125000 347.545000 167.225000 ;
      RECT 343.210000 143.100000 343.380000 145.850000 ;
      RECT 343.270000   6.340000 343.440000  16.190000 ;
      RECT 343.270000  17.340000 343.440000  27.190000 ;
      RECT 343.405000   3.925000 343.950000   4.595000 ;
      RECT 343.565000 182.950000 344.705000 196.425000 ;
      RECT 343.615000   5.815000 344.285000   5.985000 ;
      RECT 343.615000  27.400000 344.285000  27.900000 ;
      RECT 343.750000 144.010000 343.920000 144.405000 ;
      RECT 343.750000 144.405000 348.890000 144.575000 ;
      RECT 343.750000 144.575000 345.550000 145.440000 ;
      RECT 343.885000  59.635000 345.235000  59.885000 ;
      RECT 343.925000  65.035000 344.635000  65.285000 ;
      RECT 343.965000  59.595000 344.175000  59.635000 ;
      RECT 343.965000  59.885000 344.175000  59.925000 ;
      RECT 344.005000  64.995000 344.175000  65.035000 ;
      RECT 344.005000  65.285000 344.175000  65.325000 ;
      RECT 344.005000  98.970000 345.300000 104.350000 ;
      RECT 344.005000 108.170000 345.300000 113.550000 ;
      RECT 344.140000 143.300000 348.890000 143.795000 ;
      RECT 344.310000  77.110000 344.510000  80.920000 ;
      RECT 344.325000  76.400000 344.495000  77.110000 ;
      RECT 344.325000  80.920000 344.495000  81.555000 ;
      RECT 344.410000 132.010000 344.580000 141.860000 ;
      RECT 344.450000   6.340000 344.620000  16.190000 ;
      RECT 344.450000  17.340000 344.620000  27.190000 ;
      RECT 344.475000 169.005000 347.565000 169.175000 ;
      RECT 344.475000 170.565000 347.565000 170.735000 ;
      RECT 344.475000 172.125000 347.565000 172.295000 ;
      RECT 344.475000 173.685000 347.565000 173.855000 ;
      RECT 344.485000 200.645000 348.425000 203.475000 ;
      RECT 344.485000 203.475000 371.140000 204.335000 ;
      RECT 344.485000 204.335000 348.425000 215.530000 ;
      RECT 344.630000 215.530000 348.425000 215.970000 ;
      RECT 344.790000 152.320000 345.380000 152.490000 ;
      RECT 344.795000   5.820000 345.465000   5.990000 ;
      RECT 344.795000  27.400000 345.465000  27.900000 ;
      RECT 344.850000 148.350000 345.380000 148.520000 ;
      RECT 344.865000 153.765000 345.395000 153.935000 ;
      RECT 345.065000  58.960000 355.455000  59.000000 ;
      RECT 345.065000  59.000000 345.235000  59.635000 ;
      RECT 345.065000  59.885000 345.235000  60.035000 ;
      RECT 345.065000  60.035000 355.455000  62.505000 ;
      RECT 345.065000  62.505000 345.235000  63.355000 ;
      RECT 345.065000  63.355000 355.455000  63.565000 ;
      RECT 345.065000  63.565000 355.470000  66.305000 ;
      RECT 345.065000  66.305000 363.050000  68.100000 ;
      RECT 345.210000 146.610000 345.380000 147.335000 ;
      RECT 345.210000 147.335000 345.740000 147.505000 ;
      RECT 345.210000 147.675000 345.380000 148.350000 ;
      RECT 345.210000 148.520000 345.380000 149.025000 ;
      RECT 345.210000 149.335000 345.920000 149.505000 ;
      RECT 345.210000 149.505000 345.380000 149.780000 ;
      RECT 345.210000 149.780000 345.405000 150.310000 ;
      RECT 345.210000 150.310000 345.380000 150.870000 ;
      RECT 345.210000 151.960000 345.380000 152.320000 ;
      RECT 345.210000 152.490000 345.380000 152.630000 ;
      RECT 345.210000 153.240000 345.380000 153.765000 ;
      RECT 345.210000 154.870000 345.920000 155.540000 ;
      RECT 345.210000 155.540000 345.380000 157.580000 ;
      RECT 345.300000  46.875000 346.795000  51.195000 ;
      RECT 345.300000  51.195000 353.860000  54.460000 ;
      RECT 345.440000 151.455000 345.970000 151.625000 ;
      RECT 345.470000 177.450000 346.320000 184.190000 ;
      RECT 345.470000 184.190000 348.425000 200.645000 ;
      RECT 345.480000   3.925000 346.135000   4.595000 ;
      RECT 345.570000  77.050000 345.775000  80.250000 ;
      RECT 345.605000  76.400000 345.775000  77.050000 ;
      RECT 345.605000  80.250000 345.775000  81.150000 ;
      RECT 345.630000   6.340000 345.800000  16.190000 ;
      RECT 345.630000  17.340000 345.800000  27.190000 ;
      RECT 345.750000 145.285000 346.340000 145.455000 ;
      RECT 345.750000 145.455000 345.970000 146.960000 ;
      RECT 345.750000 147.840000 345.920000 149.335000 ;
      RECT 345.750000 149.850000 345.920000 150.575000 ;
      RECT 345.750000 150.575000 348.850000 150.745000 ;
      RECT 345.750000 151.200000 345.920000 151.455000 ;
      RECT 345.750000 151.625000 345.920000 154.590000 ;
      RECT 345.750000 156.300000 345.920000 157.250000 ;
      RECT 345.750000 157.250000 346.280000 157.420000 ;
      RECT 345.750000 157.420000 345.920000 157.650000 ;
      RECT 345.830000  81.610000 346.540000  81.780000 ;
      RECT 345.955000  59.795000 346.125000  60.035000 ;
      RECT 345.985000  80.880000 346.155000  81.610000 ;
      RECT 346.140000 145.725000 348.975000 145.895000 ;
      RECT 346.140000 146.605000 348.850000 146.775000 ;
      RECT 346.140000 147.485000 348.850000 147.655000 ;
      RECT 346.140000 148.365000 349.790000 148.535000 ;
      RECT 346.140000 149.245000 348.850000 149.415000 ;
      RECT 346.140000 149.795000 348.850000 149.965000 ;
      RECT 346.140000 151.455000 348.850000 151.625000 ;
      RECT 346.140000 152.335000 349.790000 152.505000 ;
      RECT 346.140000 153.215000 349.140000 153.385000 ;
      RECT 346.140000 153.765000 348.920000 153.935000 ;
      RECT 346.140000 154.645000 349.790000 154.815000 ;
      RECT 346.140000 155.525000 349.150000 155.695000 ;
      RECT 346.180000  59.435000 354.460000  59.605000 ;
      RECT 346.185000 156.075000 349.180000 156.245000 ;
      RECT 346.315000  59.390000 354.400000  59.435000 ;
      RECT 346.370000  77.110000 346.570000  80.650000 ;
      RECT 346.385000  76.400000 346.555000  77.110000 ;
      RECT 346.385000  80.650000 346.555000  81.150000 ;
      RECT 346.470000 156.855000 349.180000 157.025000 ;
      RECT 346.470000 157.635000 349.180000 157.805000 ;
      RECT 346.530000  85.710000 346.700000  95.560000 ;
      RECT 346.530000 116.960000 346.700000 126.810000 ;
      RECT 346.635000   5.415000 346.805000  28.375000 ;
      RECT 346.690000 132.010000 346.860000 141.970000 ;
      RECT 346.705000  99.140000 346.875000 103.890000 ;
      RECT 346.705000 108.340000 346.875000 113.090000 ;
      RECT 346.755000  85.370000 350.755000  85.540000 ;
      RECT 346.755000  95.920000 350.755000  96.090000 ;
      RECT 346.755000 116.430000 350.755000 116.600000 ;
      RECT 346.755000 126.980000 350.755000 127.150000 ;
      RECT 346.870000  85.540000 350.640000  95.920000 ;
      RECT 346.930000  98.800000 350.930000  98.970000 ;
      RECT 346.930000 104.350000 350.930000 104.520000 ;
      RECT 346.930000 108.000000 350.930000 108.170000 ;
      RECT 346.930000 113.550000 350.930000 113.720000 ;
      RECT 346.950000  77.110000 347.150000  80.650000 ;
      RECT 346.965000  76.050000 347.135000  77.110000 ;
      RECT 346.965000  80.650000 347.135000  82.020000 ;
      RECT 346.965000 163.625000 347.545000 164.015000 ;
      RECT 346.965000 165.785000 347.545000 166.175000 ;
      RECT 346.965000 178.435000 347.495000 178.605000 ;
      RECT 347.000000 116.600000 350.640000 126.980000 ;
      RECT 347.085000 176.430000 347.255000 178.435000 ;
      RECT 347.085000 178.605000 347.255000 183.390000 ;
      RECT 347.155000   6.305000 347.325000   6.500000 ;
      RECT 347.155000   6.500000 347.440000   9.840000 ;
      RECT 347.155000   9.840000 347.325000  23.580000 ;
      RECT 347.155000  23.580000 347.440000  26.920000 ;
      RECT 347.155000  26.920000 347.325000  27.115000 ;
      RECT 347.335000   3.925000 348.020000   4.595000 ;
      RECT 347.395000 168.825000 347.565000 169.005000 ;
      RECT 347.395000 169.175000 347.565000 169.355000 ;
      RECT 347.395000 170.385000 347.565000 170.565000 ;
      RECT 347.395000 170.735000 347.565000 170.915000 ;
      RECT 347.395000 171.945000 347.565000 172.125000 ;
      RECT 347.395000 172.295000 347.565000 172.475000 ;
      RECT 347.395000 173.505000 347.565000 173.685000 ;
      RECT 347.395000 173.855000 347.565000 174.465000 ;
      RECT 347.395000 174.465000 351.015000 174.635000 ;
      RECT 347.425000 168.075000 351.015000 168.245000 ;
      RECT 347.575000 215.970000 348.425000 225.590000 ;
      RECT 347.575000 225.590000 371.140000 226.440000 ;
      RECT 347.575000 226.440000 348.425000 248.525000 ;
      RECT 347.575000 248.525000 364.855000 249.375000 ;
      RECT 347.575000 249.375000 348.425000 252.535000 ;
      RECT 347.665000 177.270000 347.835000 179.980000 ;
      RECT 347.665000 180.740000 347.835000 183.450000 ;
      RECT 347.695000  44.015000 348.225000  44.185000 ;
      RECT 347.695000  44.640000 348.225000  44.810000 ;
      RECT 347.695000  45.270000 348.225000  45.440000 ;
      RECT 347.705000  43.945000 348.215000  44.015000 ;
      RECT 347.705000  44.185000 348.215000  44.275000 ;
      RECT 347.705000  44.575000 348.215000  44.640000 ;
      RECT 347.705000  44.810000 348.215000  44.905000 ;
      RECT 347.705000  45.205000 348.215000  45.270000 ;
      RECT 347.705000  45.440000 348.215000  45.535000 ;
      RECT 347.735000 168.580000 347.905000 170.540000 ;
      RECT 347.735000 170.540000 352.415000 170.740000 ;
      RECT 347.735000 170.740000 347.905000 171.290000 ;
      RECT 347.735000 171.570000 347.905000 174.080000 ;
      RECT 347.735000 174.080000 351.685000 174.280000 ;
      RECT 347.815000 162.900000 348.085000 163.570000 ;
      RECT 347.815000 163.570000 347.985000 164.100000 ;
      RECT 347.815000 165.410000 348.085000 166.080000 ;
      RECT 347.875000   5.945000 350.585000   6.115000 ;
      RECT 347.875000  10.225000 350.585000  10.395000 ;
      RECT 347.875000  11.505000 350.585000  11.675000 ;
      RECT 347.875000  12.785000 350.585000  12.955000 ;
      RECT 347.875000  14.065000 350.585000  14.235000 ;
      RECT 347.875000  15.345000 350.585000  15.515000 ;
      RECT 347.875000  16.625000 350.585000  16.795000 ;
      RECT 347.875000  17.905000 350.585000  18.075000 ;
      RECT 347.875000  19.185000 350.585000  19.355000 ;
      RECT 347.875000  20.465000 350.585000  20.635000 ;
      RECT 347.875000  21.745000 350.585000  21.915000 ;
      RECT 347.875000  23.025000 350.585000  23.195000 ;
      RECT 347.875000  27.305000 350.585000  27.475000 ;
      RECT 347.890000 176.600000 354.400000 176.770000 ;
      RECT 347.890000 176.770000 352.930000 176.800000 ;
      RECT 347.890000 183.620000 354.400000 183.790000 ;
      RECT 347.895000  75.120000 348.750000  82.955000 ;
      RECT 348.080000  47.935000 354.305000  48.105000 ;
      RECT 348.080000  48.105000 348.250000  48.825000 ;
      RECT 348.080000  49.185000 348.250000  49.955000 ;
      RECT 348.080000  49.955000 354.305000  50.125000 ;
      RECT 348.195000  50.125000 354.305000  50.135000 ;
      RECT 348.285000  98.970000 349.580000 104.350000 ;
      RECT 348.285000 108.170000 349.580000 113.550000 ;
      RECT 348.305000 162.845000 351.015000 163.015000 ;
      RECT 348.305000 163.625000 351.015000 163.795000 ;
      RECT 348.305000 164.305000 352.545000 164.575000 ;
      RECT 348.305000 165.185000 351.015000 165.355000 ;
      RECT 348.305000 165.830000 356.575000 166.070000 ;
      RECT 348.305000 166.070000 351.015000 166.135000 ;
      RECT 348.305000 166.515000 351.015000 166.580000 ;
      RECT 348.305000 166.580000 356.575000 166.785000 ;
      RECT 348.305000 167.295000 351.015000 167.465000 ;
      RECT 348.305000 168.855000 351.015000 169.025000 ;
      RECT 348.305000 169.635000 351.325000 169.970000 ;
      RECT 348.305000 170.140000 355.775000 170.310000 ;
      RECT 348.305000 170.310000 351.015000 170.355000 ;
      RECT 348.305000 171.065000 351.015000 171.235000 ;
      RECT 348.305000 173.585000 351.015000 173.755000 ;
      RECT 348.445000 177.270000 348.615000 180.150000 ;
      RECT 348.445000 180.150000 351.735000 180.570000 ;
      RECT 348.445000 180.570000 348.615000 183.450000 ;
      RECT 348.600000 171.555000 349.005000 171.885000 ;
      RECT 348.600000 171.885000 348.770000 172.935000 ;
      RECT 348.600000 172.935000 349.005000 173.265000 ;
      RECT 348.790000  47.905000 354.305000  47.935000 ;
      RECT 348.790000  48.415000 353.540000  48.585000 ;
      RECT 348.790000  48.945000 353.540000  49.115000 ;
      RECT 348.790000  49.465000 353.495000  49.475000 ;
      RECT 348.790000  49.475000 353.540000  49.645000 ;
      RECT 348.940000 172.415000 349.610000 172.575000 ;
      RECT 348.940000 172.575000 351.300000 172.745000 ;
      RECT 348.970000 132.010000 349.140000 141.860000 ;
      RECT 349.100000   2.335000 349.630000   2.505000 ;
      RECT 349.110000   2.235000 349.620000   2.335000 ;
      RECT 349.110000   2.505000 349.620000   2.905000 ;
      RECT 349.185000 184.215000 362.055000 186.105000 ;
      RECT 349.185000 186.105000 385.370000 186.695000 ;
      RECT 349.185000 186.695000 353.925000 192.515000 ;
      RECT 349.185000 192.515000 355.960000 195.580000 ;
      RECT 349.185000 195.580000 385.370000 202.215000 ;
      RECT 349.185000 202.215000 443.295000 202.710000 ;
      RECT 349.185000 205.100000 369.515000 205.120000 ;
      RECT 349.185000 205.120000 369.520000 206.330000 ;
      RECT 349.185000 206.330000 352.875000 217.345000 ;
      RECT 349.185000 217.345000 352.475000 223.550000 ;
      RECT 349.185000 223.550000 369.515000 224.820000 ;
      RECT 349.185000 250.140000 382.945000 253.385000 ;
      RECT 349.225000 177.270000 349.395000 179.980000 ;
      RECT 349.225000 180.740000 349.395000 183.450000 ;
      RECT 349.375000   3.925000 350.150000   4.595000 ;
      RECT 349.440000 205.070000 352.875000 205.100000 ;
      RECT 349.505000 171.235000 349.675000 171.655000 ;
      RECT 349.520000 227.595000 362.855000 228.345000 ;
      RECT 349.520000 228.345000 350.270000 246.620000 ;
      RECT 349.520000 246.620000 362.855000 247.375000 ;
      RECT 349.620000 142.950000 356.680000 143.120000 ;
      RECT 349.620000 143.120000 349.790000 148.365000 ;
      RECT 349.620000 148.535000 349.790000 152.335000 ;
      RECT 349.620000 152.505000 349.790000 154.645000 ;
      RECT 349.620000 154.815000 349.790000 158.215000 ;
      RECT 349.990000 173.165000 350.160000 173.585000 ;
      RECT 350.005000 177.270000 350.175000 180.150000 ;
      RECT 350.005000 180.570000 350.175000 183.450000 ;
      RECT 350.145000  31.485000 350.315000  32.155000 ;
      RECT 350.145000  32.665000 350.315000  33.335000 ;
      RECT 350.145000  33.845000 350.315000  34.515000 ;
      RECT 350.145000  35.025000 350.315000  35.695000 ;
      RECT 350.235000  59.795000 350.405000  60.035000 ;
      RECT 350.380000 172.935000 354.870000 173.060000 ;
      RECT 350.380000 173.060000 351.815000 173.265000 ;
      RECT 350.385000  14.955000 350.975000  15.125000 ;
      RECT 350.385000  15.735000 350.975000  15.905000 ;
      RECT 350.385000  17.515000 350.975000  17.685000 ;
      RECT 350.385000  18.295000 350.975000  18.465000 ;
      RECT 350.390000 172.075000 351.060000 172.405000 ;
      RECT 350.440000 164.815000 352.895000 164.985000 ;
      RECT 350.535000 147.070000 351.425000 147.600000 ;
      RECT 350.535000 148.365000 351.425000 149.940000 ;
      RECT 350.535000 150.570000 351.425000 151.610000 ;
      RECT 350.535000 152.350000 351.425000 154.015000 ;
      RECT 350.555000 143.885000 358.295000 145.100000 ;
      RECT 350.555000 145.100000 351.405000 147.070000 ;
      RECT 350.555000 147.600000 351.405000 148.365000 ;
      RECT 350.555000 149.940000 351.405000 150.570000 ;
      RECT 350.555000 151.610000 351.405000 152.350000 ;
      RECT 350.555000 154.015000 351.405000 159.150000 ;
      RECT 350.650000 171.555000 351.815000 171.885000 ;
      RECT 350.735000 166.785000 356.575000 166.795000 ;
      RECT 350.740000 167.665000 352.895000 167.835000 ;
      RECT 350.785000 177.270000 350.955000 179.980000 ;
      RECT 350.785000 180.740000 350.955000 183.450000 ;
      RECT 350.805000   6.305000 350.975000  14.955000 ;
      RECT 350.805000  15.125000 350.975000  15.735000 ;
      RECT 350.805000  15.905000 350.975000  17.515000 ;
      RECT 350.805000  17.685000 350.975000  18.295000 ;
      RECT 350.805000  18.465000 350.975000  27.115000 ;
      RECT 350.810000  85.710000 352.130000  95.620000 ;
      RECT 350.810000 116.900000 352.130000 126.810000 ;
      RECT 350.985000  99.140000 351.155000 103.890000 ;
      RECT 350.985000 108.340000 351.155000 113.090000 ;
      RECT 351.025000  31.485000 351.195000  32.155000 ;
      RECT 351.025000  32.665000 351.195000  33.335000 ;
      RECT 351.025000  33.845000 351.195000  34.515000 ;
      RECT 351.025000  35.025000 351.195000  35.695000 ;
      RECT 351.085000 229.105000 361.380000 229.275000 ;
      RECT 351.085000 229.275000 351.260000 245.690000 ;
      RECT 351.085000 245.690000 361.380000 245.865000 ;
      RECT 351.130000   3.925000 351.825000   4.595000 ;
      RECT 351.210000  98.800000 355.210000  98.970000 ;
      RECT 351.210000 104.350000 355.210000 104.520000 ;
      RECT 351.210000 108.000000 355.210000 108.170000 ;
      RECT 351.210000 113.550000 355.210000 113.720000 ;
      RECT 351.250000 132.010000 351.420000 141.970000 ;
      RECT 351.485000 163.965000 352.155000 164.135000 ;
      RECT 351.485000 166.990000 352.415000 167.160000 ;
      RECT 351.485000 168.515000 352.155000 168.685000 ;
      RECT 351.485000 169.160000 352.415000 169.330000 ;
      RECT 351.485000 170.915000 351.815000 171.285000 ;
      RECT 351.485000 171.285000 354.590000 171.455000 ;
      RECT 351.485000 171.455000 351.815000 171.555000 ;
      RECT 351.485000 172.890000 354.870000 172.935000 ;
      RECT 351.485000 173.265000 351.815000 173.850000 ;
      RECT 351.485000 174.280000 351.685000 174.405000 ;
      RECT 351.485000 174.405000 368.960000 174.605000 ;
      RECT 351.525000   5.930000 353.970000   5.945000 ;
      RECT 351.525000   5.945000 354.235000   6.115000 ;
      RECT 351.525000   6.115000 353.970000  10.225000 ;
      RECT 351.525000  10.225000 354.235000  10.395000 ;
      RECT 351.525000  10.395000 353.970000  11.505000 ;
      RECT 351.525000  11.505000 354.235000  11.675000 ;
      RECT 351.525000  11.675000 353.970000  12.785000 ;
      RECT 351.525000  12.785000 354.235000  12.955000 ;
      RECT 351.525000  14.065000 354.235000  14.235000 ;
      RECT 351.525000  15.345000 354.235000  15.515000 ;
      RECT 351.525000  16.625000 354.235000  16.795000 ;
      RECT 351.525000  17.905000 354.235000  18.075000 ;
      RECT 351.525000  19.185000 354.235000  19.355000 ;
      RECT 351.525000  20.465000 354.235000  20.635000 ;
      RECT 351.525000  21.745000 354.235000  21.915000 ;
      RECT 351.525000  21.915000 353.910000  23.025000 ;
      RECT 351.525000  23.025000 354.235000  23.195000 ;
      RECT 351.525000  23.195000 353.910000  27.305000 ;
      RECT 351.525000  27.305000 354.235000  27.475000 ;
      RECT 351.565000 169.635000 351.945000 169.970000 ;
      RECT 351.565000 177.270000 351.735000 180.150000 ;
      RECT 351.565000 180.570000 351.735000 183.450000 ;
      RECT 351.570000 230.095000 351.740000 245.125000 ;
      RECT 351.595000  31.155000 361.485000  31.325000 ;
      RECT 351.595000  32.335000 361.485000  32.505000 ;
      RECT 351.595000  33.515000 361.485000  33.685000 ;
      RECT 351.595000  34.695000 361.485000  34.865000 ;
      RECT 351.595000  35.875000 361.485000  36.045000 ;
      RECT 351.700000  73.985000 354.110000  74.155000 ;
      RECT 351.700000  74.155000 351.870000  80.160000 ;
      RECT 351.700000  80.160000 354.110000  80.360000 ;
      RECT 351.710000 229.695000 353.160000 229.865000 ;
      RECT 351.855000 174.020000 370.250000 174.220000 ;
      RECT 351.955000 162.445000 369.460000 162.645000 ;
      RECT 351.955000 162.645000 352.155000 163.965000 ;
      RECT 351.965000 168.155000 352.135000 168.515000 ;
      RECT 352.180000  74.405000 352.350000  79.155000 ;
      RECT 352.185000  85.370000 356.185000  85.540000 ;
      RECT 352.185000  95.920000 356.185000  96.090000 ;
      RECT 352.185000 116.430000 356.185000 116.600000 ;
      RECT 352.185000 126.980000 356.185000 127.150000 ;
      RECT 352.245000 166.965000 352.415000 166.990000 ;
      RECT 352.245000 167.160000 352.415000 167.495000 ;
      RECT 352.245000 168.930000 352.415000 169.160000 ;
      RECT 352.245000 169.330000 352.415000 169.595000 ;
      RECT 352.245000 170.740000 352.415000 171.115000 ;
      RECT 352.245000 173.260000 363.520000 173.460000 ;
      RECT 352.245000 173.460000 352.415000 173.790000 ;
      RECT 352.300000  85.540000 356.070000  95.920000 ;
      RECT 352.300000 116.600000 356.070000 126.980000 ;
      RECT 352.345000 177.270000 352.515000 179.980000 ;
      RECT 352.345000 180.740000 352.515000 183.450000 ;
      RECT 352.350000 230.175000 352.520000 245.125000 ;
      RECT 352.475000  79.665000 353.285000  79.835000 ;
      RECT 352.535000 168.020000 352.865000 168.575000 ;
      RECT 352.565000  98.970000 353.860000 104.350000 ;
      RECT 352.565000 108.170000 353.860000 113.550000 ;
      RECT 352.565000 163.175000 352.895000 163.730000 ;
      RECT 352.565000 166.240000 360.260000 166.410000 ;
      RECT 352.725000 164.985000 352.895000 165.090000 ;
      RECT 352.725000 165.090000 356.970000 165.260000 ;
      RECT 352.725000 167.390000 356.970000 167.560000 ;
      RECT 352.725000 167.560000 352.895000 167.665000 ;
      RECT 352.870000 130.030000 355.585000 130.200000 ;
      RECT 352.870000 130.910000 355.585000 131.080000 ;
      RECT 352.895000 177.270000 353.065000 179.980000 ;
      RECT 352.895000 180.740000 353.065000 183.450000 ;
      RECT 353.065000 163.120000 356.025000 163.290000 ;
      RECT 353.065000 163.900000 355.775000 164.070000 ;
      RECT 353.065000 164.680000 356.025000 164.850000 ;
      RECT 353.065000 165.460000 355.775000 165.630000 ;
      RECT 353.065000 167.020000 355.775000 167.190000 ;
      RECT 353.065000 167.800000 356.025000 167.970000 ;
      RECT 353.065000 168.580000 355.775000 168.750000 ;
      RECT 353.065000 169.360000 356.025000 169.530000 ;
      RECT 353.065000 170.920000 356.025000 171.090000 ;
      RECT 353.065000 171.700000 355.775000 171.870000 ;
      RECT 353.065000 172.480000 356.025000 172.650000 ;
      RECT 353.130000 230.095000 353.300000 245.125000 ;
      RECT 353.170000   3.925000 356.475000   4.595000 ;
      RECT 353.265000 163.885000 353.795000 163.900000 ;
      RECT 353.325000 207.860000 367.365000 208.335000 ;
      RECT 353.325000 208.335000 367.555000 209.185000 ;
      RECT 353.325000 209.185000 354.515000 213.440000 ;
      RECT 353.325000 213.440000 367.555000 213.950000 ;
      RECT 353.325000 213.950000 354.515000 218.195000 ;
      RECT 353.325000 218.195000 354.705000 218.200000 ;
      RECT 353.325000 218.200000 367.555000 219.330000 ;
      RECT 353.325000 219.330000 367.525000 219.390000 ;
      RECT 353.335000 173.630000 356.045000 173.800000 ;
      RECT 353.460000  74.405000 353.630000  79.155000 ;
      RECT 353.530000 132.010000 353.700000 141.860000 ;
      RECT 353.610000 229.275000 353.780000 245.690000 ;
      RECT 353.650000  54.670000 353.860000  58.790000 ;
      RECT 353.675000 177.270000 353.845000 183.450000 ;
      RECT 353.760000  48.640000 353.930000  49.420000 ;
      RECT 353.800000  45.835000 355.510000  46.165000 ;
      RECT 353.910000  43.280000 363.370000  43.610000 ;
      RECT 353.910000  43.610000 354.590000  44.275000 ;
      RECT 353.920000  44.575000 354.590000  45.535000 ;
      RECT 353.940000  74.155000 354.110000  80.160000 ;
      RECT 354.035000  14.955000 354.625000  15.125000 ;
      RECT 354.035000  15.735000 354.625000  15.905000 ;
      RECT 354.035000  17.515000 354.625000  17.685000 ;
      RECT 354.035000  18.295000 354.625000  18.465000 ;
      RECT 354.090000 230.095000 354.260000 245.125000 ;
      RECT 354.130000  48.105000 354.305000  49.955000 ;
      RECT 354.230000 229.695000 355.680000 229.865000 ;
      RECT 354.280000 163.460000 357.440000 163.730000 ;
      RECT 354.280000 168.920000 357.440000 169.190000 ;
      RECT 354.355000 147.710000 369.515000 147.880000 ;
      RECT 354.355000 147.880000 354.525000 159.775000 ;
      RECT 354.355000 159.775000 369.515000 159.945000 ;
      RECT 354.415000 147.690000 369.515000 147.710000 ;
      RECT 354.455000   6.305000 354.625000  10.035000 ;
      RECT 354.455000  13.175000 354.625000  14.955000 ;
      RECT 354.455000  15.125000 354.625000  15.735000 ;
      RECT 354.455000  15.905000 354.625000  17.515000 ;
      RECT 354.455000  17.685000 354.625000  18.295000 ;
      RECT 354.455000  18.465000 354.625000  27.115000 ;
      RECT 354.455000 177.270000 354.625000 179.980000 ;
      RECT 354.455000 180.740000 354.625000 183.450000 ;
      RECT 354.515000  59.795000 354.685000  60.035000 ;
      RECT 354.675000  73.725000 355.955000  76.640000 ;
      RECT 354.675000  76.640000 356.795000  78.760000 ;
      RECT 354.675000  78.760000 366.875000  78.930000 ;
      RECT 354.675000  78.930000 366.815000  79.190000 ;
      RECT 354.675000  79.190000 366.875000  79.595000 ;
      RECT 354.795000 178.435000 355.325000 178.605000 ;
      RECT 354.870000 230.175000 355.040000 245.125000 ;
      RECT 354.925000 214.380000 355.095000 217.340000 ;
      RECT 354.935000 148.790000 355.105000 151.500000 ;
      RECT 354.935000 152.010000 355.105000 154.720000 ;
      RECT 354.935000 155.975000 355.105000 156.345000 ;
      RECT 354.935000 156.345000 355.465000 156.875000 ;
      RECT 354.935000 156.875000 355.105000 158.880000 ;
      RECT 355.010000 155.270000 361.120000 155.440000 ;
      RECT 355.035000 176.430000 355.205000 178.435000 ;
      RECT 355.035000 178.605000 355.205000 183.390000 ;
      RECT 355.050000  43.980000 364.060000  44.145000 ;
      RECT 355.050000  44.145000 363.915000  44.150000 ;
      RECT 355.050000  44.150000 355.510000  45.835000 ;
      RECT 355.050000  46.165000 355.510000  46.705000 ;
      RECT 355.105000  79.595000 366.875000  82.420000 ;
      RECT 355.150000 217.560000 357.430000 217.730000 ;
      RECT 355.155000 148.070000 367.385000 148.240000 ;
      RECT 355.160000 159.100000 356.850000 159.270000 ;
      RECT 355.175000   5.945000 357.885000   6.115000 ;
      RECT 355.175000  10.225000 357.885000  10.395000 ;
      RECT 355.175000  11.505000 357.885000  11.675000 ;
      RECT 355.175000  12.785000 357.885000  12.955000 ;
      RECT 355.175000  14.065000 357.885000  14.235000 ;
      RECT 355.175000  15.345000 357.885000  15.515000 ;
      RECT 355.175000  16.625000 357.885000  16.795000 ;
      RECT 355.175000  17.905000 357.885000  18.075000 ;
      RECT 355.175000  19.185000 357.885000  19.355000 ;
      RECT 355.175000  20.465000 357.885000  20.635000 ;
      RECT 355.175000  21.745000 357.885000  21.915000 ;
      RECT 355.175000  23.025000 357.885000  23.195000 ;
      RECT 355.175000  27.305000 357.885000  27.475000 ;
      RECT 355.245000  59.000000 355.455000  60.035000 ;
      RECT 355.245000  62.505000 355.455000  63.355000 ;
      RECT 355.265000  99.140000 355.435000 103.890000 ;
      RECT 355.265000 108.340000 355.435000 113.090000 ;
      RECT 355.585000  98.800000 356.215000  98.970000 ;
      RECT 355.585000 104.350000 356.215000 104.520000 ;
      RECT 355.585000 108.000000 356.215000 108.170000 ;
      RECT 355.585000 113.550000 356.215000 113.720000 ;
      RECT 355.625000 130.400000 356.255000 130.570000 ;
      RECT 355.650000 230.095000 355.820000 245.125000 ;
      RECT 355.665000  98.970000 355.835000 104.350000 ;
      RECT 355.665000 108.170000 355.835000 113.550000 ;
      RECT 355.715000 148.630000 355.885000 151.500000 ;
      RECT 355.715000 151.670000 360.565000 151.840000 ;
      RECT 355.715000 151.840000 355.885000 154.735000 ;
      RECT 355.810000 132.010000 355.980000 141.970000 ;
      RECT 356.045000  98.970000 356.215000 101.080000 ;
      RECT 356.045000 101.080000 356.225000 101.970000 ;
      RECT 356.045000 101.970000 356.215000 104.350000 ;
      RECT 356.045000 108.170000 356.215000 110.280000 ;
      RECT 356.045000 110.280000 356.225000 111.170000 ;
      RECT 356.045000 111.170000 356.215000 113.550000 ;
      RECT 356.085000 130.240000 356.255000 130.400000 ;
      RECT 356.085000 130.570000 356.255000 130.910000 ;
      RECT 356.085000 177.155000 356.255000 178.205000 ;
      RECT 356.085000 178.435000 356.255000 178.765000 ;
      RECT 356.085000 179.385000 356.255000 179.715000 ;
      RECT 356.085000 179.885000 356.255000 182.595000 ;
      RECT 356.130000 229.275000 356.300000 245.690000 ;
      RECT 356.205000 214.630000 356.375000 217.340000 ;
      RECT 356.215000 155.830000 358.145000 156.000000 ;
      RECT 356.215000 156.000000 356.385000 158.880000 ;
      RECT 356.220000 190.940000 356.805000 191.110000 ;
      RECT 356.240000  85.710000 357.090000  89.620000 ;
      RECT 356.240000  89.620000 357.130000  94.495000 ;
      RECT 356.240000  94.495000 357.090000  95.620000 ;
      RECT 356.240000 116.900000 357.090000 118.025000 ;
      RECT 356.240000 118.025000 357.130000 122.900000 ;
      RECT 356.240000 122.900000 357.090000 126.810000 ;
      RECT 356.245000 165.560000 358.690000 165.830000 ;
      RECT 356.245000 166.795000 356.575000 166.820000 ;
      RECT 356.245000 166.820000 358.690000 167.090000 ;
      RECT 356.325000 172.415000 357.410000 172.560000 ;
      RECT 356.325000 172.560000 357.580000 172.745000 ;
      RECT 356.355000 176.655000 356.865000 176.985000 ;
      RECT 356.355000 183.065000 356.865000 183.395000 ;
      RECT 356.375000 217.730000 357.370000 217.735000 ;
      RECT 356.425000 176.985000 356.795000 183.065000 ;
      RECT 356.495000 148.790000 356.665000 151.500000 ;
      RECT 356.495000 152.010000 356.665000 154.720000 ;
      RECT 356.510000 129.620000 356.680000 131.490000 ;
      RECT 356.510000 131.660000 356.680000 142.950000 ;
      RECT 356.610000 230.095000 356.780000 245.125000 ;
      RECT 356.625000  73.910000 366.875000  74.080000 ;
      RECT 356.625000  74.080000 356.795000  75.580000 ;
      RECT 356.625000  98.560000 356.795000 104.760000 ;
      RECT 356.625000 107.760000 356.795000 113.960000 ;
      RECT 356.635000 190.360000 356.805000 190.940000 ;
      RECT 356.635000 191.110000 356.805000 191.370000 ;
      RECT 356.635000 192.220000 356.805000 193.230000 ;
      RECT 356.640000 164.425000 356.970000 165.090000 ;
      RECT 356.640000 167.560000 356.970000 168.225000 ;
      RECT 356.750000 229.695000 358.200000 229.865000 ;
      RECT 356.780000 169.850000 357.110000 169.920000 ;
      RECT 356.780000 169.920000 363.520000 170.290000 ;
      RECT 356.780000 170.290000 357.110000 170.360000 ;
      RECT 356.780000 170.730000 357.110000 170.800000 ;
      RECT 356.780000 170.800000 363.860000 171.170000 ;
      RECT 356.780000 171.170000 357.110000 171.240000 ;
      RECT 356.780000 171.610000 357.110000 171.680000 ;
      RECT 356.780000 171.680000 363.520000 171.820000 ;
      RECT 356.780000 171.820000 366.710000 171.990000 ;
      RECT 356.780000 171.990000 363.520000 172.050000 ;
      RECT 356.780000 172.050000 357.110000 172.120000 ;
      RECT 356.780000 173.040000 357.110000 173.110000 ;
      RECT 356.780000 173.110000 363.520000 173.260000 ;
      RECT 356.780000 173.460000 363.520000 173.480000 ;
      RECT 356.780000 173.480000 357.110000 173.550000 ;
      RECT 356.860000 191.620000 360.860000 191.790000 ;
      RECT 356.860000 193.480000 360.860000 193.650000 ;
      RECT 356.885000  46.800000 363.165000  46.970000 ;
      RECT 356.885000  46.970000 357.055000  50.370000 ;
      RECT 356.885000  50.370000 360.030000  50.540000 ;
      RECT 356.885000  50.540000 357.055000  53.175000 ;
      RECT 356.885000  53.175000 364.905000  53.265000 ;
      RECT 356.885000  53.265000 364.875000  53.345000 ;
      RECT 356.920000  95.620000 357.090000  95.730000 ;
      RECT 356.920000 116.790000 357.090000 116.900000 ;
      RECT 356.965000 177.155000 357.135000 182.900000 ;
      RECT 357.060000 219.390000 367.525000 219.455000 ;
      RECT 357.095000 156.170000 357.265000 159.045000 ;
      RECT 357.095000 159.045000 357.625000 159.575000 ;
      RECT 357.110000 163.450000 357.440000 163.460000 ;
      RECT 357.110000 163.730000 357.440000 163.960000 ;
      RECT 357.110000 166.070000 360.260000 166.240000 ;
      RECT 357.110000 166.410000 360.260000 166.580000 ;
      RECT 357.110000 168.690000 357.440000 168.920000 ;
      RECT 357.110000 169.190000 357.440000 169.200000 ;
      RECT 357.155000 209.680000 357.325000 210.690000 ;
      RECT 357.155000 212.185000 357.325000 212.915000 ;
      RECT 357.205000  74.590000 357.375000  75.600000 ;
      RECT 357.205000  76.650000 357.375000  77.660000 ;
      RECT 357.235000 176.655000 358.625000 176.985000 ;
      RECT 357.235000 183.065000 358.625000 183.395000 ;
      RECT 357.275000 148.630000 357.445000 151.500000 ;
      RECT 357.275000 151.840000 357.445000 154.735000 ;
      RECT 357.275000 169.500000 363.860000 169.670000 ;
      RECT 357.275000 169.670000 363.020000 169.750000 ;
      RECT 357.275000 171.340000 362.895000 171.510000 ;
      RECT 357.275000 172.745000 357.580000 172.770000 ;
      RECT 357.275000 172.770000 363.020000 172.940000 ;
      RECT 357.305000 176.985000 357.675000 183.065000 ;
      RECT 357.310000 211.785000 357.980000 211.955000 ;
      RECT 357.340000  56.030000 363.035000  56.200000 ;
      RECT 357.340000  56.200000 357.510000  64.455000 ;
      RECT 357.340000  64.455000 363.035000  64.625000 ;
      RECT 357.380000 210.910000 358.860000 211.080000 ;
      RECT 357.390000 230.175000 357.560000 245.125000 ;
      RECT 357.445000 128.205000 358.295000 143.885000 ;
      RECT 357.485000 214.380000 357.655000 217.340000 ;
      RECT 357.510000  48.245000 357.680000  49.740000 ;
      RECT 357.580000 170.460000 360.290000 170.630000 ;
      RECT 357.580000 172.220000 360.290000 172.390000 ;
      RECT 357.580000 173.650000 360.290000 173.820000 ;
      RECT 357.710000 217.560000 359.990000 217.730000 ;
      RECT 357.735000  47.675000 360.515000  47.845000 ;
      RECT 357.845000 177.155000 358.015000 178.205000 ;
      RECT 357.845000 178.435000 358.015000 178.765000 ;
      RECT 357.845000 179.385000 358.015000 179.715000 ;
      RECT 357.845000 179.885000 358.015000 182.595000 ;
      RECT 357.970000 164.015000 358.140000 165.025000 ;
      RECT 357.975000 156.000000 358.145000 158.880000 ;
      RECT 357.980000   6.500000 358.275000   9.840000 ;
      RECT 357.980000  23.580000 358.275000  26.920000 ;
      RECT 358.005000   3.925000 358.515000   4.595000 ;
      RECT 358.005000   6.305000 358.275000   6.500000 ;
      RECT 358.005000   9.840000 358.275000   9.915000 ;
      RECT 358.025000   2.235000 358.535000   2.905000 ;
      RECT 358.035000 209.680000 358.205000 210.690000 ;
      RECT 358.035000 212.245000 358.205000 213.115000 ;
      RECT 358.050000 217.730000 358.815000 217.735000 ;
      RECT 358.055000 148.790000 358.225000 151.500000 ;
      RECT 358.055000 152.010000 358.225000 154.720000 ;
      RECT 358.105000   9.915000 358.275000  10.035000 ;
      RECT 358.105000  10.605000 358.275000  12.565000 ;
      RECT 358.105000  13.165000 358.275000  20.525000 ;
      RECT 358.105000  21.155000 358.275000  21.575000 ;
      RECT 358.105000  21.575000 358.285000  22.110000 ;
      RECT 358.105000  22.110000 358.275000  22.505000 ;
      RECT 358.105000  23.385000 358.275000  23.580000 ;
      RECT 358.105000  26.920000 358.275000  27.115000 ;
      RECT 358.170000 230.095000 358.340000 245.125000 ;
      RECT 358.185000 176.985000 358.555000 183.065000 ;
      RECT 358.200000 159.100000 361.590000 159.270000 ;
      RECT 358.250000  57.920000 358.480000  63.485000 ;
      RECT 358.250000  63.485000 359.440000  63.515000 ;
      RECT 358.250000  63.515000 362.110000  63.685000 ;
      RECT 358.250000  63.685000 359.440000  63.715000 ;
      RECT 358.260000 211.785000 358.930000 211.955000 ;
      RECT 358.280000  56.945000 362.110000  57.175000 ;
      RECT 358.280000  57.175000 358.450000  57.920000 ;
      RECT 358.315000 158.675000 358.845000 159.100000 ;
      RECT 358.360000 163.450000 358.690000 165.560000 ;
      RECT 358.360000 167.090000 358.690000 169.200000 ;
      RECT 358.430000  84.825000 358.600000  96.855000 ;
      RECT 358.430000  97.145000 358.600000 106.160000 ;
      RECT 358.430000 106.360000 358.600000 115.375000 ;
      RECT 358.430000 115.675000 358.600000 127.885000 ;
      RECT 358.485000  74.590000 358.655000  77.660000 ;
      RECT 358.505000  15.485000 358.705000  16.910000 ;
      RECT 358.525000   5.415000 358.705000  15.485000 ;
      RECT 358.525000  16.910000 358.705000  28.375000 ;
      RECT 358.650000 229.275000 358.820000 245.690000 ;
      RECT 358.725000 177.155000 358.895000 182.900000 ;
      RECT 358.760000  57.980000 358.930000  62.830000 ;
      RECT 358.765000 214.630000 358.935000 217.340000 ;
      RECT 358.825000  75.820000 360.875000  75.990000 ;
      RECT 358.835000 148.630000 359.005000 151.500000 ;
      RECT 358.835000 151.840000 359.005000 154.735000 ;
      RECT 358.895000 156.455000 359.425000 156.985000 ;
      RECT 358.915000 209.680000 359.085000 210.690000 ;
      RECT 358.915000 212.245000 359.085000 213.115000 ;
      RECT 358.995000 176.655000 359.505000 176.985000 ;
      RECT 358.995000 183.065000 359.505000 183.395000 ;
      RECT 359.045000  50.540000 360.030000  50.820000 ;
      RECT 359.060000 134.865000 372.360000 141.545000 ;
      RECT 359.065000 176.985000 359.435000 183.065000 ;
      RECT 359.105000  76.620000 359.275000  77.970000 ;
      RECT 359.130000 230.095000 359.300000 245.125000 ;
      RECT 359.150000  57.400000 359.820000  57.570000 ;
      RECT 359.220000  57.390000 359.750000  57.400000 ;
      RECT 359.250000 163.270000 360.160000 164.105000 ;
      RECT 359.250000 164.105000 359.630000 164.690000 ;
      RECT 359.250000 165.100000 362.280000 165.270000 ;
      RECT 359.250000 165.980000 360.260000 166.070000 ;
      RECT 359.250000 166.580000 360.260000 167.030000 ;
      RECT 359.250000 167.030000 359.630000 167.740000 ;
      RECT 359.250000 167.980000 362.340000 168.150000 ;
      RECT 359.250000 168.150000 360.590000 168.320000 ;
      RECT 359.250000 168.670000 360.250000 169.030000 ;
      RECT 359.250000 169.030000 360.260000 169.200000 ;
      RECT 359.255000 156.170000 359.425000 156.455000 ;
      RECT 359.255000 156.985000 359.425000 158.880000 ;
      RECT 359.270000 229.695000 360.720000 229.865000 ;
      RECT 359.455000  78.350000 361.485000  78.520000 ;
      RECT 359.605000 177.155000 359.775000 178.205000 ;
      RECT 359.605000 178.435000 359.775000 178.765000 ;
      RECT 359.605000 179.385000 359.775000 179.715000 ;
      RECT 359.605000 179.885000 359.775000 182.595000 ;
      RECT 359.615000 148.790000 359.785000 151.500000 ;
      RECT 359.615000 152.010000 359.785000 154.720000 ;
      RECT 359.705000  51.305000 360.030000  52.535000 ;
      RECT 359.710000 209.185000 360.220000 213.440000 ;
      RECT 359.765000  74.590000 359.935000  75.600000 ;
      RECT 359.790000  48.245000 359.960000  49.740000 ;
      RECT 359.805000 156.170000 359.975000 158.880000 ;
      RECT 359.830000 164.360000 363.050000 164.530000 ;
      RECT 359.830000 164.530000 360.160000 164.720000 ;
      RECT 359.830000 167.385000 363.020000 167.555000 ;
      RECT 359.830000 167.555000 360.160000 167.810000 ;
      RECT 359.860000  50.820000 360.030000  51.305000 ;
      RECT 359.860000  52.535000 360.030000  53.095000 ;
      RECT 359.860000  53.095000 364.905000  53.175000 ;
      RECT 359.880000   0.930000 360.060000  28.185000 ;
      RECT 359.880000  28.185000 363.565000  28.365000 ;
      RECT 359.910000 230.175000 360.080000 245.125000 ;
      RECT 359.970000  86.645000 360.860000  88.205000 ;
      RECT 359.970000  89.825000 360.860000  94.985000 ;
      RECT 359.970000  97.085000 360.860000  99.415000 ;
      RECT 359.970000 103.775000 360.860000 108.215000 ;
      RECT 359.970000 112.835000 360.860000 115.480000 ;
      RECT 359.970000 117.405000 360.860000 122.700000 ;
      RECT 359.970000 125.500000 360.860000 127.655000 ;
      RECT 359.970000 128.425000 360.860000 129.725000 ;
      RECT 359.970000 130.805000 360.860000 134.385000 ;
      RECT 359.990000  84.410000 360.840000  86.645000 ;
      RECT 359.990000  88.205000 360.840000  89.825000 ;
      RECT 359.990000  94.985000 360.840000  97.085000 ;
      RECT 359.990000  99.415000 360.840000 103.775000 ;
      RECT 359.990000 108.215000 360.840000 112.835000 ;
      RECT 359.990000 115.480000 360.840000 117.405000 ;
      RECT 359.990000 122.700000 360.840000 125.500000 ;
      RECT 359.990000 127.655000 360.840000 128.425000 ;
      RECT 359.990000 129.725000 360.840000 130.805000 ;
      RECT 359.990000 134.385000 360.840000 134.865000 ;
      RECT 360.040000  58.080000 360.210000  62.830000 ;
      RECT 360.045000 214.380000 360.215000 217.340000 ;
      RECT 360.155000 177.155000 360.325000 182.900000 ;
      RECT 360.265000  74.590000 361.215000  74.760000 ;
      RECT 360.270000 217.560000 362.550000 217.730000 ;
      RECT 360.330000 217.730000 361.325000 217.735000 ;
      RECT 360.355000  50.575000 360.525000  51.925000 ;
      RECT 360.385000  52.230000 360.995000  52.400000 ;
      RECT 360.385000  76.620000 361.215000  76.790000 ;
      RECT 360.385000  76.790000 360.555000  77.970000 ;
      RECT 360.395000 148.630000 360.565000 151.500000 ;
      RECT 360.395000 151.840000 360.565000 154.735000 ;
      RECT 360.420000 168.320000 360.590000 168.540000 ;
      RECT 360.425000 176.655000 360.935000 176.985000 ;
      RECT 360.425000 183.065000 360.935000 183.395000 ;
      RECT 360.430000  57.400000 361.100000  57.570000 ;
      RECT 360.460000 170.460000 360.790000 170.630000 ;
      RECT 360.460000 173.650000 360.790000 173.820000 ;
      RECT 360.495000 176.985000 360.865000 183.065000 ;
      RECT 360.500000  57.390000 361.030000  57.400000 ;
      RECT 360.510000 163.530000 361.090000 163.705000 ;
      RECT 360.510000 163.705000 363.690000 163.875000 ;
      RECT 360.510000 163.875000 361.090000 164.060000 ;
      RECT 360.570000  48.245000 360.740000  49.595000 ;
      RECT 360.640000 164.530000 361.310000 164.890000 ;
      RECT 360.640000 167.555000 361.310000 167.670000 ;
      RECT 360.650000 187.400000 360.820000 188.070000 ;
      RECT 360.650000 188.350000 360.820000 189.020000 ;
      RECT 360.665000  52.195000 360.995000  52.230000 ;
      RECT 360.665000  52.400000 360.995000  52.845000 ;
      RECT 360.685000 155.945000 360.855000 158.880000 ;
      RECT 360.690000 230.095000 360.860000 245.125000 ;
      RECT 360.705000  75.120000 360.875000  75.820000 ;
      RECT 360.750000 165.270000 361.090000 165.720000 ;
      RECT 360.750000 165.720000 360.920000 167.145000 ;
      RECT 360.760000   2.965000 379.105000   3.135000 ;
      RECT 360.760000   3.135000 374.905000   3.665000 ;
      RECT 360.760000   3.665000 361.460000  13.725000 ;
      RECT 360.760000  13.725000 374.905000  14.425000 ;
      RECT 360.760000  16.045000 374.905000  16.245000 ;
      RECT 360.760000  16.245000 379.105000  16.415000 ;
      RECT 360.760000  16.415000 374.650000  16.745000 ;
      RECT 360.760000  16.745000 361.460000  26.805000 ;
      RECT 360.760000  26.805000 374.650000  27.505000 ;
      RECT 360.795000  47.675000 361.465000  47.845000 ;
      RECT 360.915000 190.360000 361.085000 191.370000 ;
      RECT 360.915000 192.220000 361.085000 193.230000 ;
      RECT 360.960000  47.845000 361.130000  48.780000 ;
      RECT 361.015000  77.070000 361.185000  78.350000 ;
      RECT 361.035000 177.155000 361.205000 178.205000 ;
      RECT 361.035000 178.435000 361.205000 178.765000 ;
      RECT 361.035000 179.385000 361.205000 179.715000 ;
      RECT 361.035000 179.885000 361.205000 182.595000 ;
      RECT 361.040000 187.245000 363.965000 187.415000 ;
      RECT 361.040000 188.125000 364.000000 188.295000 ;
      RECT 361.040000 189.005000 363.750000 189.175000 ;
      RECT 361.045000  74.760000 361.215000  75.820000 ;
      RECT 361.045000  75.820000 362.115000  75.990000 ;
      RECT 361.045000  75.990000 361.215000  76.620000 ;
      RECT 361.120000 168.320000 362.990000 168.490000 ;
      RECT 361.135000  50.575000 361.305000  51.135000 ;
      RECT 361.135000  51.135000 361.325000  51.925000 ;
      RECT 361.140000 191.620000 369.140000 191.790000 ;
      RECT 361.140000 193.480000 369.140000 193.650000 ;
      RECT 361.150000 166.305000 361.320000 166.820000 ;
      RECT 361.150000 166.820000 363.690000 166.990000 ;
      RECT 361.155000  51.925000 361.325000  52.025000 ;
      RECT 361.170000 229.275000 361.380000 245.690000 ;
      RECT 361.175000 148.790000 361.345000 151.500000 ;
      RECT 361.175000 152.010000 361.345000 154.735000 ;
      RECT 361.200000 172.220000 363.020000 172.390000 ;
      RECT 361.210000 170.460000 361.785000 170.630000 ;
      RECT 361.210000 173.650000 361.740000 173.820000 ;
      RECT 361.285000 176.690000 361.815000 176.860000 ;
      RECT 361.290000  63.485000 362.110000  63.515000 ;
      RECT 361.290000  63.685000 362.110000  63.715000 ;
      RECT 361.305000 176.655000 361.815000 176.690000 ;
      RECT 361.305000 176.860000 361.815000 176.985000 ;
      RECT 361.305000 183.065000 361.815000 183.395000 ;
      RECT 361.320000  57.980000 361.490000  62.830000 ;
      RECT 361.325000 214.630000 361.495000 217.340000 ;
      RECT 361.350000  48.100000 361.520000  49.595000 ;
      RECT 361.375000 176.985000 361.745000 183.065000 ;
      RECT 361.445000  52.195000 361.775000  52.845000 ;
      RECT 361.490000 165.470000 362.990000 165.780000 ;
      RECT 361.490000 165.780000 361.740000 166.440000 ;
      RECT 361.565000 156.170000 361.735000 158.880000 ;
      RECT 361.575000  50.005000 363.420000  50.175000 ;
      RECT 361.595000 209.800000 361.765000 212.510000 ;
      RECT 361.635000  50.000000 363.340000  50.005000 ;
      RECT 361.645000  74.080000 361.815000  75.580000 ;
      RECT 361.665000  76.620000 361.835000  77.970000 ;
      RECT 361.715000 117.400000 361.915000 125.365000 ;
      RECT 361.715000 125.365000 371.155000 125.415000 ;
      RECT 361.715000 125.415000 363.940000 126.035000 ;
      RECT 361.715000 126.035000 363.910000 127.040000 ;
      RECT 361.715000 127.040000 363.940000 127.705000 ;
      RECT 361.715000 127.705000 371.155000 127.755000 ;
      RECT 361.715000 127.755000 361.915000 133.100000 ;
      RECT 361.720000 103.825000 361.915000 104.365000 ;
      RECT 361.720000 104.365000 363.445000 105.115000 ;
      RECT 361.720000 105.115000 361.915000 107.090000 ;
      RECT 361.720000 107.090000 363.445000 107.840000 ;
      RECT 361.720000 107.840000 361.915000 108.450000 ;
      RECT 361.725000 152.010000 361.895000 154.720000 ;
      RECT 361.735000  31.485000 361.905000  32.155000 ;
      RECT 361.735000  32.665000 361.905000  33.335000 ;
      RECT 361.735000  33.845000 361.905000  34.515000 ;
      RECT 361.735000  35.025000 361.905000  35.695000 ;
      RECT 361.745000  84.375000 371.155000  84.545000 ;
      RECT 361.745000  84.545000 361.915000 103.825000 ;
      RECT 361.745000 108.450000 361.915000 117.400000 ;
      RECT 361.745000 133.100000 361.915000 133.775000 ;
      RECT 361.745000 133.775000 371.155000 133.945000 ;
      RECT 361.760000 159.100000 362.290000 159.270000 ;
      RECT 361.820000 212.730000 363.300000 212.900000 ;
      RECT 361.880000  57.175000 362.110000  63.485000 ;
      RECT 361.880000 155.270000 362.550000 155.440000 ;
      RECT 361.905000 155.440000 362.115000 159.100000 ;
      RECT 361.905000 159.270000 362.115000 159.440000 ;
      RECT 361.915000  50.575000 362.085000  51.925000 ;
      RECT 361.915000 177.155000 362.085000 179.320000 ;
      RECT 361.915000 179.320000 362.340000 179.850000 ;
      RECT 361.915000 179.850000 362.085000 182.900000 ;
      RECT 361.945000  52.230000 362.555000  52.400000 ;
      RECT 361.950000 164.700000 362.340000 164.870000 ;
      RECT 361.950000 164.870000 362.280000 165.100000 ;
      RECT 361.955000 148.630000 362.125000 151.500000 ;
      RECT 361.955000 170.460000 363.020000 170.630000 ;
      RECT 361.970000 173.650000 363.020000 173.820000 ;
      RECT 361.985000  75.120000 362.455000  75.650000 ;
      RECT 362.000000 163.270000 363.050000 163.440000 ;
      RECT 362.000000 166.150000 363.020000 166.320000 ;
      RECT 362.000000 169.030000 362.890000 169.200000 ;
      RECT 362.010000 165.980000 363.020000 166.150000 ;
      RECT 362.010000 166.320000 363.020000 166.510000 ;
      RECT 362.010000 167.200000 363.020000 167.385000 ;
      RECT 362.010000 167.750000 362.340000 167.980000 ;
      RECT 362.015000  78.350000 364.045000  78.520000 ;
      RECT 362.040000 164.150000 363.050000 164.360000 ;
      RECT 362.105000  85.420000 362.275000  86.400000 ;
      RECT 362.105000 105.820000 362.275000 106.490000 ;
      RECT 362.105000 228.345000 362.855000 246.620000 ;
      RECT 362.130000  48.245000 362.300000  49.595000 ;
      RECT 362.170000 176.655000 363.120000 176.985000 ;
      RECT 362.220000   4.425000 366.595000   5.135000 ;
      RECT 362.220000   5.135000 362.920000  12.265000 ;
      RECT 362.220000  12.265000 366.595000  12.965000 ;
      RECT 362.220000  17.505000 366.595000  18.205000 ;
      RECT 362.220000  18.205000 362.920000  25.335000 ;
      RECT 362.220000  25.335000 366.595000  26.045000 ;
      RECT 362.225000  52.195000 362.555000  52.230000 ;
      RECT 362.225000  52.400000 362.555000  52.845000 ;
      RECT 362.225000  87.565000 362.395000  94.355000 ;
      RECT 362.225000  99.615000 362.950000  99.785000 ;
      RECT 362.225000  99.785000 362.395000 103.265000 ;
      RECT 362.225000 103.265000 362.950000 103.435000 ;
      RECT 362.225000 108.815000 362.395000 112.465000 ;
      RECT 362.225000 112.465000 362.950000 112.635000 ;
      RECT 362.225000 117.835000 362.395000 124.625000 ;
      RECT 362.225000 128.155000 362.395000 132.905000 ;
      RECT 362.285000  74.560000 362.455000  74.590000 ;
      RECT 362.285000  74.590000 363.235000  74.760000 ;
      RECT 362.285000  74.760000 362.455000  75.120000 ;
      RECT 362.285000  75.650000 362.455000  76.620000 ;
      RECT 362.285000  76.620000 363.115000  76.790000 ;
      RECT 362.315000  77.070000 362.485000  78.350000 ;
      RECT 362.360000  30.425000 362.530000  36.580000 ;
      RECT 362.360000  72.420000 372.185000  72.730000 ;
      RECT 362.445000 155.945000 362.615000 158.880000 ;
      RECT 362.450000  87.175000 370.450000  87.345000 ;
      RECT 362.450000  94.825000 370.450000  94.995000 ;
      RECT 362.450000 117.195000 370.450000 117.365000 ;
      RECT 362.450000 124.845000 370.450000 125.015000 ;
      RECT 362.450000 133.415000 363.120000 133.585000 ;
      RECT 362.465000 181.885000 363.885000 182.265000 ;
      RECT 362.465000 182.265000 363.300000 182.795000 ;
      RECT 362.465000 184.635000 362.635000 185.685000 ;
      RECT 362.475000 209.800000 362.645000 212.510000 ;
      RECT 362.490000 133.405000 363.060000 133.415000 ;
      RECT 362.495000  85.175000 365.205000  85.345000 ;
      RECT 362.495000  86.455000 365.205000  86.625000 ;
      RECT 362.510000 177.155000 362.680000 178.595000 ;
      RECT 362.510000 179.625000 362.710000 180.825000 ;
      RECT 362.510000 180.825000 362.680000 180.975000 ;
      RECT 362.540000 179.575000 362.710000 179.625000 ;
      RECT 362.565000  87.345000 370.305000  94.825000 ;
      RECT 362.565000 100.795000 363.175000 100.965000 ;
      RECT 362.565000 109.995000 363.175000 110.165000 ;
      RECT 362.565000 117.365000 370.305000 124.845000 ;
      RECT 362.605000 152.010000 362.775000 154.720000 ;
      RECT 362.605000 214.380000 362.775000 217.340000 ;
      RECT 362.615000 105.675000 363.285000 105.850000 ;
      RECT 362.615000 106.460000 363.285000 106.630000 ;
      RECT 362.645000  75.820000 364.675000  75.990000 ;
      RECT 362.695000  48.245000 362.865000  49.595000 ;
      RECT 362.695000  50.575000 362.865000  51.140000 ;
      RECT 362.695000  51.140000 362.885000  51.925000 ;
      RECT 362.700000  40.760000 363.370000  41.720000 ;
      RECT 362.700000  42.020000 363.370000  42.980000 ;
      RECT 362.715000  51.925000 362.885000  52.025000 ;
      RECT 362.725000 183.145000 363.255000 183.725000 ;
      RECT 362.735000 148.790000 362.905000 151.500000 ;
      RECT 362.735000 179.035000 363.900000 179.205000 ;
      RECT 362.795000 155.270000 363.465000 155.440000 ;
      RECT 362.820000 164.730000 362.990000 165.470000 ;
      RECT 362.820000 167.780000 362.990000 168.320000 ;
      RECT 362.830000 217.560000 365.110000 217.730000 ;
      RECT 362.850000 176.985000 363.120000 179.035000 ;
      RECT 362.865000  56.200000 363.035000  64.455000 ;
      RECT 362.900000 183.725000 363.070000 185.625000 ;
      RECT 362.945000  76.790000 363.115000  77.970000 ;
      RECT 362.995000  45.925000 364.905000  46.095000 ;
      RECT 362.995000  46.095000 363.165000  46.800000 ;
      RECT 363.005000  52.195000 363.335000  52.845000 ;
      RECT 363.005000 100.005000 363.175000 100.795000 ;
      RECT 363.005000 100.965000 363.175000 102.715000 ;
      RECT 363.005000 109.205000 363.175000 109.995000 ;
      RECT 363.005000 110.165000 363.175000 111.915000 ;
      RECT 363.035000  95.425000 363.985000  95.595000 ;
      RECT 363.035000  95.595000 363.205000  99.075000 ;
      RECT 363.035000  99.075000 363.985000  99.245000 ;
      RECT 363.035000 113.005000 363.985000 113.175000 ;
      RECT 363.035000 113.175000 363.205000 116.655000 ;
      RECT 363.035000 116.655000 363.985000 116.825000 ;
      RECT 363.105000 128.155000 363.275000 132.905000 ;
      RECT 363.190000 169.840000 363.520000 169.920000 ;
      RECT 363.190000 170.290000 363.520000 170.370000 ;
      RECT 363.190000 170.730000 363.860000 170.800000 ;
      RECT 363.190000 171.170000 363.860000 171.240000 ;
      RECT 363.190000 171.610000 363.520000 171.680000 ;
      RECT 363.190000 172.050000 363.520000 172.120000 ;
      RECT 363.190000 173.040000 363.520000 173.110000 ;
      RECT 363.190000 173.480000 363.520000 173.550000 ;
      RECT 363.235000 217.730000 364.230000 217.735000 ;
      RECT 363.290000 177.785000 365.100000 177.955000 ;
      RECT 363.290000 177.955000 363.460000 178.455000 ;
      RECT 363.290000 179.625000 363.460000 181.145000 ;
      RECT 363.290000 181.145000 365.020000 181.315000 ;
      RECT 363.295000 155.440000 363.465000 155.700000 ;
      RECT 363.295000 155.700000 363.925000 155.870000 ;
      RECT 363.325000 156.170000 363.495000 158.880000 ;
      RECT 363.330000 133.415000 370.090000 133.585000 ;
      RECT 363.345000  99.615000 364.115000  99.785000 ;
      RECT 363.345000 103.265000 364.115000 103.435000 ;
      RECT 363.345000 108.815000 364.115000 108.985000 ;
      RECT 363.345000 112.465000 364.115000 112.635000 ;
      RECT 363.345000 184.675000 363.725000 185.685000 ;
      RECT 363.355000 209.800000 363.525000 212.510000 ;
      RECT 363.385000  28.365000 363.565000  37.515000 ;
      RECT 363.390000 133.405000 370.090000 133.415000 ;
      RECT 363.395000   6.000000 363.935000  11.395000 ;
      RECT 363.395000  19.075000 363.935000  24.470000 ;
      RECT 363.425000  99.785000 364.035000  99.815000 ;
      RECT 363.425000 108.985000 364.035000 109.015000 ;
      RECT 363.475000  46.445000 363.645000  47.795000 ;
      RECT 363.475000  48.245000 363.645000  49.595000 ;
      RECT 363.475000  50.575000 363.645000  51.925000 ;
      RECT 363.485000 152.010000 363.655000 154.720000 ;
      RECT 363.515000 148.630000 363.685000 151.500000 ;
      RECT 363.520000 163.875000 363.690000 164.890000 ;
      RECT 363.520000 164.890000 370.275000 165.060000 ;
      RECT 363.520000 166.990000 363.690000 168.020000 ;
      RECT 363.520000 168.020000 364.360000 168.090000 ;
      RECT 363.520000 168.090000 370.770000 168.190000 ;
      RECT 363.555000 182.465000 363.915000 182.795000 ;
      RECT 363.555000 182.795000 363.725000 183.275000 ;
      RECT 363.555000 183.275000 364.085000 183.945000 ;
      RECT 363.555000 183.945000 363.725000 184.675000 ;
      RECT 363.565000  74.590000 363.735000  75.600000 ;
      RECT 363.580000 212.730000 364.250000 212.900000 ;
      RECT 363.690000 169.670000 363.860000 169.850000 ;
      RECT 363.690000 169.850000 364.360000 169.920000 ;
      RECT 363.690000 169.920000 370.770000 170.290000 ;
      RECT 363.690000 170.290000 364.360000 170.360000 ;
      RECT 363.690000 171.240000 363.860000 171.410000 ;
      RECT 363.690000 171.410000 366.710000 171.580000 ;
      RECT 363.700000  50.005000 364.370000  50.175000 ;
      RECT 363.710000 125.185000 370.075000 125.215000 ;
      RECT 363.710000 125.215000 371.155000 125.365000 ;
      RECT 363.710000 127.755000 371.155000 127.905000 ;
      RECT 363.710000 127.905000 370.075000 127.935000 ;
      RECT 363.710000 155.105000 364.720000 155.440000 ;
      RECT 363.740000   5.420000 365.065000   5.830000 ;
      RECT 363.740000  24.640000 365.065000  25.050000 ;
      RECT 363.745000  39.745000 364.060000  43.980000 ;
      RECT 363.755000 155.870000 363.925000 156.845000 ;
      RECT 363.765000 173.025000 364.360000 173.110000 ;
      RECT 363.765000 173.110000 371.125000 173.480000 ;
      RECT 363.765000 173.480000 364.360000 173.555000 ;
      RECT 363.770000 104.675000 363.940000 104.850000 ;
      RECT 363.770000 104.850000 369.590000 105.120000 ;
      RECT 363.770000 105.120000 363.940000 105.630000 ;
      RECT 363.770000 105.630000 369.590000 105.900000 ;
      RECT 363.770000 105.900000 363.940000 106.410000 ;
      RECT 363.770000 106.410000 369.590000 106.680000 ;
      RECT 363.770000 106.680000 363.940000 107.190000 ;
      RECT 363.770000 107.190000 369.590000 107.460000 ;
      RECT 363.770000 107.460000 363.940000 107.575000 ;
      RECT 363.785000  52.335000 364.115000  52.845000 ;
      RECT 363.815000  50.175000 364.080000  52.335000 ;
      RECT 363.815000  95.595000 363.985000  99.075000 ;
      RECT 363.815000 113.175000 363.985000 116.655000 ;
      RECT 363.855000  30.295000 365.110000  30.465000 ;
      RECT 363.855000  30.665000 365.470000  30.835000 ;
      RECT 363.885000 214.630000 364.055000 217.340000 ;
      RECT 363.895000 184.585000 364.465000 184.915000 ;
      RECT 363.895000 184.915000 364.065000 184.975000 ;
      RECT 363.925000 185.455000 364.975000 185.625000 ;
      RECT 363.985000 128.135000 364.155000 132.905000 ;
      RECT 364.005000 226.440000 371.140000 226.450000 ;
      RECT 364.005000 226.450000 364.855000 248.525000 ;
      RECT 364.030000 163.330000 364.360000 163.400000 ;
      RECT 364.030000 163.400000 370.770000 163.770000 ;
      RECT 364.030000 163.770000 365.580000 163.840000 ;
      RECT 364.030000 164.210000 364.360000 164.280000 ;
      RECT 364.030000 164.280000 370.770000 164.650000 ;
      RECT 364.030000 164.650000 364.360000 164.720000 ;
      RECT 364.030000 165.060000 364.360000 165.710000 ;
      RECT 364.030000 165.710000 370.770000 166.080000 ;
      RECT 364.030000 166.080000 364.360000 166.150000 ;
      RECT 364.030000 166.520000 364.360000 166.590000 ;
      RECT 364.030000 166.590000 370.770000 166.960000 ;
      RECT 364.030000 166.960000 364.360000 167.030000 ;
      RECT 364.030000 168.190000 370.770000 168.460000 ;
      RECT 364.030000 168.460000 364.360000 168.530000 ;
      RECT 364.030000 168.900000 364.360000 168.970000 ;
      RECT 364.030000 168.970000 370.770000 169.340000 ;
      RECT 364.030000 169.340000 364.360000 169.410000 ;
      RECT 364.030000 170.730000 364.360000 170.800000 ;
      RECT 364.030000 170.800000 370.770000 171.170000 ;
      RECT 364.030000 171.170000 364.360000 171.240000 ;
      RECT 364.030000 172.160000 364.360000 172.230000 ;
      RECT 364.030000 172.230000 370.770000 172.600000 ;
      RECT 364.030000 172.600000 364.360000 172.670000 ;
      RECT 364.070000 178.125000 364.240000 178.965000 ;
      RECT 364.070000 178.965000 365.595000 179.455000 ;
      RECT 364.070000 179.455000 364.240000 180.975000 ;
      RECT 364.155000  95.425000 364.925000  95.595000 ;
      RECT 364.155000  99.075000 368.765000  99.245000 ;
      RECT 364.155000 113.005000 368.765000 113.175000 ;
      RECT 364.155000 116.655000 364.925000 116.825000 ;
      RECT 364.160000 104.510000 369.130000 104.680000 ;
      RECT 364.160000 105.290000 369.120000 105.460000 ;
      RECT 364.160000 106.070000 369.130000 106.240000 ;
      RECT 364.160000 106.850000 369.120000 107.020000 ;
      RECT 364.160000 107.630000 369.130000 107.800000 ;
      RECT 364.190000 164.190000 364.360000 164.210000 ;
      RECT 364.225000  76.620000 364.395000  77.970000 ;
      RECT 364.235000  99.045000 364.845000  99.075000 ;
      RECT 364.235000 113.175000 364.845000 113.205000 ;
      RECT 364.235000 209.800000 364.405000 212.510000 ;
      RECT 364.255000  46.445000 364.425000  47.795000 ;
      RECT 364.255000  48.245000 364.425000  49.595000 ;
      RECT 364.255000  50.575000 364.425000  51.925000 ;
      RECT 364.285000  99.615000 365.395000  99.785000 ;
      RECT 364.285000  99.785000 364.455000 103.265000 ;
      RECT 364.285000 103.265000 365.390000 103.435000 ;
      RECT 364.285000 108.815000 365.395000 108.985000 ;
      RECT 364.285000 108.985000 364.455000 112.465000 ;
      RECT 364.285000 112.465000 365.390000 112.635000 ;
      RECT 364.295000 148.790000 364.465000 151.500000 ;
      RECT 364.295000 181.885000 364.465000 183.385000 ;
      RECT 364.295000 183.385000 366.340000 183.555000 ;
      RECT 364.295000 183.555000 364.915000 183.725000 ;
      RECT 364.295000 183.725000 364.465000 184.585000 ;
      RECT 364.365000 152.010000 364.535000 154.865000 ;
      RECT 364.450000 125.695000 369.200000 125.865000 ;
      RECT 364.450000 126.475000 369.200000 126.645000 ;
      RECT 364.450000 127.255000 369.200000 127.425000 ;
      RECT 364.455000  95.595000 364.625000  99.045000 ;
      RECT 364.455000 113.205000 364.625000 116.655000 ;
      RECT 364.530000 126.645000 369.120000 126.650000 ;
      RECT 364.530000 163.060000 370.275000 163.230000 ;
      RECT 364.530000 163.840000 365.580000 163.940000 ;
      RECT 364.530000 163.940000 366.140000 164.110000 ;
      RECT 364.530000 164.820000 370.275000 164.890000 ;
      RECT 364.530000 165.370000 370.275000 165.540000 ;
      RECT 364.530000 166.250000 366.140000 166.420000 ;
      RECT 364.530000 167.130000 370.275000 167.300000 ;
      RECT 364.530000 167.680000 366.140000 167.850000 ;
      RECT 364.530000 168.630000 369.000000 168.800000 ;
      RECT 364.530000 169.580000 366.140000 169.750000 ;
      RECT 364.530000 171.340000 366.710000 171.410000 ;
      RECT 364.530000 171.990000 366.710000 172.060000 ;
      RECT 364.530000 173.650000 366.140000 173.820000 ;
      RECT 364.550000 155.440000 364.720000 158.880000 ;
      RECT 364.565000 142.760000 368.865000 142.930000 ;
      RECT 364.565000 142.930000 364.735000 144.580000 ;
      RECT 364.565000 144.580000 368.865000 144.750000 ;
      RECT 364.655000 170.460000 370.275000 170.630000 ;
      RECT 364.655000 172.770000 370.275000 172.940000 ;
      RECT 364.665000 184.125000 365.635000 184.375000 ;
      RECT 364.665000 184.375000 364.975000 185.455000 ;
      RECT 364.705000 159.100000 365.375000 159.270000 ;
      RECT 364.735000  46.095000 364.905000  53.095000 ;
      RECT 364.790000  56.665000 372.355000  56.835000 ;
      RECT 364.790000  56.835000 364.960000  70.255000 ;
      RECT 364.790000  70.255000 372.355000  70.425000 ;
      RECT 364.845000  74.590000 365.015000  77.660000 ;
      RECT 364.850000 179.625000 365.020000 181.145000 ;
      RECT 364.865000 128.155000 365.035000 132.905000 ;
      RECT 364.870000   6.000000 365.410000  11.395000 ;
      RECT 364.870000  19.075000 365.410000  24.470000 ;
      RECT 364.930000 177.955000 365.100000 178.455000 ;
      RECT 364.940000  28.980000 368.250000  29.150000 ;
      RECT 364.940000  29.150000 365.110000  30.295000 ;
      RECT 364.985000 143.270000 365.515000 143.440000 ;
      RECT 364.985000 143.440000 365.155000 144.135000 ;
      RECT 365.005000 209.185000 367.555000 213.440000 ;
      RECT 365.075000 148.630000 365.245000 151.500000 ;
      RECT 365.095000  95.485000 365.265000  98.855000 ;
      RECT 365.095000 113.725000 365.265000 116.765000 ;
      RECT 365.165000 214.380000 365.335000 217.340000 ;
      RECT 365.175000 181.885000 366.935000 182.265000 ;
      RECT 365.175000 182.265000 366.225000 182.895000 ;
      RECT 365.175000 184.645000 365.705000 185.655000 ;
      RECT 365.245000 152.010000 365.415000 154.720000 ;
      RECT 365.300000  29.320000 367.460000  29.490000 ;
      RECT 365.300000  29.490000 365.470000  30.665000 ;
      RECT 365.315000 187.220000 365.485000 187.325000 ;
      RECT 365.315000 187.325000 365.885000 187.495000 ;
      RECT 365.315000 187.495000 365.485000 187.550000 ;
      RECT 365.345000 184.635000 365.515000 184.645000 ;
      RECT 365.430000 156.170000 365.600000 158.880000 ;
      RECT 365.435000  95.425000 366.205000  95.595000 ;
      RECT 365.435000 116.655000 366.205000 116.825000 ;
      RECT 365.435000 177.785000 366.615000 177.955000 ;
      RECT 365.435000 177.955000 365.620000 178.625000 ;
      RECT 365.435000 178.625000 365.935000 178.795000 ;
      RECT 365.470000 155.270000 368.860000 155.440000 ;
      RECT 365.480000 187.770000 369.630000 187.940000 ;
      RECT 365.515000  99.045000 366.125000  99.075000 ;
      RECT 365.515000 113.175000 366.125000 113.205000 ;
      RECT 365.560000 102.485000 365.735000 102.715000 ;
      RECT 365.560000 102.715000 365.730000 103.375000 ;
      RECT 365.560000 111.685000 365.735000 111.915000 ;
      RECT 365.560000 111.915000 365.730000 112.465000 ;
      RECT 365.560000 112.465000 366.675000 112.635000 ;
      RECT 365.565000  99.615000 366.675000  99.785000 ;
      RECT 365.565000  99.785000 365.735000 102.485000 ;
      RECT 365.565000 108.815000 366.675000 108.985000 ;
      RECT 365.565000 108.985000 365.735000 111.685000 ;
      RECT 365.565000 188.455000 365.735000 189.410000 ;
      RECT 365.625000 227.215000 382.945000 250.140000 ;
      RECT 365.655000 183.785000 366.185000 183.955000 ;
      RECT 365.670000  29.675000 375.340000  29.845000 ;
      RECT 365.670000  29.845000 365.840000  30.350000 ;
      RECT 365.670000  30.350000 365.965000  37.025000 ;
      RECT 365.670000  37.025000 365.840000  39.135000 ;
      RECT 365.670000  39.135000 365.965000  41.605000 ;
      RECT 365.670000  41.605000 375.340000  41.775000 ;
      RECT 365.670000  41.775000 365.965000  51.935000 ;
      RECT 365.670000  51.935000 365.840000  52.565000 ;
      RECT 365.670000  52.565000 365.965000  53.095000 ;
      RECT 365.670000  53.095000 374.155000  53.265000 ;
      RECT 365.705000 143.240000 368.455000 143.410000 ;
      RECT 365.705000 143.670000 368.415000 143.840000 ;
      RECT 365.705000 144.100000 368.455000 144.270000 ;
      RECT 365.735000  95.595000 365.905000  99.045000 ;
      RECT 365.735000 113.205000 365.905000 116.655000 ;
      RECT 365.745000 128.135000 365.915000 132.905000 ;
      RECT 365.765000 178.795000 365.935000 179.300000 ;
      RECT 365.765000 179.300000 366.005000 180.975000 ;
      RECT 365.790000 178.125000 366.275000 178.455000 ;
      RECT 365.790000 189.630000 367.790000 189.800000 ;
      RECT 365.825000  84.545000 371.155000  86.190000 ;
      RECT 365.850000 189.800000 367.720000 189.810000 ;
      RECT 365.855000 148.790000 366.025000 151.500000 ;
      RECT 365.860000 213.950000 367.555000 218.200000 ;
      RECT 365.895000   5.135000 366.595000  12.265000 ;
      RECT 365.895000  18.205000 366.595000  25.335000 ;
      RECT 365.905000 103.265000 366.675000 103.435000 ;
      RECT 366.015000 183.955000 366.185000 185.625000 ;
      RECT 366.105000 178.455000 366.275000 178.855000 ;
      RECT 366.105000 178.855000 366.415000 179.130000 ;
      RECT 366.125000  74.590000 366.295000  75.600000 ;
      RECT 366.125000  76.650000 366.295000  77.660000 ;
      RECT 366.125000 152.010000 366.295000 154.890000 ;
      RECT 366.125000 154.890000 368.060000 155.015000 ;
      RECT 366.125000 155.015000 368.055000 155.060000 ;
      RECT 366.175000 179.130000 366.415000 179.965000 ;
      RECT 366.175000 179.965000 366.525000 180.975000 ;
      RECT 366.250000  57.685000 366.420000  62.535000 ;
      RECT 366.250000  64.050000 366.420000  68.900000 ;
      RECT 366.265000  30.195000 366.435000  32.905000 ;
      RECT 366.265000  38.545000 366.435000  41.255000 ;
      RECT 366.345000  34.025000 366.515000  36.775000 ;
      RECT 366.350000 158.740000 366.880000 159.270000 ;
      RECT 366.375000  96.145000 366.545000  98.855000 ;
      RECT 366.375000 113.725000 366.545000 116.435000 ;
      RECT 366.395000 184.645000 366.750000 185.655000 ;
      RECT 366.405000  42.415000 366.575000  52.305000 ;
      RECT 366.420000  33.455000 367.090000  33.625000 ;
      RECT 366.420000  37.825000 367.090000  37.995000 ;
      RECT 366.445000 177.675000 366.615000 177.785000 ;
      RECT 366.445000 177.955000 366.615000 178.685000 ;
      RECT 366.560000 166.250000 367.090000 166.420000 ;
      RECT 366.560000 167.680000 367.090000 167.850000 ;
      RECT 366.560000 169.580000 367.090000 169.750000 ;
      RECT 366.560000 173.650000 367.090000 173.820000 ;
      RECT 366.570000  37.285000 367.570000  37.455000 ;
      RECT 366.580000 182.465000 367.005000 182.795000 ;
      RECT 366.580000 182.795000 366.750000 183.275000 ;
      RECT 366.580000 183.275000 366.865000 183.945000 ;
      RECT 366.580000 183.945000 366.750000 184.645000 ;
      RECT 366.585000 178.855000 367.095000 179.185000 ;
      RECT 366.620000  63.270000 367.290000  63.440000 ;
      RECT 366.625000 128.155000 366.795000 132.905000 ;
      RECT 366.630000  42.025000 367.415000  42.195000 ;
      RECT 366.630000  52.675000 367.415000  52.845000 ;
      RECT 366.635000 148.630000 366.805000 151.500000 ;
      RECT 366.650000 179.185000 366.845000 179.795000 ;
      RECT 366.650000 179.795000 366.860000 179.815000 ;
      RECT 366.650000 179.815000 366.870000 179.835000 ;
      RECT 366.650000 179.835000 366.885000 179.845000 ;
      RECT 366.665000 179.845000 366.890000 179.865000 ;
      RECT 366.675000 179.865000 366.890000 179.885000 ;
      RECT 366.695000 179.885000 366.890000 179.895000 ;
      RECT 366.695000 179.895000 367.885000 180.360000 ;
      RECT 366.705000  74.080000 366.875000  75.580000 ;
      RECT 366.705000  76.640000 366.875000  78.760000 ;
      RECT 366.710000 155.440000 366.880000 158.740000 ;
      RECT 366.715000  95.425000 367.485000  95.595000 ;
      RECT 366.715000 116.655000 367.485000 116.825000 ;
      RECT 366.760000 163.940000 367.090000 164.110000 ;
      RECT 366.800000  99.045000 367.410000  99.075000 ;
      RECT 366.800000 113.175000 367.410000 113.205000 ;
      RECT 366.805000  42.195000 367.355000  42.495000 ;
      RECT 366.845000  99.615000 367.955000  99.785000 ;
      RECT 366.845000  99.785000 367.015000 103.265000 ;
      RECT 366.845000 103.265000 367.955000 103.435000 ;
      RECT 366.845000 108.815000 367.955000 108.985000 ;
      RECT 366.845000 108.985000 367.015000 112.465000 ;
      RECT 366.845000 112.465000 367.955000 112.635000 ;
      RECT 367.005000 152.010000 367.175000 154.720000 ;
      RECT 367.015000 179.395000 367.525000 179.725000 ;
      RECT 367.020000  95.595000 367.190000  99.045000 ;
      RECT 367.020000 113.205000 367.190000 116.655000 ;
      RECT 367.135000 180.360000 367.885000 180.975000 ;
      RECT 367.145000  30.195000 367.315000  32.905000 ;
      RECT 367.145000  38.545000 367.315000  39.040000 ;
      RECT 367.145000  39.040000 367.320000  41.130000 ;
      RECT 367.145000  41.130000 367.315000  41.605000 ;
      RECT 367.225000 177.675000 367.525000 178.685000 ;
      RECT 367.260000 163.940000 369.970000 164.110000 ;
      RECT 367.260000 166.250000 369.970000 166.420000 ;
      RECT 367.260000 167.680000 370.275000 167.850000 ;
      RECT 367.260000 169.580000 369.970000 169.750000 ;
      RECT 367.260000 171.340000 369.970000 171.430000 ;
      RECT 367.260000 171.430000 371.935000 171.990000 ;
      RECT 367.260000 171.990000 369.970000 172.060000 ;
      RECT 367.260000 173.650000 369.970000 173.820000 ;
      RECT 367.265000 159.100000 367.935000 159.270000 ;
      RECT 367.265000 178.685000 367.525000 179.395000 ;
      RECT 367.300000 186.950000 367.830000 187.120000 ;
      RECT 367.355000   3.665000 368.055000  13.725000 ;
      RECT 367.355000  16.745000 368.055000  26.805000 ;
      RECT 367.365000 159.270000 367.895000 159.285000 ;
      RECT 367.370000  33.455000 368.850000  33.625000 ;
      RECT 367.370000  37.825000 368.850000  37.995000 ;
      RECT 367.415000 148.630000 367.585000 151.500000 ;
      RECT 367.485000  73.910000 369.875000  74.080000 ;
      RECT 367.485000  74.080000 367.655000  80.160000 ;
      RECT 367.485000  80.160000 369.875000  80.330000 ;
      RECT 367.505000 128.135000 367.675000 132.905000 ;
      RECT 367.515000 181.365000 371.945000 185.455000 ;
      RECT 367.530000  57.685000 367.700000  62.535000 ;
      RECT 367.530000  64.050000 367.700000  68.900000 ;
      RECT 367.540000 187.120000 367.820000 187.555000 ;
      RECT 367.585000  42.025000 368.710000  42.195000 ;
      RECT 367.585000  42.195000 367.755000  52.675000 ;
      RECT 367.585000  52.675000 368.710000  52.845000 ;
      RECT 367.625000  34.025000 367.795000  36.735000 ;
      RECT 367.655000  95.485000 367.825000  98.855000 ;
      RECT 367.655000 113.725000 367.825000 116.765000 ;
      RECT 367.680000 189.160000 368.210000 189.330000 ;
      RECT 367.715000 179.455000 367.885000 179.895000 ;
      RECT 367.720000  29.150000 368.250000  29.490000 ;
      RECT 367.725000 177.695000 371.945000 178.695000 ;
      RECT 367.800000 185.455000 371.945000 185.835000 ;
      RECT 367.800000 185.835000 385.370000 186.105000 ;
      RECT 367.825000  79.690000 369.050000  79.860000 ;
      RECT 367.845000 189.080000 368.015000 189.160000 ;
      RECT 367.845000 189.330000 368.015000 189.410000 ;
      RECT 367.850000  37.285000 368.850000  37.455000 ;
      RECT 367.885000 152.010000 368.055000 152.890000 ;
      RECT 367.885000 152.890000 368.060000 154.890000 ;
      RECT 367.900000  63.270000 369.850000  63.440000 ;
      RECT 367.920000  57.265000 368.590000  57.435000 ;
      RECT 367.920000  69.340000 368.590000  69.510000 ;
      RECT 367.980000 194.230000 368.150000 194.900000 ;
      RECT 367.990000 156.170000 368.160000 158.880000 ;
      RECT 367.995000  95.425000 368.765000  95.595000 ;
      RECT 367.995000 116.655000 368.765000 116.825000 ;
      RECT 368.025000  30.195000 368.260000  33.065000 ;
      RECT 368.025000  38.385000 368.290000  41.255000 ;
      RECT 368.065000  74.510000 368.235000  79.470000 ;
      RECT 368.075000  99.045000 368.685000  99.075000 ;
      RECT 368.075000 113.175000 368.685000 113.205000 ;
      RECT 368.125000  99.615000 369.235000  99.785000 ;
      RECT 368.125000  99.785000 368.295000 103.265000 ;
      RECT 368.125000 103.265000 369.235000 103.435000 ;
      RECT 368.125000 108.815000 369.235000 108.985000 ;
      RECT 368.125000 108.985000 368.295000 112.465000 ;
      RECT 368.125000 112.465000 369.235000 112.635000 ;
      RECT 368.225000 176.430000 371.945000 177.695000 ;
      RECT 368.225000 178.695000 371.945000 181.365000 ;
      RECT 368.295000  95.595000 368.465000  99.045000 ;
      RECT 368.295000 113.205000 368.465000 116.655000 ;
      RECT 368.315000 206.330000 369.520000 223.340000 ;
      RECT 368.315000 223.340000 369.515000 223.550000 ;
      RECT 368.370000 194.005000 369.380000 194.175000 ;
      RECT 368.370000 194.885000 369.380000 195.055000 ;
      RECT 368.385000 128.155000 368.555000 132.905000 ;
      RECT 368.480000 194.175000 369.325000 194.180000 ;
      RECT 368.545000  99.785000 369.155000  99.815000 ;
      RECT 368.545000 108.985000 369.155000 109.015000 ;
      RECT 368.595000  74.720000 368.765000  79.470000 ;
      RECT 368.695000 142.930000 368.865000 144.580000 ;
      RECT 368.765000  42.415000 368.935000  52.305000 ;
      RECT 368.765000 152.010000 368.935000 154.720000 ;
      RECT 368.805000 187.220000 370.045000 187.550000 ;
      RECT 368.810000  57.685000 368.980000  62.535000 ;
      RECT 368.810000  64.050000 368.980000  68.900000 ;
      RECT 368.815000   4.425000 373.190000   5.135000 ;
      RECT 368.815000   5.135000 369.515000  12.265000 ;
      RECT 368.815000  12.265000 373.190000  12.965000 ;
      RECT 368.815000  17.505000 373.190000  18.205000 ;
      RECT 368.815000  18.205000 369.515000  25.335000 ;
      RECT 368.815000  25.335000 373.190000  26.045000 ;
      RECT 368.870000 162.645000 369.460000 162.860000 ;
      RECT 368.905000  29.845000 375.340000  29.880000 ;
      RECT 368.905000  29.880000 369.670000  32.905000 ;
      RECT 368.905000  34.025000 369.670000  35.050000 ;
      RECT 368.905000  35.050000 375.340000  36.400000 ;
      RECT 368.905000  36.400000 369.670000  36.775000 ;
      RECT 368.905000  38.545000 369.670000  41.570000 ;
      RECT 368.905000  41.570000 375.340000  41.605000 ;
      RECT 368.935000  95.425000 369.885000  95.595000 ;
      RECT 368.935000  95.595000 369.105000  99.075000 ;
      RECT 368.935000  99.075000 369.885000  99.245000 ;
      RECT 368.935000 113.725000 369.105000 116.435000 ;
      RECT 368.990000  42.025000 370.115000  42.195000 ;
      RECT 368.990000  52.675000 370.115000  52.845000 ;
      RECT 369.125000  74.510000 369.295000  79.470000 ;
      RECT 369.160000 113.005000 369.985000 113.175000 ;
      RECT 369.160000 116.655000 369.830000 116.825000 ;
      RECT 369.195000 190.360000 369.365000 191.370000 ;
      RECT 369.195000 192.220000 369.365000 193.230000 ;
      RECT 369.200000  57.265000 369.870000  57.435000 ;
      RECT 369.200000  69.340000 369.870000  69.510000 ;
      RECT 369.265000 128.135000 369.435000 132.905000 ;
      RECT 369.345000 147.880000 369.515000 159.775000 ;
      RECT 369.375000 113.175000 369.545000 116.655000 ;
      RECT 369.405000  99.615000 370.355000  99.785000 ;
      RECT 369.405000  99.785000 369.575000 103.265000 ;
      RECT 369.405000 103.265000 370.355000 103.435000 ;
      RECT 369.405000 109.205000 369.575000 111.915000 ;
      RECT 369.420000 104.730000 369.590000 104.850000 ;
      RECT 369.420000 105.120000 369.590000 105.630000 ;
      RECT 369.420000 105.900000 369.590000 106.410000 ;
      RECT 369.420000 106.680000 369.590000 107.190000 ;
      RECT 369.420000 107.460000 369.590000 107.570000 ;
      RECT 369.420000 125.920000 369.590000 127.200000 ;
      RECT 369.500000  32.905000 369.670000  34.025000 ;
      RECT 369.500000  36.775000 369.670000  38.545000 ;
      RECT 369.630000 108.815000 370.300000 108.985000 ;
      RECT 369.705000  74.080000 369.875000  80.160000 ;
      RECT 369.715000  95.595000 369.885000  99.075000 ;
      RECT 369.715000 113.725000 369.885000 116.435000 ;
      RECT 369.750000 190.495000 370.000000 193.230000 ;
      RECT 369.775000 193.230000 369.945000 195.580000 ;
      RECT 369.815000 104.255000 371.155000 107.995000 ;
      RECT 369.815000 108.535000 369.985000 108.815000 ;
      RECT 369.815000 108.985000 369.985000 113.005000 ;
      RECT 369.845000 125.415000 371.155000 127.705000 ;
      RECT 369.945000  42.195000 370.115000  52.675000 ;
      RECT 370.000000   6.000000 370.540000  11.395000 ;
      RECT 370.000000  19.075000 370.540000  24.470000 ;
      RECT 370.090000  57.685000 370.260000  62.535000 ;
      RECT 370.090000  64.050000 370.260000  68.900000 ;
      RECT 370.145000 128.155000 370.315000 132.905000 ;
      RECT 370.185000  99.785000 370.355000 103.265000 ;
      RECT 370.185000 109.205000 370.355000 111.915000 ;
      RECT 370.280000 204.335000 371.140000 225.590000 ;
      RECT 370.330000 141.545000 372.360000 161.195000 ;
      RECT 370.345000   5.420000 371.670000   5.830000 ;
      RECT 370.345000  24.640000 371.670000  25.050000 ;
      RECT 370.435000  30.645000 374.405000  30.815000 ;
      RECT 370.435000  30.815000 370.605000  34.085000 ;
      RECT 370.440000 163.330000 370.770000 163.400000 ;
      RECT 370.440000 163.770000 370.770000 163.840000 ;
      RECT 370.440000 164.210000 370.770000 164.280000 ;
      RECT 370.440000 164.650000 370.770000 164.720000 ;
      RECT 370.440000 165.640000 370.770000 165.710000 ;
      RECT 370.440000 166.080000 370.770000 166.150000 ;
      RECT 370.440000 166.520000 370.770000 166.590000 ;
      RECT 370.440000 166.960000 370.770000 167.030000 ;
      RECT 370.440000 168.020000 370.770000 168.090000 ;
      RECT 370.440000 168.460000 370.770000 168.530000 ;
      RECT 370.440000 168.900000 370.770000 168.970000 ;
      RECT 370.440000 169.340000 370.770000 169.410000 ;
      RECT 370.440000 169.850000 370.770000 169.920000 ;
      RECT 370.440000 170.290000 370.770000 170.360000 ;
      RECT 370.440000 170.730000 370.770000 170.800000 ;
      RECT 370.440000 171.170000 370.770000 171.260000 ;
      RECT 370.440000 172.160000 370.770000 172.230000 ;
      RECT 370.440000 172.600000 370.770000 172.690000 ;
      RECT 370.440000 173.040000 371.125000 173.110000 ;
      RECT 370.440000 173.480000 371.125000 173.550000 ;
      RECT 370.460000  63.270000 371.130000  63.440000 ;
      RECT 370.475000  88.310000 370.675000  93.725000 ;
      RECT 370.475000 118.465000 370.675000 123.880000 ;
      RECT 370.490000  40.635000 374.405000  40.805000 ;
      RECT 370.505000  87.565000 370.675000  88.310000 ;
      RECT 370.505000  93.725000 370.675000  94.355000 ;
      RECT 370.505000 117.835000 370.675000 118.465000 ;
      RECT 370.505000 123.880000 370.675000 124.625000 ;
      RECT 370.530000 186.695000 385.370000 195.580000 ;
      RECT 370.665000  41.775000 371.675000  53.095000 ;
      RECT 370.915000  31.065000 371.085000  33.775000 ;
      RECT 370.915000  37.675000 371.085000  40.385000 ;
      RECT 370.940000 165.425000 371.935000 171.430000 ;
      RECT 370.940000 171.990000 371.935000 172.100000 ;
      RECT 370.955000 173.020000 371.125000 173.040000 ;
      RECT 370.985000  86.190000 371.155000 104.255000 ;
      RECT 370.985000 107.995000 371.155000 125.215000 ;
      RECT 370.985000 127.905000 371.155000 133.775000 ;
      RECT 371.040000 173.750000 371.945000 174.835000 ;
      RECT 371.230000 162.215000 372.360000 164.565000 ;
      RECT 371.275000  34.325000 372.285000  34.345000 ;
      RECT 371.275000  34.345000 373.960000  34.515000 ;
      RECT 371.275000  36.935000 373.960000  37.105000 ;
      RECT 371.275000  37.105000 372.285000  37.125000 ;
      RECT 371.325000 172.935000 371.945000 173.750000 ;
      RECT 371.370000  57.685000 371.540000  62.535000 ;
      RECT 371.370000  64.050000 371.540000  68.900000 ;
      RECT 371.425000 165.335000 371.935000 165.425000 ;
      RECT 371.475000   6.000000 372.015000  11.395000 ;
      RECT 371.475000  19.075000 372.015000  24.470000 ;
      RECT 371.695000  31.065000 371.865000  33.775000 ;
      RECT 371.695000  37.675000 371.865000  40.385000 ;
      RECT 371.945000 202.710000 443.295000 206.365000 ;
      RECT 371.945000 206.365000 387.620000 211.275000 ;
      RECT 371.945000 211.275000 443.295000 214.880000 ;
      RECT 371.945000 214.880000 382.945000 227.215000 ;
      RECT 372.185000  56.835000 372.355000  70.255000 ;
      RECT 372.225000  42.025000 373.350000  42.195000 ;
      RECT 372.225000  42.195000 372.395000  52.675000 ;
      RECT 372.225000  52.675000 373.350000  52.845000 ;
      RECT 372.475000  31.065000 372.645000  33.775000 ;
      RECT 372.475000  37.675000 372.645000  40.385000 ;
      RECT 372.490000   5.135000 373.190000  12.265000 ;
      RECT 372.490000  18.205000 373.190000  25.335000 ;
      RECT 372.765000  82.505000 372.995000 184.540000 ;
      RECT 372.765000 184.540000 382.225000 184.770000 ;
      RECT 372.795000  53.700000 374.905000  53.870000 ;
      RECT 372.795000  53.870000 372.965000  82.505000 ;
      RECT 372.865000  34.325000 373.535000  34.345000 ;
      RECT 372.865000  37.105000 373.535000  37.125000 ;
      RECT 373.405000  42.415000 373.575000  52.305000 ;
      RECT 373.525000  56.710000 373.855000  58.300000 ;
      RECT 373.755000  31.065000 373.925000  33.775000 ;
      RECT 373.755000  37.675000 373.925000  40.385000 ;
      RECT 373.950000   3.665000 374.905000  13.725000 ;
      RECT 373.950000  16.745000 374.650000  26.805000 ;
      RECT 373.985000  41.775000 374.320000  42.710000 ;
      RECT 373.985000  42.710000 374.155000  53.095000 ;
      RECT 374.215000  54.165000 374.865000  56.710000 ;
      RECT 374.235000  30.815000 374.405000  34.085000 ;
      RECT 374.235000  37.365000 374.405000  40.635000 ;
      RECT 374.335000  56.710000 374.865000  58.050000 ;
      RECT 374.735000  14.425000 374.905000  16.045000 ;
      RECT 374.735000  42.790000 375.695000  42.960000 ;
      RECT 374.735000  42.960000 374.905000  53.700000 ;
      RECT 375.170000  29.880000 375.340000  35.050000 ;
      RECT 375.170000  36.400000 375.340000  41.570000 ;
      RECT 375.285000  17.350000 377.305000  18.100000 ;
      RECT 375.285000  27.930000 377.305000  28.680000 ;
      RECT 375.465000  43.425000 375.795000  44.015000 ;
      RECT 375.465000 182.950000 375.795000 183.555000 ;
      RECT 375.525000  41.725000 382.225000  41.895000 ;
      RECT 375.525000  41.895000 375.695000  42.790000 ;
      RECT 375.665000   3.905000 378.175000   4.075000 ;
      RECT 375.665000   4.075000 375.835000  15.315000 ;
      RECT 375.665000  15.315000 378.175000  15.485000 ;
      RECT 376.060000  14.905000 377.370000  15.075000 ;
      RECT 376.245000   4.675000 376.415000  14.525000 ;
      RECT 376.275000 182.950000 376.605000 183.550000 ;
      RECT 376.470000   4.315000 377.370000   4.485000 ;
      RECT 376.585000   4.485000 377.255000  14.905000 ;
      RECT 377.085000 182.950000 377.415000 183.550000 ;
      RECT 377.425000   4.675000 377.595000  14.565000 ;
      RECT 377.895000 182.950000 378.225000 183.550000 ;
      RECT 378.005000   4.075000 378.175000  15.315000 ;
      RECT 378.325000  41.695000 382.225000  41.725000 ;
      RECT 378.325000  41.895000 382.225000  41.925000 ;
      RECT 378.705000 182.950000 379.035000 183.550000 ;
      RECT 378.935000   3.135000 379.105000  16.245000 ;
      RECT 379.515000 136.140000 379.845000 136.730000 ;
      RECT 379.515000 182.950000 379.845000 183.540000 ;
      RECT 380.100000   0.415000 385.640000   8.500000 ;
      RECT 380.100000   8.500000 400.380000   9.250000 ;
      RECT 380.100000   9.250000 386.090000  41.120000 ;
      RECT 380.325000  65.275000 380.655000  65.865000 ;
      RECT 381.135000  65.275000 381.550000  65.865000 ;
      RECT 381.995000  41.925000 382.225000 184.540000 ;
      RECT 382.770000  41.120000 386.090000 134.915000 ;
      RECT 382.770000 134.915000 383.970000 148.030000 ;
      RECT 382.770000 148.030000 385.370000 185.835000 ;
      RECT 384.150000 216.230000 444.600000 217.090000 ;
      RECT 384.150000 217.090000 385.010000 240.090000 ;
      RECT 384.150000 240.090000 408.075000 240.120000 ;
      RECT 384.150000 240.120000 420.680000 240.290000 ;
      RECT 384.775000 136.240000 384.955000 146.960000 ;
      RECT 384.775000 146.960000 396.285000 147.140000 ;
      RECT 385.000000 240.290000 408.075000 240.320000 ;
      RECT 385.720000 134.915000 386.090000 146.015000 ;
      RECT 385.720000 146.015000 395.340000 146.325000 ;
      RECT 386.070000 218.170000 439.970000 218.340000 ;
      RECT 386.070000 218.340000 386.240000 228.475000 ;
      RECT 386.070000 228.475000 439.970000 228.645000 ;
      RECT 386.070000 228.645000 386.240000 238.890000 ;
      RECT 386.070000 238.890000 420.055000 239.055000 ;
      RECT 386.070000 239.055000 413.105000 239.060000 ;
      RECT 386.205000 147.140000 386.385000 199.940000 ;
      RECT 386.205000 199.940000 428.415000 200.145000 ;
      RECT 386.270000   9.660000 386.600000  10.310000 ;
      RECT 386.270000  27.735000 386.600000  29.785000 ;
      RECT 386.270000  47.580000 386.600000  48.230000 ;
      RECT 386.270000  48.610000 386.600000  49.260000 ;
      RECT 386.270000  67.055000 386.600000  67.705000 ;
      RECT 386.270000  68.085000 386.600000  68.735000 ;
      RECT 386.270000  86.530000 386.600000  87.180000 ;
      RECT 386.270000  87.560000 386.600000  88.210000 ;
      RECT 386.270000 106.005000 386.600000 106.655000 ;
      RECT 386.270000 107.035000 386.600000 107.685000 ;
      RECT 386.270000 125.480000 386.600000 126.130000 ;
      RECT 386.270000 126.510000 386.600000 127.160000 ;
      RECT 386.270000 144.955000 386.600000 145.605000 ;
      RECT 386.440000 246.700000 387.060000 252.915000 ;
      RECT 386.440000 252.915000 415.045000 253.535000 ;
      RECT 386.575000   0.300000 477.515000   1.970000 ;
      RECT 386.680000 222.890000 387.535000 223.900000 ;
      RECT 386.680000 233.220000 387.535000 234.230000 ;
      RECT 386.770000 214.880000 443.295000 215.425000 ;
      RECT 386.820000 224.560000 387.085000 225.770000 ;
      RECT 386.820000 225.770000 389.445000 226.020000 ;
      RECT 386.820000 231.100000 389.445000 231.350000 ;
      RECT 386.820000 231.350000 387.085000 232.560000 ;
      RECT 386.900000   9.660000 387.230000  10.310000 ;
      RECT 386.900000  27.735000 387.230000  29.785000 ;
      RECT 386.900000  47.580000 387.230000  48.230000 ;
      RECT 386.900000  48.610000 387.230000  49.260000 ;
      RECT 386.900000  67.055000 387.230000  67.705000 ;
      RECT 386.900000  68.085000 387.230000  68.735000 ;
      RECT 386.900000  86.530000 387.230000  87.180000 ;
      RECT 386.900000  87.560000 387.230000  88.210000 ;
      RECT 386.900000 106.005000 387.230000 106.655000 ;
      RECT 386.900000 107.035000 387.230000 107.685000 ;
      RECT 386.900000 125.480000 387.230000 126.130000 ;
      RECT 386.900000 126.510000 387.230000 127.160000 ;
      RECT 386.900000 144.955000 387.230000 145.605000 ;
      RECT 387.050000 226.570000 387.560000 227.580000 ;
      RECT 387.050000 229.540000 387.560000 230.550000 ;
      RECT 387.085000 224.150000 390.345000 224.320000 ;
      RECT 387.085000 232.800000 390.345000 232.970000 ;
      RECT 387.150000 147.725000 391.730000 148.085000 ;
      RECT 387.150000 148.085000 387.330000 198.900000 ;
      RECT 387.150000 198.900000 391.730000 199.200000 ;
      RECT 387.345000 248.605000 387.875000 248.775000 ;
      RECT 387.345000 248.775000 387.735000 252.275000 ;
      RECT 387.410000 245.925000 388.080000 248.415000 ;
      RECT 387.465000 235.700000 387.635000 238.410000 ;
      RECT 387.530000   9.660000 387.860000  10.310000 ;
      RECT 387.530000  27.735000 387.860000  29.785000 ;
      RECT 387.530000  47.580000 387.860000  48.230000 ;
      RECT 387.530000  48.610000 387.860000  49.260000 ;
      RECT 387.530000  67.055000 387.860000  67.705000 ;
      RECT 387.530000  68.085000 387.860000  68.735000 ;
      RECT 387.530000  86.530000 387.860000  87.180000 ;
      RECT 387.530000  87.560000 387.860000  88.210000 ;
      RECT 387.530000 106.005000 387.860000 106.655000 ;
      RECT 387.530000 107.035000 387.860000 107.685000 ;
      RECT 387.530000 125.480000 387.860000 126.130000 ;
      RECT 387.530000 126.510000 387.860000 127.160000 ;
      RECT 387.530000 144.955000 387.860000 145.605000 ;
      RECT 387.615000 227.830000 389.055000 228.000000 ;
      RECT 387.615000 229.120000 389.055000 229.290000 ;
      RECT 387.665000 234.980000 388.565000 235.120000 ;
      RECT 387.665000 235.120000 388.335000 235.150000 ;
      RECT 387.700000 148.495000 388.030000 149.145000 ;
      RECT 387.700000 157.540000 388.030000 158.190000 ;
      RECT 387.700000 158.570000 388.030000 159.220000 ;
      RECT 387.700000 167.615000 388.030000 168.265000 ;
      RECT 387.700000 168.645000 388.030000 169.295000 ;
      RECT 387.700000 177.690000 388.030000 178.340000 ;
      RECT 387.700000 178.720000 388.030000 179.370000 ;
      RECT 387.700000 187.765000 388.030000 188.415000 ;
      RECT 387.700000 188.795000 388.030000 189.445000 ;
      RECT 387.700000 197.840000 388.030000 198.490000 ;
      RECT 387.765000 226.020000 388.045000 227.590000 ;
      RECT 387.765000 229.530000 388.045000 231.100000 ;
      RECT 387.820000 218.710000 387.990000 221.420000 ;
      RECT 387.875000 222.890000 388.405000 223.900000 ;
      RECT 387.875000 224.570000 388.405000 225.580000 ;
      RECT 387.875000 231.540000 388.405000 232.550000 ;
      RECT 387.875000 233.220000 388.405000 234.230000 ;
      RECT 387.920000 249.565000 388.850000 252.425000 ;
      RECT 388.020000 221.970000 388.690000 222.000000 ;
      RECT 388.020000 222.000000 388.920000 222.140000 ;
      RECT 388.035000 234.950000 388.565000 234.980000 ;
      RECT 388.150000   4.470000 393.020000   4.650000 ;
      RECT 388.150000   4.650000 388.330000   8.125000 ;
      RECT 388.150000   8.125000 425.580000   8.180000 ;
      RECT 388.150000   8.180000 401.325000   8.305000 ;
      RECT 388.160000   9.660000 388.490000  10.310000 ;
      RECT 388.160000  27.735000 388.490000  29.785000 ;
      RECT 388.160000  47.580000 388.490000  48.230000 ;
      RECT 388.160000  48.610000 388.490000  49.260000 ;
      RECT 388.160000  67.055000 388.490000  67.705000 ;
      RECT 388.160000  68.085000 388.490000  68.735000 ;
      RECT 388.160000  86.530000 388.490000  87.180000 ;
      RECT 388.160000  87.560000 388.490000  88.210000 ;
      RECT 388.160000 106.005000 388.490000 106.655000 ;
      RECT 388.160000 107.035000 388.490000 107.685000 ;
      RECT 388.160000 125.480000 388.490000 126.130000 ;
      RECT 388.160000 126.510000 388.490000 127.160000 ;
      RECT 388.160000 144.955000 388.490000 145.605000 ;
      RECT 388.250000 226.570000 388.420000 227.580000 ;
      RECT 388.250000 229.540000 388.420000 230.550000 ;
      RECT 388.330000 148.495000 388.660000 149.145000 ;
      RECT 388.330000 157.540000 388.660000 158.190000 ;
      RECT 388.330000 158.570000 388.660000 159.220000 ;
      RECT 388.330000 167.615000 388.660000 168.265000 ;
      RECT 388.330000 168.645000 388.660000 169.295000 ;
      RECT 388.330000 177.690000 388.660000 178.340000 ;
      RECT 388.330000 178.720000 388.660000 179.370000 ;
      RECT 388.330000 187.765000 388.660000 188.415000 ;
      RECT 388.330000 188.795000 388.660000 189.445000 ;
      RECT 388.330000 197.840000 388.660000 198.490000 ;
      RECT 388.345000 235.700000 388.515000 238.410000 ;
      RECT 388.390000 222.140000 388.920000 222.170000 ;
      RECT 388.420000 207.340000 388.590000 210.050000 ;
      RECT 388.420000 241.395000 388.590000 244.105000 ;
      RECT 388.615000 206.950000 389.285000 207.120000 ;
      RECT 388.615000 244.325000 389.285000 244.495000 ;
      RECT 388.625000 226.020000 388.905000 227.590000 ;
      RECT 388.625000 229.530000 388.905000 231.100000 ;
      RECT 388.700000 218.710000 388.870000 221.420000 ;
      RECT 388.740000   4.950000 388.910000   5.960000 ;
      RECT 388.740000   6.620000 388.910000   7.630000 ;
      RECT 388.785000 246.265000 391.150000 246.775000 ;
      RECT 388.790000   9.660000 389.120000  10.310000 ;
      RECT 388.790000  27.735000 389.120000  29.785000 ;
      RECT 388.790000  47.580000 389.120000  48.230000 ;
      RECT 388.790000  48.610000 389.120000  49.260000 ;
      RECT 388.790000  67.055000 389.120000  67.705000 ;
      RECT 388.790000  68.085000 389.120000  68.735000 ;
      RECT 388.790000  86.530000 389.120000  87.180000 ;
      RECT 388.790000  87.560000 389.120000  88.210000 ;
      RECT 388.790000 106.005000 389.120000 106.655000 ;
      RECT 388.790000 107.035000 389.120000 107.685000 ;
      RECT 388.790000 125.480000 389.120000 126.130000 ;
      RECT 388.790000 126.510000 389.120000 127.160000 ;
      RECT 388.790000 144.955000 389.120000 145.605000 ;
      RECT 388.905000 248.995000 390.285000 249.165000 ;
      RECT 388.920000 246.775000 389.185000 248.075000 ;
      RECT 388.960000 148.495000 389.290000 149.145000 ;
      RECT 388.960000 157.540000 389.290000 158.190000 ;
      RECT 388.960000 158.570000 389.290000 159.220000 ;
      RECT 388.960000 167.615000 389.290000 168.265000 ;
      RECT 388.960000 168.645000 389.290000 169.295000 ;
      RECT 388.960000 177.690000 389.290000 178.340000 ;
      RECT 388.960000 178.720000 389.290000 179.370000 ;
      RECT 388.960000 187.765000 389.290000 188.415000 ;
      RECT 388.960000 188.795000 389.290000 189.445000 ;
      RECT 388.960000 197.840000 389.290000 198.490000 ;
      RECT 388.965000   6.220000 394.955000   6.390000 ;
      RECT 389.040000 222.890000 389.570000 223.900000 ;
      RECT 389.040000 233.220000 389.570000 234.230000 ;
      RECT 389.110000 226.570000 389.620000 227.580000 ;
      RECT 389.110000 229.540000 389.620000 230.550000 ;
      RECT 389.165000 224.560000 389.445000 225.770000 ;
      RECT 389.165000 231.350000 389.445000 232.560000 ;
      RECT 389.240000 249.475000 389.850000 252.915000 ;
      RECT 389.245000 248.605000 389.775000 248.775000 ;
      RECT 389.300000 207.340000 390.620000 210.110000 ;
      RECT 389.300000 241.335000 390.620000 244.105000 ;
      RECT 389.365000 247.065000 389.645000 248.605000 ;
      RECT 389.420000   9.660000 389.750000  10.310000 ;
      RECT 389.420000  27.735000 389.750000  29.785000 ;
      RECT 389.420000  47.580000 389.750000  48.230000 ;
      RECT 389.420000  48.610000 389.750000  49.260000 ;
      RECT 389.420000  67.055000 389.750000  67.705000 ;
      RECT 389.420000  68.085000 389.750000  68.735000 ;
      RECT 389.420000  86.530000 389.750000  87.180000 ;
      RECT 389.420000  87.560000 389.750000  88.210000 ;
      RECT 389.420000 106.005000 389.750000 106.655000 ;
      RECT 389.420000 107.035000 389.750000 107.685000 ;
      RECT 389.420000 125.480000 389.750000 126.130000 ;
      RECT 389.420000 126.510000 389.750000 127.160000 ;
      RECT 389.420000 144.955000 389.750000 145.605000 ;
      RECT 389.590000 148.495000 389.920000 149.145000 ;
      RECT 389.590000 157.540000 389.920000 158.190000 ;
      RECT 389.590000 158.570000 389.920000 159.220000 ;
      RECT 389.590000 167.615000 389.920000 168.265000 ;
      RECT 389.590000 168.645000 389.920000 169.295000 ;
      RECT 389.590000 177.690000 389.920000 178.340000 ;
      RECT 389.590000 178.720000 389.920000 179.370000 ;
      RECT 389.590000 187.765000 389.920000 188.415000 ;
      RECT 389.590000 188.795000 389.920000 189.445000 ;
      RECT 389.590000 197.840000 389.920000 198.490000 ;
      RECT 389.620000   4.950000 389.790000   5.960000 ;
      RECT 389.620000   6.620000 389.790000   7.630000 ;
      RECT 389.805000 219.125000 390.335000 220.220000 ;
      RECT 389.830000 246.775000 390.095000 248.075000 ;
      RECT 389.855000 235.640000 390.385000 235.810000 ;
      RECT 389.965000 220.980000 390.135000 221.870000 ;
      RECT 389.965000 235.470000 390.135000 235.640000 ;
      RECT 389.965000 235.810000 390.135000 236.140000 ;
      RECT 390.050000   9.660000 390.380000  10.310000 ;
      RECT 390.050000  27.735000 390.380000  29.785000 ;
      RECT 390.050000  47.580000 390.380000  48.230000 ;
      RECT 390.050000  48.610000 390.380000  49.260000 ;
      RECT 390.050000  67.055000 390.380000  67.705000 ;
      RECT 390.050000  68.085000 390.380000  68.735000 ;
      RECT 390.050000  86.530000 390.380000  87.180000 ;
      RECT 390.050000  87.560000 390.380000  88.210000 ;
      RECT 390.050000 106.005000 390.380000 106.655000 ;
      RECT 390.050000 107.035000 390.380000 107.685000 ;
      RECT 390.050000 125.480000 390.380000 126.130000 ;
      RECT 390.050000 126.510000 390.380000 127.160000 ;
      RECT 390.050000 144.955000 390.380000 145.605000 ;
      RECT 390.165000 236.900000 390.335000 238.260000 ;
      RECT 390.220000 148.495000 390.550000 149.145000 ;
      RECT 390.220000 157.540000 390.550000 158.190000 ;
      RECT 390.220000 158.570000 390.550000 159.220000 ;
      RECT 390.220000 167.615000 390.550000 168.265000 ;
      RECT 390.220000 168.645000 390.550000 169.295000 ;
      RECT 390.220000 177.690000 390.550000 178.340000 ;
      RECT 390.220000 178.720000 390.550000 179.370000 ;
      RECT 390.220000 187.765000 390.550000 188.415000 ;
      RECT 390.220000 188.795000 390.550000 189.445000 ;
      RECT 390.220000 197.840000 390.550000 198.490000 ;
      RECT 390.220000 222.890000 390.750000 223.900000 ;
      RECT 390.220000 224.570000 390.750000 225.580000 ;
      RECT 390.220000 231.540000 390.750000 232.550000 ;
      RECT 390.220000 233.220000 390.750000 234.230000 ;
      RECT 390.240000 249.565000 391.170000 252.425000 ;
      RECT 390.340000 247.065000 390.510000 248.075000 ;
      RECT 390.355000 220.470000 391.025000 220.640000 ;
      RECT 390.355000 236.480000 391.025000 236.650000 ;
      RECT 390.500000   4.950000 390.670000   5.960000 ;
      RECT 390.500000   6.620000 390.670000   7.630000 ;
      RECT 390.625000 218.520000 391.215000 218.690000 ;
      RECT 390.625000 238.530000 391.215000 238.700000 ;
      RECT 390.650000 210.325000 392.850000 210.995000 ;
      RECT 390.650000 240.675000 392.850000 240.845000 ;
      RECT 390.670000 218.690000 391.215000 220.220000 ;
      RECT 390.670000 236.900000 391.215000 238.530000 ;
      RECT 390.680000   9.660000 391.010000  10.310000 ;
      RECT 390.680000  27.735000 391.010000  31.070000 ;
      RECT 390.680000  47.580000 391.010000  48.230000 ;
      RECT 390.680000  48.610000 391.010000  49.260000 ;
      RECT 390.680000  67.055000 391.010000  67.705000 ;
      RECT 390.680000  68.085000 391.010000  68.735000 ;
      RECT 390.680000  86.530000 391.010000  87.180000 ;
      RECT 390.680000  87.560000 391.010000  88.210000 ;
      RECT 390.680000 106.005000 391.010000 106.655000 ;
      RECT 390.680000 107.035000 391.010000 107.685000 ;
      RECT 390.680000 125.480000 391.010000 126.130000 ;
      RECT 390.680000 126.510000 391.010000 127.160000 ;
      RECT 390.680000 144.955000 391.010000 145.605000 ;
      RECT 390.735000 248.605000 391.405000 248.775000 ;
      RECT 390.745000 246.775000 391.010000 248.075000 ;
      RECT 390.825000 207.540000 391.130000 210.325000 ;
      RECT 390.825000 240.845000 392.850000 241.215000 ;
      RECT 390.825000 241.215000 391.130000 243.905000 ;
      RECT 390.850000 148.495000 391.180000 149.145000 ;
      RECT 390.850000 157.540000 391.180000 158.190000 ;
      RECT 390.850000 158.570000 391.180000 159.220000 ;
      RECT 390.850000 167.615000 391.180000 168.265000 ;
      RECT 390.850000 168.645000 391.180000 169.295000 ;
      RECT 390.850000 177.690000 391.180000 178.340000 ;
      RECT 390.850000 178.720000 391.180000 179.370000 ;
      RECT 390.850000 187.765000 391.180000 188.415000 ;
      RECT 390.850000 188.795000 391.180000 189.445000 ;
      RECT 390.850000 197.840000 391.180000 198.490000 ;
      RECT 390.885000 236.070000 391.415000 236.240000 ;
      RECT 390.895000 226.570000 391.405000 227.580000 ;
      RECT 390.895000 229.540000 391.405000 230.550000 ;
      RECT 391.245000 220.980000 391.415000 221.650000 ;
      RECT 391.245000 235.470000 391.415000 236.070000 ;
      RECT 391.310000   9.660000 391.640000  10.310000 ;
      RECT 391.310000  27.735000 391.640000  29.885000 ;
      RECT 391.310000  47.580000 391.640000  48.230000 ;
      RECT 391.310000  48.610000 391.640000  49.260000 ;
      RECT 391.310000  67.055000 391.640000  67.705000 ;
      RECT 391.310000  68.085000 391.640000  68.735000 ;
      RECT 391.310000  86.530000 391.640000  87.180000 ;
      RECT 391.310000  87.560000 391.640000  88.210000 ;
      RECT 391.310000 106.005000 391.640000 106.655000 ;
      RECT 391.310000 119.155000 391.640000 119.805000 ;
      RECT 391.310000 125.480000 391.640000 126.130000 ;
      RECT 391.310000 126.510000 391.640000 127.160000 ;
      RECT 391.310000 144.955000 391.640000 145.605000 ;
      RECT 391.330000 207.340000 391.500000 210.050000 ;
      RECT 391.330000 241.395000 391.500000 244.105000 ;
      RECT 391.380000   4.950000 391.550000   5.960000 ;
      RECT 391.380000   6.620000 391.550000   7.630000 ;
      RECT 391.415000 218.520000 392.005000 218.690000 ;
      RECT 391.415000 218.690000 391.790000 220.080000 ;
      RECT 391.415000 220.080000 392.025000 220.580000 ;
      RECT 391.415000 220.580000 392.390000 220.790000 ;
      RECT 391.415000 236.420000 392.390000 236.540000 ;
      RECT 391.415000 236.540000 392.025000 237.040000 ;
      RECT 391.415000 237.040000 391.790000 238.530000 ;
      RECT 391.415000 238.530000 392.005000 238.700000 ;
      RECT 391.460000 227.830000 392.900000 228.000000 ;
      RECT 391.460000 229.120000 392.900000 229.290000 ;
      RECT 391.460000 249.565000 391.840000 252.275000 ;
      RECT 391.550000 148.085000 391.730000 198.900000 ;
      RECT 391.585000 247.405000 391.840000 249.565000 ;
      RECT 391.665000 226.270000 391.835000 227.580000 ;
      RECT 391.665000 229.540000 391.835000 230.850000 ;
      RECT 391.670000 220.790000 392.390000 221.650000 ;
      RECT 391.670000 235.470000 392.390000 236.420000 ;
      RECT 391.825000 222.650000 391.995000 225.360000 ;
      RECT 391.825000 231.760000 391.995000 234.470000 ;
      RECT 391.940000   9.660000 392.270000  10.310000 ;
      RECT 391.940000  27.735000 392.270000  29.885000 ;
      RECT 391.940000  47.580000 392.270000  48.230000 ;
      RECT 391.940000  48.610000 392.270000  49.260000 ;
      RECT 391.940000  67.055000 392.270000  67.705000 ;
      RECT 391.940000  68.085000 392.270000  68.735000 ;
      RECT 391.940000  86.530000 392.270000  87.180000 ;
      RECT 391.940000  87.560000 392.270000  88.210000 ;
      RECT 391.940000 106.005000 392.270000 106.655000 ;
      RECT 391.940000 107.035000 392.270000 107.685000 ;
      RECT 391.940000 125.480000 392.270000 126.130000 ;
      RECT 391.940000 126.510000 392.270000 127.160000 ;
      RECT 391.940000 144.955000 392.270000 145.605000 ;
      RECT 391.990000 219.185000 392.520000 219.880000 ;
      RECT 391.990000 237.240000 392.160000 238.260000 ;
      RECT 392.020000 248.605000 392.550000 248.775000 ;
      RECT 392.020000 248.775000 392.410000 252.275000 ;
      RECT 392.050000 225.910000 394.190000 226.080000 ;
      RECT 392.050000 231.040000 394.190000 231.210000 ;
      RECT 392.085000 245.095000 395.570000 245.765000 ;
      RECT 392.085000 245.765000 392.755000 248.415000 ;
      RECT 392.095000 226.570000 392.265000 227.600000 ;
      RECT 392.095000 229.520000 392.265000 230.550000 ;
      RECT 392.180000 207.440000 392.850000 207.610000 ;
      RECT 392.180000 208.220000 392.910000 209.540000 ;
      RECT 392.180000 210.150000 392.850000 210.325000 ;
      RECT 392.180000 241.215000 392.850000 241.295000 ;
      RECT 392.180000 241.905000 392.910000 243.225000 ;
      RECT 392.180000 243.835000 392.850000 244.495000 ;
      RECT 392.215000 220.220000 393.215000 220.390000 ;
      RECT 392.215000 236.730000 393.215000 236.900000 ;
      RECT 392.260000   4.950000 392.430000   5.960000 ;
      RECT 392.260000   6.620000 392.430000   7.630000 ;
      RECT 392.345000 222.630000 392.875000 222.800000 ;
      RECT 392.345000 234.320000 392.875000 234.490000 ;
      RECT 392.495000 147.140000 392.675000 147.710000 ;
      RECT 392.495000 147.710000 406.805000 147.890000 ;
      RECT 392.525000 226.270000 392.695000 227.580000 ;
      RECT 392.525000 229.540000 392.695000 230.850000 ;
      RECT 392.570000   9.660000 392.900000  10.310000 ;
      RECT 392.570000  27.735000 392.900000  29.885000 ;
      RECT 392.570000  47.580000 392.900000  48.230000 ;
      RECT 392.570000  48.610000 392.900000  49.260000 ;
      RECT 392.570000  67.055000 392.900000  67.705000 ;
      RECT 392.570000  68.085000 392.900000  68.735000 ;
      RECT 392.570000  86.530000 392.900000  87.180000 ;
      RECT 392.570000  87.560000 392.900000  88.210000 ;
      RECT 392.570000 106.005000 392.900000 106.655000 ;
      RECT 392.570000 119.155000 392.900000 119.805000 ;
      RECT 392.570000 125.620000 392.900000 126.130000 ;
      RECT 392.570000 126.510000 392.900000 127.160000 ;
      RECT 392.570000 144.955000 392.900000 145.605000 ;
      RECT 392.595000 249.565000 393.525000 252.425000 ;
      RECT 392.650000 125.540000 392.820000 125.620000 ;
      RECT 392.705000 222.800000 392.875000 225.360000 ;
      RECT 392.705000 231.760000 392.875000 234.320000 ;
      RECT 392.760000 207.855000 393.360000 208.025000 ;
      RECT 392.760000 243.420000 393.360000 243.590000 ;
      RECT 392.840000   4.650000 393.020000   5.790000 ;
      RECT 392.840000   5.790000 402.640000   5.970000 ;
      RECT 392.910000 155.160000 393.080000 155.420000 ;
      RECT 392.910000 155.420000 395.015000 155.750000 ;
      RECT 392.955000 226.570000 393.465000 227.580000 ;
      RECT 392.955000 229.540000 393.465000 230.550000 ;
      RECT 393.100000 220.640000 393.270000 221.650000 ;
      RECT 393.100000 235.470000 393.270000 236.480000 ;
      RECT 393.140000   6.620000 393.310000   7.630000 ;
      RECT 393.185000 219.210000 394.645000 219.880000 ;
      RECT 393.185000 237.240000 394.645000 237.910000 ;
      RECT 393.190000 207.585000 393.360000 207.855000 ;
      RECT 393.190000 208.025000 393.360000 208.255000 ;
      RECT 393.190000 209.515000 393.360000 209.680000 ;
      RECT 393.190000 209.680000 394.210000 209.850000 ;
      RECT 393.190000 209.850000 393.360000 210.185000 ;
      RECT 393.190000 241.260000 393.360000 241.595000 ;
      RECT 393.190000 241.595000 394.210000 241.765000 ;
      RECT 393.190000 241.765000 393.360000 241.930000 ;
      RECT 393.190000 243.190000 393.360000 243.420000 ;
      RECT 393.190000 243.590000 393.360000 243.860000 ;
      RECT 393.200000   9.660000 393.530000  10.310000 ;
      RECT 393.200000  27.735000 393.530000  29.885000 ;
      RECT 393.200000  47.720000 393.530000  49.260000 ;
      RECT 393.200000  67.055000 393.530000  67.705000 ;
      RECT 393.200000  68.085000 393.530000  68.735000 ;
      RECT 393.200000  86.530000 393.530000  87.180000 ;
      RECT 393.200000  87.560000 393.530000  88.210000 ;
      RECT 393.200000 106.005000 393.530000 106.655000 ;
      RECT 393.200000 107.035000 393.530000 107.685000 ;
      RECT 393.200000 125.480000 393.530000 126.130000 ;
      RECT 393.200000 126.510000 393.530000 127.160000 ;
      RECT 393.200000 144.955000 393.530000 145.605000 ;
      RECT 393.365000 222.650000 393.535000 225.360000 ;
      RECT 393.365000 231.760000 393.535000 234.470000 ;
      RECT 393.445000 147.890000 393.625000 154.950000 ;
      RECT 393.445000 155.920000 419.985000 156.100000 ;
      RECT 393.445000 156.100000 393.625000 182.010000 ;
      RECT 393.445000 182.010000 428.475000 182.190000 ;
      RECT 393.445000 182.190000 393.625000 199.580000 ;
      RECT 393.445000 199.580000 393.675000 199.940000 ;
      RECT 393.450000 154.950000 393.620000 155.230000 ;
      RECT 393.460000 246.265000 395.825000 246.775000 ;
      RECT 393.560000 207.410000 394.210000 209.680000 ;
      RECT 393.560000 241.765000 394.210000 244.495000 ;
      RECT 393.580000 248.995000 394.960000 249.165000 ;
      RECT 393.595000 246.775000 393.860000 248.075000 ;
      RECT 393.830000   9.660000 394.160000  10.310000 ;
      RECT 393.830000  27.560000 394.160000  29.885000 ;
      RECT 393.830000  33.580000 394.160000  35.640000 ;
      RECT 393.830000  47.170000 394.160000  48.230000 ;
      RECT 393.830000  48.610000 394.160000  49.260000 ;
      RECT 393.830000  67.055000 394.160000  67.705000 ;
      RECT 393.830000  68.085000 394.160000  68.735000 ;
      RECT 393.830000  86.530000 394.160000  87.180000 ;
      RECT 393.830000  87.560000 394.160000  88.210000 ;
      RECT 393.830000 106.005000 394.160000 106.655000 ;
      RECT 393.830000 119.155000 394.160000 119.805000 ;
      RECT 393.830000 125.480000 394.160000 126.130000 ;
      RECT 393.830000 126.510000 394.160000 127.160000 ;
      RECT 393.830000 144.955000 394.160000 145.605000 ;
      RECT 393.915000 249.475000 394.525000 252.915000 ;
      RECT 393.920000 248.605000 394.450000 248.775000 ;
      RECT 394.020000   6.620000 394.190000   7.630000 ;
      RECT 394.040000 247.065000 394.320000 248.605000 ;
      RECT 394.200000 148.240000 394.370000 155.230000 ;
      RECT 394.245000 222.650000 394.415000 225.360000 ;
      RECT 394.245000 231.760000 394.415000 234.470000 ;
      RECT 394.390000 156.865000 405.860000 157.045000 ;
      RECT 394.390000 157.045000 395.150000 162.575000 ;
      RECT 394.390000 162.575000 395.625000 162.905000 ;
      RECT 394.390000 162.905000 395.150000 168.535000 ;
      RECT 394.390000 168.535000 395.625000 168.865000 ;
      RECT 394.390000 168.865000 395.150000 174.495000 ;
      RECT 394.390000 174.495000 395.625000 174.825000 ;
      RECT 394.390000 174.825000 395.150000 180.455000 ;
      RECT 394.390000 180.455000 395.625000 180.785000 ;
      RECT 394.390000 180.785000 395.150000 180.955000 ;
      RECT 394.390000 180.955000 405.860000 181.135000 ;
      RECT 394.390000 182.955000 427.470000 183.135000 ;
      RECT 394.390000 183.135000 394.570000 189.290000 ;
      RECT 394.390000 189.290000 427.470000 189.470000 ;
      RECT 394.460000   9.660000 394.790000  10.680000 ;
      RECT 394.460000  27.735000 394.790000  29.855000 ;
      RECT 394.460000  33.580000 394.790000  35.640000 ;
      RECT 394.460000  48.610000 394.790000  49.260000 ;
      RECT 394.460000  67.055000 394.790000  67.705000 ;
      RECT 394.460000  68.085000 394.790000  68.735000 ;
      RECT 394.460000  86.530000 394.790000  87.180000 ;
      RECT 394.460000  87.560000 394.790000  88.210000 ;
      RECT 394.460000 106.005000 394.790000 106.655000 ;
      RECT 394.460000 107.035000 394.790000 107.685000 ;
      RECT 394.460000 125.480000 394.790000 126.130000 ;
      RECT 394.460000 126.510000 394.790000 127.160000 ;
      RECT 394.460000 144.955000 394.790000 145.605000 ;
      RECT 394.505000 246.775000 394.770000 248.075000 ;
      RECT 394.610000 189.470000 394.790000 199.020000 ;
      RECT 394.610000 199.020000 427.470000 199.200000 ;
      RECT 394.640000 206.365000 395.490000 211.275000 ;
      RECT 394.900000   6.620000 395.070000   7.630000 ;
      RECT 394.900000 243.845000 395.570000 245.095000 ;
      RECT 394.915000 249.565000 395.845000 252.425000 ;
      RECT 394.980000 183.610000 395.150000 188.370000 ;
      RECT 395.015000 247.065000 395.185000 248.075000 ;
      RECT 395.025000 218.340000 395.195000 228.475000 ;
      RECT 395.025000 228.645000 395.195000 238.890000 ;
      RECT 395.030000 190.240000 395.365000 193.970000 ;
      RECT 395.030000 194.520000 395.365000 198.250000 ;
      RECT 395.090000   9.660000 395.420000  10.680000 ;
      RECT 395.090000  27.560000 395.420000  29.855000 ;
      RECT 395.090000  33.580000 395.420000  35.075000 ;
      RECT 395.125000   6.220000 396.655000   6.390000 ;
      RECT 395.160000  35.485000 396.180000  35.665000 ;
      RECT 395.160000  35.665000 395.340000 146.015000 ;
      RECT 395.180000   2.640000 401.930000   2.820000 ;
      RECT 395.180000   2.820000 395.360000   4.845000 ;
      RECT 395.180000   4.845000 401.930000   5.025000 ;
      RECT 395.205000 188.870000 396.685000 189.040000 ;
      RECT 395.410000 248.605000 396.080000 248.775000 ;
      RECT 395.420000 246.775000 395.685000 248.075000 ;
      RECT 395.480000 148.220000 395.650000 155.230000 ;
      RECT 395.560000 189.470000 426.710000 190.050000 ;
      RECT 395.560000 190.050000 415.820000 194.160000 ;
      RECT 395.560000 194.160000 426.710000 194.330000 ;
      RECT 395.560000 194.330000 405.395000 198.440000 ;
      RECT 395.560000 198.440000 426.710000 199.020000 ;
      RECT 395.575000 219.210000 397.035000 219.880000 ;
      RECT 395.575000 237.240000 397.035000 237.910000 ;
      RECT 395.690000 188.530000 396.220000 188.870000 ;
      RECT 395.720000   9.660000 396.050000  10.680000 ;
      RECT 395.720000  27.735000 396.050000  29.855000 ;
      RECT 395.720000  33.580000 396.050000  35.075000 ;
      RECT 395.760000 157.395000 395.930000 162.245000 ;
      RECT 395.760000 163.355000 395.930000 168.205000 ;
      RECT 395.760000 169.315000 395.930000 174.165000 ;
      RECT 395.760000 175.275000 395.930000 180.125000 ;
      RECT 395.770000   3.170000 395.940000   4.195000 ;
      RECT 395.805000 222.650000 395.975000 225.360000 ;
      RECT 395.805000 231.760000 395.975000 234.470000 ;
      RECT 395.860000 183.610000 396.030000 188.360000 ;
      RECT 395.865000   4.425000 396.545000   4.595000 ;
      RECT 395.940000 155.420000 397.470000 155.750000 ;
      RECT 396.010000 207.410000 396.660000 209.680000 ;
      RECT 396.010000 209.680000 397.030000 209.850000 ;
      RECT 396.010000 241.595000 397.030000 241.765000 ;
      RECT 396.010000 241.765000 396.660000 244.495000 ;
      RECT 396.030000 225.910000 398.170000 226.080000 ;
      RECT 396.030000 231.040000 398.170000 231.210000 ;
      RECT 396.105000  38.145000 418.880000  38.465000 ;
      RECT 396.105000  38.465000 396.285000 121.735000 ;
      RECT 396.105000 121.735000 419.985000 121.915000 ;
      RECT 396.105000 121.915000 396.285000 145.535000 ;
      RECT 396.105000 145.535000 397.305000 145.715000 ;
      RECT 396.105000 145.715000 396.285000 146.960000 ;
      RECT 396.105000 147.140000 396.285000 147.710000 ;
      RECT 396.135000 249.565000 396.515000 252.275000 ;
      RECT 396.180000   6.620000 396.350000   7.630000 ;
      RECT 396.200000 162.575000 399.770000 162.905000 ;
      RECT 396.200000 168.535000 399.770000 168.865000 ;
      RECT 396.200000 174.495000 399.770000 174.825000 ;
      RECT 396.200000 180.455000 399.770000 180.785000 ;
      RECT 396.260000 247.405000 396.515000 249.565000 ;
      RECT 396.350000   9.660000 396.680000  10.680000 ;
      RECT 396.350000  27.560000 396.680000  29.855000 ;
      RECT 396.350000  33.580000 396.680000  35.890000 ;
      RECT 396.350000  35.890000 396.910000  36.060000 ;
      RECT 396.460000 147.345000 399.870000 147.515000 ;
      RECT 396.515000 146.115000 397.045000 147.145000 ;
      RECT 396.635000 145.115000 397.305000 145.285000 ;
      RECT 396.685000 222.650000 396.855000 225.360000 ;
      RECT 396.685000 231.760000 396.855000 234.470000 ;
      RECT 396.695000 122.165000 397.420000 122.335000 ;
      RECT 396.695000 122.335000 396.865000 129.815000 ;
      RECT 396.695000 129.815000 397.420000 129.985000 ;
      RECT 396.695000 129.985000 396.865000 137.465000 ;
      RECT 396.695000 137.465000 397.420000 137.635000 ;
      RECT 396.695000 137.635000 396.865000 145.115000 ;
      RECT 396.695000 248.605000 397.225000 248.775000 ;
      RECT 396.695000 248.775000 397.085000 252.275000 ;
      RECT 396.715000   4.425000 398.955000   4.595000 ;
      RECT 396.730000   6.620000 396.900000   7.630000 ;
      RECT 396.740000 183.610000 396.910000 188.370000 ;
      RECT 396.755000 226.570000 397.265000 227.580000 ;
      RECT 396.755000 229.540000 397.265000 230.550000 ;
      RECT 396.760000 244.710000 397.430000 248.415000 ;
      RECT 396.850000   3.170000 397.020000   4.180000 ;
      RECT 396.850000  35.485000 400.380000  35.665000 ;
      RECT 396.860000 207.585000 397.030000 207.855000 ;
      RECT 396.860000 207.855000 397.460000 208.025000 ;
      RECT 396.860000 208.025000 397.030000 208.255000 ;
      RECT 396.860000 209.515000 397.030000 209.680000 ;
      RECT 396.860000 209.850000 397.030000 210.185000 ;
      RECT 396.860000 241.260000 397.030000 241.595000 ;
      RECT 396.860000 241.765000 397.030000 241.930000 ;
      RECT 396.860000 243.190000 397.030000 243.420000 ;
      RECT 396.860000 243.420000 397.460000 243.590000 ;
      RECT 396.860000 243.590000 397.030000 243.860000 ;
      RECT 396.950000 220.640000 397.120000 221.650000 ;
      RECT 396.950000 235.470000 397.120000 236.480000 ;
      RECT 396.955000   6.220000 398.955000   6.390000 ;
      RECT 396.980000   9.660000 397.310000  10.280000 ;
      RECT 396.980000  27.735000 397.310000  29.855000 ;
      RECT 396.980000  33.580000 397.310000  35.075000 ;
      RECT 397.005000 220.220000 398.005000 220.390000 ;
      RECT 397.005000 236.730000 398.005000 236.900000 ;
      RECT 397.030000 188.870000 406.760000 189.040000 ;
      RECT 397.070000   6.390000 398.840000   6.760000 ;
      RECT 397.205000  38.965000 418.885000  39.145000 ;
      RECT 397.205000  39.145000 397.385000  63.005000 ;
      RECT 397.205000  63.005000 425.725000  63.185000 ;
      RECT 397.205000  63.185000 397.385000 109.660000 ;
      RECT 397.205000 109.660000 397.990000 121.735000 ;
      RECT 397.270000 249.565000 398.200000 252.425000 ;
      RECT 397.310000 208.220000 398.040000 209.540000 ;
      RECT 397.310000 241.905000 398.040000 243.225000 ;
      RECT 397.320000 227.830000 398.760000 228.000000 ;
      RECT 397.320000 229.120000 398.760000 229.290000 ;
      RECT 397.345000 222.630000 397.875000 222.800000 ;
      RECT 397.345000 222.800000 397.515000 225.360000 ;
      RECT 397.345000 231.760000 397.515000 234.320000 ;
      RECT 397.345000 234.320000 397.875000 234.490000 ;
      RECT 397.370000 207.440000 398.040000 207.610000 ;
      RECT 397.370000 210.150000 398.040000 210.325000 ;
      RECT 397.370000 210.325000 399.570000 210.995000 ;
      RECT 397.370000 240.675000 399.570000 240.845000 ;
      RECT 397.370000 240.845000 399.395000 241.215000 ;
      RECT 397.370000 241.215000 398.040000 241.295000 ;
      RECT 397.370000 243.835000 398.040000 244.495000 ;
      RECT 397.475000 122.555000 397.645000 129.565000 ;
      RECT 397.475000 130.205000 397.645000 137.215000 ;
      RECT 397.475000 137.855000 397.645000 144.645000 ;
      RECT 397.475000 144.815000 397.645000 145.530000 ;
      RECT 397.475000 145.530000 398.765000 145.700000 ;
      RECT 397.475000 145.700000 397.645000 147.125000 ;
      RECT 397.525000 226.270000 397.695000 227.580000 ;
      RECT 397.525000 229.540000 397.695000 230.850000 ;
      RECT 397.610000   9.660000 397.940000  10.280000 ;
      RECT 397.610000  27.560000 397.940000  29.855000 ;
      RECT 397.610000  33.580000 397.940000  35.075000 ;
      RECT 397.700000 219.185000 398.230000 219.880000 ;
      RECT 397.760000 148.240000 397.930000 155.230000 ;
      RECT 397.830000 220.580000 398.805000 220.790000 ;
      RECT 397.830000 220.790000 398.550000 221.650000 ;
      RECT 397.830000 235.470000 398.550000 236.420000 ;
      RECT 397.830000 236.420000 398.805000 236.540000 ;
      RECT 397.855000 122.165000 399.545000 122.335000 ;
      RECT 397.855000 129.815000 399.545000 129.985000 ;
      RECT 397.855000 144.890000 399.545000 145.285000 ;
      RECT 397.895000 146.115000 398.425000 147.145000 ;
      RECT 397.930000   3.170000 398.100000   4.195000 ;
      RECT 397.955000 226.570000 398.125000 227.600000 ;
      RECT 397.955000 229.520000 398.125000 230.550000 ;
      RECT 398.020000 183.610000 398.190000 188.360000 ;
      RECT 398.060000 237.240000 398.230000 238.260000 ;
      RECT 398.135000 246.265000 400.500000 246.775000 ;
      RECT 398.150000  39.910000 417.940000  40.090000 ;
      RECT 398.150000  40.090000 398.330000  62.060000 ;
      RECT 398.150000  62.060000 417.940000  62.240000 ;
      RECT 398.150000  63.950000 400.560000  64.130000 ;
      RECT 398.150000  64.130000 398.330000  75.235000 ;
      RECT 398.150000  75.235000 400.290000  75.415000 ;
      RECT 398.150000  75.415000 398.330000  86.330000 ;
      RECT 398.150000  86.330000 400.290000  86.510000 ;
      RECT 398.150000  86.510000 398.330000  97.430000 ;
      RECT 398.150000  97.430000 400.290000  97.610000 ;
      RECT 398.150000  97.610000 398.330000 108.715000 ;
      RECT 398.150000 108.715000 424.780000 108.895000 ;
      RECT 398.165000 109.115000 398.755000 109.435000 ;
      RECT 398.165000 109.435000 398.590000 110.595000 ;
      RECT 398.195000 220.080000 398.805000 220.580000 ;
      RECT 398.195000 236.540000 398.805000 237.040000 ;
      RECT 398.215000 218.520000 398.805000 218.690000 ;
      RECT 398.215000 238.530000 398.805000 238.700000 ;
      RECT 398.220000 155.420000 399.750000 155.750000 ;
      RECT 398.225000 222.650000 398.395000 225.360000 ;
      RECT 398.225000 231.760000 398.395000 234.470000 ;
      RECT 398.240000   9.660000 398.570000  10.280000 ;
      RECT 398.240000  27.735000 398.570000  29.855000 ;
      RECT 398.240000  33.580000 398.570000  35.075000 ;
      RECT 398.255000 248.995000 399.635000 249.165000 ;
      RECT 398.270000 246.775000 398.535000 248.075000 ;
      RECT 398.385000 226.270000 398.555000 227.580000 ;
      RECT 398.385000 229.540000 398.555000 230.850000 ;
      RECT 398.430000 218.690000 398.805000 220.080000 ;
      RECT 398.430000 237.040000 398.805000 238.530000 ;
      RECT 398.590000 249.475000 399.200000 252.915000 ;
      RECT 398.595000 145.700000 398.765000 146.115000 ;
      RECT 398.595000 146.115000 399.205000 147.125000 ;
      RECT 398.595000 248.605000 399.125000 248.775000 ;
      RECT 398.715000 247.065000 398.995000 248.605000 ;
      RECT 398.720000 207.340000 398.890000 210.050000 ;
      RECT 398.720000 241.395000 398.890000 244.105000 ;
      RECT 398.740000  40.920000 398.910000  50.770000 ;
      RECT 398.740000  51.380000 398.910000  61.230000 ;
      RECT 398.740000  64.770000 398.910000  74.660000 ;
      RECT 398.740000  75.840000 398.910000  85.730000 ;
      RECT 398.740000  86.965000 398.910000  96.855000 ;
      RECT 398.740000  98.035000 398.910000 107.925000 ;
      RECT 398.760000 110.605000 398.940000 120.970000 ;
      RECT 398.765000 109.660000 407.190000 109.840000 ;
      RECT 398.765000 110.405000 398.935000 110.605000 ;
      RECT 398.805000 220.980000 398.975000 221.650000 ;
      RECT 398.805000 235.470000 398.975000 236.070000 ;
      RECT 398.805000 236.070000 399.335000 236.240000 ;
      RECT 398.815000 226.570000 399.325000 227.580000 ;
      RECT 398.815000 229.540000 399.325000 230.550000 ;
      RECT 398.870000   9.660000 399.200000  10.310000 ;
      RECT 398.870000  27.295000 399.200000  29.855000 ;
      RECT 398.870000  33.580000 399.200000  35.075000 ;
      RECT 398.945000 145.535000 419.985000 145.715000 ;
      RECT 399.005000 218.520000 399.595000 218.690000 ;
      RECT 399.005000 218.690000 399.550000 220.220000 ;
      RECT 399.005000 236.900000 399.550000 238.530000 ;
      RECT 399.005000 238.530000 399.595000 238.700000 ;
      RECT 399.010000   3.170000 399.180000   4.180000 ;
      RECT 399.010000   6.620000 399.180000   7.630000 ;
      RECT 399.090000 207.540000 399.395000 210.325000 ;
      RECT 399.090000 241.215000 399.395000 243.905000 ;
      RECT 399.100000  40.330000 402.830000  40.340000 ;
      RECT 399.100000  40.340000 407.110000  40.745000 ;
      RECT 399.100000  61.405000 407.110000  61.810000 ;
      RECT 399.100000  64.380000 402.830000  64.550000 ;
      RECT 399.100000 108.295000 402.830000 108.465000 ;
      RECT 399.180000 246.775000 399.445000 248.075000 ;
      RECT 399.195000 220.470000 399.865000 220.640000 ;
      RECT 399.195000 236.480000 399.865000 236.650000 ;
      RECT 399.235000   4.425000 401.115000   4.595000 ;
      RECT 399.235000   6.220000 401.235000   6.390000 ;
      RECT 399.300000 183.610000 399.470000 188.370000 ;
      RECT 399.350000 110.765000 399.520000 120.655000 ;
      RECT 399.470000 222.890000 400.000000 223.900000 ;
      RECT 399.470000 224.570000 400.000000 225.580000 ;
      RECT 399.470000 231.540000 400.000000 232.550000 ;
      RECT 399.470000 233.220000 400.000000 234.230000 ;
      RECT 399.500000   9.660000 399.830000  10.310000 ;
      RECT 399.500000  27.735000 399.830000  29.855000 ;
      RECT 399.500000  33.580000 399.830000  35.075000 ;
      RECT 399.590000 249.565000 400.520000 252.425000 ;
      RECT 399.600000 207.340000 400.920000 210.110000 ;
      RECT 399.600000 241.335000 400.920000 244.105000 ;
      RECT 399.635000 146.115000 400.165000 147.145000 ;
      RECT 399.690000 110.375000 406.260000 110.545000 ;
      RECT 399.690000 121.025000 400.360000 121.195000 ;
      RECT 399.690000 247.065000 399.860000 248.075000 ;
      RECT 399.755000 122.555000 399.925000 129.565000 ;
      RECT 399.755000 130.205000 399.925000 137.215000 ;
      RECT 399.755000 137.855000 399.925000 144.645000 ;
      RECT 399.835000 235.640000 400.365000 235.810000 ;
      RECT 399.875000 224.150000 403.135000 224.320000 ;
      RECT 399.875000 232.800000 403.135000 232.970000 ;
      RECT 399.885000 219.125000 400.415000 220.220000 ;
      RECT 399.885000 236.900000 400.055000 238.260000 ;
      RECT 400.040000 148.220000 400.210000 155.230000 ;
      RECT 400.040000 157.395000 400.210000 162.245000 ;
      RECT 400.040000 163.355000 400.210000 168.205000 ;
      RECT 400.040000 169.315000 400.210000 174.165000 ;
      RECT 400.040000 175.275000 400.210000 180.125000 ;
      RECT 400.085000 220.980000 400.255000 221.870000 ;
      RECT 400.085000 235.470000 400.255000 235.640000 ;
      RECT 400.085000 235.810000 400.255000 236.140000 ;
      RECT 400.085000 248.605000 400.755000 248.775000 ;
      RECT 400.090000   3.170000 400.260000   4.195000 ;
      RECT 400.095000 246.775000 400.360000 248.075000 ;
      RECT 400.135000 122.165000 401.825000 122.335000 ;
      RECT 400.135000 129.815000 401.825000 129.985000 ;
      RECT 400.135000 144.890000 401.825000 145.285000 ;
      RECT 400.200000   9.250000 400.380000  35.485000 ;
      RECT 400.460000  75.235000 401.470000  75.405000 ;
      RECT 400.460000  86.330000 401.470000  86.500000 ;
      RECT 400.460000  97.430000 401.470000  97.600000 ;
      RECT 400.480000 162.575000 404.050000 162.905000 ;
      RECT 400.480000 168.535000 404.050000 168.865000 ;
      RECT 400.480000 174.495000 404.050000 174.825000 ;
      RECT 400.480000 180.455000 404.050000 180.785000 ;
      RECT 400.500000 155.420000 402.030000 155.750000 ;
      RECT 400.530000 110.545000 400.700000 120.655000 ;
      RECT 400.580000 183.610000 400.750000 188.360000 ;
      RECT 400.600000   3.605000 400.830000   4.425000 ;
      RECT 400.600000 226.570000 401.110000 227.580000 ;
      RECT 400.600000 229.540000 401.110000 230.550000 ;
      RECT 400.650000 222.890000 401.180000 223.900000 ;
      RECT 400.650000 233.220000 401.180000 234.230000 ;
      RECT 400.730000  63.505000 401.260000  64.380000 ;
      RECT 400.775000 224.560000 401.055000 225.770000 ;
      RECT 400.775000 225.770000 403.400000 226.020000 ;
      RECT 400.775000 231.100000 403.400000 231.350000 ;
      RECT 400.775000 231.350000 401.055000 232.560000 ;
      RECT 400.810000 249.565000 401.190000 252.275000 ;
      RECT 400.870000 121.025000 401.540000 121.195000 ;
      RECT 400.935000 206.950000 401.605000 207.120000 ;
      RECT 400.935000 244.325000 401.605000 244.495000 ;
      RECT 400.935000 247.405000 401.190000 249.565000 ;
      RECT 401.145000   8.010000 425.580000   8.125000 ;
      RECT 401.145000   8.305000 401.325000  12.285000 ;
      RECT 401.165000 227.830000 402.605000 228.000000 ;
      RECT 401.165000 229.120000 402.605000 229.290000 ;
      RECT 401.170000   3.170000 401.340000   4.180000 ;
      RECT 401.290000   6.620000 401.460000   7.630000 ;
      RECT 401.300000 222.000000 402.200000 222.140000 ;
      RECT 401.300000 222.140000 401.830000 222.170000 ;
      RECT 401.315000 226.020000 401.595000 227.590000 ;
      RECT 401.315000 229.530000 401.595000 231.100000 ;
      RECT 401.350000 218.710000 401.520000 221.420000 ;
      RECT 401.370000 248.605000 401.900000 248.775000 ;
      RECT 401.370000 248.775000 401.760000 252.275000 ;
      RECT 401.430000  63.950000 405.340000  64.130000 ;
      RECT 401.435000 244.695000 402.105000 248.415000 ;
      RECT 401.530000 221.970000 402.200000 222.000000 ;
      RECT 401.630000 207.340000 401.800000 210.050000 ;
      RECT 401.630000 241.395000 401.800000 244.105000 ;
      RECT 401.640000  75.235000 404.570000  75.415000 ;
      RECT 401.640000  86.330000 404.570000  86.510000 ;
      RECT 401.640000  97.430000 404.570000  97.610000 ;
      RECT 401.655000 234.950000 402.185000 234.980000 ;
      RECT 401.655000 234.980000 402.555000 235.120000 ;
      RECT 401.705000 235.700000 401.875000 238.410000 ;
      RECT 401.710000 110.765000 401.880000 120.655000 ;
      RECT 401.750000   2.820000 401.930000   4.845000 ;
      RECT 401.800000 226.570000 401.970000 227.580000 ;
      RECT 401.800000 229.540000 401.970000 230.550000 ;
      RECT 401.815000 222.890000 402.345000 223.900000 ;
      RECT 401.815000 224.570000 402.345000 225.580000 ;
      RECT 401.815000 231.540000 402.345000 232.550000 ;
      RECT 401.815000 233.220000 402.345000 234.230000 ;
      RECT 401.860000 183.610000 402.030000 188.370000 ;
      RECT 401.885000 235.120000 402.555000 235.150000 ;
      RECT 401.945000 249.565000 402.875000 252.425000 ;
      RECT 402.035000 122.555000 402.205000 129.565000 ;
      RECT 402.035000 130.205000 402.205000 137.215000 ;
      RECT 402.035000 137.855000 402.205000 144.645000 ;
      RECT 402.050000 121.025000 402.720000 121.195000 ;
      RECT 402.090000  29.290000 412.720000  29.470000 ;
      RECT 402.090000  29.470000 402.270000  35.490000 ;
      RECT 402.090000  35.490000 411.535000  35.670000 ;
      RECT 402.175000 226.020000 402.455000 227.590000 ;
      RECT 402.175000 229.530000 402.455000 231.100000 ;
      RECT 402.230000 218.710000 402.400000 221.420000 ;
      RECT 402.320000 148.240000 402.490000 155.230000 ;
      RECT 402.415000 122.165000 404.105000 122.335000 ;
      RECT 402.415000 129.815000 404.105000 129.985000 ;
      RECT 402.415000 144.890000 404.105000 145.285000 ;
      RECT 402.460000   5.970000 402.640000   8.010000 ;
      RECT 402.460000   8.180000 402.630000  12.170000 ;
      RECT 402.460000  12.780000 402.630000  15.700000 ;
      RECT 402.460000  15.700000 438.335000  15.870000 ;
      RECT 402.460000  15.870000 402.630000  16.435000 ;
      RECT 402.460000  16.605000 405.310000  16.775000 ;
      RECT 402.460000  16.775000 402.630000  17.385000 ;
      RECT 402.460000  17.555000 402.630000  28.155000 ;
      RECT 402.460000  28.155000 444.675000  28.325000 ;
      RECT 402.585000 235.700000 402.755000 238.410000 ;
      RECT 402.660000 226.570000 403.170000 227.580000 ;
      RECT 402.660000 229.540000 403.170000 230.550000 ;
      RECT 402.680000  29.820000 402.850000  34.570000 ;
      RECT 402.685000 222.890000 403.540000 223.900000 ;
      RECT 402.685000 233.220000 403.540000 234.230000 ;
      RECT 402.700000 206.365000 405.250000 211.275000 ;
      RECT 402.780000 155.420000 404.310000 155.750000 ;
      RECT 402.810000 246.265000 405.175000 246.775000 ;
      RECT 402.850000  15.685000 442.220000  15.700000 ;
      RECT 402.860000  22.155000 403.395000  22.730000 ;
      RECT 402.890000 110.545000 403.060000 120.655000 ;
      RECT 402.925000  16.965000 403.680000  17.135000 ;
      RECT 402.925000  17.135000 403.095000  18.735000 ;
      RECT 402.925000  18.735000 403.455000  18.905000 ;
      RECT 402.925000  18.905000 403.095000  20.825000 ;
      RECT 402.925000  20.825000 403.130000  21.835000 ;
      RECT 402.930000 248.995000 404.310000 249.165000 ;
      RECT 402.945000 246.775000 403.210000 248.075000 ;
      RECT 403.000000  35.080000 408.770000  35.250000 ;
      RECT 403.020000  40.920000 403.190000  50.770000 ;
      RECT 403.020000  51.380000 403.190000  61.230000 ;
      RECT 403.020000  64.770000 403.190000  74.660000 ;
      RECT 403.020000  75.840000 403.190000  85.730000 ;
      RECT 403.020000  86.965000 403.190000  96.855000 ;
      RECT 403.020000  98.035000 403.190000 107.925000 ;
      RECT 403.040000   8.830000 403.210000  14.590000 ;
      RECT 403.120000  22.935000 403.290000  23.040000 ;
      RECT 403.120000  23.040000 404.150000  23.210000 ;
      RECT 403.120000  23.210000 403.290000  23.605000 ;
      RECT 403.135000 224.560000 403.400000 225.770000 ;
      RECT 403.135000 231.350000 403.400000 232.560000 ;
      RECT 403.140000 183.610000 403.310000 188.360000 ;
      RECT 403.230000 121.025000 403.900000 121.195000 ;
      RECT 403.265000  19.940000 403.435000  20.610000 ;
      RECT 403.265000 249.475000 403.875000 252.915000 ;
      RECT 403.270000 248.605000 403.800000 248.775000 ;
      RECT 403.305000  23.780000 404.050000  23.950000 ;
      RECT 403.305000  23.950000 403.475000  27.230000 ;
      RECT 403.305000  27.230000 407.545000  27.400000 ;
      RECT 403.310000   8.350000 403.820000   8.680000 ;
      RECT 403.310000  14.760000 403.820000  14.840000 ;
      RECT 403.310000  14.840000 403.840000  15.010000 ;
      RECT 403.310000  15.010000 403.820000  15.090000 ;
      RECT 403.380000   8.680000 403.750000  14.760000 ;
      RECT 403.380000  40.330000 407.110000  40.340000 ;
      RECT 403.380000  64.380000 407.110000  64.550000 ;
      RECT 403.380000 108.295000 407.110000 108.465000 ;
      RECT 403.390000 247.065000 403.670000 248.605000 ;
      RECT 403.420000  20.825000 403.590000  21.835000 ;
      RECT 403.450000  23.710000 403.980000  23.780000 ;
      RECT 403.460000  27.735000 404.130000  27.905000 ;
      RECT 403.460000  29.820000 403.630000  34.570000 ;
      RECT 403.630000  19.575000 404.170000  19.865000 ;
      RECT 403.630000  19.865000 403.930000  20.500000 ;
      RECT 403.630000  20.500000 404.170000  20.655000 ;
      RECT 403.640000  22.670000 404.170000  22.840000 ;
      RECT 403.760000  20.655000 404.170000  22.670000 ;
      RECT 403.855000 246.775000 404.120000 248.075000 ;
      RECT 403.880000  17.155000 404.170000  19.575000 ;
      RECT 403.920000   9.150000 404.090000  11.860000 ;
      RECT 403.920000  12.030000 404.090000  12.560000 ;
      RECT 403.920000  12.780000 404.090000  13.355000 ;
      RECT 403.920000  13.525000 404.090000  14.590000 ;
      RECT 403.980000 218.340000 404.150000 228.475000 ;
      RECT 403.980000 228.645000 404.150000 238.890000 ;
      RECT 404.070000 110.765000 404.240000 120.655000 ;
      RECT 404.100000  20.070000 404.630000  20.240000 ;
      RECT 404.185000  24.350000 404.490000  27.060000 ;
      RECT 404.190000   8.350000 404.700000   8.680000 ;
      RECT 404.190000  14.760000 404.700000  15.090000 ;
      RECT 404.240000  29.820000 404.410000  34.570000 ;
      RECT 404.260000   8.680000 404.630000  14.760000 ;
      RECT 404.265000 249.565000 405.195000 252.425000 ;
      RECT 404.315000 122.555000 404.485000 129.565000 ;
      RECT 404.315000 130.205000 404.485000 137.215000 ;
      RECT 404.315000 137.855000 404.485000 144.645000 ;
      RECT 404.320000  22.935000 404.570000  23.605000 ;
      RECT 404.320000  23.605000 404.535000  23.660000 ;
      RECT 404.320000  23.660000 404.490000  24.350000 ;
      RECT 404.320000 157.395000 404.490000 162.245000 ;
      RECT 404.320000 163.355000 404.490000 168.205000 ;
      RECT 404.320000 169.315000 404.490000 174.165000 ;
      RECT 404.320000 175.275000 404.490000 180.125000 ;
      RECT 404.340000  17.155000 404.510000  20.070000 ;
      RECT 404.340000  20.825000 404.535000  21.835000 ;
      RECT 404.365000  21.835000 404.535000  22.935000 ;
      RECT 404.365000 247.065000 404.535000 248.075000 ;
      RECT 404.410000  27.735000 405.080000  27.905000 ;
      RECT 404.410000 121.025000 405.080000 121.195000 ;
      RECT 404.420000 183.610000 404.590000 188.370000 ;
      RECT 404.590000 222.890000 405.445000 223.900000 ;
      RECT 404.590000 233.220000 405.445000 234.230000 ;
      RECT 404.600000 148.220000 404.770000 155.230000 ;
      RECT 404.625000 162.575000 406.330000 162.905000 ;
      RECT 404.625000 168.535000 405.860000 168.865000 ;
      RECT 404.625000 174.495000 405.860000 174.825000 ;
      RECT 404.625000 180.455000 405.860000 180.785000 ;
      RECT 404.660000  23.780000 405.330000  23.950000 ;
      RECT 404.695000 122.165000 406.385000 122.335000 ;
      RECT 404.695000 129.815000 406.385000 129.985000 ;
      RECT 404.695000 144.890000 406.385000 145.285000 ;
      RECT 404.730000 224.560000 404.995000 225.770000 ;
      RECT 404.730000 225.770000 407.355000 226.020000 ;
      RECT 404.730000 231.100000 407.355000 231.350000 ;
      RECT 404.730000 231.350000 404.995000 232.560000 ;
      RECT 404.740000  23.040000 405.270000  23.210000 ;
      RECT 404.740000  23.210000 405.235000  23.780000 ;
      RECT 404.740000  75.235000 405.750000  75.405000 ;
      RECT 404.740000  86.330000 405.750000  86.500000 ;
      RECT 404.740000  97.430000 405.750000  97.600000 ;
      RECT 404.760000 248.605000 405.430000 248.775000 ;
      RECT 404.770000 246.775000 405.035000 248.075000 ;
      RECT 404.800000   8.830000 404.970000  14.465000 ;
      RECT 404.800000  17.155000 404.970000  18.735000 ;
      RECT 404.800000  18.735000 405.330000  18.905000 ;
      RECT 404.800000  18.905000 404.970000  20.825000 ;
      RECT 404.800000  20.825000 405.450000  21.835000 ;
      RECT 404.960000 226.570000 405.470000 227.580000 ;
      RECT 404.960000 229.540000 405.470000 230.550000 ;
      RECT 404.995000 224.150000 408.255000 224.320000 ;
      RECT 404.995000 232.800000 408.255000 232.970000 ;
      RECT 405.010000  14.760000 405.580000  15.090000 ;
      RECT 405.020000  29.820000 405.190000  34.570000 ;
      RECT 405.065000  23.950000 405.235000  27.060000 ;
      RECT 405.070000   8.350000 405.580000   8.680000 ;
      RECT 405.100000 157.045000 405.860000 162.320000 ;
      RECT 405.100000 163.170000 405.860000 168.535000 ;
      RECT 405.100000 168.865000 405.860000 174.495000 ;
      RECT 405.100000 174.825000 405.860000 180.455000 ;
      RECT 405.100000 180.785000 405.860000 180.955000 ;
      RECT 405.140000   8.680000 405.510000  14.760000 ;
      RECT 405.140000  16.775000 405.310000  17.385000 ;
      RECT 405.235000 155.420000 406.050000 155.750000 ;
      RECT 405.250000 110.545000 405.420000 120.655000 ;
      RECT 405.280000  21.835000 405.450000  22.595000 ;
      RECT 405.280000  22.595000 407.940000  22.765000 ;
      RECT 405.290000  27.655000 408.825000  27.905000 ;
      RECT 405.375000 235.700000 405.545000 238.410000 ;
      RECT 405.485000 249.565000 405.865000 252.275000 ;
      RECT 405.500000  23.710000 406.030000  23.880000 ;
      RECT 405.510000  63.505000 406.040000  64.380000 ;
      RECT 405.525000 227.830000 406.965000 228.000000 ;
      RECT 405.525000 229.120000 406.965000 229.290000 ;
      RECT 405.575000 234.980000 406.475000 235.120000 ;
      RECT 405.575000 235.120000 406.245000 235.150000 ;
      RECT 405.590000 121.025000 406.260000 121.195000 ;
      RECT 405.610000 247.405000 405.865000 249.565000 ;
      RECT 405.620000  16.850000 405.790000  21.975000 ;
      RECT 405.620000  21.975000 406.150000  22.145000 ;
      RECT 405.630000 194.520000 405.800000 198.250000 ;
      RECT 405.675000 226.020000 405.955000 227.590000 ;
      RECT 405.675000 229.530000 405.955000 231.100000 ;
      RECT 405.680000   9.150000 405.850000  11.860000 ;
      RECT 405.680000  12.770000 405.850000  14.590000 ;
      RECT 405.680000  22.935000 405.850000  23.710000 ;
      RECT 405.680000 163.075000 405.860000 163.170000 ;
      RECT 405.700000 183.610000 405.870000 188.360000 ;
      RECT 405.730000 218.710000 405.900000 221.420000 ;
      RECT 405.785000 222.890000 406.315000 223.900000 ;
      RECT 405.785000 224.570000 406.315000 225.580000 ;
      RECT 405.785000 231.540000 406.315000 232.550000 ;
      RECT 405.785000 233.220000 406.315000 234.230000 ;
      RECT 405.800000  14.760000 406.330000  14.930000 ;
      RECT 405.800000  29.820000 405.970000  34.570000 ;
      RECT 405.880000 148.220000 406.050000 155.420000 ;
      RECT 405.890000   1.970000 477.515000   6.600000 ;
      RECT 405.920000  75.235000 408.850000  75.415000 ;
      RECT 405.920000  86.330000 408.850000  86.510000 ;
      RECT 405.920000  97.430000 408.850000  97.610000 ;
      RECT 405.930000 221.970000 406.600000 222.000000 ;
      RECT 405.930000 222.000000 406.830000 222.140000 ;
      RECT 405.945000  24.080000 406.205000  27.060000 ;
      RECT 405.945000 234.950000 406.475000 234.980000 ;
      RECT 405.960000  16.520000 408.850000  16.690000 ;
      RECT 405.960000  16.690000 406.490000  17.870000 ;
      RECT 405.960000  17.870000 406.150000  20.890000 ;
      RECT 405.960000  20.890000 407.780000  21.060000 ;
      RECT 406.020000  14.445000 406.400000  14.615000 ;
      RECT 406.020000  14.615000 406.330000  14.760000 ;
      RECT 406.045000 248.605000 406.575000 248.775000 ;
      RECT 406.045000 248.775000 406.435000 252.275000 ;
      RECT 406.110000 245.110000 406.780000 248.415000 ;
      RECT 406.160000 162.315000 406.330000 162.575000 ;
      RECT 406.160000 226.570000 406.330000 227.580000 ;
      RECT 406.160000 229.540000 406.330000 230.550000 ;
      RECT 406.210000  63.950000 409.950000  64.130000 ;
      RECT 406.230000   8.845000 406.400000  14.445000 ;
      RECT 406.255000 235.700000 406.425000 238.410000 ;
      RECT 406.280000 194.330000 415.820000 198.440000 ;
      RECT 406.300000 222.140000 406.830000 222.170000 ;
      RECT 406.320000  18.160000 406.490000  19.790000 ;
      RECT 406.320000  19.790000 406.850000  19.960000 ;
      RECT 406.320000  19.960000 406.490000  20.660000 ;
      RECT 406.320000  21.230000 406.490000  22.400000 ;
      RECT 406.330000 207.340000 406.500000 210.050000 ;
      RECT 406.330000 241.395000 406.500000 244.105000 ;
      RECT 406.405000  24.080000 406.665000  27.060000 ;
      RECT 406.430000 110.765000 406.600000 120.655000 ;
      RECT 406.500000   8.350000 407.010000   8.680000 ;
      RECT 406.500000  14.760000 407.030000  15.300000 ;
      RECT 406.525000 206.950000 407.195000 207.120000 ;
      RECT 406.525000 244.325000 407.195000 244.495000 ;
      RECT 406.535000 226.020000 406.815000 227.590000 ;
      RECT 406.535000 229.530000 406.815000 231.100000 ;
      RECT 406.570000   8.680000 406.940000  14.760000 ;
      RECT 406.580000  29.820000 406.750000  34.570000 ;
      RECT 406.590000  22.765000 407.940000  22.770000 ;
      RECT 406.595000 122.555000 406.765000 129.565000 ;
      RECT 406.595000 130.205000 406.765000 137.215000 ;
      RECT 406.595000 137.855000 406.765000 144.645000 ;
      RECT 406.610000 218.710000 406.780000 221.420000 ;
      RECT 406.620000 249.565000 407.550000 252.425000 ;
      RECT 406.625000 145.715000 406.805000 147.710000 ;
      RECT 406.625000 147.890000 406.805000 155.920000 ;
      RECT 406.625000 156.100000 406.805000 182.010000 ;
      RECT 406.750000  21.060000 406.920000  22.400000 ;
      RECT 406.800000  16.860000 407.670000  17.870000 ;
      RECT 406.800000  17.870000 407.330000  18.905000 ;
      RECT 406.820000 122.165000 407.545000 122.335000 ;
      RECT 406.820000 129.815000 407.545000 129.985000 ;
      RECT 406.820000 137.465000 407.545000 137.635000 ;
      RECT 406.820000 145.115000 407.545000 145.285000 ;
      RECT 406.950000 222.890000 407.480000 223.900000 ;
      RECT 406.950000 233.220000 407.480000 234.230000 ;
      RECT 406.980000 183.610000 407.150000 188.370000 ;
      RECT 407.010000 110.605000 407.190000 120.970000 ;
      RECT 407.015000 110.405000 407.185000 110.605000 ;
      RECT 407.020000 226.570000 407.530000 227.580000 ;
      RECT 407.020000 229.540000 407.530000 230.550000 ;
      RECT 407.075000 224.560000 407.355000 225.770000 ;
      RECT 407.075000 231.350000 407.355000 232.560000 ;
      RECT 407.110000   9.150000 407.280000  11.860000 ;
      RECT 407.110000  12.030000 407.280000  12.560000 ;
      RECT 407.110000  12.780000 407.280000  13.310000 ;
      RECT 407.110000  13.540000 407.280000  14.590000 ;
      RECT 407.175000 146.300000 407.345000 155.175000 ;
      RECT 407.180000  21.230000 407.350000  22.400000 ;
      RECT 407.195000 109.115000 408.895000 109.435000 ;
      RECT 407.210000 207.340000 408.530000 210.110000 ;
      RECT 407.210000 241.335000 408.530000 244.105000 ;
      RECT 407.300000  40.920000 407.470000  50.770000 ;
      RECT 407.300000  51.380000 407.470000  61.230000 ;
      RECT 407.300000  64.770000 407.470000  74.660000 ;
      RECT 407.300000  75.840000 407.470000  85.730000 ;
      RECT 407.300000  86.965000 407.470000  96.855000 ;
      RECT 407.300000  98.035000 407.470000 107.925000 ;
      RECT 407.340000 188.870000 407.670000 189.040000 ;
      RECT 407.360000  29.820000 407.530000  34.570000 ;
      RECT 407.360000 109.435000 407.785000 111.295000 ;
      RECT 407.375000  23.710000 407.905000  23.880000 ;
      RECT 407.375000  23.880000 407.545000  27.230000 ;
      RECT 407.375000 122.335000 407.545000 129.815000 ;
      RECT 407.375000 129.985000 407.545000 137.465000 ;
      RECT 407.375000 137.635000 407.545000 145.115000 ;
      RECT 407.380000   8.350000 407.890000   8.680000 ;
      RECT 407.380000  14.760000 407.910000  14.930000 ;
      RECT 407.380000  14.930000 407.890000  15.090000 ;
      RECT 407.420000 188.110000 407.590000 188.870000 ;
      RECT 407.450000   8.680000 407.820000  14.760000 ;
      RECT 407.485000 246.265000 409.850000 246.775000 ;
      RECT 407.500000  18.160000 407.670000  19.310000 ;
      RECT 407.500000  19.310000 410.030000  19.480000 ;
      RECT 407.500000  19.480000 407.670000  20.660000 ;
      RECT 407.570000 145.910000 413.000000 146.080000 ;
      RECT 407.570000 156.865000 419.040000 157.045000 ;
      RECT 407.570000 157.045000 408.330000 162.575000 ;
      RECT 407.570000 162.575000 408.805000 162.905000 ;
      RECT 407.570000 162.905000 408.330000 168.535000 ;
      RECT 407.570000 168.535000 408.805000 168.865000 ;
      RECT 407.570000 168.865000 408.330000 174.495000 ;
      RECT 407.570000 174.495000 408.805000 174.825000 ;
      RECT 407.570000 174.825000 408.330000 180.455000 ;
      RECT 407.570000 180.455000 408.805000 180.785000 ;
      RECT 407.570000 180.785000 408.330000 180.955000 ;
      RECT 407.570000 180.955000 419.040000 181.135000 ;
      RECT 407.605000 248.995000 408.985000 249.165000 ;
      RECT 407.610000  21.060000 407.780000  22.400000 ;
      RECT 407.620000 246.775000 407.885000 248.075000 ;
      RECT 407.660000  64.380000 411.390000  64.550000 ;
      RECT 407.660000 108.295000 411.390000 108.465000 ;
      RECT 407.665000 146.300000 408.415000 155.305000 ;
      RECT 407.715000 219.125000 408.245000 220.220000 ;
      RECT 407.765000 235.640000 408.295000 235.810000 ;
      RECT 407.780000 121.915000 408.310000 145.535000 ;
      RECT 407.860000 183.610000 408.030000 188.360000 ;
      RECT 407.875000 220.980000 408.045000 221.870000 ;
      RECT 407.875000 235.470000 408.045000 235.640000 ;
      RECT 407.875000 235.810000 408.045000 236.140000 ;
      RECT 407.940000 249.475000 408.550000 252.915000 ;
      RECT 407.945000 248.605000 408.475000 248.775000 ;
      RECT 407.955000  24.370000 408.125000  27.370000 ;
      RECT 407.955000  40.090000 408.135000  62.060000 ;
      RECT 407.955000 109.660000 408.135000 121.735000 ;
      RECT 407.990000   8.845000 408.160000  14.590000 ;
      RECT 408.020000  18.225000 408.350000  19.075000 ;
      RECT 408.040000  21.230000 408.210000  22.400000 ;
      RECT 408.065000 247.065000 408.345000 248.605000 ;
      RECT 408.075000 236.900000 408.245000 238.260000 ;
      RECT 408.100000  17.615000 408.270000  18.225000 ;
      RECT 408.130000 222.890000 408.660000 223.900000 ;
      RECT 408.130000 224.570000 408.660000 225.580000 ;
      RECT 408.130000 231.540000 408.660000 232.550000 ;
      RECT 408.130000 233.220000 408.660000 234.230000 ;
      RECT 408.140000  29.820000 408.310000  34.570000 ;
      RECT 408.175000  19.790000 408.850000  19.960000 ;
      RECT 408.250000 188.870000 412.905000 189.040000 ;
      RECT 408.260000   8.350000 409.650000   8.680000 ;
      RECT 408.260000  14.760000 409.650000  15.090000 ;
      RECT 408.265000 220.470000 408.935000 220.640000 ;
      RECT 408.265000 236.480000 408.935000 236.650000 ;
      RECT 408.295000  22.570000 409.545000  22.600000 ;
      RECT 408.295000  22.600000 409.645000  22.770000 ;
      RECT 408.295000  25.395000 408.825000  27.655000 ;
      RECT 408.305000 109.435000 408.730000 111.295000 ;
      RECT 408.330000   8.680000 408.700000  14.760000 ;
      RECT 408.470000  20.890000 410.030000  21.060000 ;
      RECT 408.470000  21.060000 408.640000  22.400000 ;
      RECT 408.530000 246.775000 408.795000 248.075000 ;
      RECT 408.535000 218.520000 409.125000 218.690000 ;
      RECT 408.535000 238.530000 409.125000 238.700000 ;
      RECT 408.545000 122.165000 409.270000 122.335000 ;
      RECT 408.545000 122.335000 408.715000 129.815000 ;
      RECT 408.545000 129.815000 409.270000 129.985000 ;
      RECT 408.545000 129.985000 408.715000 137.465000 ;
      RECT 408.545000 137.465000 409.270000 137.635000 ;
      RECT 408.545000 137.635000 408.715000 145.115000 ;
      RECT 408.545000 145.115000 409.270000 145.285000 ;
      RECT 408.560000 210.325000 410.760000 210.995000 ;
      RECT 408.560000 240.675000 410.760000 240.845000 ;
      RECT 408.580000 218.690000 409.125000 220.220000 ;
      RECT 408.580000 236.900000 409.125000 238.530000 ;
      RECT 408.620000  40.920000 408.790000  50.770000 ;
      RECT 408.620000  51.380000 408.790000  61.230000 ;
      RECT 408.680000  16.690000 408.850000  19.140000 ;
      RECT 408.680000  19.650000 408.850000  19.790000 ;
      RECT 408.680000  19.960000 408.850000  20.660000 ;
      RECT 408.735000 146.300000 408.905000 155.175000 ;
      RECT 408.735000 207.540000 409.040000 210.325000 ;
      RECT 408.735000 240.845000 410.760000 241.215000 ;
      RECT 408.735000 241.215000 409.040000 243.905000 ;
      RECT 408.795000 236.070000 409.325000 236.240000 ;
      RECT 408.805000 226.570000 409.315000 227.580000 ;
      RECT 408.805000 229.540000 409.315000 230.550000 ;
      RECT 408.870000   9.150000 409.040000  11.860000 ;
      RECT 408.870000  12.030000 409.040000  12.560000 ;
      RECT 408.870000  12.980000 409.040000  13.310000 ;
      RECT 408.870000  13.540000 409.040000  14.590000 ;
      RECT 408.900000  21.230000 409.070000  22.400000 ;
      RECT 408.900000 109.660000 417.330000 109.840000 ;
      RECT 408.900000 110.605000 409.080000 120.970000 ;
      RECT 408.920000  29.820000 409.090000  34.570000 ;
      RECT 408.940000 157.395000 409.110000 162.245000 ;
      RECT 408.940000 163.355000 409.110000 168.205000 ;
      RECT 408.940000 169.315000 409.110000 174.165000 ;
      RECT 408.940000 175.275000 409.110000 180.125000 ;
      RECT 408.940000 249.565000 409.870000 252.425000 ;
      RECT 408.980000  40.330000 412.710000  40.340000 ;
      RECT 408.980000  40.340000 416.990000  40.745000 ;
      RECT 408.980000  61.405000 416.990000  61.810000 ;
      RECT 409.020000  75.235000 410.030000  75.405000 ;
      RECT 409.020000  86.330000 410.030000  86.500000 ;
      RECT 409.020000  97.430000 410.030000  97.600000 ;
      RECT 409.040000 247.065000 409.210000 248.075000 ;
      RECT 409.140000 183.610000 409.310000 188.360000 ;
      RECT 409.155000 220.980000 409.325000 221.650000 ;
      RECT 409.155000 235.470000 409.325000 236.070000 ;
      RECT 409.210000   8.680000 409.580000  14.760000 ;
      RECT 409.210000  35.080000 410.560000  35.250000 ;
      RECT 409.240000 207.340000 409.410000 210.050000 ;
      RECT 409.240000 241.395000 409.410000 244.105000 ;
      RECT 409.300000  24.395000 409.470000  27.475000 ;
      RECT 409.325000 122.555000 409.495000 129.565000 ;
      RECT 409.325000 130.205000 409.495000 137.215000 ;
      RECT 409.325000 137.855000 409.495000 144.645000 ;
      RECT 409.325000 218.520000 409.915000 218.690000 ;
      RECT 409.325000 218.690000 409.700000 220.080000 ;
      RECT 409.325000 220.080000 409.935000 220.580000 ;
      RECT 409.325000 220.580000 410.300000 220.790000 ;
      RECT 409.325000 236.420000 410.300000 236.540000 ;
      RECT 409.325000 236.540000 409.935000 237.040000 ;
      RECT 409.325000 237.040000 409.700000 238.530000 ;
      RECT 409.325000 238.530000 409.915000 238.700000 ;
      RECT 409.330000  21.060000 409.500000  22.400000 ;
      RECT 409.370000 227.830000 410.810000 228.000000 ;
      RECT 409.370000 229.120000 410.810000 229.290000 ;
      RECT 409.380000 162.575000 412.950000 162.905000 ;
      RECT 409.380000 168.535000 412.950000 168.865000 ;
      RECT 409.380000 174.495000 412.950000 174.825000 ;
      RECT 409.380000 180.455000 412.950000 180.785000 ;
      RECT 409.435000 248.605000 410.105000 248.775000 ;
      RECT 409.445000 246.775000 409.710000 248.075000 ;
      RECT 409.490000 110.765000 409.660000 120.655000 ;
      RECT 409.500000  18.735000 410.030000  18.905000 ;
      RECT 409.515000 146.300000 410.270000 152.785000 ;
      RECT 409.515000 152.785000 409.685000 155.175000 ;
      RECT 409.575000 226.270000 409.745000 227.580000 ;
      RECT 409.575000 229.540000 409.745000 230.850000 ;
      RECT 409.580000 220.790000 410.300000 221.650000 ;
      RECT 409.580000 235.470000 410.300000 236.420000 ;
      RECT 409.625000  22.940000 410.155000  23.110000 ;
      RECT 409.625000  23.110000 409.935000  23.805000 ;
      RECT 409.625000  23.805000 410.590000  23.975000 ;
      RECT 409.705000 122.165000 411.395000 122.335000 ;
      RECT 409.705000 129.815000 411.395000 129.985000 ;
      RECT 409.705000 144.890000 411.395000 145.285000 ;
      RECT 409.735000 222.650000 409.905000 225.360000 ;
      RECT 409.735000 231.760000 409.905000 234.470000 ;
      RECT 409.750000   8.830000 409.920000  14.590000 ;
      RECT 409.760000  21.230000 409.930000  22.400000 ;
      RECT 409.765000  24.145000 409.935000  24.375000 ;
      RECT 409.765000  24.375000 410.050000  27.085000 ;
      RECT 409.800000  29.820000 409.970000  34.570000 ;
      RECT 409.830000 110.375000 416.400000 110.545000 ;
      RECT 409.830000 121.025000 410.500000 121.195000 ;
      RECT 409.860000  16.860000 410.030000  18.735000 ;
      RECT 409.860000  18.905000 410.030000  19.140000 ;
      RECT 409.860000  19.480000 410.030000  20.890000 ;
      RECT 409.900000 219.185000 410.430000 219.880000 ;
      RECT 409.900000 237.240000 410.070000 238.260000 ;
      RECT 409.960000 225.910000 412.100000 226.080000 ;
      RECT 409.960000 231.040000 412.100000 231.210000 ;
      RECT 410.005000 226.570000 410.175000 227.600000 ;
      RECT 410.005000 229.520000 410.175000 230.550000 ;
      RECT 410.020000   8.350000 410.530000   8.680000 ;
      RECT 410.020000  14.760000 410.530000  15.090000 ;
      RECT 410.090000   8.680000 410.460000  14.760000 ;
      RECT 410.090000 207.440000 410.760000 207.610000 ;
      RECT 410.090000 208.220000 410.820000 209.540000 ;
      RECT 410.090000 210.150000 410.760000 210.325000 ;
      RECT 410.090000 241.215000 410.760000 241.295000 ;
      RECT 410.090000 241.905000 410.820000 243.225000 ;
      RECT 410.090000 243.835000 410.760000 244.495000 ;
      RECT 410.105000  23.310000 410.635000  23.480000 ;
      RECT 410.105000  23.975000 410.590000  23.985000 ;
      RECT 410.105000  23.985000 410.775000  24.155000 ;
      RECT 410.105000  27.735000 412.360000  27.905000 ;
      RECT 410.120000  63.505000 410.650000  64.380000 ;
      RECT 410.125000 220.220000 411.125000 220.390000 ;
      RECT 410.125000 236.730000 411.125000 236.900000 ;
      RECT 410.160000 249.565000 410.540000 252.275000 ;
      RECT 410.200000  75.235000 414.450000  75.415000 ;
      RECT 410.200000  86.330000 414.450000  86.510000 ;
      RECT 410.200000  97.430000 414.450000  97.610000 ;
      RECT 410.220000  21.960000 410.750000  22.130000 ;
      RECT 410.220000  24.155000 410.590000  27.645000 ;
      RECT 410.220000  27.645000 412.360000  27.735000 ;
      RECT 410.255000 222.630000 410.785000 222.800000 ;
      RECT 410.255000 234.320000 410.785000 234.490000 ;
      RECT 410.285000 247.405000 410.540000 249.565000 ;
      RECT 410.325000  22.130000 410.635000  23.310000 ;
      RECT 410.420000 183.610000 410.590000 188.370000 ;
      RECT 410.435000 226.270000 410.605000 227.580000 ;
      RECT 410.435000 229.540000 410.605000 230.850000 ;
      RECT 410.440000  16.850000 410.610000  21.960000 ;
      RECT 410.615000 222.800000 410.785000 225.360000 ;
      RECT 410.615000 231.760000 410.785000 234.320000 ;
      RECT 410.630000   9.150000 410.800000  11.860000 ;
      RECT 410.630000  12.030000 410.800000  12.560000 ;
      RECT 410.630000  12.780000 410.800000  13.310000 ;
      RECT 410.630000  13.540000 410.800000  14.590000 ;
      RECT 410.670000 110.545000 410.840000 120.655000 ;
      RECT 410.670000 207.855000 411.270000 208.025000 ;
      RECT 410.670000 243.420000 411.270000 243.590000 ;
      RECT 410.680000  29.820000 410.850000  34.570000 ;
      RECT 410.720000 248.605000 411.250000 248.775000 ;
      RECT 410.720000 248.775000 411.110000 252.275000 ;
      RECT 410.760000  24.375000 410.930000  27.475000 ;
      RECT 410.785000 245.510000 411.455000 248.415000 ;
      RECT 410.805000  22.550000 411.090000  22.720000 ;
      RECT 410.805000  22.720000 410.975000  23.625000 ;
      RECT 410.805000  23.625000 411.270000  23.795000 ;
      RECT 410.820000  63.950000 413.945000  64.130000 ;
      RECT 410.865000 226.570000 411.375000 227.580000 ;
      RECT 410.865000 229.540000 411.375000 230.550000 ;
      RECT 410.880000 146.330000 411.050000 152.350000 ;
      RECT 410.880000 153.400000 411.050000 155.160000 ;
      RECT 410.880000 155.160000 411.520000 155.670000 ;
      RECT 410.900000   8.350000 411.410000   8.680000 ;
      RECT 410.900000  14.760000 411.410000  15.090000 ;
      RECT 410.905000  35.080000 411.915000  35.250000 ;
      RECT 410.920000  21.625000 411.090000  22.550000 ;
      RECT 410.970000   8.680000 411.340000  14.760000 ;
      RECT 411.010000 121.025000 411.680000 121.195000 ;
      RECT 411.010000 220.640000 411.180000 221.650000 ;
      RECT 411.010000 235.470000 411.180000 236.480000 ;
      RECT 411.095000 219.210000 412.555000 219.880000 ;
      RECT 411.095000 237.240000 412.555000 237.910000 ;
      RECT 411.100000  23.795000 411.270000  24.375000 ;
      RECT 411.100000  24.375000 411.810000  24.845000 ;
      RECT 411.100000 207.585000 411.270000 207.855000 ;
      RECT 411.100000 208.025000 411.270000 208.255000 ;
      RECT 411.100000 209.515000 411.270000 209.680000 ;
      RECT 411.100000 209.680000 412.120000 209.850000 ;
      RECT 411.100000 209.850000 411.270000 210.185000 ;
      RECT 411.100000 241.260000 411.270000 241.595000 ;
      RECT 411.100000 241.595000 412.120000 241.765000 ;
      RECT 411.100000 241.765000 411.270000 241.930000 ;
      RECT 411.100000 243.190000 411.270000 243.420000 ;
      RECT 411.100000 243.590000 411.270000 243.860000 ;
      RECT 411.145000  23.125000 411.765000  23.455000 ;
      RECT 411.275000 222.650000 411.445000 225.360000 ;
      RECT 411.275000 231.760000 411.445000 234.470000 ;
      RECT 411.295000 249.565000 412.225000 252.425000 ;
      RECT 411.370000  16.720000 414.740000  16.890000 ;
      RECT 411.370000 146.300000 412.120000 152.785000 ;
      RECT 411.410000  17.240000 411.580000  19.950000 ;
      RECT 411.440000  23.455000 411.765000  23.710000 ;
      RECT 411.440000  23.710000 412.360000  23.880000 ;
      RECT 411.470000 207.410000 412.120000 209.680000 ;
      RECT 411.470000 241.765000 412.120000 244.495000 ;
      RECT 411.510000   8.850000 411.680000  14.590000 ;
      RECT 411.530000  16.890000 414.580000  17.025000 ;
      RECT 411.580000  64.770000 411.750000  74.660000 ;
      RECT 411.580000  75.840000 411.750000  85.730000 ;
      RECT 411.580000  86.965000 411.750000  96.855000 ;
      RECT 411.580000  98.035000 411.750000 107.925000 ;
      RECT 411.605000 122.555000 411.775000 129.465000 ;
      RECT 411.605000 130.205000 411.775000 137.215000 ;
      RECT 411.605000 137.855000 411.775000 144.645000 ;
      RECT 411.640000  24.845000 411.810000  27.085000 ;
      RECT 411.660000 153.400000 411.830000 154.750000 ;
      RECT 411.700000 183.610000 411.870000 188.360000 ;
      RECT 411.705000  35.250000 411.915000  37.585000 ;
      RECT 411.705000  37.585000 412.295000  37.755000 ;
      RECT 411.780000   8.350000 413.170000   8.650000 ;
      RECT 411.780000   8.650000 412.290000   8.680000 ;
      RECT 411.780000  14.760000 412.290000  14.790000 ;
      RECT 411.780000  14.790000 413.170000  15.090000 ;
      RECT 411.800000  20.840000 411.970000  22.635000 ;
      RECT 411.815000  20.040000 412.360000  20.210000 ;
      RECT 411.850000   8.680000 412.220000  14.760000 ;
      RECT 411.850000 110.765000 412.020000 120.655000 ;
      RECT 411.905000  20.440000 412.435000  20.500000 ;
      RECT 411.905000  20.500000 412.915000  20.670000 ;
      RECT 411.960000  29.820000 412.130000  34.570000 ;
      RECT 411.970000 155.160000 412.300000 155.670000 ;
      RECT 411.980000  26.625000 412.360000  27.645000 ;
      RECT 411.985000 122.165000 413.675000 122.335000 ;
      RECT 411.985000 129.815000 413.675000 129.985000 ;
      RECT 411.985000 144.890000 413.675000 145.285000 ;
      RECT 412.020000  23.070000 412.690000  23.240000 ;
      RECT 412.050000 155.090000 412.220000 155.160000 ;
      RECT 412.085000  35.490000 412.720000  35.670000 ;
      RECT 412.090000  22.940000 412.620000  23.070000 ;
      RECT 412.155000 222.650000 412.325000 225.360000 ;
      RECT 412.155000 231.760000 412.325000 234.470000 ;
      RECT 412.160000 246.265000 414.525000 246.775000 ;
      RECT 412.190000  17.240000 412.360000  20.040000 ;
      RECT 412.190000  20.210000 412.360000  20.240000 ;
      RECT 412.190000  23.880000 412.360000  25.045000 ;
      RECT 412.190000 121.025000 412.860000 121.195000 ;
      RECT 412.235000  64.130000 412.415000  75.235000 ;
      RECT 412.235000  75.415000 412.415000  86.330000 ;
      RECT 412.235000  86.510000 412.415000  97.430000 ;
      RECT 412.235000  97.610000 412.415000 108.715000 ;
      RECT 412.280000 248.995000 413.660000 249.165000 ;
      RECT 412.290000  25.520000 413.820000  26.270000 ;
      RECT 412.295000 246.775000 412.560000 248.075000 ;
      RECT 412.320000  22.565000 412.850000  22.735000 ;
      RECT 412.390000   9.150000 412.560000  11.860000 ;
      RECT 412.390000  12.030000 412.560000  12.560000 ;
      RECT 412.390000  12.980000 412.560000  13.310000 ;
      RECT 412.390000  13.540000 412.560000  14.590000 ;
      RECT 412.440000 146.330000 412.610000 152.350000 ;
      RECT 412.440000 153.400000 412.610000 154.750000 ;
      RECT 412.530000  24.375000 413.580000  25.520000 ;
      RECT 412.530000  26.270000 413.580000  27.475000 ;
      RECT 412.540000  29.470000 412.720000  35.490000 ;
      RECT 412.575000 206.365000 413.425000 211.275000 ;
      RECT 412.615000 249.475000 413.225000 252.915000 ;
      RECT 412.620000 248.605000 413.150000 248.775000 ;
      RECT 412.660000   8.650000 413.170000   8.680000 ;
      RECT 412.660000  14.760000 413.170000  14.790000 ;
      RECT 412.680000  21.625000 412.850000  22.565000 ;
      RECT 412.730000   8.680000 413.100000  14.760000 ;
      RECT 412.740000 247.065000 413.020000 248.605000 ;
      RECT 412.750000 155.160000 413.080000 155.670000 ;
      RECT 412.830000 155.090000 413.000000 155.160000 ;
      RECT 412.900000  40.920000 413.070000  50.770000 ;
      RECT 412.900000  51.380000 413.070000  61.230000 ;
      RECT 412.900000  64.770000 413.070000  74.660000 ;
      RECT 412.900000  75.840000 413.070000  85.730000 ;
      RECT 412.900000  86.965000 413.070000  96.855000 ;
      RECT 412.900000  98.035000 413.070000 107.925000 ;
      RECT 412.930000 146.300000 413.680000 152.785000 ;
      RECT 412.935000 218.340000 413.105000 228.475000 ;
      RECT 412.935000 228.645000 415.840000 237.300000 ;
      RECT 412.935000 237.300000 420.055000 238.890000 ;
      RECT 412.970000  17.240000 413.140000  19.950000 ;
      RECT 412.980000 183.610000 413.150000 188.370000 ;
      RECT 412.980000 241.695000 418.055000 244.245000 ;
      RECT 413.030000 110.545000 413.200000 120.655000 ;
      RECT 413.195000  20.500000 414.205000  20.670000 ;
      RECT 413.205000 246.775000 413.470000 248.075000 ;
      RECT 413.220000 153.375000 413.390000 154.750000 ;
      RECT 413.220000 157.395000 413.390000 162.245000 ;
      RECT 413.220000 163.355000 413.390000 168.205000 ;
      RECT 413.220000 169.315000 413.390000 174.165000 ;
      RECT 413.220000 175.275000 413.390000 180.125000 ;
      RECT 413.260000  21.625000 413.430000  22.565000 ;
      RECT 413.260000  22.565000 413.790000  22.735000 ;
      RECT 413.260000  40.330000 416.990000  40.340000 ;
      RECT 413.260000  64.380000 416.990000  64.550000 ;
      RECT 413.260000 108.295000 416.990000 108.465000 ;
      RECT 413.270000   8.850000 413.440000  14.590000 ;
      RECT 413.280000 239.055000 420.055000 239.060000 ;
      RECT 413.370000 121.025000 414.040000 121.195000 ;
      RECT 413.370000 188.870000 414.040000 189.290000 ;
      RECT 413.420000  23.070000 414.090000  23.240000 ;
      RECT 413.485000  28.150000 444.675000  28.155000 ;
      RECT 413.485000  28.325000 413.665000  30.475000 ;
      RECT 413.485000  30.475000 414.020000  30.645000 ;
      RECT 413.485000  30.645000 413.665000  30.735000 ;
      RECT 413.485000  31.495000 413.665000  36.230000 ;
      RECT 413.485000  36.230000 432.885000  36.410000 ;
      RECT 413.485000 219.210000 414.945000 219.880000 ;
      RECT 413.490000  22.940000 414.020000  23.070000 ;
      RECT 413.530000 155.160000 413.860000 155.670000 ;
      RECT 413.540000   8.350000 414.930000   8.650000 ;
      RECT 413.540000   8.650000 414.050000   8.680000 ;
      RECT 413.540000  14.760000 414.050000  14.790000 ;
      RECT 413.540000  14.790000 414.930000  15.090000 ;
      RECT 413.610000   8.680000 413.980000  14.760000 ;
      RECT 413.610000 145.910000 419.040000 146.080000 ;
      RECT 413.610000 155.090000 413.780000 155.160000 ;
      RECT 413.615000 249.565000 414.545000 252.425000 ;
      RECT 413.660000 162.575000 417.230000 162.905000 ;
      RECT 413.660000 168.535000 417.230000 168.865000 ;
      RECT 413.660000 174.495000 417.230000 174.825000 ;
      RECT 413.660000 180.455000 417.230000 180.785000 ;
      RECT 413.675000  20.440000 414.205000  20.500000 ;
      RECT 413.715000 222.650000 413.885000 225.360000 ;
      RECT 413.715000 247.065000 413.885000 248.075000 ;
      RECT 413.750000  17.240000 413.920000  20.040000 ;
      RECT 413.750000  20.040000 414.295000  20.210000 ;
      RECT 413.750000  20.210000 413.920000  20.240000 ;
      RECT 413.750000  23.710000 414.670000  23.880000 ;
      RECT 413.750000  23.880000 413.920000  25.045000 ;
      RECT 413.750000  26.625000 414.130000  27.645000 ;
      RECT 413.750000  27.645000 415.890000  27.735000 ;
      RECT 413.750000  27.735000 416.005000  27.905000 ;
      RECT 413.855000  31.215000 414.385000  31.385000 ;
      RECT 413.855000  31.925000 414.385000  35.280000 ;
      RECT 413.885000 122.555000 414.055000 129.565000 ;
      RECT 413.885000 130.205000 414.055000 137.215000 ;
      RECT 413.885000 137.855000 414.055000 144.645000 ;
      RECT 413.910000  28.325000 444.675000  28.330000 ;
      RECT 413.920000 207.410000 414.570000 209.680000 ;
      RECT 413.920000 209.680000 414.940000 209.850000 ;
      RECT 413.940000 225.910000 416.080000 226.080000 ;
      RECT 414.000000 146.330000 414.170000 152.350000 ;
      RECT 414.000000 153.400000 414.170000 154.750000 ;
      RECT 414.075000  28.895000 414.725000  30.175000 ;
      RECT 414.110000 248.605000 414.780000 248.775000 ;
      RECT 414.120000 246.775000 414.385000 248.075000 ;
      RECT 414.140000  20.840000 414.310000  22.635000 ;
      RECT 414.150000   9.150000 414.320000  11.860000 ;
      RECT 414.150000  12.030000 414.320000  12.560000 ;
      RECT 414.150000  12.980000 414.320000  13.310000 ;
      RECT 414.150000  13.540000 414.320000  14.590000 ;
      RECT 414.155000  31.085000 414.325000  31.215000 ;
      RECT 414.155000  31.385000 414.325000  31.755000 ;
      RECT 414.185000  63.505000 414.715000  64.380000 ;
      RECT 414.210000 110.765000 414.380000 120.655000 ;
      RECT 414.260000 183.610000 414.430000 188.360000 ;
      RECT 414.265000 122.165000 415.955000 122.335000 ;
      RECT 414.265000 129.815000 415.955000 129.985000 ;
      RECT 414.265000 144.890000 415.955000 145.285000 ;
      RECT 414.300000  24.375000 415.010000  24.845000 ;
      RECT 414.300000  24.845000 414.470000  27.085000 ;
      RECT 414.310000 155.160000 414.640000 155.670000 ;
      RECT 414.345000  23.125000 414.965000  23.455000 ;
      RECT 414.345000  23.455000 414.670000  23.710000 ;
      RECT 414.390000 155.090000 414.560000 155.160000 ;
      RECT 414.420000   8.650000 414.930000   8.680000 ;
      RECT 414.420000  14.760000 414.930000  14.790000 ;
      RECT 414.490000   8.680000 414.860000  14.760000 ;
      RECT 414.490000 146.300000 415.240000 152.785000 ;
      RECT 414.495000  30.845000 415.025000  31.015000 ;
      RECT 414.500000 188.870000 417.880000 189.040000 ;
      RECT 414.530000  17.240000 414.700000  19.950000 ;
      RECT 414.550000 121.025000 415.220000 121.195000 ;
      RECT 414.555000  30.815000 415.025000  30.845000 ;
      RECT 414.555000  31.015000 415.025000  34.635000 ;
      RECT 414.595000 222.650000 414.765000 225.360000 ;
      RECT 414.620000  75.235000 415.630000  75.405000 ;
      RECT 414.620000  86.330000 415.630000  86.500000 ;
      RECT 414.620000  97.430000 415.630000  97.600000 ;
      RECT 414.665000 226.570000 415.175000 227.580000 ;
      RECT 414.770000 207.585000 414.940000 207.855000 ;
      RECT 414.770000 207.855000 415.370000 208.025000 ;
      RECT 414.770000 208.025000 414.940000 208.255000 ;
      RECT 414.770000 209.515000 414.940000 209.680000 ;
      RECT 414.770000 209.850000 414.940000 210.185000 ;
      RECT 414.780000 153.400000 414.950000 154.750000 ;
      RECT 414.835000 249.565000 415.215000 252.275000 ;
      RECT 414.840000  23.625000 415.305000  23.795000 ;
      RECT 414.840000  23.795000 415.010000  24.375000 ;
      RECT 414.860000 220.640000 415.030000 221.650000 ;
      RECT 414.915000 220.220000 415.915000 220.390000 ;
      RECT 414.960000 247.405000 415.215000 249.565000 ;
      RECT 414.990000  63.950000 417.390000  64.130000 ;
      RECT 415.020000  21.625000 415.190000  22.550000 ;
      RECT 415.020000  22.550000 415.305000  22.720000 ;
      RECT 415.030000   8.850000 415.200000  14.590000 ;
      RECT 415.090000 155.160000 415.730000 155.670000 ;
      RECT 415.135000  22.720000 415.305000  23.625000 ;
      RECT 415.180000  24.375000 415.350000  27.475000 ;
      RECT 415.195000  29.165000 415.805000  31.300000 ;
      RECT 415.195000  31.300000 416.245000  31.755000 ;
      RECT 415.195000  31.755000 415.465000  35.080000 ;
      RECT 415.195000  35.080000 416.245000  36.060000 ;
      RECT 415.220000 208.220000 415.950000 209.540000 ;
      RECT 415.230000 227.830000 416.670000 228.000000 ;
      RECT 415.255000 222.630000 415.785000 222.800000 ;
      RECT 415.255000 222.800000 415.425000 225.360000 ;
      RECT 415.280000 207.440000 415.950000 207.610000 ;
      RECT 415.280000 210.150000 415.950000 210.325000 ;
      RECT 415.280000 210.325000 417.480000 210.995000 ;
      RECT 415.295000   8.350000 416.690000   8.650000 ;
      RECT 415.295000   8.650000 415.805000   8.680000 ;
      RECT 415.300000  14.760000 415.810000  14.790000 ;
      RECT 415.300000  14.790000 416.690000  15.090000 ;
      RECT 415.335000  23.985000 416.005000  24.155000 ;
      RECT 415.360000  21.960000 415.890000  22.130000 ;
      RECT 415.370000   8.680000 415.740000  14.760000 ;
      RECT 415.390000 110.545000 415.560000 120.655000 ;
      RECT 415.435000 226.270000 415.605000 227.580000 ;
      RECT 415.475000  22.130000 415.785000  23.310000 ;
      RECT 415.475000  23.310000 416.005000  23.480000 ;
      RECT 415.500000  16.850000 415.670000  21.960000 ;
      RECT 415.520000  23.805000 416.485000  23.975000 ;
      RECT 415.520000  23.975000 416.005000  23.985000 ;
      RECT 415.520000  24.155000 415.890000  27.645000 ;
      RECT 415.540000 183.610000 415.710000 188.370000 ;
      RECT 415.560000 146.330000 415.730000 152.350000 ;
      RECT 415.560000 153.400000 415.730000 155.160000 ;
      RECT 415.610000 219.185000 416.140000 219.880000 ;
      RECT 415.635000  31.925000 415.805000  34.635000 ;
      RECT 415.730000 121.025000 416.400000 121.195000 ;
      RECT 415.740000 220.580000 416.715000 220.790000 ;
      RECT 415.740000 220.790000 416.460000 221.650000 ;
      RECT 415.800000  75.235000 417.730000  75.415000 ;
      RECT 415.800000  86.330000 417.730000  86.510000 ;
      RECT 415.800000  97.430000 417.730000  97.610000 ;
      RECT 415.865000 226.570000 416.035000 227.600000 ;
      RECT 415.910000   9.150000 416.080000  11.860000 ;
      RECT 415.910000  12.030000 416.080000  12.560000 ;
      RECT 415.910000  12.980000 416.080000  13.310000 ;
      RECT 415.910000  13.540000 416.080000  14.590000 ;
      RECT 415.955000  22.940000 416.485000  23.110000 ;
      RECT 415.975000  31.755000 416.245000  35.080000 ;
      RECT 416.060000  24.375000 416.345000  27.085000 ;
      RECT 416.075000  28.895000 416.605000  31.045000 ;
      RECT 416.080000  16.860000 416.250000  18.735000 ;
      RECT 416.080000  18.735000 416.610000  18.905000 ;
      RECT 416.080000  18.905000 416.250000  19.140000 ;
      RECT 416.080000  19.310000 418.610000  19.480000 ;
      RECT 416.080000  19.480000 416.250000  20.890000 ;
      RECT 416.080000  20.890000 417.640000  21.060000 ;
      RECT 416.105000 220.080000 416.715000 220.580000 ;
      RECT 416.125000 218.520000 416.715000 218.690000 ;
      RECT 416.135000 222.650000 416.305000 225.360000 ;
      RECT 416.165000 122.555000 416.335000 129.565000 ;
      RECT 416.165000 130.205000 416.335000 137.215000 ;
      RECT 416.165000 137.855000 416.335000 144.645000 ;
      RECT 416.175000  23.110000 416.485000  23.805000 ;
      RECT 416.175000  24.145000 416.345000  24.375000 ;
      RECT 416.180000   8.650000 416.690000   8.680000 ;
      RECT 416.180000  14.760000 416.690000  14.790000 ;
      RECT 416.180000  21.230000 416.350000  22.400000 ;
      RECT 416.250000   8.680000 416.620000  14.760000 ;
      RECT 416.280000 190.240000 416.450000 193.970000 ;
      RECT 416.280000 194.520000 416.450000 198.250000 ;
      RECT 416.295000 226.270000 416.465000 227.580000 ;
      RECT 416.340000 146.300000 417.095000 152.785000 ;
      RECT 416.340000 218.690000 416.715000 220.080000 ;
      RECT 416.400000 244.245000 418.055000 244.730000 ;
      RECT 416.400000 244.730000 419.855000 244.770000 ;
      RECT 416.400000 244.770000 420.665000 245.980000 ;
      RECT 416.400000 245.980000 419.855000 246.265000 ;
      RECT 416.415000  31.925000 417.465000  34.635000 ;
      RECT 416.465000  22.600000 417.815000  22.770000 ;
      RECT 416.545000 122.165000 418.235000 122.335000 ;
      RECT 416.545000 129.815000 418.235000 129.985000 ;
      RECT 416.545000 144.890000 418.235000 145.285000 ;
      RECT 416.565000  22.570000 417.815000  22.600000 ;
      RECT 416.570000  35.185000 417.395000  35.355000 ;
      RECT 416.570000 110.765000 416.740000 120.655000 ;
      RECT 416.610000  21.060000 416.780000  22.400000 ;
      RECT 416.630000 207.340000 416.800000 210.050000 ;
      RECT 416.640000  24.395000 416.810000  27.475000 ;
      RECT 416.715000 220.980000 416.885000 221.650000 ;
      RECT 416.725000 226.570000 417.235000 227.580000 ;
      RECT 416.790000   8.850000 416.960000  14.590000 ;
      RECT 416.805000  28.695000 418.075000  29.025000 ;
      RECT 416.820000 183.610000 416.990000 188.360000 ;
      RECT 416.870000 229.405000 444.570000 229.655000 ;
      RECT 416.880000 190.050000 426.120000 194.160000 ;
      RECT 416.880000 194.330000 426.120000 198.440000 ;
      RECT 416.910000 230.290000 417.080000 233.270000 ;
      RECT 416.915000 218.520000 417.505000 218.690000 ;
      RECT 416.915000 218.690000 417.460000 220.220000 ;
      RECT 416.925000 152.785000 417.095000 155.175000 ;
      RECT 416.965000 246.265000 419.855000 253.125000 ;
      RECT 417.000000 207.540000 417.305000 210.325000 ;
      RECT 417.040000  21.230000 417.210000  22.400000 ;
      RECT 417.060000   8.350000 417.570000   8.680000 ;
      RECT 417.060000  14.760000 417.570000  15.090000 ;
      RECT 417.105000 220.470000 417.775000 220.640000 ;
      RECT 417.130000   8.680000 417.500000  14.760000 ;
      RECT 417.135000 233.550000 420.375000 233.720000 ;
      RECT 417.150000 110.605000 417.330000 120.970000 ;
      RECT 417.180000  40.920000 417.350000  50.770000 ;
      RECT 417.180000  51.380000 417.350000  61.230000 ;
      RECT 417.180000  64.770000 417.350000  74.660000 ;
      RECT 417.180000  75.840000 417.350000  85.730000 ;
      RECT 417.180000  86.965000 417.350000  96.855000 ;
      RECT 417.180000  98.035000 417.350000 107.925000 ;
      RECT 417.225000  34.635000 417.395000  35.185000 ;
      RECT 417.260000  16.520000 420.150000  16.690000 ;
      RECT 417.260000  16.690000 417.430000  19.140000 ;
      RECT 417.260000  19.650000 417.430000  19.790000 ;
      RECT 417.260000  19.790000 417.935000  19.960000 ;
      RECT 417.260000  19.960000 417.430000  20.660000 ;
      RECT 417.285000  25.395000 417.815000  27.655000 ;
      RECT 417.285000  27.655000 420.820000  27.905000 ;
      RECT 417.295000  29.195000 417.465000  30.245000 ;
      RECT 417.295000  30.475000 417.465000  30.805000 ;
      RECT 417.295000  31.425000 417.465000  31.755000 ;
      RECT 417.335000 109.115000 417.925000 109.435000 ;
      RECT 417.380000 222.890000 417.910000 223.900000 ;
      RECT 417.380000 224.570000 417.910000 225.580000 ;
      RECT 417.470000  21.060000 417.640000  22.400000 ;
      RECT 417.500000 109.435000 417.925000 111.380000 ;
      RECT 417.500000 157.395000 417.670000 162.245000 ;
      RECT 417.500000 163.355000 417.670000 168.205000 ;
      RECT 417.500000 169.315000 417.670000 174.165000 ;
      RECT 417.500000 175.275000 417.670000 180.125000 ;
      RECT 417.510000 207.340000 418.830000 210.110000 ;
      RECT 417.560000  63.505000 418.090000  64.380000 ;
      RECT 417.560000  64.380000 419.250000  64.550000 ;
      RECT 417.560000 108.295000 419.250000 108.465000 ;
      RECT 417.565000  35.105000 418.075000  35.435000 ;
      RECT 417.635000  29.025000 418.005000  35.105000 ;
      RECT 417.670000   9.150000 417.840000  11.860000 ;
      RECT 417.670000  12.030000 417.840000  12.560000 ;
      RECT 417.670000  12.980000 417.840000  13.310000 ;
      RECT 417.670000  13.540000 417.840000  14.590000 ;
      RECT 417.705000 146.300000 417.875000 155.175000 ;
      RECT 417.760000  18.225000 418.090000  19.075000 ;
      RECT 417.760000  40.090000 417.940000  62.060000 ;
      RECT 417.785000 224.150000 421.045000 224.320000 ;
      RECT 417.790000 230.115000 417.960000 233.000000 ;
      RECT 417.795000 219.125000 418.325000 220.220000 ;
      RECT 417.805000 162.575000 419.040000 162.905000 ;
      RECT 417.805000 168.535000 419.040000 168.865000 ;
      RECT 417.805000 174.495000 419.040000 174.825000 ;
      RECT 417.805000 180.455000 419.040000 180.785000 ;
      RECT 417.840000  17.615000 418.010000  18.225000 ;
      RECT 417.900000  21.230000 418.070000  22.400000 ;
      RECT 417.900000  75.235000 418.910000  75.405000 ;
      RECT 417.900000  86.330000 418.910000  86.500000 ;
      RECT 417.900000  97.430000 418.910000  97.600000 ;
      RECT 417.940000   8.350000 418.450000   8.680000 ;
      RECT 417.940000  14.760000 418.450000  15.090000 ;
      RECT 417.985000  24.370000 418.155000  27.370000 ;
      RECT 417.995000 220.980000 418.165000 221.870000 ;
      RECT 418.010000   8.680000 418.380000  14.760000 ;
      RECT 418.095000 109.470000 418.885000 109.660000 ;
      RECT 418.095000 109.660000 425.725000 109.840000 ;
      RECT 418.095000 109.840000 418.885000 121.735000 ;
      RECT 418.100000 183.610000 418.270000 188.475000 ;
      RECT 418.170000  22.595000 420.830000  22.765000 ;
      RECT 418.170000  22.765000 419.520000  22.770000 ;
      RECT 418.175000  29.195000 418.345000  34.940000 ;
      RECT 418.195000 146.300000 418.945000 155.305000 ;
      RECT 418.205000  23.710000 418.735000  23.880000 ;
      RECT 418.260000  63.950000 419.670000  64.130000 ;
      RECT 418.270000 235.010000 418.440000 236.090000 ;
      RECT 418.280000 157.045000 419.040000 162.575000 ;
      RECT 418.280000 162.905000 419.040000 168.535000 ;
      RECT 418.280000 168.865000 419.040000 174.495000 ;
      RECT 418.280000 174.825000 419.040000 180.455000 ;
      RECT 418.280000 180.785000 419.040000 180.955000 ;
      RECT 418.330000  20.890000 420.150000  21.060000 ;
      RECT 418.330000  21.060000 418.500000  22.400000 ;
      RECT 418.440000  16.860000 419.310000  17.870000 ;
      RECT 418.440000  18.160000 418.610000  19.310000 ;
      RECT 418.440000  19.480000 418.610000  20.660000 ;
      RECT 418.440000 188.870000 425.560000 189.040000 ;
      RECT 418.445000 122.555000 418.615000 129.565000 ;
      RECT 418.445000 130.205000 418.615000 137.215000 ;
      RECT 418.445000 137.855000 418.615000 144.645000 ;
      RECT 418.450000 234.660000 419.120000 234.830000 ;
      RECT 418.510000 226.570000 419.020000 227.580000 ;
      RECT 418.520000 236.310000 419.050000 236.480000 ;
      RECT 418.550000   8.850000 418.720000  14.590000 ;
      RECT 418.560000 222.890000 419.090000 223.900000 ;
      RECT 418.565000  23.880000 418.735000  27.230000 ;
      RECT 418.565000  27.230000 422.805000  27.400000 ;
      RECT 418.630000 233.720000 418.970000 234.660000 ;
      RECT 418.630000 234.830000 418.970000 236.310000 ;
      RECT 418.670000 122.165000 419.395000 122.335000 ;
      RECT 418.670000 129.815000 419.395000 129.985000 ;
      RECT 418.670000 137.465000 419.395000 137.635000 ;
      RECT 418.670000 145.115000 419.395000 145.285000 ;
      RECT 418.670000 230.290000 418.840000 233.270000 ;
      RECT 418.685000 224.560000 418.965000 225.770000 ;
      RECT 418.685000 225.770000 421.310000 226.020000 ;
      RECT 418.705000  39.145000 418.885000  63.005000 ;
      RECT 418.710000  38.465000 418.880000  38.965000 ;
      RECT 418.725000  29.195000 418.895000  34.940000 ;
      RECT 418.760000  21.230000 418.930000  22.400000 ;
      RECT 418.780000  17.870000 419.310000  18.905000 ;
      RECT 418.820000   8.350000 420.210000   8.650000 ;
      RECT 418.820000   8.650000 419.330000   8.680000 ;
      RECT 418.820000  14.760000 419.330000  14.790000 ;
      RECT 418.820000  14.790000 420.210000  15.090000 ;
      RECT 418.845000 206.950000 419.515000 207.120000 ;
      RECT 418.890000   8.680000 419.260000  14.760000 ;
      RECT 418.995000  28.695000 422.710000  28.995000 ;
      RECT 418.995000  28.995000 420.265000  29.025000 ;
      RECT 418.995000  35.090000 420.265000  35.435000 ;
      RECT 419.065000  29.025000 419.435000  35.090000 ;
      RECT 419.075000 227.830000 420.515000 228.000000 ;
      RECT 419.080000  75.235000 420.010000  75.415000 ;
      RECT 419.080000  86.330000 420.010000  86.510000 ;
      RECT 419.080000  97.430000 420.010000  97.610000 ;
      RECT 419.100000 240.290000 420.680000 243.860000 ;
      RECT 419.150000 235.010000 419.320000 236.090000 ;
      RECT 419.190000  21.060000 419.360000  22.400000 ;
      RECT 419.210000 222.000000 420.110000 222.140000 ;
      RECT 419.210000 222.140000 419.740000 222.170000 ;
      RECT 419.225000 122.335000 419.395000 129.815000 ;
      RECT 419.225000 129.985000 419.395000 137.465000 ;
      RECT 419.225000 137.635000 419.395000 145.115000 ;
      RECT 419.225000 226.020000 419.505000 227.590000 ;
      RECT 419.260000  19.790000 419.790000  19.960000 ;
      RECT 419.260000 218.710000 419.430000 221.420000 ;
      RECT 419.265000 146.300000 419.435000 155.175000 ;
      RECT 419.380000 183.610000 419.550000 188.360000 ;
      RECT 419.430000   9.150000 419.600000  11.860000 ;
      RECT 419.430000  12.030000 419.600000  12.560000 ;
      RECT 419.430000  12.980000 419.600000  13.310000 ;
      RECT 419.430000  13.540000 419.600000  14.590000 ;
      RECT 419.440000 221.970000 420.110000 222.000000 ;
      RECT 419.445000  24.080000 419.705000  27.060000 ;
      RECT 419.460000  64.770000 419.630000  74.660000 ;
      RECT 419.460000  75.840000 419.630000  85.730000 ;
      RECT 419.460000  86.965000 419.630000  96.855000 ;
      RECT 419.460000  98.035000 419.630000 107.925000 ;
      RECT 419.540000 207.340000 419.710000 210.050000 ;
      RECT 419.550000 230.115000 419.720000 233.000000 ;
      RECT 419.605000  29.195000 419.775000  30.245000 ;
      RECT 419.605000  30.475000 419.775000  30.805000 ;
      RECT 419.605000  31.425000 419.775000  31.755000 ;
      RECT 419.605000  31.925000 419.775000  34.635000 ;
      RECT 419.620000  16.690000 420.150000  17.870000 ;
      RECT 419.620000  18.160000 419.790000  19.790000 ;
      RECT 419.620000  19.960000 419.790000  20.660000 ;
      RECT 419.620000  21.230000 419.790000  22.400000 ;
      RECT 419.700000   8.650000 420.210000   8.680000 ;
      RECT 419.700000  14.760000 420.210000  14.790000 ;
      RECT 419.710000 226.570000 419.880000 227.580000 ;
      RECT 419.725000 222.890000 420.255000 223.900000 ;
      RECT 419.725000 224.570000 420.255000 225.580000 ;
      RECT 419.770000   8.680000 420.140000  14.760000 ;
      RECT 419.805000 121.915000 419.985000 145.535000 ;
      RECT 419.805000 145.715000 419.985000 155.920000 ;
      RECT 419.805000 156.100000 419.985000 182.010000 ;
      RECT 419.840000  63.505000 420.370000  64.380000 ;
      RECT 419.840000  64.380000 421.530000  64.550000 ;
      RECT 419.840000 108.295000 421.530000 108.465000 ;
      RECT 419.905000  24.080000 420.165000  27.060000 ;
      RECT 419.945000  29.025000 420.265000  35.090000 ;
      RECT 419.960000  17.870000 420.150000  20.890000 ;
      RECT 419.960000  21.975000 420.490000  22.145000 ;
      RECT 420.080000  23.710000 420.610000  23.880000 ;
      RECT 420.085000 226.020000 420.365000 227.590000 ;
      RECT 420.140000 218.710000 420.310000 221.420000 ;
      RECT 420.180000  75.235000 421.190000  75.405000 ;
      RECT 420.180000  86.330000 421.190000  86.500000 ;
      RECT 420.180000  97.430000 421.190000  97.600000 ;
      RECT 420.260000  22.935000 420.430000  23.710000 ;
      RECT 420.310000   8.850000 420.480000  14.590000 ;
      RECT 420.320000  16.850000 420.490000  21.975000 ;
      RECT 420.430000 230.290000 420.600000 233.270000 ;
      RECT 420.465000  29.165000 420.995000  35.690000 ;
      RECT 420.540000  63.950000 421.680000  64.130000 ;
      RECT 420.570000 226.570000 421.080000 227.580000 ;
      RECT 420.580000   8.350000 421.970000   8.650000 ;
      RECT 420.580000   8.650000 421.090000   8.680000 ;
      RECT 420.580000  14.760000 421.090000  14.790000 ;
      RECT 420.580000  14.790000 421.970000  15.090000 ;
      RECT 420.595000 222.890000 421.450000 223.900000 ;
      RECT 420.630000 250.890000 454.055000 252.495000 ;
      RECT 420.630000 252.495000 465.160000 253.385000 ;
      RECT 420.650000   8.680000 421.020000  14.760000 ;
      RECT 420.660000  20.825000 421.310000  21.835000 ;
      RECT 420.660000  21.835000 420.830000  22.595000 ;
      RECT 420.660000 183.610000 420.830000 188.475000 ;
      RECT 420.750000 111.555000 427.150000 111.735000 ;
      RECT 420.750000 111.735000 420.930000 135.285000 ;
      RECT 420.750000 135.285000 427.150000 135.465000 ;
      RECT 420.750000 135.465000 423.875000 136.040000 ;
      RECT 420.750000 136.040000 420.930000 140.060000 ;
      RECT 420.750000 140.060000 423.875000 140.240000 ;
      RECT 420.750000 237.915000 420.920000 238.965000 ;
      RECT 420.750000 247.190000 420.920000 249.900000 ;
      RECT 420.780000  18.735000 421.310000  18.905000 ;
      RECT 420.780000  23.780000 421.450000  23.950000 ;
      RECT 420.800000  16.605000 426.330000  16.775000 ;
      RECT 420.800000  16.775000 420.970000  17.385000 ;
      RECT 420.815000 236.820000 449.625000 237.070000 ;
      RECT 420.840000  23.040000 421.370000  23.210000 ;
      RECT 420.875000  23.210000 421.370000  23.780000 ;
      RECT 420.875000  23.950000 421.045000  27.060000 ;
      RECT 420.930000 239.235000 421.460000 239.405000 ;
      RECT 420.985000 206.365000 422.855000 211.275000 ;
      RECT 421.020000 237.415000 421.530000 237.745000 ;
      RECT 421.020000 250.370000 421.530000 250.700000 ;
      RECT 421.030000  27.735000 421.700000  27.905000 ;
      RECT 421.045000 224.560000 421.310000 225.770000 ;
      RECT 421.065000  40.200000 423.165000  40.370000 ;
      RECT 421.065000  40.370000 421.235000  42.450000 ;
      RECT 421.065000  42.450000 421.815000  42.780000 ;
      RECT 421.065000  43.200000 421.815000  43.730000 ;
      RECT 421.065000  43.730000 421.235000  47.580000 ;
      RECT 421.065000  47.580000 445.335000  47.750000 ;
      RECT 421.090000 237.745000 421.460000 239.235000 ;
      RECT 421.090000 239.405000 421.460000 250.370000 ;
      RECT 421.140000  17.155000 421.310000  18.735000 ;
      RECT 421.140000  18.905000 421.310000  20.825000 ;
      RECT 421.180000 181.095000 423.525000 181.840000 ;
      RECT 421.190000   9.150000 421.360000  11.860000 ;
      RECT 421.190000  12.030000 421.360000  12.360000 ;
      RECT 421.190000  12.980000 421.360000  13.310000 ;
      RECT 421.190000  13.540000 421.360000  14.590000 ;
      RECT 421.265000  29.165000 421.815000  36.060000 ;
      RECT 421.310000 140.415000 441.730000 140.585000 ;
      RECT 421.310000 140.585000 421.480000 180.755000 ;
      RECT 421.310000 180.755000 430.390000 180.925000 ;
      RECT 421.335000 112.145000 421.665000 112.655000 ;
      RECT 421.335000 134.365000 421.665000 134.875000 ;
      RECT 421.340000 230.620000 421.510000 233.330000 ;
      RECT 421.340000 235.010000 421.510000 236.060000 ;
      RECT 421.355000 136.720000 421.525000 139.430000 ;
      RECT 421.360000  75.235000 422.290000  75.415000 ;
      RECT 421.360000  86.330000 422.290000  86.510000 ;
      RECT 421.360000  97.430000 422.290000  97.610000 ;
      RECT 421.415000 112.135000 421.585000 112.145000 ;
      RECT 421.415000 112.655000 421.585000 112.665000 ;
      RECT 421.415000 134.355000 421.585000 134.365000 ;
      RECT 421.415000 134.875000 421.585000 134.885000 ;
      RECT 421.460000   8.650000 421.970000   8.680000 ;
      RECT 421.460000  14.760000 421.970000  14.790000 ;
      RECT 421.480000  20.070000 422.010000  20.240000 ;
      RECT 421.520000 234.570000 422.050000 234.740000 ;
      RECT 421.530000   8.680000 421.900000  14.760000 ;
      RECT 421.530000 229.900000 422.200000 230.070000 ;
      RECT 421.540000  22.935000 421.790000  23.605000 ;
      RECT 421.575000  20.825000 421.770000  21.835000 ;
      RECT 421.575000  21.835000 421.745000  22.935000 ;
      RECT 421.575000  23.605000 421.790000  23.660000 ;
      RECT 421.600000  17.155000 421.770000  20.070000 ;
      RECT 421.610000 236.230000 422.120000 236.560000 ;
      RECT 421.620000  23.660000 421.790000  24.350000 ;
      RECT 421.620000  24.350000 421.925000  27.060000 ;
      RECT 421.630000 237.915000 421.800000 239.240000 ;
      RECT 421.630000 239.240000 422.960000 239.750000 ;
      RECT 421.630000 239.750000 421.800000 250.205000 ;
      RECT 421.645000  41.170000 421.815000  42.220000 ;
      RECT 421.645000  43.900000 421.815000  46.610000 ;
      RECT 421.645000 139.650000 422.995000 139.830000 ;
      RECT 421.680000 230.070000 422.050000 234.570000 ;
      RECT 421.680000 234.740000 422.050000 236.230000 ;
      RECT 421.740000  64.770000 421.910000  74.660000 ;
      RECT 421.740000  75.840000 421.910000  85.730000 ;
      RECT 421.740000  86.965000 421.910000  96.855000 ;
      RECT 421.740000  98.035000 421.910000 107.925000 ;
      RECT 421.850000  63.505000 422.380000  64.380000 ;
      RECT 421.850000  64.380000 423.810000  64.550000 ;
      RECT 421.890000 218.340000 422.060000 228.475000 ;
      RECT 421.915000  40.670000 422.425000  41.000000 ;
      RECT 421.915000  47.080000 422.425000  47.410000 ;
      RECT 421.940000  17.155000 422.230000  19.575000 ;
      RECT 421.940000  19.575000 422.480000  19.865000 ;
      RECT 421.940000  20.500000 422.480000  20.655000 ;
      RECT 421.940000  20.655000 422.350000  22.670000 ;
      RECT 421.940000  22.670000 422.470000  22.840000 ;
      RECT 421.940000 183.610000 422.110000 188.360000 ;
      RECT 421.960000  23.040000 422.990000  23.210000 ;
      RECT 421.980000  27.735000 422.650000  27.905000 ;
      RECT 421.985000  29.165000 422.995000  30.175000 ;
      RECT 421.985000  30.175000 422.515000  35.690000 ;
      RECT 421.985000  41.000000 422.355000  47.080000 ;
      RECT 422.035000 112.145000 422.365000 113.105000 ;
      RECT 422.035000 129.990000 422.365000 130.580000 ;
      RECT 422.040000 141.155000 422.370000 141.805000 ;
      RECT 422.040000 160.345000 422.370000 160.995000 ;
      RECT 422.040000 179.535000 422.370000 180.185000 ;
      RECT 422.060000  23.780000 422.805000  23.950000 ;
      RECT 422.070000   8.850000 422.240000  14.590000 ;
      RECT 422.120000 108.295000 423.810000 108.465000 ;
      RECT 422.130000  23.710000 422.660000  23.780000 ;
      RECT 422.180000  19.865000 422.480000  20.500000 ;
      RECT 422.220000 230.315000 422.390000 234.225000 ;
      RECT 422.220000 234.225000 423.550000 234.735000 ;
      RECT 422.220000 234.735000 422.390000 236.060000 ;
      RECT 422.235000 136.720000 422.405000 139.430000 ;
      RECT 422.250000 237.915000 422.420000 238.965000 ;
      RECT 422.250000 247.190000 422.420000 249.900000 ;
      RECT 422.335000   8.350000 423.730000   8.650000 ;
      RECT 422.335000   8.650000 422.845000   8.680000 ;
      RECT 422.340000  14.760000 422.850000  14.790000 ;
      RECT 422.340000  14.790000 423.730000  15.090000 ;
      RECT 422.410000   8.680000 422.780000  14.760000 ;
      RECT 422.430000  16.965000 423.185000  17.135000 ;
      RECT 422.460000  75.235000 423.470000  75.405000 ;
      RECT 422.460000  86.330000 423.470000  86.500000 ;
      RECT 422.460000  97.430000 423.470000  97.600000 ;
      RECT 422.500000 222.890000 423.355000 223.900000 ;
      RECT 422.520000  20.825000 422.690000  21.835000 ;
      RECT 422.520000 237.415000 423.030000 237.745000 ;
      RECT 422.520000 250.370000 423.030000 250.700000 ;
      RECT 422.525000  41.170000 422.695000  46.915000 ;
      RECT 422.550000  63.950000 424.780000  64.130000 ;
      RECT 422.590000 237.745000 422.960000 239.240000 ;
      RECT 422.590000 239.750000 422.960000 250.370000 ;
      RECT 422.635000  23.950000 422.805000  27.230000 ;
      RECT 422.640000 224.560000 422.905000 225.770000 ;
      RECT 422.640000 225.770000 425.265000 226.020000 ;
      RECT 422.655000  18.735000 423.185000  18.905000 ;
      RECT 422.675000  19.940000 422.845000  20.610000 ;
      RECT 422.685000  30.850000 422.855000  31.755000 ;
      RECT 422.685000  31.925000 423.685000  36.060000 ;
      RECT 422.715000  22.155000 423.250000  22.730000 ;
      RECT 422.735000 112.145000 423.065000 113.105000 ;
      RECT 422.735000 129.990000 423.065000 130.580000 ;
      RECT 422.820000  22.935000 422.990000  23.040000 ;
      RECT 422.820000  23.210000 422.990000  23.605000 ;
      RECT 422.840000 230.620000 423.010000 233.330000 ;
      RECT 422.840000 235.010000 423.010000 236.060000 ;
      RECT 422.850000 141.155000 423.180000 141.805000 ;
      RECT 422.850000 160.345000 423.180000 160.995000 ;
      RECT 422.850000 179.535000 423.180000 180.185000 ;
      RECT 422.870000 226.570000 423.380000 227.580000 ;
      RECT 422.905000 224.150000 426.165000 224.320000 ;
      RECT 422.950000   9.150000 423.120000  11.860000 ;
      RECT 422.950000  12.030000 423.120000  12.560000 ;
      RECT 422.950000  12.980000 423.120000  13.310000 ;
      RECT 422.950000  13.540000 423.120000  14.590000 ;
      RECT 422.980000  20.825000 423.185000  21.835000 ;
      RECT 423.015000  17.135000 423.185000  18.735000 ;
      RECT 423.015000  18.905000 423.185000  20.825000 ;
      RECT 423.030000 229.900000 423.700000 230.070000 ;
      RECT 423.075000  41.170000 423.245000  42.990000 ;
      RECT 423.075000  43.900000 423.245000  46.610000 ;
      RECT 423.100000  30.430000 423.270000  30.805000 ;
      RECT 423.110000 236.230000 423.620000 236.560000 ;
      RECT 423.115000 136.720000 423.285000 139.430000 ;
      RECT 423.130000 237.915000 423.300000 239.240000 ;
      RECT 423.130000 239.240000 424.460000 239.750000 ;
      RECT 423.130000 239.750000 423.300000 250.205000 ;
      RECT 423.180000 230.070000 423.550000 234.225000 ;
      RECT 423.180000 234.735000 423.550000 236.230000 ;
      RECT 423.220000   8.650000 423.730000   8.680000 ;
      RECT 423.220000  14.760000 423.730000  14.790000 ;
      RECT 423.220000 183.610000 423.390000 188.475000 ;
      RECT 423.290000   8.680000 423.660000  14.760000 ;
      RECT 423.335000  39.345000 423.865000  41.000000 ;
      RECT 423.345000  47.080000 423.855000  47.410000 ;
      RECT 423.375000  29.165000 424.385000  30.175000 ;
      RECT 423.415000  41.000000 423.785000  47.080000 ;
      RECT 423.435000 112.145000 423.765000 113.105000 ;
      RECT 423.435000 133.915000 423.765000 134.875000 ;
      RECT 423.435000 227.830000 424.875000 228.000000 ;
      RECT 423.480000  16.775000 423.650000  17.385000 ;
      RECT 423.480000  20.815000 423.650000  23.870000 ;
      RECT 423.515000  30.850000 423.685000  31.755000 ;
      RECT 423.585000 226.020000 423.865000 227.590000 ;
      RECT 423.640000  75.235000 424.780000  75.415000 ;
      RECT 423.640000  86.330000 424.780000  86.510000 ;
      RECT 423.640000  97.430000 424.780000  97.610000 ;
      RECT 423.640000 218.710000 423.810000 221.420000 ;
      RECT 423.660000  28.695000 427.375000  28.995000 ;
      RECT 423.660000 141.155000 423.990000 141.805000 ;
      RECT 423.660000 160.345000 423.990000 160.995000 ;
      RECT 423.660000 179.535000 423.990000 180.185000 ;
      RECT 423.695000 136.040000 423.875000 140.060000 ;
      RECT 423.695000 222.890000 424.225000 223.900000 ;
      RECT 423.695000 224.570000 424.225000 225.580000 ;
      RECT 423.720000 230.315000 423.890000 234.225000 ;
      RECT 423.720000 234.225000 425.050000 234.735000 ;
      RECT 423.720000 234.735000 423.890000 236.060000 ;
      RECT 423.750000 237.915000 423.920000 238.980000 ;
      RECT 423.750000 247.190000 423.920000 249.900000 ;
      RECT 423.830000   8.850000 424.000000  14.590000 ;
      RECT 423.840000 221.970000 424.510000 222.000000 ;
      RECT 423.840000 222.000000 424.740000 222.140000 ;
      RECT 423.855000  30.175000 424.385000  35.690000 ;
      RECT 423.880000  22.155000 424.415000  22.730000 ;
      RECT 423.945000  16.965000 424.700000  17.135000 ;
      RECT 423.945000  17.135000 424.115000  18.735000 ;
      RECT 423.945000  18.735000 424.475000  18.905000 ;
      RECT 423.945000  18.905000 424.115000  20.825000 ;
      RECT 423.945000  20.825000 424.150000  21.835000 ;
      RECT 423.955000  41.295000 424.125000  46.915000 ;
      RECT 424.020000  64.770000 424.190000  74.660000 ;
      RECT 424.020000  75.840000 424.190000  85.730000 ;
      RECT 424.020000  86.965000 424.190000  96.855000 ;
      RECT 424.020000  98.035000 424.190000 107.925000 ;
      RECT 424.020000 237.415000 424.530000 237.745000 ;
      RECT 424.020000 250.370000 424.530000 250.700000 ;
      RECT 424.035000  40.200000 424.925000  40.370000 ;
      RECT 424.070000 226.570000 424.240000 227.580000 ;
      RECT 424.090000 237.745000 424.460000 239.240000 ;
      RECT 424.090000 239.750000 424.460000 250.370000 ;
      RECT 424.100000   8.350000 424.610000   8.680000 ;
      RECT 424.100000  14.760000 424.610000  15.090000 ;
      RECT 424.135000 112.145000 424.465000 113.105000 ;
      RECT 424.135000 133.915000 424.465000 134.875000 ;
      RECT 424.140000  22.935000 424.310000  23.040000 ;
      RECT 424.140000  23.040000 425.170000  23.210000 ;
      RECT 424.140000  23.210000 424.310000  23.605000 ;
      RECT 424.170000   8.680000 424.540000  14.760000 ;
      RECT 424.210000 222.140000 424.740000 222.170000 ;
      RECT 424.225000  40.670000 425.625000  41.000000 ;
      RECT 424.225000  47.080000 424.735000  47.410000 ;
      RECT 424.240000 207.340000 424.410000 210.050000 ;
      RECT 424.285000  19.940000 424.455000  20.610000 ;
      RECT 424.295000  41.000000 424.665000  47.080000 ;
      RECT 424.325000  23.780000 425.070000  23.950000 ;
      RECT 424.325000  23.950000 424.495000  27.230000 ;
      RECT 424.325000  27.230000 428.565000  27.400000 ;
      RECT 424.340000 230.620000 424.510000 233.330000 ;
      RECT 424.340000 234.995000 424.510000 236.060000 ;
      RECT 424.435000 206.950000 425.105000 207.120000 ;
      RECT 424.440000  20.825000 424.610000  21.835000 ;
      RECT 424.445000 226.020000 424.725000 227.590000 ;
      RECT 424.470000  23.710000 425.000000  23.780000 ;
      RECT 424.470000 141.155000 424.800000 141.805000 ;
      RECT 424.470000 160.345000 424.800000 160.995000 ;
      RECT 424.470000 179.535000 424.800000 180.185000 ;
      RECT 424.480000  27.735000 425.150000  27.905000 ;
      RECT 424.500000 183.610000 424.670000 188.360000 ;
      RECT 424.520000 218.710000 424.690000 221.420000 ;
      RECT 424.530000 229.900000 425.200000 230.070000 ;
      RECT 424.555000  29.165000 425.105000  36.060000 ;
      RECT 424.600000  64.130000 424.780000  75.235000 ;
      RECT 424.600000  75.415000 424.780000  86.330000 ;
      RECT 424.600000  86.510000 424.780000  97.430000 ;
      RECT 424.600000  97.610000 424.780000 108.715000 ;
      RECT 424.610000 236.230000 425.120000 236.560000 ;
      RECT 424.630000 238.040000 424.800000 250.205000 ;
      RECT 424.650000  19.575000 425.190000  19.865000 ;
      RECT 424.650000  19.865000 424.950000  20.500000 ;
      RECT 424.650000  20.500000 425.190000  20.655000 ;
      RECT 424.660000  22.670000 425.190000  22.840000 ;
      RECT 424.680000 230.070000 425.050000 234.225000 ;
      RECT 424.680000 234.735000 425.050000 236.230000 ;
      RECT 424.710000   9.150000 424.880000  11.860000 ;
      RECT 424.710000  12.030000 424.880000  12.560000 ;
      RECT 424.710000  12.780000 424.880000  13.310000 ;
      RECT 424.710000  13.540000 424.880000  14.590000 ;
      RECT 424.750000 138.345000 424.920000 139.355000 ;
      RECT 424.780000  20.655000 425.190000  22.670000 ;
      RECT 424.805000 137.925000 425.475000 138.095000 ;
      RECT 424.835000  41.170000 425.005000  42.235000 ;
      RECT 424.835000  42.405000 425.005000  42.780000 ;
      RECT 424.835000  43.200000 425.005000  43.730000 ;
      RECT 424.835000  43.900000 425.005000  46.610000 ;
      RECT 424.835000 112.145000 425.165000 113.105000 ;
      RECT 424.835000 133.915000 425.165000 134.875000 ;
      RECT 424.860000 222.890000 425.390000 223.900000 ;
      RECT 424.895000 237.495000 425.425000 237.665000 ;
      RECT 424.900000  17.155000 425.190000  19.575000 ;
      RECT 424.900000 237.415000 425.410000 237.495000 ;
      RECT 424.900000 237.665000 425.410000 237.745000 ;
      RECT 424.900000 250.370000 425.410000 250.700000 ;
      RECT 424.930000 226.570000 425.440000 227.580000 ;
      RECT 424.970000 237.745000 425.340000 250.370000 ;
      RECT 424.985000 224.560000 425.265000 225.770000 ;
      RECT 425.095000  36.975000 425.625000  40.670000 ;
      RECT 425.105000  47.080000 425.615000  47.410000 ;
      RECT 425.120000  20.070000 425.650000  20.240000 ;
      RECT 425.120000 207.340000 426.440000 210.110000 ;
      RECT 425.175000  41.000000 425.545000  47.080000 ;
      RECT 425.205000  24.350000 425.510000  27.060000 ;
      RECT 425.220000 230.300000 425.390000 235.935000 ;
      RECT 425.280000 141.155000 425.610000 141.805000 ;
      RECT 425.280000 160.345000 425.610000 160.995000 ;
      RECT 425.280000 179.535000 425.610000 180.185000 ;
      RECT 425.340000  22.935000 425.590000  23.605000 ;
      RECT 425.340000  23.605000 425.555000  23.660000 ;
      RECT 425.340000  23.660000 425.510000  24.350000 ;
      RECT 425.360000  17.155000 425.530000  20.070000 ;
      RECT 425.360000  20.825000 425.555000  21.835000 ;
      RECT 425.375000  29.165000 425.905000  35.690000 ;
      RECT 425.385000  21.835000 425.555000  22.935000 ;
      RECT 425.405000   8.180000 425.575000  12.560000 ;
      RECT 425.405000  13.080000 426.340000  14.600000 ;
      RECT 425.405000  14.600000 430.360000  15.685000 ;
      RECT 425.410000 229.900000 426.080000 230.070000 ;
      RECT 425.430000  27.735000 426.100000  27.905000 ;
      RECT 425.485000 236.310000 426.015000 236.480000 ;
      RECT 425.490000 236.230000 426.000000 236.310000 ;
      RECT 425.490000 236.480000 426.000000 236.560000 ;
      RECT 425.510000 237.915000 425.680000 239.240000 ;
      RECT 425.510000 239.240000 426.840000 239.750000 ;
      RECT 425.510000 247.190000 425.680000 249.900000 ;
      RECT 425.530000 138.345000 425.700000 139.355000 ;
      RECT 425.535000 112.145000 425.865000 113.105000 ;
      RECT 425.535000 134.365000 425.865000 134.875000 ;
      RECT 425.545000  48.420000 445.335000  48.600000 ;
      RECT 425.545000  48.600000 425.725000  63.005000 ;
      RECT 425.545000  63.185000 425.725000 109.660000 ;
      RECT 425.555000 133.915000 425.865000 134.365000 ;
      RECT 425.560000 230.070000 425.930000 236.230000 ;
      RECT 425.625000 219.125000 426.155000 220.220000 ;
      RECT 425.680000  23.780000 426.350000  23.950000 ;
      RECT 425.715000  41.295000 425.885000  46.915000 ;
      RECT 425.760000  23.040000 426.290000  23.210000 ;
      RECT 425.760000  23.210000 426.255000  23.780000 ;
      RECT 425.780000 183.610000 425.950000 188.475000 ;
      RECT 425.785000 220.980000 425.955000 221.870000 ;
      RECT 425.820000  17.155000 425.990000  18.735000 ;
      RECT 425.820000  18.735000 426.350000  18.905000 ;
      RECT 425.820000  18.905000 425.990000  20.825000 ;
      RECT 425.820000  20.825000 426.470000  21.835000 ;
      RECT 425.975000  38.175000 426.505000  41.000000 ;
      RECT 425.985000  47.080000 426.495000  47.410000 ;
      RECT 426.005000 188.870000 427.100000 189.040000 ;
      RECT 426.040000 222.890000 426.570000 223.900000 ;
      RECT 426.040000 224.570000 426.570000 225.580000 ;
      RECT 426.055000  41.000000 426.425000  47.080000 ;
      RECT 426.085000  23.950000 426.255000  27.060000 ;
      RECT 426.090000 141.155000 426.420000 141.805000 ;
      RECT 426.090000 160.345000 426.420000 160.995000 ;
      RECT 426.090000 179.535000 426.420000 180.185000 ;
      RECT 426.100000 230.620000 426.270000 233.330000 ;
      RECT 426.100000 234.570000 426.270000 236.060000 ;
      RECT 426.105000  28.995000 427.375000  29.025000 ;
      RECT 426.105000  29.025000 426.425000  35.105000 ;
      RECT 426.105000  35.105000 427.375000  35.435000 ;
      RECT 426.130000 237.915000 426.300000 238.965000 ;
      RECT 426.130000 247.190000 426.300000 249.900000 ;
      RECT 426.160000  16.775000 426.330000  17.385000 ;
      RECT 426.175000 220.470000 426.845000 220.640000 ;
      RECT 426.235000 112.145000 426.565000 113.105000 ;
      RECT 426.235000 133.910000 426.565000 134.875000 ;
      RECT 426.300000  21.835000 426.470000  22.595000 ;
      RECT 426.300000  22.595000 428.960000  22.765000 ;
      RECT 426.310000  27.655000 429.845000  27.905000 ;
      RECT 426.400000 237.415000 426.910000 237.745000 ;
      RECT 426.400000 250.370000 426.910000 250.700000 ;
      RECT 426.445000 218.520000 427.035000 218.690000 ;
      RECT 426.470000 210.325000 428.670000 210.995000 ;
      RECT 426.470000 237.745000 426.840000 239.240000 ;
      RECT 426.470000 239.750000 426.840000 250.370000 ;
      RECT 426.490000 218.690000 427.035000 220.220000 ;
      RECT 426.520000  23.710000 427.050000  23.880000 ;
      RECT 426.560000 183.610000 426.730000 188.475000 ;
      RECT 426.595000  29.195000 426.765000  30.245000 ;
      RECT 426.595000  30.475000 426.765000  30.805000 ;
      RECT 426.595000  31.425000 426.765000  31.755000 ;
      RECT 426.595000  31.925000 426.765000  34.635000 ;
      RECT 426.595000  41.170000 426.765000  42.990000 ;
      RECT 426.595000  43.900000 426.765000  46.610000 ;
      RECT 426.640000  16.850000 426.810000  21.975000 ;
      RECT 426.640000  21.975000 427.170000  22.145000 ;
      RECT 426.645000 207.540000 426.950000 210.325000 ;
      RECT 426.690000  40.200000 427.220000  40.370000 ;
      RECT 426.700000  22.935000 426.870000  23.710000 ;
      RECT 426.715000 226.570000 427.225000 227.580000 ;
      RECT 426.720000 230.620000 426.890000 233.330000 ;
      RECT 426.720000 234.995000 426.890000 236.060000 ;
      RECT 426.725000 190.240000 427.050000 193.970000 ;
      RECT 426.725000 194.520000 427.050000 198.250000 ;
      RECT 426.900000 141.155000 427.230000 141.805000 ;
      RECT 426.900000 160.345000 427.230000 160.995000 ;
      RECT 426.900000 179.535000 427.230000 180.185000 ;
      RECT 426.900000 234.010000 427.430000 234.180000 ;
      RECT 426.910000 229.900000 427.580000 230.070000 ;
      RECT 426.930000 188.110000 427.100000 188.870000 ;
      RECT 426.935000  29.025000 427.305000  35.105000 ;
      RECT 426.955000 137.765000 433.185000 137.945000 ;
      RECT 426.955000 137.945000 427.135000 139.995000 ;
      RECT 426.955000 139.995000 433.185000 140.175000 ;
      RECT 426.965000  24.080000 427.225000  27.060000 ;
      RECT 426.970000   8.420000 438.355000   8.930000 ;
      RECT 426.970000   8.930000 427.500000  12.090000 ;
      RECT 426.970000  12.090000 428.380000  13.125000 ;
      RECT 426.970000  13.125000 429.100000  13.540000 ;
      RECT 426.970000  13.540000 430.360000  14.600000 ;
      RECT 426.970000 111.735000 427.150000 135.285000 ;
      RECT 426.980000  16.520000 429.870000  16.690000 ;
      RECT 426.980000  16.690000 427.510000  17.870000 ;
      RECT 426.980000  17.870000 427.170000  20.890000 ;
      RECT 426.980000  20.890000 428.800000  21.060000 ;
      RECT 426.990000 236.230000 427.500000 236.560000 ;
      RECT 427.010000 237.915000 427.180000 250.220000 ;
      RECT 427.060000 230.070000 427.430000 234.010000 ;
      RECT 427.060000 234.180000 427.430000 236.230000 ;
      RECT 427.065000 220.980000 427.235000 221.650000 ;
      RECT 427.145000  41.170000 427.315000  42.990000 ;
      RECT 427.145000  43.900000 427.315000  46.610000 ;
      RECT 427.150000 207.340000 427.320000 210.050000 ;
      RECT 427.235000 218.520000 427.825000 218.690000 ;
      RECT 427.235000 218.690000 427.610000 220.080000 ;
      RECT 427.235000 220.080000 427.845000 220.580000 ;
      RECT 427.235000 220.580000 428.210000 220.790000 ;
      RECT 427.280000 227.830000 428.720000 228.000000 ;
      RECT 427.290000 183.135000 427.470000 189.290000 ;
      RECT 427.290000 189.470000 427.470000 199.020000 ;
      RECT 427.325000 138.635000 427.830000 139.305000 ;
      RECT 427.340000  18.160000 427.510000  19.790000 ;
      RECT 427.340000  19.790000 427.870000  19.960000 ;
      RECT 427.340000  19.960000 427.510000  20.660000 ;
      RECT 427.340000  21.230000 427.510000  22.400000 ;
      RECT 427.405000  39.375000 427.935000  41.000000 ;
      RECT 427.415000  47.080000 427.925000  47.410000 ;
      RECT 427.425000  24.080000 427.685000  27.060000 ;
      RECT 427.475000  29.195000 427.645000  34.940000 ;
      RECT 427.485000  41.000000 427.855000  47.080000 ;
      RECT 427.485000 226.270000 427.655000 227.580000 ;
      RECT 427.490000 220.790000 428.210000 221.650000 ;
      RECT 427.600000 230.315000 427.770000 235.935000 ;
      RECT 427.610000  22.765000 428.960000  22.770000 ;
      RECT 427.630000 237.915000 427.800000 238.980000 ;
      RECT 427.630000 247.190000 427.800000 249.900000 ;
      RECT 427.645000 222.650000 427.815000 225.360000 ;
      RECT 427.710000 141.155000 428.040000 141.805000 ;
      RECT 427.710000 160.345000 428.040000 160.995000 ;
      RECT 427.710000 179.535000 428.040000 180.185000 ;
      RECT 427.770000  21.060000 427.940000  22.400000 ;
      RECT 427.790000 229.900000 428.460000 230.070000 ;
      RECT 427.810000 219.185000 428.340000 219.880000 ;
      RECT 427.810000 239.795000 428.340000 239.965000 ;
      RECT 427.820000  16.860000 428.690000  17.870000 ;
      RECT 427.820000  17.870000 428.350000  18.905000 ;
      RECT 427.870000 225.910000 430.010000 226.080000 ;
      RECT 427.870000 236.230000 428.380000 236.560000 ;
      RECT 427.900000 237.415000 428.410000 237.745000 ;
      RECT 427.900000 250.370000 428.410000 250.700000 ;
      RECT 427.915000 226.570000 428.085000 227.600000 ;
      RECT 427.940000 230.070000 428.310000 236.230000 ;
      RECT 427.970000 237.745000 428.340000 239.795000 ;
      RECT 427.970000 239.965000 428.340000 250.370000 ;
      RECT 428.000000 207.440000 428.670000 207.610000 ;
      RECT 428.000000 208.220000 428.730000 209.540000 ;
      RECT 428.000000 210.150000 428.670000 210.325000 ;
      RECT 428.005000 138.355000 433.185000 138.525000 ;
      RECT 428.005000 138.885000 432.755000 139.055000 ;
      RECT 428.005000 139.415000 433.185000 139.585000 ;
      RECT 428.025000  29.195000 428.195000  34.940000 ;
      RECT 428.025000  41.295000 428.195000  46.915000 ;
      RECT 428.035000 220.220000 429.035000 220.390000 ;
      RECT 428.090000   9.490000 436.730000   9.710000 ;
      RECT 428.135000  40.200000 429.025000  40.370000 ;
      RECT 428.165000 222.630000 428.695000 222.800000 ;
      RECT 428.200000  21.230000 428.370000  22.400000 ;
      RECT 428.210000   9.960000 428.380000  11.015000 ;
      RECT 428.235000 182.190000 428.475000 182.415000 ;
      RECT 428.235000 182.415000 428.480000 188.345000 ;
      RECT 428.235000 188.345000 428.415000 199.940000 ;
      RECT 428.255000   9.180000 436.705000   9.490000 ;
      RECT 428.295000  28.695000 432.010000  28.995000 ;
      RECT 428.295000  28.995000 429.565000  29.025000 ;
      RECT 428.295000  35.105000 429.565000  35.435000 ;
      RECT 428.295000  40.670000 428.805000  41.000000 ;
      RECT 428.295000  47.080000 428.805000  47.410000 ;
      RECT 428.345000 226.270000 428.515000 227.580000 ;
      RECT 428.365000  29.025000 428.735000  35.090000 ;
      RECT 428.365000  35.090000 429.565000  35.105000 ;
      RECT 428.365000  41.000000 428.735000  47.080000 ;
      RECT 428.395000  23.710000 428.925000  23.880000 ;
      RECT 428.395000  23.880000 428.565000  27.230000 ;
      RECT 428.480000 230.620000 428.650000 233.330000 ;
      RECT 428.480000 234.225000 429.810000 234.735000 ;
      RECT 428.480000 234.735000 428.650000 236.060000 ;
      RECT 428.510000 238.040000 428.680000 250.205000 ;
      RECT 428.520000  18.160000 428.690000  19.310000 ;
      RECT 428.520000  19.310000 431.050000  19.480000 ;
      RECT 428.520000  19.480000 428.690000  20.660000 ;
      RECT 428.520000 141.155000 428.850000 141.805000 ;
      RECT 428.520000 160.345000 428.850000 160.995000 ;
      RECT 428.520000 179.535000 428.850000 180.185000 ;
      RECT 428.525000 222.800000 428.695000 225.360000 ;
      RECT 428.580000 207.855000 429.180000 208.025000 ;
      RECT 428.630000  21.060000 428.800000  22.400000 ;
      RECT 428.775000 226.570000 429.285000 227.580000 ;
      RECT 428.780000 237.415000 429.290000 237.745000 ;
      RECT 428.780000 250.370000 429.290000 250.700000 ;
      RECT 428.850000 237.745000 429.220000 250.370000 ;
      RECT 428.905000  29.195000 429.075000  30.245000 ;
      RECT 428.905000  30.475000 429.075000  30.805000 ;
      RECT 428.905000  31.425000 429.075000  31.755000 ;
      RECT 428.905000  31.925000 429.075000  34.635000 ;
      RECT 428.905000  41.170000 429.075000  42.235000 ;
      RECT 428.905000  42.405000 429.075000  42.780000 ;
      RECT 428.905000  43.200000 429.075000  43.730000 ;
      RECT 428.905000  43.900000 429.075000  46.610000 ;
      RECT 428.920000 220.640000 429.090000 221.650000 ;
      RECT 428.975000  24.370000 429.145000  27.370000 ;
      RECT 429.005000 219.210000 430.465000 219.880000 ;
      RECT 429.010000 207.585000 429.180000 207.855000 ;
      RECT 429.010000 208.025000 429.180000 208.255000 ;
      RECT 429.010000 209.515000 429.180000 209.680000 ;
      RECT 429.010000 209.680000 430.030000 209.850000 ;
      RECT 429.010000 209.850000 429.180000 210.185000 ;
      RECT 429.040000  18.225000 429.370000  19.075000 ;
      RECT 429.060000  21.230000 429.230000  22.400000 ;
      RECT 429.100000 230.620000 429.270000 233.330000 ;
      RECT 429.100000 235.010000 429.270000 236.060000 ;
      RECT 429.120000  17.615000 429.290000  18.225000 ;
      RECT 429.155000 135.640000 437.515000 135.670000 ;
      RECT 429.155000 135.670000 444.415000 135.840000 ;
      RECT 429.155000 135.840000 437.515000 135.870000 ;
      RECT 429.185000  49.370000 442.555000  49.540000 ;
      RECT 429.185000  49.540000 429.355000 135.640000 ;
      RECT 429.185000 222.650000 429.355000 225.360000 ;
      RECT 429.195000  19.790000 429.870000  19.960000 ;
      RECT 429.235000  38.575000 429.765000  41.000000 ;
      RECT 429.245000  29.025000 429.565000  35.090000 ;
      RECT 429.245000  47.080000 429.755000  47.410000 ;
      RECT 429.290000 229.900000 429.960000 230.070000 ;
      RECT 429.315000  22.570000 430.565000  22.600000 ;
      RECT 429.315000  22.600000 430.665000  22.770000 ;
      RECT 429.315000  25.395000 429.845000  27.655000 ;
      RECT 429.315000  41.000000 429.685000  47.080000 ;
      RECT 429.330000 141.155000 429.660000 141.805000 ;
      RECT 429.330000 160.345000 429.660000 160.995000 ;
      RECT 429.330000 179.535000 429.660000 180.185000 ;
      RECT 429.370000 236.230000 429.880000 236.560000 ;
      RECT 429.380000 207.410000 430.030000 209.680000 ;
      RECT 429.390000 237.915000 429.560000 239.240000 ;
      RECT 429.390000 239.240000 430.720000 239.750000 ;
      RECT 429.390000 247.190000 429.560000 249.900000 ;
      RECT 429.440000 230.070000 429.810000 234.225000 ;
      RECT 429.440000 234.735000 429.810000 236.230000 ;
      RECT 429.490000   9.960000 429.660000  13.100000 ;
      RECT 429.490000  20.890000 431.050000  21.060000 ;
      RECT 429.490000  21.060000 429.660000  22.400000 ;
      RECT 429.595000  49.850000 430.125000  50.020000 ;
      RECT 429.700000  16.690000 429.870000  19.140000 ;
      RECT 429.700000  19.650000 429.870000  19.790000 ;
      RECT 429.700000  19.960000 429.870000  20.660000 ;
      RECT 429.710000  56.485000 430.040000  57.175000 ;
      RECT 429.710000  63.640000 430.040000  64.330000 ;
      RECT 429.710000  70.795000 430.040000  71.485000 ;
      RECT 429.710000  77.950000 430.040000  78.640000 ;
      RECT 429.710000  85.105000 430.040000  85.795000 ;
      RECT 429.710000  92.260000 430.040000  92.950000 ;
      RECT 429.710000  99.415000 430.040000 100.105000 ;
      RECT 429.710000 106.570000 430.040000 107.260000 ;
      RECT 429.710000 113.725000 430.040000 114.415000 ;
      RECT 429.710000 120.880000 430.040000 121.570000 ;
      RECT 429.710000 128.035000 430.040000 128.725000 ;
      RECT 429.710000 135.190000 430.810000 135.360000 ;
      RECT 429.765000  29.165000 430.295000  34.635000 ;
      RECT 429.830000  11.450000 431.860000  11.620000 ;
      RECT 429.830000  13.140000 430.360000  13.540000 ;
      RECT 429.855000  41.170000 430.025000  45.640000 ;
      RECT 429.920000  21.230000 430.090000  22.400000 ;
      RECT 429.980000 230.315000 430.150000 234.225000 ;
      RECT 429.980000 234.225000 431.310000 234.735000 ;
      RECT 429.980000 234.735000 430.150000 236.060000 ;
      RECT 430.010000 237.915000 430.180000 238.965000 ;
      RECT 430.010000 247.190000 430.180000 249.900000 ;
      RECT 430.065000 222.650000 430.235000 225.360000 ;
      RECT 430.115000  38.575000 430.645000  41.000000 ;
      RECT 430.125000  47.080000 430.635000  47.410000 ;
      RECT 430.140000 141.155000 430.470000 141.805000 ;
      RECT 430.140000 160.345000 430.470000 160.995000 ;
      RECT 430.140000 179.535000 430.470000 180.185000 ;
      RECT 430.195000  41.000000 430.565000  47.080000 ;
      RECT 430.220000 180.925000 430.390000 199.940000 ;
      RECT 430.220000 199.940000 441.730000 200.115000 ;
      RECT 430.280000 237.415000 430.790000 237.745000 ;
      RECT 430.280000 250.370000 430.790000 250.700000 ;
      RECT 430.320000  24.395000 430.490000  27.475000 ;
      RECT 430.350000  21.060000 430.520000  22.400000 ;
      RECT 430.350000 237.745000 430.720000 239.240000 ;
      RECT 430.350000 239.750000 430.720000 250.370000 ;
      RECT 430.385000  92.780000 430.915000  92.950000 ;
      RECT 430.480000  49.850000 431.580000  50.020000 ;
      RECT 430.480000  56.485000 430.810000  57.175000 ;
      RECT 430.480000  63.640000 430.810000  64.330000 ;
      RECT 430.480000  70.795000 430.810000  71.485000 ;
      RECT 430.480000  77.950000 430.810000  78.640000 ;
      RECT 430.480000  85.105000 430.810000  85.795000 ;
      RECT 430.480000  92.260000 430.810000  92.780000 ;
      RECT 430.480000  99.415000 430.810000 100.105000 ;
      RECT 430.480000 106.570000 430.810000 107.260000 ;
      RECT 430.480000 113.725000 430.810000 114.415000 ;
      RECT 430.480000 120.880000 430.810000 121.570000 ;
      RECT 430.480000 128.035000 430.810000 128.725000 ;
      RECT 430.485000 206.365000 431.335000 211.275000 ;
      RECT 430.520000  18.735000 431.050000  18.905000 ;
      RECT 430.565000  29.165000 431.115000  36.060000 ;
      RECT 430.600000 230.620000 430.770000 233.330000 ;
      RECT 430.600000 234.995000 430.770000 236.060000 ;
      RECT 430.645000  22.940000 431.175000  23.110000 ;
      RECT 430.645000  23.110000 430.955000  23.805000 ;
      RECT 430.645000  23.805000 431.610000  23.975000 ;
      RECT 430.770000   9.960000 430.940000  11.015000 ;
      RECT 430.770000  12.020000 430.940000  14.730000 ;
      RECT 430.780000  21.230000 430.950000  22.400000 ;
      RECT 430.785000  24.145000 430.955000  24.375000 ;
      RECT 430.785000  24.375000 431.070000  27.085000 ;
      RECT 430.790000 229.900000 431.460000 230.070000 ;
      RECT 430.805000  41.170000 430.975000  42.220000 ;
      RECT 430.805000  42.450000 431.525000  42.780000 ;
      RECT 430.805000  43.400000 431.525000  43.730000 ;
      RECT 430.805000  43.900000 430.975000  46.915000 ;
      RECT 430.815000  40.170000 432.385000  40.370000 ;
      RECT 430.845000 218.340000 431.015000 228.475000 ;
      RECT 430.870000 236.230000 431.380000 236.560000 ;
      RECT 430.880000  16.860000 431.050000  18.735000 ;
      RECT 430.880000  18.905000 431.050000  19.140000 ;
      RECT 430.880000  19.480000 431.050000  20.890000 ;
      RECT 430.890000 237.915000 431.060000 239.240000 ;
      RECT 430.890000 239.240000 433.720000 239.750000 ;
      RECT 430.890000 239.750000 431.060000 250.205000 ;
      RECT 430.940000 230.070000 431.310000 234.225000 ;
      RECT 430.940000 234.735000 431.310000 236.230000 ;
      RECT 430.950000 141.155000 431.280000 141.805000 ;
      RECT 430.950000 160.345000 431.280000 160.995000 ;
      RECT 430.950000 179.535000 431.280000 180.185000 ;
      RECT 430.950000 198.725000 431.280000 199.375000 ;
      RECT 431.125000  23.310000 431.655000  23.480000 ;
      RECT 431.125000  23.975000 431.610000  23.985000 ;
      RECT 431.125000  23.985000 431.795000  24.155000 ;
      RECT 431.125000  27.735000 433.380000  27.905000 ;
      RECT 431.145000  92.085000 432.435000  92.470000 ;
      RECT 431.145000  92.470000 431.665000  93.080000 ;
      RECT 431.165000  70.745000 431.665000  71.185000 ;
      RECT 431.165000  71.185000 433.890000  71.810000 ;
      RECT 431.185000  15.285000 431.855000  15.455000 ;
      RECT 431.240000  21.960000 431.770000  22.130000 ;
      RECT 431.240000  24.155000 431.610000  27.645000 ;
      RECT 431.240000  27.645000 433.380000  27.735000 ;
      RECT 431.245000  14.760000 431.775000  15.285000 ;
      RECT 431.250000  56.485000 431.580000  57.175000 ;
      RECT 431.250000  63.640000 431.580000  64.330000 ;
      RECT 431.250000  77.950000 433.890000  78.640000 ;
      RECT 431.250000  84.800000 433.890000  85.395000 ;
      RECT 431.250000  85.395000 432.350000  85.795000 ;
      RECT 431.250000  99.415000 431.580000 100.105000 ;
      RECT 431.250000 106.570000 431.580000 106.740000 ;
      RECT 431.250000 107.090000 431.580000 107.260000 ;
      RECT 431.250000 113.725000 431.580000 114.415000 ;
      RECT 431.250000 120.880000 431.580000 121.570000 ;
      RECT 431.250000 128.035000 431.580000 128.725000 ;
      RECT 431.250000 135.190000 432.350000 135.360000 ;
      RECT 431.285000  29.165000 432.295000  30.175000 ;
      RECT 431.285000  30.175000 431.815000  34.635000 ;
      RECT 431.335000 106.740000 431.505000 107.090000 ;
      RECT 431.345000  22.130000 431.655000  23.310000 ;
      RECT 431.355000  41.170000 431.525000  42.220000 ;
      RECT 431.355000  43.900000 431.525000  46.915000 ;
      RECT 431.395000 219.210000 432.855000 219.880000 ;
      RECT 431.460000  16.850000 431.630000  21.960000 ;
      RECT 431.480000 230.315000 431.650000 235.935000 ;
      RECT 431.625000 222.650000 431.795000 225.360000 ;
      RECT 431.670000 229.900000 432.340000 230.070000 ;
      RECT 431.695000  40.670000 432.205000  41.000000 ;
      RECT 431.695000  47.080000 432.205000  47.410000 ;
      RECT 431.735000 236.310000 432.265000 236.480000 ;
      RECT 431.750000 236.230000 432.260000 236.310000 ;
      RECT 431.750000 236.480000 432.260000 236.560000 ;
      RECT 431.760000 141.155000 432.090000 141.805000 ;
      RECT 431.760000 160.345000 432.090000 160.995000 ;
      RECT 431.760000 179.535000 432.090000 180.185000 ;
      RECT 431.760000 198.725000 432.090000 199.375000 ;
      RECT 431.765000  41.000000 432.135000  47.080000 ;
      RECT 431.780000  24.375000 431.950000  27.475000 ;
      RECT 431.820000 230.070000 432.190000 236.230000 ;
      RECT 431.825000  22.550000 432.110000  22.720000 ;
      RECT 431.825000  22.720000 431.995000  23.625000 ;
      RECT 431.825000  23.625000 432.290000  23.795000 ;
      RECT 431.830000 207.410000 432.480000 209.680000 ;
      RECT 431.830000 209.680000 432.850000 209.850000 ;
      RECT 431.850000 225.910000 433.990000 226.080000 ;
      RECT 431.900000  11.820000 432.430000  11.990000 ;
      RECT 431.915000  49.850000 432.445000  50.020000 ;
      RECT 431.935000  92.740000 432.435000  97.165000 ;
      RECT 431.935000  97.165000 433.205000  97.610000 ;
      RECT 431.935000  99.415000 432.435000  99.895000 ;
      RECT 431.935000  99.895000 433.205000 100.145000 ;
      RECT 431.935000 106.570000 433.205000 107.260000 ;
      RECT 431.935000 113.610000 433.205000 114.065000 ;
      RECT 431.935000 114.065000 432.435000 114.415000 ;
      RECT 431.940000  21.625000 432.110000  22.550000 ;
      RECT 431.985000  30.850000 432.155000  31.755000 ;
      RECT 431.985000  31.925000 432.515000  36.060000 ;
      RECT 432.020000  56.485000 432.350000  57.175000 ;
      RECT 432.020000  63.640000 432.350000  64.330000 ;
      RECT 432.020000  70.495000 433.120000  71.005000 ;
      RECT 432.020000 120.880000 432.350000 121.570000 ;
      RECT 432.020000 128.035000 432.350000 128.725000 ;
      RECT 432.050000   9.960000 432.220000  11.820000 ;
      RECT 432.050000  11.990000 432.220000  14.730000 ;
      RECT 432.120000  23.795000 432.290000  24.375000 ;
      RECT 432.120000  24.375000 432.830000  24.845000 ;
      RECT 432.165000  23.125000 432.785000  23.455000 ;
      RECT 432.305000  41.170000 432.475000  45.640000 ;
      RECT 432.350000  30.475000 432.885000  30.645000 ;
      RECT 432.360000 230.620000 432.530000 233.330000 ;
      RECT 432.360000 234.570000 432.530000 236.060000 ;
      RECT 432.390000  16.720000 435.760000  16.890000 ;
      RECT 432.420000  11.450000 432.950000  11.620000 ;
      RECT 432.430000  17.240000 432.600000  19.950000 ;
      RECT 432.460000  23.455000 432.785000  23.710000 ;
      RECT 432.460000  23.710000 433.380000  23.880000 ;
      RECT 432.505000 222.650000 432.675000 225.360000 ;
      RECT 432.550000  16.890000 435.600000  17.025000 ;
      RECT 432.565000  37.775000 433.095000  41.000000 ;
      RECT 432.570000 141.155000 432.900000 141.805000 ;
      RECT 432.570000 160.345000 432.900000 160.995000 ;
      RECT 432.570000 179.535000 432.900000 180.185000 ;
      RECT 432.570000 198.725000 432.900000 199.375000 ;
      RECT 432.575000  47.080000 433.085000  47.410000 ;
      RECT 432.575000 226.570000 433.085000 227.580000 ;
      RECT 432.600000   9.960000 432.770000  11.450000 ;
      RECT 432.600000  11.620000 432.770000  14.730000 ;
      RECT 432.645000  41.000000 433.015000  47.080000 ;
      RECT 432.660000  24.845000 432.830000  27.085000 ;
      RECT 432.680000 207.585000 432.850000 207.855000 ;
      RECT 432.680000 207.855000 433.280000 208.025000 ;
      RECT 432.680000 208.025000 432.850000 208.255000 ;
      RECT 432.680000 209.515000 432.850000 209.680000 ;
      RECT 432.680000 209.850000 432.850000 210.185000 ;
      RECT 432.705000  28.330000 444.675000  28.335000 ;
      RECT 432.705000  28.335000 432.885000  30.475000 ;
      RECT 432.705000  30.645000 432.885000  30.735000 ;
      RECT 432.705000  31.495000 432.885000  36.230000 ;
      RECT 432.705000  97.610000 433.205000  99.625000 ;
      RECT 432.705000 114.970000 433.205000 135.640000 ;
      RECT 432.770000 220.640000 432.940000 221.650000 ;
      RECT 432.790000  49.790000 433.890000  50.300000 ;
      RECT 432.790000  56.485000 433.120000  57.175000 ;
      RECT 432.790000  63.640000 433.120000  64.330000 ;
      RECT 432.790000  85.585000 433.890000  85.925000 ;
      RECT 432.790000  92.260000 433.120000  92.950000 ;
      RECT 432.820000  20.840000 432.990000  22.635000 ;
      RECT 432.825000 220.220000 433.825000 220.390000 ;
      RECT 432.835000  20.040000 433.380000  20.210000 ;
      RECT 432.925000  20.440000 433.455000  20.500000 ;
      RECT 432.925000  20.500000 433.935000  20.670000 ;
      RECT 432.945000  15.280000 433.615000  15.450000 ;
      RECT 432.980000 230.620000 433.150000 233.330000 ;
      RECT 432.980000 234.995000 433.150000 236.060000 ;
      RECT 433.000000  26.625000 433.380000  27.645000 ;
      RECT 433.005000  15.130000 433.535000  15.280000 ;
      RECT 433.005000 137.945000 433.185000 138.355000 ;
      RECT 433.005000 138.525000 433.185000 139.415000 ;
      RECT 433.005000 139.585000 433.185000 139.995000 ;
      RECT 433.010000 237.915000 433.180000 238.980000 ;
      RECT 433.010000 247.190000 433.180000 249.900000 ;
      RECT 433.040000  23.070000 433.710000  23.240000 ;
      RECT 433.110000  22.940000 433.640000  23.070000 ;
      RECT 433.130000 208.220000 433.860000 209.540000 ;
      RECT 433.140000 227.830000 434.580000 228.000000 ;
      RECT 433.160000 234.010000 433.690000 234.180000 ;
      RECT 433.165000 222.630000 433.695000 222.800000 ;
      RECT 433.165000 222.800000 433.335000 225.360000 ;
      RECT 433.170000 229.900000 433.840000 230.070000 ;
      RECT 433.190000 207.440000 433.860000 207.610000 ;
      RECT 433.190000 210.150000 433.860000 210.325000 ;
      RECT 433.190000 210.325000 435.390000 210.995000 ;
      RECT 433.210000  17.240000 433.380000  20.040000 ;
      RECT 433.210000  20.210000 433.380000  20.240000 ;
      RECT 433.210000  23.880000 433.380000  25.045000 ;
      RECT 433.250000 236.230000 433.760000 236.560000 ;
      RECT 433.255000  41.170000 433.425000  42.235000 ;
      RECT 433.255000  42.405000 433.425000  42.780000 ;
      RECT 433.255000  43.400000 433.425000  43.730000 ;
      RECT 433.255000  43.900000 433.425000  46.610000 ;
      RECT 433.265000  40.200000 434.225000  40.370000 ;
      RECT 433.280000 237.415000 433.790000 237.745000 ;
      RECT 433.280000 250.370000 433.790000 250.700000 ;
      RECT 433.300000  11.450000 434.990000  11.620000 ;
      RECT 433.310000  25.520000 434.840000  26.270000 ;
      RECT 433.320000 230.070000 433.690000 234.010000 ;
      RECT 433.320000 234.180000 433.690000 236.230000 ;
      RECT 433.340000  22.565000 433.870000  22.735000 ;
      RECT 433.345000 226.270000 433.515000 227.580000 ;
      RECT 433.350000 237.745000 433.720000 239.240000 ;
      RECT 433.350000 239.750000 433.720000 250.370000 ;
      RECT 433.380000 141.155000 433.710000 141.805000 ;
      RECT 433.380000 160.345000 433.710000 160.995000 ;
      RECT 433.380000 179.535000 433.710000 180.185000 ;
      RECT 433.380000 198.725000 433.710000 199.375000 ;
      RECT 433.520000 219.185000 434.050000 219.880000 ;
      RECT 433.525000  40.670000 434.035000  41.000000 ;
      RECT 433.525000  47.080000 434.035000  47.410000 ;
      RECT 433.550000  24.375000 434.600000  25.520000 ;
      RECT 433.550000  26.270000 434.600000  27.475000 ;
      RECT 433.560000  56.485000 433.890000  57.175000 ;
      RECT 433.560000  63.640000 433.890000  64.330000 ;
      RECT 433.560000  70.495000 434.660000  71.005000 ;
      RECT 433.560000  92.260000 433.890000  92.950000 ;
      RECT 433.560000  99.415000 433.890000 100.105000 ;
      RECT 433.560000 106.570000 433.890000 107.260000 ;
      RECT 433.560000 113.725000 433.890000 114.415000 ;
      RECT 433.560000 120.880000 433.890000 121.570000 ;
      RECT 433.560000 128.035000 433.890000 128.725000 ;
      RECT 433.560000 134.945000 434.660000 135.400000 ;
      RECT 433.595000  41.000000 433.965000  47.080000 ;
      RECT 433.650000 220.580000 434.625000 220.790000 ;
      RECT 433.650000 220.790000 434.370000 221.650000 ;
      RECT 433.700000  21.625000 433.870000  22.565000 ;
      RECT 433.775000 226.570000 433.945000 227.600000 ;
      RECT 433.860000 230.315000 434.030000 235.935000 ;
      RECT 433.880000   9.960000 434.050000  11.015000 ;
      RECT 433.880000  12.020000 434.050000  14.730000 ;
      RECT 433.890000 238.040000 434.060000 250.205000 ;
      RECT 433.980000 136.685000 444.415000 139.805000 ;
      RECT 433.990000  17.240000 434.160000  19.950000 ;
      RECT 434.015000 220.080000 434.625000 220.580000 ;
      RECT 434.035000 218.520000 434.625000 218.690000 ;
      RECT 434.045000 222.650000 434.215000 225.360000 ;
      RECT 434.050000 229.900000 434.720000 230.070000 ;
      RECT 434.130000 236.230000 434.640000 236.560000 ;
      RECT 434.135000  41.295000 434.305000  46.915000 ;
      RECT 434.145000 237.495000 434.675000 237.665000 ;
      RECT 434.160000 237.415000 434.670000 237.495000 ;
      RECT 434.160000 237.665000 434.670000 237.745000 ;
      RECT 434.160000 250.370000 434.670000 250.700000 ;
      RECT 434.190000 141.155000 434.520000 141.805000 ;
      RECT 434.190000 160.345000 434.520000 160.995000 ;
      RECT 434.190000 179.535000 434.520000 180.185000 ;
      RECT 434.190000 198.725000 434.520000 199.375000 ;
      RECT 434.200000 230.070000 434.570000 236.230000 ;
      RECT 434.205000 226.270000 434.375000 227.580000 ;
      RECT 434.210000  71.315000 434.740000  71.485000 ;
      RECT 434.215000  20.500000 435.225000  20.670000 ;
      RECT 434.225000 120.880000 434.755000 121.050000 ;
      RECT 434.230000 237.745000 434.600000 250.370000 ;
      RECT 434.250000 218.690000 434.625000 220.080000 ;
      RECT 434.280000  21.625000 434.450000  22.565000 ;
      RECT 434.280000  22.565000 434.810000  22.735000 ;
      RECT 434.330000  49.785000 435.430000  50.295000 ;
      RECT 434.330000  56.485000 434.660000  57.175000 ;
      RECT 434.330000  63.640000 434.660000  64.330000 ;
      RECT 434.330000  77.950000 434.660000  78.640000 ;
      RECT 434.330000  85.105000 434.660000  85.795000 ;
      RECT 434.330000  92.260000 434.660000  92.950000 ;
      RECT 434.330000  99.415000 434.660000 100.105000 ;
      RECT 434.330000 106.570000 434.660000 107.260000 ;
      RECT 434.330000 113.725000 434.660000 114.415000 ;
      RECT 434.330000 121.050000 434.660000 121.570000 ;
      RECT 434.330000 128.035000 434.660000 128.725000 ;
      RECT 434.395000  39.375000 434.925000  41.000000 ;
      RECT 434.405000  47.080000 434.915000  47.410000 ;
      RECT 434.440000  23.070000 435.110000  23.240000 ;
      RECT 434.460000  13.140000 434.990000  13.340000 ;
      RECT 434.460000  13.340000 438.335000  13.565000 ;
      RECT 434.460000  13.565000 443.200000  15.625000 ;
      RECT 434.460000  15.625000 442.220000  15.685000 ;
      RECT 434.475000  41.000000 434.845000  47.080000 ;
      RECT 434.510000  22.940000 435.040000  23.070000 ;
      RECT 434.540000 207.340000 434.710000 210.050000 ;
      RECT 434.625000 220.980000 434.795000 221.650000 ;
      RECT 434.635000 226.570000 435.145000 227.580000 ;
      RECT 434.695000  20.440000 435.225000  20.500000 ;
      RECT 434.740000 230.620000 434.910000 233.330000 ;
      RECT 434.740000 234.225000 436.070000 234.735000 ;
      RECT 434.740000 234.735000 434.910000 236.060000 ;
      RECT 434.770000  17.240000 434.940000  20.040000 ;
      RECT 434.770000  20.040000 435.315000  20.210000 ;
      RECT 434.770000  20.210000 434.940000  20.240000 ;
      RECT 434.770000  23.710000 435.690000  23.880000 ;
      RECT 434.770000  23.880000 434.940000  25.045000 ;
      RECT 434.770000  26.625000 435.150000  27.645000 ;
      RECT 434.770000  27.645000 436.910000  27.735000 ;
      RECT 434.770000  27.735000 437.025000  27.905000 ;
      RECT 434.770000 237.915000 434.940000 239.240000 ;
      RECT 434.770000 239.240000 436.100000 239.750000 ;
      RECT 434.770000 247.190000 434.940000 249.900000 ;
      RECT 434.825000 218.520000 435.415000 218.690000 ;
      RECT 434.825000 218.690000 435.370000 220.220000 ;
      RECT 434.910000 207.540000 435.215000 210.325000 ;
      RECT 434.985000  92.260000 435.515000  92.430000 ;
      RECT 435.000000 141.155000 435.330000 141.805000 ;
      RECT 435.000000 160.345000 435.330000 160.995000 ;
      RECT 435.000000 179.535000 435.330000 180.185000 ;
      RECT 435.000000 198.725000 435.330000 199.375000 ;
      RECT 435.015000  41.170000 435.185000  42.990000 ;
      RECT 435.015000  43.900000 435.185000  46.610000 ;
      RECT 435.015000  93.535000 435.515000 135.640000 ;
      RECT 435.015000 220.470000 435.685000 220.640000 ;
      RECT 435.095000  40.200000 435.655000  40.370000 ;
      RECT 435.100000  56.485000 435.430000  57.175000 ;
      RECT 435.100000  63.640000 435.430000  64.330000 ;
      RECT 435.100000  70.795000 435.430000  71.485000 ;
      RECT 435.100000  77.950000 435.430000  78.640000 ;
      RECT 435.100000  85.105000 435.430000  85.795000 ;
      RECT 435.160000   9.960000 435.330000  12.540000 ;
      RECT 435.160000  12.540000 435.740000  12.710000 ;
      RECT 435.160000  12.710000 435.330000  13.100000 ;
      RECT 435.160000  20.840000 435.330000  22.635000 ;
      RECT 435.290000 222.890000 435.820000 223.900000 ;
      RECT 435.290000 224.570000 435.820000 225.580000 ;
      RECT 435.320000  24.375000 436.030000  24.845000 ;
      RECT 435.320000  24.845000 435.490000  27.085000 ;
      RECT 435.360000 230.620000 435.530000 233.330000 ;
      RECT 435.360000 235.010000 435.530000 236.060000 ;
      RECT 435.365000  23.125000 435.985000  23.455000 ;
      RECT 435.365000  23.455000 435.690000  23.710000 ;
      RECT 435.390000 237.915000 435.560000 238.965000 ;
      RECT 435.390000 247.190000 435.560000 249.900000 ;
      RECT 435.420000 207.340000 436.740000 210.110000 ;
      RECT 435.535000  28.335000 441.625000  28.690000 ;
      RECT 435.535000  28.690000 435.715000  30.475000 ;
      RECT 435.535000  30.475000 436.070000  30.645000 ;
      RECT 435.535000  30.645000 435.715000  30.790000 ;
      RECT 435.550000  17.240000 435.720000  19.950000 ;
      RECT 435.550000 229.900000 436.220000 230.070000 ;
      RECT 435.565000  41.170000 435.735000  43.350000 ;
      RECT 435.565000  43.900000 435.735000  46.610000 ;
      RECT 435.630000 236.230000 436.140000 236.560000 ;
      RECT 435.645000  31.945000 435.815000  35.315000 ;
      RECT 435.645000  35.315000 441.255000  35.485000 ;
      RECT 435.660000 237.415000 436.170000 237.745000 ;
      RECT 435.660000 250.370000 436.170000 250.700000 ;
      RECT 435.695000 224.150000 438.955000 224.320000 ;
      RECT 435.700000 230.070000 436.070000 234.225000 ;
      RECT 435.700000 234.735000 436.070000 236.230000 ;
      RECT 435.705000 219.125000 436.235000 220.220000 ;
      RECT 435.730000 237.745000 436.100000 239.240000 ;
      RECT 435.730000 239.750000 436.100000 250.370000 ;
      RECT 435.740000  13.140000 438.355000  13.280000 ;
      RECT 435.740000  13.280000 438.335000  13.340000 ;
      RECT 435.755000  49.950000 435.985000  66.660000 ;
      RECT 435.785000  49.540000 435.955000  49.950000 ;
      RECT 435.785000  66.660000 435.955000 135.640000 ;
      RECT 435.810000 141.155000 436.140000 141.805000 ;
      RECT 435.810000 160.345000 436.140000 160.995000 ;
      RECT 435.810000 179.535000 436.140000 180.185000 ;
      RECT 435.810000 198.725000 436.140000 199.375000 ;
      RECT 435.825000  38.145000 436.355000  41.000000 ;
      RECT 435.835000  47.080000 436.345000  47.410000 ;
      RECT 435.860000  23.625000 436.325000  23.795000 ;
      RECT 435.860000  23.795000 436.030000  24.375000 ;
      RECT 435.905000  41.000000 436.275000  47.080000 ;
      RECT 435.905000 220.980000 436.075000 221.870000 ;
      RECT 436.040000  21.625000 436.210000  22.550000 ;
      RECT 436.040000  22.550000 436.325000  22.720000 ;
      RECT 436.125000  29.165000 436.295000  30.245000 ;
      RECT 436.125000  32.255000 436.295000  34.965000 ;
      RECT 436.155000  22.720000 436.325000  23.625000 ;
      RECT 436.200000  24.375000 436.370000  27.475000 ;
      RECT 436.225000  92.260000 436.755000  92.430000 ;
      RECT 436.225000  93.535000 436.725000 135.640000 ;
      RECT 436.240000 230.315000 436.410000 234.225000 ;
      RECT 436.240000 234.225000 437.570000 234.735000 ;
      RECT 436.240000 234.735000 436.410000 236.060000 ;
      RECT 436.270000 237.915000 436.440000 250.205000 ;
      RECT 436.310000  49.785000 437.410000  50.295000 ;
      RECT 436.310000  56.485000 436.640000  57.175000 ;
      RECT 436.310000  63.640000 436.640000  64.330000 ;
      RECT 436.310000  70.795000 436.640000  71.485000 ;
      RECT 436.310000  77.950000 436.640000  78.640000 ;
      RECT 436.310000  85.105000 436.640000  85.795000 ;
      RECT 436.355000  23.985000 437.025000  24.155000 ;
      RECT 436.380000  21.960000 436.910000  22.130000 ;
      RECT 436.420000 226.570000 436.930000 227.580000 ;
      RECT 436.440000   9.960000 436.610000  11.015000 ;
      RECT 436.440000  12.090000 436.610000  13.140000 ;
      RECT 436.445000  41.295000 436.615000  46.915000 ;
      RECT 436.470000 222.890000 437.000000 223.900000 ;
      RECT 436.495000  22.130000 436.805000  23.310000 ;
      RECT 436.495000  23.310000 437.025000  23.480000 ;
      RECT 436.520000  16.850000 436.690000  21.960000 ;
      RECT 436.540000  23.805000 437.505000  23.975000 ;
      RECT 436.540000  23.975000 437.025000  23.985000 ;
      RECT 436.540000  24.155000 436.910000  27.645000 ;
      RECT 436.585000  29.165000 436.755000  34.965000 ;
      RECT 436.595000 224.560000 436.875000 225.770000 ;
      RECT 436.595000 225.770000 439.220000 226.020000 ;
      RECT 436.620000 141.155000 436.950000 141.805000 ;
      RECT 436.620000 160.345000 436.950000 160.995000 ;
      RECT 436.620000 179.535000 436.950000 180.185000 ;
      RECT 436.620000 198.725000 436.950000 199.375000 ;
      RECT 436.705000  38.575000 437.235000  41.000000 ;
      RECT 436.715000  47.080000 437.225000  47.410000 ;
      RECT 436.755000 206.950000 437.425000 207.120000 ;
      RECT 436.785000  41.000000 437.155000  47.080000 ;
      RECT 436.860000 230.620000 437.030000 233.330000 ;
      RECT 436.860000 234.995000 437.030000 236.060000 ;
      RECT 436.890000 237.915000 437.060000 238.980000 ;
      RECT 436.890000 247.190000 437.060000 249.900000 ;
      RECT 436.925000  30.600000 439.075000  30.770000 ;
      RECT 436.975000  22.940000 437.505000  23.110000 ;
      RECT 436.985000 120.880000 437.515000 121.050000 ;
      RECT 436.985000 227.830000 438.425000 228.000000 ;
      RECT 437.000000  71.315000 437.530000  71.485000 ;
      RECT 437.045000  29.165000 437.215000  30.245000 ;
      RECT 437.045000  32.255000 437.215000  34.965000 ;
      RECT 437.050000 229.900000 437.720000 230.070000 ;
      RECT 437.070000 239.795000 437.600000 239.965000 ;
      RECT 437.080000  24.375000 437.365000  27.085000 ;
      RECT 437.080000  56.485000 437.410000  57.175000 ;
      RECT 437.080000  63.640000 437.410000  64.330000 ;
      RECT 437.080000  70.495000 438.180000  71.005000 ;
      RECT 437.080000  77.950000 437.410000  78.640000 ;
      RECT 437.080000  85.105000 437.410000  85.795000 ;
      RECT 437.080000  92.260000 437.410000  92.950000 ;
      RECT 437.080000  99.415000 437.410000 100.105000 ;
      RECT 437.080000 106.570000 437.410000 107.260000 ;
      RECT 437.080000 113.725000 437.410000 114.415000 ;
      RECT 437.080000 121.050000 437.410000 121.570000 ;
      RECT 437.080000 128.035000 437.410000 128.725000 ;
      RECT 437.080000 134.945000 438.180000 135.400000 ;
      RECT 437.100000  16.860000 437.270000  18.735000 ;
      RECT 437.100000  18.735000 437.630000  18.905000 ;
      RECT 437.100000  18.905000 437.270000  19.140000 ;
      RECT 437.100000  19.310000 439.630000  19.480000 ;
      RECT 437.100000  19.480000 437.270000  20.890000 ;
      RECT 437.100000  20.890000 438.660000  21.060000 ;
      RECT 437.120000 222.000000 438.020000 222.140000 ;
      RECT 437.120000 222.140000 437.650000 222.170000 ;
      RECT 437.130000 236.230000 437.640000 236.560000 ;
      RECT 437.135000 226.020000 437.415000 227.590000 ;
      RECT 437.160000 237.415000 437.670000 237.745000 ;
      RECT 437.160000 250.370000 437.670000 250.700000 ;
      RECT 437.170000 218.710000 437.340000 221.420000 ;
      RECT 437.195000  23.110000 437.505000  23.805000 ;
      RECT 437.195000  24.145000 437.365000  24.375000 ;
      RECT 437.200000  21.230000 437.370000  22.400000 ;
      RECT 437.200000 230.070000 437.570000 234.225000 ;
      RECT 437.200000 234.735000 437.570000 236.230000 ;
      RECT 437.230000 237.745000 437.600000 239.795000 ;
      RECT 437.230000 239.965000 437.600000 250.370000 ;
      RECT 437.325000  41.170000 437.495000  42.235000 ;
      RECT 437.325000  42.405000 437.495000  42.780000 ;
      RECT 437.325000  43.200000 437.495000  43.730000 ;
      RECT 437.325000  43.900000 437.495000  46.610000 ;
      RECT 437.350000 221.970000 438.020000 222.000000 ;
      RECT 437.405000  40.200000 440.605000  40.370000 ;
      RECT 437.430000 141.155000 437.760000 141.805000 ;
      RECT 437.430000 160.345000 437.760000 160.995000 ;
      RECT 437.430000 179.535000 437.760000 180.185000 ;
      RECT 437.430000 198.725000 437.760000 199.375000 ;
      RECT 437.450000 207.340000 437.620000 210.050000 ;
      RECT 437.465000   8.930000 438.355000   9.310000 ;
      RECT 437.465000  11.275000 438.355000  12.165000 ;
      RECT 437.465000  13.110000 438.355000  13.140000 ;
      RECT 437.485000   9.310000 438.335000  11.275000 ;
      RECT 437.485000  12.165000 438.335000  13.110000 ;
      RECT 437.485000  22.600000 438.835000  22.770000 ;
      RECT 437.525000  31.945000 437.695000  35.315000 ;
      RECT 437.585000  22.570000 438.835000  22.600000 ;
      RECT 437.595000  40.670000 438.105000  41.000000 ;
      RECT 437.595000  47.080000 438.105000  47.410000 ;
      RECT 437.620000 226.570000 437.790000 227.580000 ;
      RECT 437.630000  21.060000 437.800000  22.400000 ;
      RECT 437.635000 222.890000 438.165000 223.900000 ;
      RECT 437.635000 224.570000 438.165000 225.580000 ;
      RECT 437.660000  24.395000 437.830000  27.475000 ;
      RECT 437.665000  41.000000 438.035000  47.080000 ;
      RECT 437.740000 230.315000 437.910000 235.935000 ;
      RECT 437.745000  29.165000 437.915000  30.245000 ;
      RECT 437.770000 238.040000 437.940000 250.205000 ;
      RECT 437.850000  49.790000 438.950000  50.300000 ;
      RECT 437.850000  56.485000 438.180000  57.175000 ;
      RECT 437.850000  63.640000 438.180000  64.330000 ;
      RECT 437.850000  71.185000 440.575000  71.810000 ;
      RECT 437.850000  77.950000 440.490000  78.640000 ;
      RECT 437.850000  84.800000 440.490000  85.395000 ;
      RECT 437.850000  85.585000 438.950000  85.925000 ;
      RECT 437.850000  92.260000 438.180000  92.950000 ;
      RECT 437.850000  99.415000 438.180000 100.105000 ;
      RECT 437.850000 106.570000 438.180000 107.260000 ;
      RECT 437.850000 113.725000 438.180000 114.415000 ;
      RECT 437.850000 120.880000 438.180000 121.570000 ;
      RECT 437.850000 128.035000 438.180000 128.725000 ;
      RECT 437.930000 229.900000 438.600000 230.070000 ;
      RECT 437.945000  30.940000 438.355000  31.470000 ;
      RECT 437.995000 226.020000 438.275000 227.590000 ;
      RECT 438.000000 236.310000 438.530000 236.480000 ;
      RECT 438.010000 236.230000 438.520000 236.310000 ;
      RECT 438.010000 236.480000 438.520000 236.560000 ;
      RECT 438.025000  33.575000 438.335000  34.965000 ;
      RECT 438.040000 237.415000 438.550000 237.745000 ;
      RECT 438.040000 250.370000 438.550000 250.700000 ;
      RECT 438.050000 218.710000 438.220000 221.420000 ;
      RECT 438.060000  21.230000 438.230000  22.400000 ;
      RECT 438.080000 230.070000 438.450000 236.230000 ;
      RECT 438.105000  32.635000 439.075000  33.305000 ;
      RECT 438.110000 237.745000 438.480000 250.370000 ;
      RECT 438.205000  41.170000 438.375000  46.910000 ;
      RECT 438.240000 141.155000 438.570000 141.805000 ;
      RECT 438.240000 160.345000 438.570000 160.995000 ;
      RECT 438.240000 179.535000 438.570000 180.185000 ;
      RECT 438.240000 198.725000 438.570000 199.375000 ;
      RECT 438.280000  16.520000 441.170000  16.690000 ;
      RECT 438.280000  16.690000 438.450000  19.140000 ;
      RECT 438.280000  19.650000 438.450000  19.790000 ;
      RECT 438.280000  19.790000 438.955000  19.960000 ;
      RECT 438.280000  19.960000 438.450000  20.660000 ;
      RECT 438.305000  25.395000 438.835000  27.655000 ;
      RECT 438.305000  27.655000 441.840000  27.905000 ;
      RECT 438.475000  40.670000 438.985000  41.000000 ;
      RECT 438.475000  47.080000 438.985000  47.410000 ;
      RECT 438.480000 226.570000 438.990000 227.580000 ;
      RECT 438.490000  21.060000 438.660000  22.400000 ;
      RECT 438.505000 222.890000 439.360000 223.900000 ;
      RECT 438.525000  29.165000 439.075000  30.600000 ;
      RECT 438.525000  30.770000 439.075000  32.635000 ;
      RECT 438.525000  33.305000 439.075000  33.985000 ;
      RECT 438.525000  33.985000 439.535000  34.155000 ;
      RECT 438.535000  97.165000 439.805000  97.610000 ;
      RECT 438.535000  97.610000 439.035000  99.625000 ;
      RECT 438.535000  99.895000 439.805000 100.145000 ;
      RECT 438.535000 106.570000 439.805000 107.260000 ;
      RECT 438.535000 113.610000 439.805000 114.065000 ;
      RECT 438.535000 114.970000 439.035000 135.640000 ;
      RECT 438.535000 135.640000 444.415000 135.670000 ;
      RECT 438.545000  41.000000 438.915000  47.080000 ;
      RECT 438.620000  56.485000 438.950000  57.175000 ;
      RECT 438.620000  63.640000 438.950000  64.330000 ;
      RECT 438.620000  70.495000 439.720000  71.005000 ;
      RECT 438.620000  92.260000 438.950000  92.950000 ;
      RECT 438.620000 135.840000 444.415000 135.870000 ;
      RECT 438.620000 230.620000 438.790000 233.330000 ;
      RECT 438.620000 234.570000 438.790000 236.060000 ;
      RECT 438.650000 237.915000 438.820000 239.240000 ;
      RECT 438.650000 239.240000 439.980000 239.750000 ;
      RECT 438.650000 247.190000 438.820000 249.900000 ;
      RECT 438.730000   9.540000 439.260000   9.710000 ;
      RECT 438.780000  18.225000 439.110000  19.075000 ;
      RECT 438.860000  17.615000 439.030000  18.225000 ;
      RECT 438.920000  21.230000 439.090000  22.400000 ;
      RECT 438.955000 224.560000 439.220000 225.770000 ;
      RECT 439.005000  24.370000 439.175000  27.370000 ;
      RECT 439.050000 141.155000 439.380000 141.805000 ;
      RECT 439.050000 160.345000 439.380000 160.995000 ;
      RECT 439.050000 179.535000 439.380000 180.185000 ;
      RECT 439.050000 198.725000 439.380000 199.375000 ;
      RECT 439.085000  41.170000 439.255000  42.220000 ;
      RECT 439.085000  42.450000 439.255000  42.780000 ;
      RECT 439.085000  43.400000 439.255000  43.730000 ;
      RECT 439.085000  43.900000 439.255000  46.610000 ;
      RECT 439.090000   8.010000 443.200000   8.880000 ;
      RECT 439.090000   8.880000 439.260000   9.540000 ;
      RECT 439.090000   9.710000 439.260000  10.560000 ;
      RECT 439.090000  10.560000 439.380000  10.730000 ;
      RECT 439.090000  10.730000 439.810000  11.060000 ;
      RECT 439.090000  11.230000 439.810000  11.560000 ;
      RECT 439.090000  11.560000 439.260000  12.750000 ;
      RECT 439.130000 206.365000 443.295000 211.275000 ;
      RECT 439.190000  22.595000 441.850000  22.765000 ;
      RECT 439.190000  22.765000 440.540000  22.770000 ;
      RECT 439.225000  23.710000 439.755000  23.880000 ;
      RECT 439.240000 230.620000 439.410000 233.330000 ;
      RECT 439.240000 234.995000 439.410000 236.060000 ;
      RECT 439.245000  33.445000 440.255000  33.615000 ;
      RECT 439.270000 237.915000 439.440000 238.965000 ;
      RECT 439.270000 247.190000 439.440000 249.900000 ;
      RECT 439.295000  49.850000 439.825000  50.020000 ;
      RECT 439.305000  29.165000 439.475000  30.245000 ;
      RECT 439.305000  92.085000 440.595000  92.470000 ;
      RECT 439.305000  92.740000 439.805000  97.165000 ;
      RECT 439.305000  99.415000 439.805000  99.895000 ;
      RECT 439.305000 114.065000 439.805000 114.415000 ;
      RECT 439.350000  20.890000 441.170000  21.060000 ;
      RECT 439.350000  21.060000 439.520000  22.400000 ;
      RECT 439.355000  40.670000 439.865000  41.000000 ;
      RECT 439.355000  47.080000 439.865000  47.410000 ;
      RECT 439.390000  56.485000 439.720000  57.175000 ;
      RECT 439.390000  63.640000 439.720000  64.330000 ;
      RECT 439.390000  85.395000 440.490000  85.795000 ;
      RECT 439.390000 120.880000 439.720000 121.570000 ;
      RECT 439.390000 128.035000 439.720000 128.725000 ;
      RECT 439.390000 135.190000 440.490000 135.360000 ;
      RECT 439.425000  41.000000 439.795000  47.080000 ;
      RECT 439.430000 229.900000 440.100000 230.070000 ;
      RECT 439.460000  16.860000 440.330000  17.870000 ;
      RECT 439.460000  18.160000 439.630000  19.310000 ;
      RECT 439.460000  19.480000 439.630000  20.660000 ;
      RECT 439.475000 236.310000 440.020000 236.480000 ;
      RECT 439.510000 236.230000 440.020000 236.310000 ;
      RECT 439.510000 236.480000 440.020000 236.560000 ;
      RECT 439.525000  40.570000 439.695000  40.670000 ;
      RECT 439.540000 237.415000 440.050000 237.745000 ;
      RECT 439.540000 250.370000 440.050000 250.700000 ;
      RECT 439.580000 230.070000 439.950000 236.230000 ;
      RECT 439.585000  23.880000 439.755000  27.230000 ;
      RECT 439.585000  27.230000 443.825000  27.400000 ;
      RECT 439.610000 237.745000 439.980000 239.240000 ;
      RECT 439.610000 239.750000 439.980000 250.370000 ;
      RECT 439.640000   9.550000 439.810000  10.560000 ;
      RECT 439.640000  11.730000 439.810000  12.740000 ;
      RECT 439.705000  29.165000 440.255000  33.445000 ;
      RECT 439.705000  33.615000 440.255000  34.295000 ;
      RECT 439.705000  34.295000 440.675000  34.965000 ;
      RECT 439.780000  21.230000 439.950000  22.400000 ;
      RECT 439.800000  17.870000 440.330000  18.905000 ;
      RECT 439.800000 218.340000 439.970000 228.475000 ;
      RECT 439.860000 141.155000 440.190000 141.805000 ;
      RECT 439.860000 160.345000 440.190000 160.995000 ;
      RECT 439.860000 179.535000 440.190000 180.185000 ;
      RECT 439.860000 198.725000 440.190000 199.375000 ;
      RECT 439.965000  41.170000 440.135000  46.915000 ;
      RECT 439.980000   9.050000 440.150000  13.240000 ;
      RECT 440.075000  70.745000 440.575000  71.185000 ;
      RECT 440.075000  92.470000 440.595000  93.080000 ;
      RECT 440.120000 230.315000 440.290000 235.935000 ;
      RECT 440.150000 237.915000 440.320000 239.240000 ;
      RECT 440.150000 239.240000 442.985000 239.750000 ;
      RECT 440.150000 239.750000 440.320000 250.205000 ;
      RECT 440.160000  49.850000 441.260000  50.020000 ;
      RECT 440.160000  56.485000 440.490000  57.175000 ;
      RECT 440.160000  63.640000 440.490000  64.330000 ;
      RECT 440.160000  99.415000 440.490000 100.105000 ;
      RECT 440.160000 106.570000 440.490000 106.740000 ;
      RECT 440.160000 107.090000 440.490000 107.260000 ;
      RECT 440.160000 113.725000 440.490000 114.415000 ;
      RECT 440.160000 120.880000 440.490000 121.570000 ;
      RECT 440.160000 128.035000 440.490000 128.725000 ;
      RECT 440.210000  21.060000 440.380000  22.400000 ;
      RECT 440.235000 106.740000 440.405000 107.090000 ;
      RECT 440.280000  19.790000 440.810000  19.960000 ;
      RECT 440.310000 229.900000 440.980000 230.070000 ;
      RECT 440.350000   9.050000 440.520000  13.240000 ;
      RECT 440.390000 236.230000 440.900000 236.560000 ;
      RECT 440.425000  30.940000 440.755000  31.470000 ;
      RECT 440.445000  32.555000 440.765000  34.025000 ;
      RECT 440.460000 230.070000 440.830000 233.875000 ;
      RECT 440.460000 233.875000 441.060000 234.045000 ;
      RECT 440.460000 234.045000 440.830000 236.230000 ;
      RECT 440.465000  24.080000 440.725000  27.060000 ;
      RECT 440.515000  41.170000 440.685000  42.235000 ;
      RECT 440.515000  42.405000 440.685000  42.780000 ;
      RECT 440.515000  43.200000 440.685000  43.730000 ;
      RECT 440.515000  43.900000 440.685000  46.610000 ;
      RECT 440.640000  16.690000 441.170000  17.870000 ;
      RECT 440.640000  18.160000 440.810000  19.790000 ;
      RECT 440.640000  19.960000 440.810000  20.660000 ;
      RECT 440.640000  21.230000 440.810000  22.400000 ;
      RECT 440.670000 141.155000 441.000000 141.805000 ;
      RECT 440.670000 160.345000 441.000000 160.995000 ;
      RECT 440.670000 179.535000 441.000000 180.185000 ;
      RECT 440.670000 198.725000 441.000000 199.375000 ;
      RECT 440.720000   9.050000 441.570000   9.380000 ;
      RECT 440.720000   9.380000 440.890000  12.910000 ;
      RECT 440.720000  12.910000 441.570000  13.240000 ;
      RECT 440.775000  36.975000 441.305000  41.000000 ;
      RECT 440.785000  47.080000 441.295000  47.410000 ;
      RECT 440.825000  92.780000 441.355000  92.950000 ;
      RECT 440.855000  41.000000 441.225000  47.080000 ;
      RECT 440.865000  29.165000 441.035000  30.245000 ;
      RECT 440.925000  24.080000 441.185000  27.060000 ;
      RECT 440.930000  56.485000 441.260000  57.175000 ;
      RECT 440.930000  63.640000 441.260000  64.330000 ;
      RECT 440.930000  70.795000 441.260000  71.485000 ;
      RECT 440.930000  77.950000 441.260000  78.640000 ;
      RECT 440.930000  85.105000 441.260000  85.795000 ;
      RECT 440.930000  92.260000 441.260000  92.780000 ;
      RECT 440.930000  99.415000 441.260000 100.105000 ;
      RECT 440.930000 106.570000 441.260000 107.260000 ;
      RECT 440.930000 113.725000 441.260000 114.415000 ;
      RECT 440.930000 120.880000 441.260000 121.570000 ;
      RECT 440.930000 128.035000 441.260000 128.725000 ;
      RECT 440.930000 135.190000 442.030000 135.360000 ;
      RECT 440.980000  17.870000 441.170000  20.890000 ;
      RECT 440.980000  21.975000 441.510000  22.145000 ;
      RECT 441.000000 230.620000 441.170000 233.330000 ;
      RECT 441.000000 234.225000 442.330000 234.735000 ;
      RECT 441.000000 234.735000 441.170000 236.060000 ;
      RECT 441.020000 217.090000 441.250000 229.405000 ;
      RECT 441.060000   9.550000 441.230000  10.560000 ;
      RECT 441.060000  10.730000 441.230000  11.060000 ;
      RECT 441.060000  11.230000 441.230000  11.560000 ;
      RECT 441.060000  11.730000 441.230000  12.740000 ;
      RECT 441.085000  31.945000 441.255000  35.315000 ;
      RECT 441.095000  30.475000 441.625000  30.645000 ;
      RECT 441.100000  23.710000 441.630000  23.880000 ;
      RECT 441.280000  22.935000 441.450000  23.710000 ;
      RECT 441.340000  16.850000 441.510000  21.975000 ;
      RECT 441.395000  41.295000 441.565000  46.915000 ;
      RECT 441.400000   9.380000 441.570000  12.910000 ;
      RECT 441.445000  28.690000 441.625000  30.475000 ;
      RECT 441.445000  30.645000 441.625000  30.790000 ;
      RECT 441.560000 140.585000 441.730000 199.940000 ;
      RECT 441.615000  49.850000 442.145000  50.020000 ;
      RECT 441.620000 230.620000 441.790000 233.330000 ;
      RECT 441.620000 235.010000 441.790000 236.060000 ;
      RECT 441.655000  38.565000 442.185000  41.000000 ;
      RECT 441.665000  47.080000 442.175000  47.410000 ;
      RECT 441.680000  20.825000 442.330000  21.835000 ;
      RECT 441.680000  21.835000 441.850000  22.595000 ;
      RECT 441.700000  56.485000 442.030000  57.175000 ;
      RECT 441.700000  63.640000 442.030000  64.330000 ;
      RECT 441.700000  70.795000 442.030000  71.485000 ;
      RECT 441.700000  77.950000 442.030000  78.640000 ;
      RECT 441.700000  85.105000 442.030000  85.795000 ;
      RECT 441.700000  92.260000 442.030000  92.950000 ;
      RECT 441.700000  99.415000 442.030000 100.105000 ;
      RECT 441.700000 106.570000 442.030000 107.260000 ;
      RECT 441.700000 113.725000 442.030000 114.415000 ;
      RECT 441.700000 120.880000 442.030000 121.570000 ;
      RECT 441.700000 128.035000 442.030000 128.725000 ;
      RECT 441.735000  41.000000 442.105000  47.080000 ;
      RECT 441.770000   9.050000 441.940000  13.240000 ;
      RECT 441.800000  18.735000 442.330000  18.905000 ;
      RECT 441.800000  23.780000 442.470000  23.950000 ;
      RECT 441.810000 229.900000 442.480000 230.070000 ;
      RECT 441.820000  16.605000 444.670000  16.775000 ;
      RECT 441.820000  16.775000 441.990000  17.385000 ;
      RECT 441.860000  23.040000 442.390000  23.210000 ;
      RECT 441.890000 236.230000 442.400000 236.560000 ;
      RECT 441.895000  23.210000 442.390000  23.780000 ;
      RECT 441.895000  23.950000 442.065000  27.060000 ;
      RECT 441.925000 215.425000 443.295000 215.440000 ;
      RECT 441.960000 230.070000 442.330000 234.225000 ;
      RECT 441.960000 234.735000 442.330000 236.230000 ;
      RECT 442.010000  27.735000 442.720000  27.905000 ;
      RECT 442.140000   9.050000 442.310000  13.240000 ;
      RECT 442.150000 139.805000 444.415000 185.105000 ;
      RECT 442.150000 185.105000 466.740000 190.715000 ;
      RECT 442.150000 190.715000 443.295000 202.215000 ;
      RECT 442.160000  17.155000 442.330000  18.735000 ;
      RECT 442.160000  18.905000 442.330000  20.825000 ;
      RECT 442.275000  41.170000 442.445000  43.350000 ;
      RECT 442.275000  43.900000 442.445000  46.610000 ;
      RECT 442.275000 237.915000 442.445000 238.980000 ;
      RECT 442.275000 247.190000 442.445000 249.900000 ;
      RECT 442.355000  40.200000 442.915000  40.370000 ;
      RECT 442.385000  49.540000 442.555000  61.065000 ;
      RECT 442.385000  61.065000 450.130000  88.065000 ;
      RECT 442.385000  88.065000 444.415000 135.640000 ;
      RECT 442.385000 218.755000 442.555000 223.505000 ;
      RECT 442.385000 223.505000 444.835000 228.605000 ;
      RECT 442.480000   9.550000 442.650000  10.560000 ;
      RECT 442.480000  10.730000 443.200000  11.060000 ;
      RECT 442.480000  11.230000 443.200000  11.560000 ;
      RECT 442.480000  11.730000 442.650000  12.740000 ;
      RECT 442.500000  20.070000 443.030000  20.240000 ;
      RECT 442.500000 230.315000 443.005000 236.060000 ;
      RECT 442.545000 237.415000 443.055000 237.745000 ;
      RECT 442.545000 250.370000 443.055000 250.700000 ;
      RECT 442.560000  22.935000 442.810000  23.605000 ;
      RECT 442.595000  20.825000 442.790000  21.835000 ;
      RECT 442.595000  21.835000 442.765000  22.935000 ;
      RECT 442.595000  23.605000 442.810000  23.660000 ;
      RECT 442.610000 218.175000 444.610000 218.345000 ;
      RECT 442.615000 237.745000 442.985000 239.240000 ;
      RECT 442.615000 239.750000 442.985000 250.370000 ;
      RECT 442.620000  17.155000 442.790000  20.070000 ;
      RECT 442.640000  23.660000 442.810000  24.350000 ;
      RECT 442.640000  24.350000 442.945000  27.060000 ;
      RECT 442.655000 230.005000 443.185000 230.175000 ;
      RECT 442.655000 230.175000 443.005000 230.315000 ;
      RECT 442.705000 136.615000 444.415000 136.685000 ;
      RECT 442.725000 136.270000 444.415000 136.615000 ;
      RECT 442.745000 135.870000 444.415000 136.270000 ;
      RECT 442.820000   9.540000 443.350000   9.710000 ;
      RECT 442.825000  41.170000 442.995000  42.990000 ;
      RECT 442.825000  43.900000 442.995000  46.610000 ;
      RECT 442.960000  17.155000 443.250000  19.575000 ;
      RECT 442.960000  19.575000 443.500000  19.865000 ;
      RECT 442.960000  20.500000 443.500000  20.655000 ;
      RECT 442.960000  20.655000 443.370000  22.670000 ;
      RECT 442.960000  22.670000 443.490000  22.840000 ;
      RECT 442.980000  23.040000 444.010000  23.210000 ;
      RECT 443.000000  27.735000 443.670000  27.905000 ;
      RECT 443.030000   8.880000 443.200000   9.540000 ;
      RECT 443.030000   9.710000 443.200000  10.730000 ;
      RECT 443.030000  11.560000 443.200000  12.750000 ;
      RECT 443.080000  23.780000 443.825000  23.950000 ;
      RECT 443.085000  38.965000 443.615000  41.000000 ;
      RECT 443.095000  47.080000 443.605000  47.410000 ;
      RECT 443.125000 218.345000 444.065000 222.180000 ;
      RECT 443.150000  23.710000 443.680000  23.780000 ;
      RECT 443.155000 238.040000 443.325000 250.205000 ;
      RECT 443.165000  41.000000 443.535000  47.080000 ;
      RECT 443.200000  19.865000 443.500000  20.500000 ;
      RECT 443.225000  53.325000 444.350000  53.370000 ;
      RECT 443.225000  53.370000 447.595000  53.540000 ;
      RECT 443.225000  53.540000 444.350000  53.585000 ;
      RECT 443.225000  53.585000 443.485000  56.940000 ;
      RECT 443.225000  58.505000 443.485000  59.970000 ;
      RECT 443.225000  59.970000 444.350000  60.015000 ;
      RECT 443.225000  60.015000 447.595000  60.185000 ;
      RECT 443.225000  60.185000 444.350000  60.230000 ;
      RECT 443.270000  56.940000 443.440000  58.505000 ;
      RECT 443.415000 237.495000 443.945000 237.665000 ;
      RECT 443.425000 237.415000 443.935000 237.495000 ;
      RECT 443.425000 237.665000 443.935000 237.745000 ;
      RECT 443.425000 250.370000 443.935000 250.700000 ;
      RECT 443.450000  16.965000 444.205000  17.135000 ;
      RECT 443.495000 237.745000 443.865000 250.370000 ;
      RECT 443.540000  20.825000 443.710000  21.835000 ;
      RECT 443.655000  23.950000 443.825000  27.230000 ;
      RECT 443.670000  19.075000 443.840000  19.770000 ;
      RECT 443.675000  18.735000 444.205000  18.905000 ;
      RECT 443.695000  19.940000 443.865000  20.610000 ;
      RECT 443.705000  41.295000 443.875000  46.915000 ;
      RECT 443.710000 192.100000 458.545000 193.220000 ;
      RECT 443.710000 193.220000 444.600000 198.880000 ;
      RECT 443.710000 198.880000 444.570000 209.620000 ;
      RECT 443.710000 209.620000 444.600000 211.910000 ;
      RECT 443.710000 211.910000 444.570000 215.230000 ;
      RECT 443.710000 215.230000 444.600000 216.230000 ;
      RECT 443.735000  22.155000 444.270000  22.730000 ;
      RECT 443.785000  40.170000 445.335000  40.370000 ;
      RECT 443.840000  22.935000 444.010000  23.040000 ;
      RECT 443.840000  23.210000 444.010000  23.605000 ;
      RECT 443.975000  40.670000 444.485000  41.000000 ;
      RECT 443.975000  47.080000 444.485000  47.410000 ;
      RECT 444.000000  20.825000 444.205000  21.835000 ;
      RECT 444.030000  54.740000 446.830000  54.910000 ;
      RECT 444.030000  56.300000 446.830000  56.470000 ;
      RECT 444.030000  57.860000 446.830000  58.030000 ;
      RECT 444.030000  59.420000 446.830000  59.590000 ;
      RECT 444.035000  17.135000 444.205000  18.735000 ;
      RECT 444.035000  18.905000 444.205000  20.825000 ;
      RECT 444.035000 237.915000 444.205000 239.240000 ;
      RECT 444.035000 239.240000 445.365000 239.750000 ;
      RECT 444.035000 247.190000 444.205000 249.900000 ;
      RECT 444.045000  41.000000 444.415000  47.080000 ;
      RECT 444.120000  53.960000 446.830000  54.130000 ;
      RECT 444.120000  55.520000 446.830000  55.690000 ;
      RECT 444.120000  57.080000 446.830000  57.250000 ;
      RECT 444.120000  58.640000 446.830000  58.810000 ;
      RECT 444.370000 232.320000 444.600000 234.950000 ;
      RECT 444.370000 234.950000 470.480000 235.180000 ;
      RECT 444.400000 229.655000 444.570000 232.320000 ;
      RECT 444.495000  22.835000 444.675000  28.150000 ;
      RECT 444.500000  16.775000 444.670000  17.385000 ;
      RECT 444.500000  20.815000 444.670000  22.835000 ;
      RECT 444.510000   6.600000 477.515000  11.235000 ;
      RECT 444.585000  41.170000 444.755000  42.235000 ;
      RECT 444.585000  42.405000 446.350000  42.780000 ;
      RECT 444.585000  43.400000 445.335000  43.730000 ;
      RECT 444.585000  43.900000 444.755000  46.610000 ;
      RECT 444.655000 237.915000 444.825000 238.965000 ;
      RECT 444.655000 247.190000 444.825000 249.900000 ;
      RECT 444.665000 218.755000 444.835000 223.505000 ;
      RECT 444.860000  61.055000 450.130000  61.065000 ;
      RECT 444.925000 237.415000 445.435000 237.745000 ;
      RECT 444.925000 250.370000 445.435000 250.700000 ;
      RECT 444.955000  40.370000 445.335000  41.740000 ;
      RECT 444.955000  41.740000 446.350000  42.405000 ;
      RECT 444.995000 237.745000 445.365000 239.240000 ;
      RECT 444.995000 239.750000 445.365000 250.370000 ;
      RECT 445.155000  48.600000 445.335000  51.285000 ;
      RECT 445.160000  43.730000 445.335000  47.075000 ;
      RECT 445.165000  47.075000 445.335000  47.580000 ;
      RECT 445.200000  54.130000 446.810000  54.230000 ;
      RECT 445.320000  11.235000 477.515000  11.240000 ;
      RECT 445.320000  11.240000 447.420000  24.755000 ;
      RECT 445.320000  24.755000 477.515000  29.000000 ;
      RECT 445.320000  29.000000 450.130000  39.285000 ;
      RECT 445.425000 113.455000 446.290000 145.465000 ;
      RECT 445.425000 145.465000 462.110000 146.460000 ;
      RECT 445.425000 146.460000 446.290000 182.820000 ;
      RECT 445.425000 182.820000 462.110000 183.680000 ;
      RECT 445.425000 183.680000 447.490000 183.685000 ;
      RECT 445.430000  89.195000 462.110000  90.055000 ;
      RECT 445.430000  90.055000 446.290000 113.455000 ;
      RECT 445.535000 237.915000 445.705000 239.235000 ;
      RECT 445.535000 239.235000 446.065000 239.405000 ;
      RECT 445.535000 239.405000 445.705000 250.205000 ;
      RECT 445.625000 199.915000 466.450000 200.145000 ;
      RECT 445.625000 201.280000 445.855000 206.125000 ;
      RECT 445.625000 209.620000 445.855000 211.185000 ;
      RECT 445.625000 211.185000 466.450000 211.415000 ;
      RECT 445.625000 211.415000 445.855000 211.910000 ;
      RECT 445.625000 215.230000 445.855000 219.275000 ;
      RECT 445.625000 222.440000 466.450000 222.670000 ;
      RECT 445.625000 222.670000 445.855000 229.450000 ;
      RECT 445.625000 232.320000 445.855000 233.700000 ;
      RECT 445.625000 233.700000 466.450000 233.930000 ;
      RECT 445.655000 200.145000 445.825000 201.280000 ;
      RECT 445.655000 206.125000 445.825000 209.620000 ;
      RECT 445.655000 211.910000 445.825000 215.230000 ;
      RECT 445.655000 219.275000 445.825000 222.440000 ;
      RECT 445.655000 229.450000 445.825000 232.320000 ;
      RECT 445.980000 194.525000 446.150000 198.525000 ;
      RECT 446.155000 237.915000 446.325000 238.980000 ;
      RECT 446.155000 247.190000 446.325000 249.900000 ;
      RECT 446.265000 200.695000 446.435000 210.545000 ;
      RECT 446.265000 211.940000 446.435000 221.790000 ;
      RECT 446.265000 223.200000 446.435000 233.050000 ;
      RECT 446.345000 237.495000 446.935000 237.665000 ;
      RECT 446.425000 237.415000 446.935000 237.495000 ;
      RECT 446.425000 237.665000 446.935000 237.745000 ;
      RECT 446.425000 250.370000 446.935000 250.700000 ;
      RECT 446.490000 210.765000 450.490000 210.935000 ;
      RECT 446.490000 222.010000 450.490000 222.180000 ;
      RECT 446.490000 233.270000 450.490000 233.440000 ;
      RECT 446.495000 237.745000 446.865000 250.370000 ;
      RECT 446.560000 194.300000 456.410000 194.470000 ;
      RECT 446.560000 198.580000 456.410000 198.750000 ;
      RECT 447.010000  54.185000 447.180000  59.445000 ;
      RECT 447.035000 238.040000 447.205000 250.205000 ;
      RECT 447.165000  97.235000 447.495000  97.305000 ;
      RECT 447.165000  97.305000 460.845000  97.675000 ;
      RECT 447.165000  97.675000 447.495000  97.745000 ;
      RECT 447.165000  98.115000 447.495000  98.185000 ;
      RECT 447.165000  98.185000 460.845000  98.555000 ;
      RECT 447.165000  98.555000 447.495000  98.625000 ;
      RECT 447.165000 110.745000 447.495000 110.815000 ;
      RECT 447.165000 110.815000 460.845000 111.185000 ;
      RECT 447.165000 111.185000 447.495000 111.255000 ;
      RECT 447.165000 111.625000 447.495000 111.695000 ;
      RECT 447.165000 111.695000 460.845000 112.065000 ;
      RECT 447.165000 112.065000 447.495000 112.135000 ;
      RECT 447.165000 124.255000 447.495000 124.325000 ;
      RECT 447.165000 124.325000 460.845000 124.695000 ;
      RECT 447.165000 124.695000 447.495000 124.765000 ;
      RECT 447.165000 125.135000 447.495000 125.205000 ;
      RECT 447.165000 125.205000 460.845000 125.575000 ;
      RECT 447.165000 125.575000 447.495000 125.645000 ;
      RECT 447.165000 137.765000 447.495000 137.835000 ;
      RECT 447.165000 137.835000 460.845000 138.205000 ;
      RECT 447.165000 138.205000 447.495000 138.275000 ;
      RECT 447.165000 138.645000 447.495000 138.715000 ;
      RECT 447.165000 138.715000 460.845000 139.085000 ;
      RECT 447.165000 139.085000 447.495000 139.155000 ;
      RECT 447.215000  91.770000 447.385000  95.390000 ;
      RECT 447.215000  97.215000 447.385000  97.235000 ;
      RECT 447.215000  98.625000 447.385000  98.645000 ;
      RECT 447.215000 100.470000 447.385000 104.090000 ;
      RECT 447.215000 105.280000 447.385000 108.900000 ;
      RECT 447.215000 110.725000 447.385000 110.745000 ;
      RECT 447.215000 112.135000 447.385000 112.155000 ;
      RECT 447.215000 113.980000 447.385000 117.600000 ;
      RECT 447.215000 118.790000 447.385000 122.410000 ;
      RECT 447.215000 124.235000 447.385000 124.255000 ;
      RECT 447.215000 125.645000 447.385000 125.665000 ;
      RECT 447.215000 127.490000 447.385000 131.110000 ;
      RECT 447.215000 132.300000 447.385000 135.920000 ;
      RECT 447.215000 137.745000 447.385000 137.765000 ;
      RECT 447.215000 139.155000 447.385000 139.175000 ;
      RECT 447.215000 141.000000 447.385000 144.620000 ;
      RECT 447.295000 237.495000 447.825000 237.665000 ;
      RECT 447.305000 237.415000 447.815000 237.495000 ;
      RECT 447.305000 237.665000 447.815000 237.745000 ;
      RECT 447.305000 250.370000 447.815000 250.700000 ;
      RECT 447.375000 237.745000 447.745000 246.105000 ;
      RECT 447.375000 246.105000 447.905000 246.275000 ;
      RECT 447.375000 246.275000 447.745000 250.370000 ;
      RECT 447.425000  53.540000 447.595000  60.015000 ;
      RECT 447.665000  96.965000 460.350000  97.135000 ;
      RECT 447.665000  97.845000 448.715000  98.015000 ;
      RECT 447.665000  98.725000 460.350000  98.895000 ;
      RECT 447.665000 110.475000 460.350000 110.645000 ;
      RECT 447.665000 111.355000 448.715000 111.525000 ;
      RECT 447.665000 112.235000 460.350000 112.405000 ;
      RECT 447.665000 123.985000 460.350000 124.155000 ;
      RECT 447.665000 124.865000 448.715000 125.035000 ;
      RECT 447.665000 125.745000 460.350000 125.915000 ;
      RECT 447.665000 137.495000 460.350000 137.665000 ;
      RECT 447.665000 138.375000 448.715000 138.545000 ;
      RECT 447.665000 139.255000 460.350000 139.425000 ;
      RECT 447.710000  39.285000 450.130000  52.425000 ;
      RECT 447.725000  24.750000 477.515000  24.755000 ;
      RECT 447.755000  96.230000 449.145000  96.400000 ;
      RECT 447.755000  99.460000 449.145000  99.630000 ;
      RECT 447.755000 109.740000 449.145000 109.910000 ;
      RECT 447.755000 112.970000 449.145000 113.140000 ;
      RECT 447.755000 123.250000 449.145000 123.420000 ;
      RECT 447.755000 126.480000 449.145000 126.650000 ;
      RECT 447.755000 136.760000 449.145000 136.930000 ;
      RECT 447.755000 139.990000 449.145000 140.160000 ;
      RECT 447.765000  91.345000 460.045000  91.915000 ;
      RECT 447.765000  92.125000 460.045000  92.695000 ;
      RECT 447.765000  92.905000 460.045000  93.475000 ;
      RECT 447.765000  93.685000 460.045000  94.255000 ;
      RECT 447.765000  94.465000 460.045000  95.035000 ;
      RECT 447.765000  95.245000 460.045000  95.815000 ;
      RECT 447.765000 100.045000 460.045000 100.615000 ;
      RECT 447.765000 100.825000 460.045000 101.395000 ;
      RECT 447.765000 101.605000 460.045000 102.175000 ;
      RECT 447.765000 102.385000 460.045000 102.955000 ;
      RECT 447.765000 103.165000 460.045000 103.735000 ;
      RECT 447.765000 103.945000 460.045000 104.515000 ;
      RECT 447.765000 104.855000 460.045000 105.425000 ;
      RECT 447.765000 105.635000 460.045000 106.205000 ;
      RECT 447.765000 106.415000 460.045000 106.985000 ;
      RECT 447.765000 107.195000 460.045000 107.765000 ;
      RECT 447.765000 107.975000 460.045000 108.545000 ;
      RECT 447.765000 108.755000 460.045000 109.325000 ;
      RECT 447.765000 113.555000 460.045000 114.125000 ;
      RECT 447.765000 114.335000 460.045000 114.905000 ;
      RECT 447.765000 115.115000 460.045000 115.685000 ;
      RECT 447.765000 115.895000 460.045000 116.465000 ;
      RECT 447.765000 116.675000 460.045000 117.245000 ;
      RECT 447.765000 117.455000 460.045000 118.025000 ;
      RECT 447.765000 118.365000 460.045000 118.935000 ;
      RECT 447.765000 119.145000 460.045000 119.715000 ;
      RECT 447.765000 119.925000 460.045000 120.495000 ;
      RECT 447.765000 120.705000 460.045000 121.275000 ;
      RECT 447.765000 121.485000 460.045000 122.055000 ;
      RECT 447.765000 122.265000 460.045000 122.835000 ;
      RECT 447.765000 127.065000 460.045000 127.635000 ;
      RECT 447.765000 127.845000 460.045000 128.415000 ;
      RECT 447.765000 128.625000 460.045000 129.195000 ;
      RECT 447.765000 129.405000 460.045000 129.975000 ;
      RECT 447.765000 130.185000 460.045000 130.755000 ;
      RECT 447.765000 130.965000 460.045000 131.535000 ;
      RECT 447.765000 131.875000 460.045000 132.445000 ;
      RECT 447.765000 132.655000 460.045000 133.225000 ;
      RECT 447.765000 133.435000 460.045000 134.005000 ;
      RECT 447.765000 134.215000 460.045000 134.785000 ;
      RECT 447.765000 134.995000 460.045000 135.565000 ;
      RECT 447.765000 135.775000 460.045000 136.345000 ;
      RECT 447.765000 140.575000 460.045000 141.145000 ;
      RECT 447.765000 141.355000 460.045000 141.925000 ;
      RECT 447.765000 142.135000 460.045000 142.705000 ;
      RECT 447.765000 142.915000 460.045000 143.485000 ;
      RECT 447.765000 143.695000 460.045000 144.265000 ;
      RECT 447.765000 144.475000 460.045000 145.045000 ;
      RECT 447.915000 237.915000 448.085000 239.240000 ;
      RECT 447.915000 239.240000 449.245000 239.750000 ;
      RECT 447.915000 247.190000 448.085000 249.900000 ;
      RECT 448.085000  15.745000 448.615000  15.915000 ;
      RECT 448.150000  13.335000 451.050000  13.585000 ;
      RECT 448.150000  17.370000 451.040000  17.925000 ;
      RECT 448.150000  17.925000 451.220000  18.175000 ;
      RECT 448.160000  13.585000 451.040000  14.040000 ;
      RECT 448.160000  17.200000 451.040000  17.370000 ;
      RECT 448.275000  14.040000 448.605000  15.335000 ;
      RECT 448.285000  15.505000 448.615000  15.745000 ;
      RECT 448.285000  15.915000 448.615000  15.985000 ;
      RECT 448.295000  16.155000 448.545000  17.200000 ;
      RECT 448.340000 146.920000 448.510000 181.625000 ;
      RECT 448.535000 237.915000 448.705000 238.965000 ;
      RECT 448.535000 247.190000 448.705000 249.900000 ;
      RECT 448.600000  52.425000 450.130000  61.055000 ;
      RECT 448.725000  16.155000 448.975000  16.935000 ;
      RECT 448.805000  14.395000 449.895000  15.335000 ;
      RECT 448.805000  15.335000 448.975000  16.155000 ;
      RECT 448.805000 237.415000 449.315000 237.745000 ;
      RECT 448.805000 250.370000 449.315000 250.700000 ;
      RECT 448.865000 146.880000 458.585000 147.145000 ;
      RECT 448.865000 147.800000 449.875000 147.970000 ;
      RECT 448.865000 148.680000 449.875000 148.850000 ;
      RECT 448.865000 149.560000 449.875000 149.730000 ;
      RECT 448.865000 150.385000 458.585000 150.650000 ;
      RECT 448.865000 151.310000 458.585000 151.575000 ;
      RECT 448.865000 152.230000 449.875000 152.400000 ;
      RECT 448.865000 153.110000 449.875000 153.280000 ;
      RECT 448.865000 153.990000 449.875000 154.160000 ;
      RECT 448.865000 154.815000 458.585000 155.080000 ;
      RECT 448.865000 155.740000 458.585000 156.005000 ;
      RECT 448.865000 156.660000 449.875000 156.830000 ;
      RECT 448.865000 157.540000 449.875000 157.710000 ;
      RECT 448.865000 158.420000 449.875000 158.590000 ;
      RECT 448.865000 159.245000 458.585000 159.510000 ;
      RECT 448.865000 160.170000 458.585000 160.435000 ;
      RECT 448.865000 161.090000 449.875000 161.260000 ;
      RECT 448.865000 161.970000 449.875000 162.140000 ;
      RECT 448.865000 162.850000 449.875000 163.020000 ;
      RECT 448.865000 163.675000 458.585000 163.940000 ;
      RECT 448.865000 164.600000 458.585000 164.865000 ;
      RECT 448.865000 165.520000 449.875000 165.690000 ;
      RECT 448.865000 166.400000 449.875000 166.570000 ;
      RECT 448.865000 167.280000 449.875000 167.450000 ;
      RECT 448.865000 168.105000 458.585000 168.370000 ;
      RECT 448.865000 169.030000 458.585000 169.295000 ;
      RECT 448.865000 169.950000 449.875000 170.120000 ;
      RECT 448.865000 170.830000 449.875000 171.000000 ;
      RECT 448.865000 171.710000 449.875000 171.880000 ;
      RECT 448.865000 172.535000 458.585000 172.800000 ;
      RECT 448.865000 173.460000 458.585000 173.725000 ;
      RECT 448.865000 174.380000 449.875000 174.550000 ;
      RECT 448.865000 175.260000 449.875000 175.430000 ;
      RECT 448.865000 176.140000 449.875000 176.310000 ;
      RECT 448.865000 176.965000 458.585000 177.230000 ;
      RECT 448.865000 177.890000 458.585000 178.155000 ;
      RECT 448.865000 178.810000 449.875000 178.980000 ;
      RECT 448.865000 179.690000 449.875000 179.860000 ;
      RECT 448.865000 180.570000 449.875000 180.740000 ;
      RECT 448.865000 181.395000 458.585000 181.660000 ;
      RECT 448.875000 237.745000 449.245000 239.240000 ;
      RECT 448.875000 239.750000 449.245000 250.370000 ;
      RECT 448.945000  97.845000 449.275000  98.015000 ;
      RECT 448.945000 111.355000 449.275000 111.525000 ;
      RECT 448.945000 124.865000 449.275000 125.035000 ;
      RECT 448.945000 138.375000 449.275000 138.545000 ;
      RECT 449.145000  14.305000 449.895000  14.395000 ;
      RECT 449.145000  15.505000 449.475000  15.985000 ;
      RECT 449.155000  16.155000 449.485000  17.200000 ;
      RECT 449.415000 237.915000 449.585000 250.205000 ;
      RECT 449.655000  15.335000 449.895000  15.505000 ;
      RECT 449.655000  15.505000 450.415000  15.985000 ;
      RECT 449.985000 244.735000 467.055000 246.035000 ;
      RECT 450.085000  14.040000 450.415000  15.335000 ;
      RECT 450.085000  16.155000 450.415000  17.200000 ;
      RECT 450.085000 240.120000 450.255000 242.390000 ;
      RECT 450.085000 242.390000 470.480000 244.115000 ;
      RECT 450.270000 237.965000 450.440000 238.075000 ;
      RECT 450.270000 238.075000 450.445000 238.965000 ;
      RECT 450.270000 238.965000 450.440000 238.975000 ;
      RECT 450.320000 148.060000 454.305000 148.590000 ;
      RECT 450.320000 148.965000 454.735000 149.495000 ;
      RECT 450.320000 149.675000 455.165000 150.205000 ;
      RECT 450.320000 152.490000 455.595000 153.020000 ;
      RECT 450.320000 153.395000 454.735000 153.925000 ;
      RECT 450.320000 154.105000 455.165000 154.635000 ;
      RECT 450.320000 156.920000 454.305000 157.450000 ;
      RECT 450.320000 157.825000 456.025000 158.355000 ;
      RECT 450.320000 158.535000 455.165000 159.065000 ;
      RECT 450.320000 161.350000 455.595000 161.880000 ;
      RECT 450.320000 162.255000 456.025000 162.785000 ;
      RECT 450.320000 162.965000 455.165000 163.495000 ;
      RECT 450.320000 165.780000 454.305000 166.310000 ;
      RECT 450.320000 166.685000 454.735000 167.215000 ;
      RECT 450.320000 167.395000 456.455000 167.925000 ;
      RECT 450.320000 170.210000 455.595000 170.740000 ;
      RECT 450.320000 171.115000 454.735000 171.645000 ;
      RECT 450.320000 171.825000 456.455000 172.355000 ;
      RECT 450.320000 174.640000 454.305000 175.170000 ;
      RECT 450.320000 175.545000 456.025000 176.075000 ;
      RECT 450.320000 176.255000 456.455000 176.785000 ;
      RECT 450.320000 179.070000 455.595000 179.600000 ;
      RECT 450.320000 179.975000 456.025000 180.505000 ;
      RECT 450.320000 180.685000 456.455000 181.215000 ;
      RECT 450.325000 247.250000 450.495000 250.230000 ;
      RECT 450.460000 237.545000 451.130000 237.715000 ;
      RECT 450.545000 200.695000 450.715000 210.545000 ;
      RECT 450.545000 211.940000 450.715000 221.790000 ;
      RECT 450.545000 223.200000 450.715000 233.050000 ;
      RECT 450.550000 246.265000 461.585000 246.970000 ;
      RECT 450.585000  14.305000 450.915000  16.935000 ;
      RECT 450.640000 240.720000 451.220000 242.390000 ;
      RECT 450.770000 210.765000 465.610000 210.935000 ;
      RECT 450.770000 222.010000 465.610000 222.180000 ;
      RECT 450.770000 233.270000 465.610000 233.440000 ;
      RECT 451.060000 240.300000 452.660000 240.470000 ;
      RECT 451.150000 237.965000 451.320000 238.975000 ;
      RECT 451.205000 247.520000 451.375000 250.230000 ;
      RECT 451.400000  62.475000 460.915000  62.975000 ;
      RECT 451.400000  62.975000 452.620000  78.420000 ;
      RECT 451.400000  78.420000 460.915000  78.920000 ;
      RECT 451.400000  78.920000 452.620000  86.845000 ;
      RECT 451.400000  86.845000 460.915000  89.195000 ;
      RECT 451.835000 237.935000 452.005000 239.210000 ;
      RECT 451.835000 240.720000 452.005000 241.730000 ;
      RECT 451.900000  30.235000 464.800000  30.405000 ;
      RECT 451.900000  30.405000 452.070000  46.485000 ;
      RECT 451.900000  46.485000 460.685000  46.655000 ;
      RECT 451.900000  46.655000 452.070000  62.475000 ;
      RECT 452.085000 247.250000 452.255000 250.230000 ;
      RECT 452.715000 236.365000 455.320000 238.945000 ;
      RECT 452.715000 240.720000 454.605000 242.390000 ;
      RECT 452.965000 247.520000 453.135000 250.230000 ;
      RECT 453.170000  48.385000 453.340000  53.135000 ;
      RECT 453.170000  56.125000 453.340000  60.875000 ;
      RECT 453.170000  64.575000 453.340000  69.325000 ;
      RECT 453.170000  72.085000 453.340000  76.835000 ;
      RECT 453.170000  80.535000 453.340000  85.285000 ;
      RECT 453.220000  31.915000 453.390000  36.665000 ;
      RECT 453.220000  38.695000 453.390000  43.445000 ;
      RECT 453.220000  53.485000 456.360000  53.655000 ;
      RECT 453.220000  55.605000 456.360000  55.775000 ;
      RECT 453.220000  69.675000 456.360000  69.845000 ;
      RECT 453.220000  71.565000 456.360000  71.735000 ;
      RECT 453.220000  85.635000 456.360000  85.805000 ;
      RECT 453.240000  47.705000 453.910000  47.875000 ;
      RECT 453.240000  61.385000 453.910000  61.555000 ;
      RECT 453.240000  63.895000 453.910000  64.065000 ;
      RECT 453.240000  77.345000 453.910000  77.515000 ;
      RECT 453.240000  79.855000 453.910000  80.025000 ;
      RECT 453.395000  47.000000 459.095000  47.370000 ;
      RECT 453.395000  47.370000 453.765000  47.705000 ;
      RECT 453.395000  61.555000 453.765000  61.890000 ;
      RECT 453.395000  61.890000 459.095000  62.260000 ;
      RECT 453.395000  63.190000 459.095000  63.560000 ;
      RECT 453.395000  63.560000 453.765000  63.895000 ;
      RECT 453.395000  77.515000 453.765000  77.850000 ;
      RECT 453.395000  77.850000 459.095000  78.220000 ;
      RECT 453.395000  79.150000 459.095000  79.520000 ;
      RECT 453.395000  79.520000 453.765000  79.855000 ;
      RECT 453.445000  30.785000 456.740000  30.955000 ;
      RECT 453.445000  30.955000 454.925000  31.405000 ;
      RECT 453.445000  43.955000 454.925000  44.355000 ;
      RECT 453.445000  44.355000 457.145000  44.525000 ;
      RECT 453.755000  48.415000 454.315000  48.735000 ;
      RECT 453.755000  60.525000 454.315000  60.845000 ;
      RECT 453.755000  64.605000 454.315000  64.925000 ;
      RECT 453.755000  76.485000 454.315000  76.805000 ;
      RECT 453.755000  80.565000 454.315000  80.885000 ;
      RECT 453.845000 247.250000 454.015000 250.230000 ;
      RECT 453.950000  48.385000 454.120000  48.415000 ;
      RECT 453.950000  48.735000 454.120000  53.135000 ;
      RECT 453.950000  56.125000 454.120000  60.525000 ;
      RECT 453.950000  60.845000 454.120000  60.875000 ;
      RECT 453.950000  64.575000 454.120000  64.605000 ;
      RECT 453.950000  64.925000 454.120000  69.325000 ;
      RECT 453.950000  72.085000 454.120000  76.485000 ;
      RECT 453.950000  76.805000 454.120000  76.835000 ;
      RECT 453.950000  80.535000 454.120000  80.565000 ;
      RECT 453.950000  80.885000 454.120000  85.285000 ;
      RECT 454.075000  12.275000 454.585000  15.045000 ;
      RECT 454.100000  31.915000 454.270000  36.665000 ;
      RECT 454.100000  38.695000 454.270000  43.445000 ;
      RECT 454.415000  49.575000 454.980000  49.895000 ;
      RECT 454.415000  59.365000 454.980000  59.685000 ;
      RECT 454.415000  65.765000 454.980000  66.085000 ;
      RECT 454.415000  75.325000 454.980000  75.645000 ;
      RECT 454.415000  81.725000 454.980000  82.045000 ;
      RECT 454.420000 240.300000 456.140000 240.470000 ;
      RECT 454.570000  48.385000 454.740000  49.575000 ;
      RECT 454.570000  49.895000 454.740000  53.135000 ;
      RECT 454.570000  56.125000 454.740000  59.365000 ;
      RECT 454.570000  59.685000 454.740000  60.875000 ;
      RECT 454.570000  64.575000 454.740000  65.765000 ;
      RECT 454.570000  66.085000 454.740000  69.325000 ;
      RECT 454.570000  72.085000 454.740000  75.325000 ;
      RECT 454.570000  75.645000 454.740000  76.835000 ;
      RECT 454.570000  80.535000 454.740000  81.725000 ;
      RECT 454.570000  82.045000 454.740000  85.285000 ;
      RECT 454.600000 250.310000 456.530000 250.480000 ;
      RECT 454.600000 250.480000 455.055000 251.030000 ;
      RECT 454.615000  21.090000 455.070000  21.640000 ;
      RECT 454.615000  21.640000 456.545000  21.810000 ;
      RECT 454.615000  44.710000 456.545000  44.880000 ;
      RECT 454.615000  44.880000 455.070000  45.430000 ;
      RECT 454.625000  47.705000 455.295000  47.875000 ;
      RECT 454.625000  61.385000 455.295000  61.555000 ;
      RECT 454.625000  63.895000 455.295000  64.065000 ;
      RECT 454.625000  77.345000 455.295000  77.515000 ;
      RECT 454.625000  79.855000 455.295000  80.025000 ;
      RECT 454.640000  15.535000 457.880000  15.705000 ;
      RECT 454.825000 200.695000 454.995000 210.545000 ;
      RECT 454.825000 211.940000 454.995000 221.790000 ;
      RECT 454.825000 223.200000 454.995000 233.050000 ;
      RECT 454.910000 251.380000 456.860000 251.730000 ;
      RECT 454.925000  20.390000 456.875000  20.740000 ;
      RECT 454.925000  45.780000 456.875000  46.130000 ;
      RECT 454.980000  31.915000 455.150000  36.665000 ;
      RECT 454.980000  38.695000 455.150000  43.445000 ;
      RECT 455.145000  48.415000 455.705000  48.735000 ;
      RECT 455.145000  60.525000 455.705000  60.845000 ;
      RECT 455.145000  64.605000 455.705000  64.925000 ;
      RECT 455.145000  76.485000 455.705000  76.805000 ;
      RECT 455.145000  80.565000 455.705000  80.885000 ;
      RECT 455.205000  31.235000 456.685000  31.405000 ;
      RECT 455.205000  43.955000 456.685000  44.125000 ;
      RECT 455.295000  12.275000 455.465000  14.985000 ;
      RECT 455.315000 240.720000 455.485000 241.730000 ;
      RECT 455.350000  48.385000 455.520000  48.415000 ;
      RECT 455.350000  48.735000 455.520000  53.135000 ;
      RECT 455.350000  56.125000 455.520000  60.525000 ;
      RECT 455.350000  60.845000 455.520000  60.875000 ;
      RECT 455.350000  64.575000 455.520000  64.605000 ;
      RECT 455.350000  64.925000 455.520000  69.325000 ;
      RECT 455.350000  72.085000 455.520000  76.485000 ;
      RECT 455.350000  76.805000 455.520000  76.835000 ;
      RECT 455.350000  80.535000 455.520000  80.565000 ;
      RECT 455.350000  80.885000 455.520000  85.285000 ;
      RECT 455.575000  47.705000 456.245000  47.875000 ;
      RECT 455.575000  61.385000 456.245000  61.555000 ;
      RECT 455.575000  63.895000 456.245000  64.065000 ;
      RECT 455.575000  77.345000 456.245000  77.515000 ;
      RECT 455.575000  79.855000 456.245000  80.025000 ;
      RECT 455.635000 250.665000 455.805000 251.195000 ;
      RECT 455.650000  20.925000 455.820000  21.455000 ;
      RECT 455.650000  45.065000 455.820000  45.595000 ;
      RECT 455.860000  31.915000 456.030000  36.665000 ;
      RECT 455.860000  38.695000 456.030000  43.445000 ;
      RECT 455.940000  48.995000 456.475000  49.315000 ;
      RECT 455.940000  59.945000 456.475000  60.265000 ;
      RECT 455.940000  65.185000 456.475000  65.505000 ;
      RECT 455.940000  75.905000 456.475000  76.225000 ;
      RECT 455.940000  81.145000 456.475000  81.465000 ;
      RECT 455.955000 240.720000 456.535000 242.390000 ;
      RECT 456.030000 237.935000 456.200000 238.945000 ;
      RECT 456.130000  48.385000 456.300000  48.995000 ;
      RECT 456.130000  49.315000 456.300000  53.135000 ;
      RECT 456.130000  56.125000 456.300000  59.945000 ;
      RECT 456.130000  60.265000 456.300000  60.875000 ;
      RECT 456.130000  64.575000 456.300000  65.185000 ;
      RECT 456.130000  65.505000 456.300000  69.325000 ;
      RECT 456.130000  72.085000 456.300000  75.905000 ;
      RECT 456.130000  76.225000 456.300000  76.835000 ;
      RECT 456.130000  80.535000 456.300000  81.145000 ;
      RECT 456.130000  81.465000 456.300000  85.285000 ;
      RECT 456.175000  12.275000 456.345000  14.985000 ;
      RECT 456.325000 250.700000 456.860000 251.380000 ;
      RECT 456.340000  16.735000 456.510000  19.445000 ;
      RECT 456.340000  20.740000 456.875000  21.420000 ;
      RECT 456.340000  45.100000 456.875000  45.780000 ;
      RECT 456.675000 147.360000 457.345000 147.530000 ;
      RECT 456.675000 151.790000 457.345000 151.960000 ;
      RECT 456.675000 156.220000 457.345000 156.390000 ;
      RECT 456.675000 160.650000 457.345000 160.820000 ;
      RECT 456.675000 165.080000 457.345000 165.250000 ;
      RECT 456.675000 169.510000 457.345000 169.680000 ;
      RECT 456.675000 173.940000 457.345000 174.110000 ;
      RECT 456.675000 178.370000 457.345000 178.540000 ;
      RECT 456.695000 148.625000 458.575000 148.905000 ;
      RECT 456.695000 153.055000 458.575000 153.335000 ;
      RECT 456.695000 157.485000 458.575000 157.765000 ;
      RECT 456.695000 161.915000 458.575000 162.195000 ;
      RECT 456.695000 166.345000 458.575000 166.625000 ;
      RECT 456.695000 170.775000 458.575000 171.055000 ;
      RECT 456.695000 175.205000 458.575000 175.485000 ;
      RECT 456.695000 179.635000 458.575000 179.915000 ;
      RECT 456.740000  31.855000 457.250000  36.665000 ;
      RECT 456.740000  38.695000 457.250000  43.505000 ;
      RECT 456.965000 241.810000 465.080000 241.995000 ;
      RECT 456.965000 241.995000 457.495000 242.085000 ;
      RECT 457.025000  96.205000 462.110000  96.375000 ;
      RECT 457.025000  99.485000 462.110000  99.655000 ;
      RECT 457.025000 109.715000 462.110000 109.885000 ;
      RECT 457.025000 112.995000 462.110000 113.165000 ;
      RECT 457.025000 123.225000 462.110000 123.395000 ;
      RECT 457.025000 126.505000 462.110000 126.675000 ;
      RECT 457.025000 136.735000 462.110000 136.905000 ;
      RECT 457.025000 140.015000 462.110000 140.185000 ;
      RECT 457.030000  47.675000 457.200000  47.705000 ;
      RECT 457.030000  47.705000 457.655000  47.875000 ;
      RECT 457.030000  47.875000 457.200000  52.855000 ;
      RECT 457.030000  52.855000 457.655000  53.865000 ;
      RECT 457.030000  55.395000 457.655000  56.405000 ;
      RECT 457.030000  56.405000 457.200000  61.385000 ;
      RECT 457.030000  61.385000 457.655000  61.555000 ;
      RECT 457.030000  61.555000 457.200000  61.585000 ;
      RECT 457.030000  63.865000 457.200000  63.895000 ;
      RECT 457.030000  63.895000 457.655000  64.065000 ;
      RECT 457.030000  64.065000 457.200000  69.045000 ;
      RECT 457.030000  69.045000 457.655000  70.055000 ;
      RECT 457.030000  71.355000 457.655000  72.365000 ;
      RECT 457.030000  72.365000 457.200000  77.345000 ;
      RECT 457.030000  77.345000 457.655000  77.515000 ;
      RECT 457.030000  77.515000 457.200000  77.545000 ;
      RECT 457.030000  79.825000 457.200000  79.855000 ;
      RECT 457.030000  79.855000 457.655000  80.025000 ;
      RECT 457.030000  80.025000 457.200000  85.005000 ;
      RECT 457.030000  85.005000 457.655000  86.015000 ;
      RECT 457.045000 236.190000 457.215000 238.900000 ;
      RECT 457.055000  12.275000 457.225000  14.985000 ;
      RECT 457.060000 241.450000 463.320000 241.620000 ;
      RECT 457.085000 250.780000 458.500000 251.080000 ;
      RECT 457.100000  21.040000 458.515000  21.340000 ;
      RECT 457.100000  45.180000 458.515000  45.480000 ;
      RECT 457.220000  18.195000 457.940000  19.445000 ;
      RECT 457.240000 239.450000 457.910000 239.620000 ;
      RECT 457.335000  97.845000 460.045000  98.015000 ;
      RECT 457.335000 111.355000 460.045000 111.525000 ;
      RECT 457.335000 124.865000 460.045000 125.035000 ;
      RECT 457.335000 138.375000 460.045000 138.545000 ;
      RECT 457.385000  96.165000 462.110000  96.205000 ;
      RECT 457.385000  96.375000 462.110000  96.415000 ;
      RECT 457.385000  99.445000 462.110000  99.485000 ;
      RECT 457.385000  99.655000 462.110000  99.695000 ;
      RECT 457.385000 109.675000 462.110000 109.715000 ;
      RECT 457.385000 109.885000 462.110000 109.925000 ;
      RECT 457.385000 112.955000 462.110000 112.995000 ;
      RECT 457.385000 113.165000 462.110000 113.205000 ;
      RECT 457.385000 123.185000 462.110000 123.225000 ;
      RECT 457.385000 123.395000 462.110000 123.435000 ;
      RECT 457.385000 126.465000 462.110000 126.505000 ;
      RECT 457.385000 126.675000 462.110000 126.715000 ;
      RECT 457.385000 136.695000 462.110000 136.735000 ;
      RECT 457.385000 136.905000 462.110000 136.945000 ;
      RECT 457.385000 139.975000 462.110000 140.015000 ;
      RECT 457.385000 140.185000 462.110000 140.225000 ;
      RECT 457.485000  50.590000 457.655000  51.640000 ;
      RECT 457.485000  57.620000 457.655000  58.670000 ;
      RECT 457.485000  66.780000 457.655000  67.830000 ;
      RECT 457.485000  73.580000 457.655000  74.630000 ;
      RECT 457.485000  82.740000 457.655000  83.790000 ;
      RECT 457.565000 147.745000 459.345000 148.025000 ;
      RECT 457.565000 149.505000 459.345000 149.785000 ;
      RECT 457.565000 152.175000 459.345000 152.455000 ;
      RECT 457.565000 153.935000 459.345000 154.215000 ;
      RECT 457.565000 156.605000 459.345000 156.885000 ;
      RECT 457.565000 158.365000 459.345000 158.645000 ;
      RECT 457.565000 161.035000 459.345000 161.315000 ;
      RECT 457.565000 162.795000 459.345000 163.075000 ;
      RECT 457.565000 165.465000 459.345000 165.745000 ;
      RECT 457.565000 167.225000 459.345000 167.505000 ;
      RECT 457.565000 169.895000 459.345000 170.175000 ;
      RECT 457.565000 171.655000 459.345000 171.935000 ;
      RECT 457.565000 174.325000 459.345000 174.605000 ;
      RECT 457.565000 176.085000 459.345000 176.365000 ;
      RECT 457.565000 178.755000 459.345000 179.035000 ;
      RECT 457.565000 180.515000 459.345000 180.795000 ;
      RECT 457.585000 193.220000 458.545000 197.915000 ;
      RECT 457.585000 197.915000 470.480000 198.880000 ;
      RECT 457.755000  50.090000 458.265000  50.420000 ;
      RECT 457.755000  54.035000 458.265000  54.365000 ;
      RECT 457.755000  54.895000 458.265000  55.225000 ;
      RECT 457.755000  58.840000 458.265000  59.170000 ;
      RECT 457.755000  66.280000 458.265000  66.610000 ;
      RECT 457.755000  70.225000 458.265000  70.555000 ;
      RECT 457.755000  70.855000 458.265000  71.185000 ;
      RECT 457.755000  74.800000 458.265000  75.130000 ;
      RECT 457.755000  82.240000 458.265000  82.570000 ;
      RECT 457.755000  86.185000 458.265000  86.515000 ;
      RECT 457.825000  50.420000 458.195000  51.895000 ;
      RECT 457.825000  51.895000 458.355000  52.065000 ;
      RECT 457.825000  52.290000 458.355000  52.460000 ;
      RECT 457.825000  52.460000 458.195000  54.035000 ;
      RECT 457.825000  55.225000 458.195000  56.800000 ;
      RECT 457.825000  56.800000 458.355000  56.970000 ;
      RECT 457.825000  57.195000 458.355000  57.365000 ;
      RECT 457.825000  57.365000 458.195000  58.840000 ;
      RECT 457.825000  66.610000 458.195000  68.085000 ;
      RECT 457.825000  68.085000 458.355000  68.255000 ;
      RECT 457.825000  68.480000 458.355000  68.650000 ;
      RECT 457.825000  68.650000 458.195000  70.225000 ;
      RECT 457.825000  71.185000 458.195000  72.760000 ;
      RECT 457.825000  72.760000 458.355000  72.930000 ;
      RECT 457.825000  73.155000 458.355000  73.325000 ;
      RECT 457.825000  73.325000 458.195000  74.800000 ;
      RECT 457.825000  82.570000 458.195000  84.045000 ;
      RECT 457.825000  84.045000 458.355000  84.215000 ;
      RECT 457.825000  84.440000 458.355000  84.610000 ;
      RECT 457.825000  84.610000 458.195000  86.185000 ;
      RECT 457.925000 236.190000 458.435000 236.395000 ;
      RECT 457.925000 236.395000 459.245000 238.960000 ;
      RECT 457.935000  12.275000 459.255000  15.045000 ;
      RECT 458.365000  50.590000 458.535000  51.600000 ;
      RECT 458.365000  52.815000 458.535000  53.865000 ;
      RECT 458.365000  55.395000 458.535000  56.445000 ;
      RECT 458.365000  57.660000 458.535000  58.670000 ;
      RECT 458.365000  66.780000 458.535000  67.790000 ;
      RECT 458.365000  69.005000 458.535000  70.055000 ;
      RECT 458.365000  71.355000 458.535000  72.405000 ;
      RECT 458.365000  73.620000 458.535000  74.630000 ;
      RECT 458.365000  82.740000 458.535000  83.750000 ;
      RECT 458.365000  84.965000 458.535000  86.015000 ;
      RECT 458.635000  50.090000 459.145000  50.420000 ;
      RECT 458.635000  54.035000 460.175000  54.365000 ;
      RECT 458.635000  54.895000 460.175000  55.225000 ;
      RECT 458.635000  58.840000 459.145000  59.170000 ;
      RECT 458.635000  66.280000 459.145000  66.610000 ;
      RECT 458.635000  70.225000 460.175000  70.555000 ;
      RECT 458.635000  70.855000 460.175000  71.185000 ;
      RECT 458.635000  74.800000 459.145000  75.130000 ;
      RECT 458.635000  82.240000 459.145000  82.570000 ;
      RECT 458.635000  86.185000 460.175000  86.515000 ;
      RECT 458.725000  47.370000 459.095000  50.090000 ;
      RECT 458.725000  59.170000 459.095000  61.890000 ;
      RECT 458.725000  63.560000 459.095000  66.280000 ;
      RECT 458.725000  75.130000 459.095000  77.850000 ;
      RECT 458.725000  79.520000 459.095000  82.240000 ;
      RECT 458.735000 236.190000 459.245000 236.395000 ;
      RECT 458.885000  51.895000 459.415000  52.065000 ;
      RECT 458.885000  52.290000 459.415000  52.460000 ;
      RECT 458.885000  56.800000 459.415000  56.970000 ;
      RECT 458.885000  57.195000 459.415000  57.365000 ;
      RECT 458.885000  68.085000 459.415000  68.255000 ;
      RECT 458.885000  68.480000 459.415000  68.650000 ;
      RECT 458.885000  72.760000 459.415000  72.930000 ;
      RECT 458.885000  73.155000 459.415000  73.325000 ;
      RECT 458.885000  84.045000 459.415000  84.215000 ;
      RECT 458.885000  84.440000 459.415000  84.610000 ;
      RECT 458.900000 249.430000 459.070000 252.140000 ;
      RECT 458.905000 248.710000 460.605000 248.880000 ;
      RECT 459.095000 146.730000 459.345000 147.745000 ;
      RECT 459.095000 148.025000 459.345000 149.505000 ;
      RECT 459.095000 149.785000 459.345000 150.800000 ;
      RECT 459.095000 151.160000 459.345000 152.175000 ;
      RECT 459.095000 152.455000 459.345000 153.935000 ;
      RECT 459.095000 154.215000 459.345000 155.230000 ;
      RECT 459.095000 155.590000 459.345000 156.605000 ;
      RECT 459.095000 156.885000 459.345000 158.365000 ;
      RECT 459.095000 158.645000 459.345000 159.660000 ;
      RECT 459.095000 160.020000 459.345000 161.035000 ;
      RECT 459.095000 161.315000 459.345000 162.795000 ;
      RECT 459.095000 163.075000 459.345000 164.090000 ;
      RECT 459.095000 164.450000 459.345000 165.465000 ;
      RECT 459.095000 165.745000 459.345000 167.225000 ;
      RECT 459.095000 167.505000 459.345000 168.520000 ;
      RECT 459.095000 168.880000 459.345000 169.895000 ;
      RECT 459.095000 170.175000 459.345000 171.655000 ;
      RECT 459.095000 171.935000 459.345000 172.950000 ;
      RECT 459.095000 173.310000 459.345000 174.325000 ;
      RECT 459.095000 174.605000 459.345000 176.085000 ;
      RECT 459.095000 176.365000 459.345000 177.380000 ;
      RECT 459.095000 177.740000 459.345000 178.755000 ;
      RECT 459.095000 179.035000 459.345000 180.515000 ;
      RECT 459.095000 180.795000 459.345000 181.810000 ;
      RECT 459.105000 200.695000 459.275000 210.545000 ;
      RECT 459.105000 211.940000 459.275000 221.790000 ;
      RECT 459.105000 223.200000 459.275000 233.050000 ;
      RECT 459.190000  15.535000 460.790000  15.705000 ;
      RECT 459.245000  50.590000 459.415000  51.895000 ;
      RECT 459.245000  52.460000 459.415000  53.865000 ;
      RECT 459.245000  55.395000 459.415000  56.800000 ;
      RECT 459.245000  57.365000 459.415000  58.670000 ;
      RECT 459.245000  66.780000 459.415000  68.085000 ;
      RECT 459.245000  68.650000 459.415000  70.055000 ;
      RECT 459.245000  71.355000 459.415000  72.760000 ;
      RECT 459.245000  73.325000 459.415000  74.630000 ;
      RECT 459.245000  82.740000 459.415000  84.045000 ;
      RECT 459.245000  84.610000 459.415000  86.015000 ;
      RECT 459.250000  16.735000 459.420000  19.445000 ;
      RECT 459.275000 239.450000 459.945000 239.620000 ;
      RECT 459.645000  47.175000 460.175000  47.345000 ;
      RECT 459.645000  61.915000 460.175000  62.085000 ;
      RECT 459.645000  63.365000 460.175000  63.535000 ;
      RECT 459.645000  77.875000 460.175000  78.045000 ;
      RECT 459.645000  79.325000 460.175000  79.495000 ;
      RECT 459.780000 249.430000 459.950000 252.140000 ;
      RECT 459.805000  47.170000 460.175000  47.175000 ;
      RECT 459.805000  47.345000 460.175000  54.035000 ;
      RECT 459.805000  55.225000 460.175000  61.915000 ;
      RECT 459.805000  62.085000 460.175000  62.090000 ;
      RECT 459.805000  63.360000 460.175000  63.365000 ;
      RECT 459.805000  63.535000 460.175000  70.225000 ;
      RECT 459.805000  71.185000 460.175000  77.875000 ;
      RECT 459.805000  78.045000 460.175000  78.050000 ;
      RECT 459.805000  79.320000 460.175000  79.325000 ;
      RECT 459.805000  79.495000 460.175000  86.185000 ;
      RECT 459.955000 236.190000 460.125000 238.900000 ;
      RECT 459.965000  12.275000 460.135000  14.985000 ;
      RECT 460.090000 190.715000 466.740000 196.790000 ;
      RECT 460.130000  16.675000 460.640000  18.195000 ;
      RECT 460.130000  18.195000 460.850000  19.445000 ;
      RECT 460.515000  46.655000 460.685000  62.470000 ;
      RECT 460.515000  62.470000 460.915000  62.475000 ;
      RECT 460.515000  62.975000 460.915000  78.420000 ;
      RECT 460.515000  78.920000 460.915000  86.845000 ;
      RECT 460.515000  97.235000 460.845000  97.305000 ;
      RECT 460.515000  97.675000 460.845000  97.745000 ;
      RECT 460.515000  98.115000 460.845000  98.185000 ;
      RECT 460.515000  98.555000 460.845000  98.625000 ;
      RECT 460.515000 110.745000 460.845000 110.815000 ;
      RECT 460.515000 111.185000 460.845000 111.255000 ;
      RECT 460.515000 111.625000 460.845000 111.695000 ;
      RECT 460.515000 112.065000 460.845000 112.135000 ;
      RECT 460.515000 124.255000 460.845000 124.325000 ;
      RECT 460.515000 124.695000 460.845000 124.765000 ;
      RECT 460.515000 125.135000 460.845000 125.205000 ;
      RECT 460.515000 125.575000 460.845000 125.645000 ;
      RECT 460.515000 137.765000 460.845000 137.835000 ;
      RECT 460.515000 138.205000 460.845000 138.275000 ;
      RECT 460.515000 138.645000 460.845000 138.715000 ;
      RECT 460.515000 139.085000 460.845000 139.155000 ;
      RECT 460.595000  91.770000 460.765000  95.390000 ;
      RECT 460.595000 100.470000 460.765000 104.090000 ;
      RECT 460.595000 105.280000 460.765000 108.900000 ;
      RECT 460.595000 113.980000 460.765000 117.600000 ;
      RECT 460.595000 118.790000 460.765000 122.410000 ;
      RECT 460.595000 127.490000 460.765000 131.110000 ;
      RECT 460.595000 132.300000 460.765000 135.920000 ;
      RECT 460.595000 141.000000 460.765000 144.620000 ;
      RECT 460.660000 249.370000 462.550000 252.140000 ;
      RECT 460.840000  32.985000 461.010000  33.235000 ;
      RECT 460.840000  33.235000 463.230000  33.405000 ;
      RECT 460.840000  33.405000 461.010000  33.515000 ;
      RECT 460.845000  12.275000 462.735000  15.045000 ;
      RECT 461.180000  47.605000 461.350000  48.120000 ;
      RECT 461.180000  48.120000 461.445000  51.135000 ;
      RECT 461.180000  58.125000 461.445000  61.140000 ;
      RECT 461.180000  61.140000 461.350000  61.655000 ;
      RECT 461.180000  63.795000 461.350000  64.310000 ;
      RECT 461.180000  64.310000 461.445000  67.325000 ;
      RECT 461.180000  74.085000 461.445000  77.100000 ;
      RECT 461.180000  77.100000 461.350000  77.615000 ;
      RECT 461.180000  79.755000 461.350000  80.270000 ;
      RECT 461.180000  80.270000 461.445000  83.285000 ;
      RECT 461.250000  90.055000 462.110000  96.165000 ;
      RECT 461.250000  96.415000 462.110000  99.445000 ;
      RECT 461.250000  99.695000 462.110000 109.675000 ;
      RECT 461.250000 109.925000 462.110000 112.955000 ;
      RECT 461.250000 113.205000 462.110000 123.185000 ;
      RECT 461.250000 123.435000 462.110000 126.465000 ;
      RECT 461.250000 126.715000 462.110000 136.695000 ;
      RECT 461.250000 136.945000 462.110000 139.975000 ;
      RECT 461.250000 140.225000 462.110000 145.465000 ;
      RECT 461.250000 146.460000 462.110000 182.820000 ;
      RECT 461.470000 249.250000 461.720000 249.370000 ;
      RECT 461.545000  47.625000 462.055000  47.955000 ;
      RECT 461.545000  61.305000 462.055000  61.635000 ;
      RECT 461.545000  63.815000 462.055000  64.145000 ;
      RECT 461.545000  77.265000 462.055000  77.595000 ;
      RECT 461.545000  79.775000 462.055000  80.105000 ;
      RECT 461.615000  47.955000 461.985000  52.290000 ;
      RECT 461.615000  52.290000 462.145000  52.460000 ;
      RECT 461.615000  56.800000 462.145000  56.970000 ;
      RECT 461.615000  56.970000 461.985000  61.305000 ;
      RECT 461.615000  64.145000 461.985000  68.480000 ;
      RECT 461.615000  68.480000 462.145000  68.650000 ;
      RECT 461.615000  72.760000 462.145000  72.930000 ;
      RECT 461.615000  72.930000 461.985000  77.265000 ;
      RECT 461.615000  80.105000 461.985000  84.440000 ;
      RECT 461.615000  84.440000 462.145000  84.610000 ;
      RECT 461.620000  20.655000 462.570000  21.905000 ;
      RECT 461.620000  44.615000 462.570000  45.865000 ;
      RECT 461.620000 236.190000 461.790000 240.940000 ;
      RECT 461.655000  15.045000 461.905000  15.165000 ;
      RECT 461.845000  35.415000 462.565000  36.665000 ;
      RECT 461.845000  38.695000 462.565000  39.945000 ;
      RECT 462.055000  21.905000 462.565000  23.425000 ;
      RECT 462.055000  33.895000 462.565000  35.415000 ;
      RECT 462.055000  37.215000 462.565000  38.695000 ;
      RECT 462.055000  39.945000 462.565000  39.985000 ;
      RECT 462.055000  43.095000 462.565000  44.615000 ;
      RECT 462.155000  48.425000 462.325000  51.135000 ;
      RECT 462.155000  58.125000 462.325000  60.835000 ;
      RECT 462.155000  64.615000 462.325000  67.325000 ;
      RECT 462.155000  74.085000 462.325000  76.795000 ;
      RECT 462.155000  80.575000 462.325000  83.285000 ;
      RECT 462.400000 248.710000 464.085000 248.880000 ;
      RECT 462.415000  23.915000 464.100000  24.085000 ;
      RECT 462.415000  42.435000 464.100000  42.605000 ;
      RECT 462.425000  47.625000 462.935000  47.705000 ;
      RECT 462.425000  47.705000 462.955000  47.875000 ;
      RECT 462.425000  47.875000 462.935000  47.955000 ;
      RECT 462.425000  61.305000 462.935000  61.385000 ;
      RECT 462.425000  61.385000 462.955000  61.555000 ;
      RECT 462.425000  61.555000 462.935000  61.635000 ;
      RECT 462.425000  63.815000 462.935000  63.895000 ;
      RECT 462.425000  63.895000 462.955000  64.065000 ;
      RECT 462.425000  64.065000 462.935000  64.145000 ;
      RECT 462.425000  77.265000 462.935000  77.345000 ;
      RECT 462.425000  77.345000 462.955000  77.515000 ;
      RECT 462.425000  77.515000 462.935000  77.595000 ;
      RECT 462.425000  79.775000 462.935000  79.855000 ;
      RECT 462.425000  79.855000 462.955000  80.025000 ;
      RECT 462.425000  80.025000 462.935000  80.105000 ;
      RECT 462.500000 236.190000 462.670000 240.940000 ;
      RECT 462.550000  15.535000 464.270000  15.705000 ;
      RECT 462.730000  18.195000 463.450000  19.445000 ;
      RECT 462.940000  16.675000 463.450000  18.195000 ;
      RECT 463.035000  48.120000 463.205000  52.290000 ;
      RECT 463.035000  52.290000 463.565000  52.460000 ;
      RECT 463.035000  56.800000 463.565000  56.970000 ;
      RECT 463.035000  56.970000 463.205000  61.140000 ;
      RECT 463.035000  64.310000 463.205000  68.480000 ;
      RECT 463.035000  68.480000 463.565000  68.650000 ;
      RECT 463.035000  72.760000 463.565000  72.930000 ;
      RECT 463.035000  72.930000 463.205000  77.100000 ;
      RECT 463.035000  80.270000 463.205000  84.440000 ;
      RECT 463.035000  84.440000 463.565000  84.610000 ;
      RECT 463.220000  87.055000 466.740000 185.105000 ;
      RECT 463.260000 249.430000 463.430000 252.140000 ;
      RECT 463.275000  20.655000 463.445000  23.365000 ;
      RECT 463.275000  33.955000 463.445000  36.665000 ;
      RECT 463.275000  37.215000 463.445000  39.925000 ;
      RECT 463.275000  43.155000 463.445000  45.865000 ;
      RECT 463.380000 236.190000 463.550000 240.940000 ;
      RECT 463.385000 200.695000 463.555000 210.545000 ;
      RECT 463.385000 211.940000 463.555000 221.790000 ;
      RECT 463.385000 223.200000 463.555000 233.050000 ;
      RECT 463.445000  12.275000 463.615000  14.985000 ;
      RECT 463.600000 241.450000 465.080000 241.810000 ;
      RECT 464.140000 249.430000 464.310000 252.140000 ;
      RECT 464.155000  20.655000 464.325000  23.365000 ;
      RECT 464.155000  43.095000 464.800000  45.865000 ;
      RECT 464.160000  16.735000 464.330000  19.445000 ;
      RECT 464.260000 236.190000 464.430000 240.940000 ;
      RECT 464.325000  12.275000 464.495000  14.985000 ;
      RECT 464.360000  46.880000 467.360000  47.345000 ;
      RECT 464.360000  47.345000 466.130000  87.055000 ;
      RECT 464.630000  30.405000 464.800000  43.095000 ;
      RECT 464.720000 247.445000 465.160000 252.495000 ;
      RECT 465.140000 236.190000 465.650000 241.000000 ;
      RECT 465.560000  29.000000 477.515000  45.815000 ;
      RECT 465.560000  45.815000 467.360000  46.880000 ;
      RECT 465.665000 200.695000 465.835000 210.545000 ;
      RECT 465.665000 211.940000 465.835000 221.790000 ;
      RECT 465.665000 223.200000 465.835000 233.050000 ;
      RECT 466.045000 246.035000 467.055000 253.445000 ;
      RECT 466.220000 200.145000 466.450000 211.185000 ;
      RECT 466.220000 211.415000 466.450000 222.440000 ;
      RECT 466.220000 222.670000 466.450000 233.700000 ;
      RECT 466.845000  47.705000 467.375000  47.875000 ;
      RECT 466.845000  61.385000 467.375000  61.555000 ;
      RECT 466.845000  63.895000 467.375000  64.065000 ;
      RECT 466.845000  77.345000 467.375000  77.515000 ;
      RECT 466.845000  79.855000 467.375000  80.025000 ;
      RECT 466.925000  51.500000 467.455000  51.670000 ;
      RECT 466.925000  57.590000 467.455000  57.760000 ;
      RECT 466.925000  67.690000 467.455000  67.860000 ;
      RECT 466.925000  73.550000 467.455000  73.720000 ;
      RECT 466.925000  83.650000 467.455000  83.820000 ;
      RECT 467.085000   0.130000 477.515000   0.300000 ;
      RECT 467.085000  11.240000 477.515000  24.750000 ;
      RECT 467.205000  47.875000 467.375000  48.120000 ;
      RECT 467.205000  48.120000 467.455000  51.500000 ;
      RECT 467.205000  57.760000 467.455000  61.140000 ;
      RECT 467.205000  61.140000 467.375000  61.385000 ;
      RECT 467.205000  64.065000 467.375000  64.310000 ;
      RECT 467.205000  64.310000 467.455000  67.690000 ;
      RECT 467.205000  73.720000 467.455000  77.100000 ;
      RECT 467.205000  77.100000 467.375000  77.345000 ;
      RECT 467.205000  80.025000 467.375000  80.270000 ;
      RECT 467.205000  80.270000 467.455000  83.650000 ;
      RECT 467.245000  52.225000 469.100000  52.475000 ;
      RECT 467.245000  56.785000 469.100000  57.035000 ;
      RECT 467.245000  68.415000 469.100000  68.665000 ;
      RECT 467.245000  72.745000 469.100000  72.995000 ;
      RECT 467.245000  84.375000 469.100000  84.625000 ;
      RECT 467.450000 198.880000 470.480000 234.950000 ;
      RECT 467.480000 235.180000 470.480000 242.390000 ;
      RECT 467.555000  47.625000 468.065000  47.955000 ;
      RECT 467.555000  61.305000 468.065000  61.635000 ;
      RECT 467.555000  63.815000 468.065000  64.145000 ;
      RECT 467.555000  77.265000 468.065000  77.595000 ;
      RECT 467.555000  79.775000 468.065000  80.105000 ;
      RECT 467.625000  47.955000 467.995000  51.950000 ;
      RECT 467.625000  57.310000 467.995000  61.305000 ;
      RECT 467.625000  64.145000 467.995000  68.140000 ;
      RECT 467.625000  73.270000 467.995000  77.265000 ;
      RECT 467.625000  80.105000 467.995000  84.100000 ;
      RECT 467.820000 244.115000 470.480000 253.385000 ;
      RECT 467.850000  88.840000 470.480000 197.915000 ;
      RECT 467.980000  88.770000 470.480000  88.840000 ;
      RECT 468.165000  48.235000 468.615000  52.225000 ;
      RECT 468.165000  57.035000 468.615000  61.025000 ;
      RECT 468.165000  64.425000 468.615000  68.415000 ;
      RECT 468.165000  72.995000 468.615000  76.985000 ;
      RECT 468.165000  80.385000 468.615000  84.375000 ;
      RECT 468.415000  46.665000 468.945000  47.705000 ;
      RECT 468.415000  61.555000 468.945000  62.595000 ;
      RECT 468.415000  62.855000 468.945000  63.895000 ;
      RECT 468.415000  77.515000 468.945000  78.555000 ;
      RECT 468.415000  78.815000 468.945000  79.855000 ;
      RECT 468.435000  47.705000 468.945000  47.955000 ;
      RECT 468.435000  61.305000 468.945000  61.555000 ;
      RECT 468.435000  63.895000 468.945000  64.145000 ;
      RECT 468.435000  77.265000 468.945000  77.515000 ;
      RECT 468.435000  79.855000 468.945000  80.105000 ;
      RECT 468.850000  52.475000 469.100000  53.485000 ;
      RECT 468.850000  53.485000 471.420000  53.735000 ;
      RECT 468.850000  55.525000 471.420000  55.775000 ;
      RECT 468.850000  55.775000 469.100000  56.785000 ;
      RECT 468.850000  68.665000 469.100000  69.675000 ;
      RECT 468.850000  69.675000 471.420000  69.925000 ;
      RECT 468.850000  71.485000 471.420000  71.735000 ;
      RECT 468.850000  71.735000 469.100000  72.745000 ;
      RECT 468.850000  84.625000 469.100000  85.635000 ;
      RECT 468.850000  85.635000 471.420000  85.885000 ;
      RECT 469.045000  48.120000 469.215000  51.950000 ;
      RECT 469.045000  57.310000 469.215000  61.140000 ;
      RECT 469.045000  64.310000 469.215000  68.140000 ;
      RECT 469.045000  73.270000 469.215000  77.100000 ;
      RECT 469.045000  80.270000 469.215000  84.100000 ;
      RECT 469.485000  48.995000 470.045000  49.315000 ;
      RECT 469.485000  59.945000 470.045000  60.265000 ;
      RECT 469.485000  65.185000 470.045000  65.505000 ;
      RECT 469.485000  75.905000 470.045000  76.225000 ;
      RECT 469.485000  81.145000 470.045000  81.465000 ;
      RECT 469.650000  48.385000 469.820000  48.995000 ;
      RECT 469.650000  49.315000 469.820000  53.135000 ;
      RECT 469.650000  56.125000 469.820000  59.945000 ;
      RECT 469.650000  60.265000 469.820000  60.875000 ;
      RECT 469.650000  64.575000 469.820000  65.185000 ;
      RECT 469.650000  65.505000 469.820000  69.325000 ;
      RECT 469.650000  72.085000 469.820000  75.905000 ;
      RECT 469.650000  76.225000 469.820000  76.835000 ;
      RECT 469.650000  80.535000 469.820000  81.145000 ;
      RECT 469.650000  81.465000 469.820000  85.285000 ;
      RECT 469.705000  47.705000 470.375000  47.875000 ;
      RECT 469.705000  61.385000 470.375000  61.555000 ;
      RECT 469.705000  63.895000 470.375000  64.065000 ;
      RECT 469.705000  77.345000 470.375000  77.515000 ;
      RECT 469.705000  79.855000 470.375000  80.025000 ;
      RECT 470.200000  48.415000 470.760000  48.735000 ;
      RECT 470.200000  60.525000 470.760000  60.845000 ;
      RECT 470.200000  64.605000 470.760000  64.925000 ;
      RECT 470.200000  76.485000 470.760000  76.805000 ;
      RECT 470.200000  80.565000 470.760000  80.885000 ;
      RECT 470.430000  48.385000 470.600000  48.415000 ;
      RECT 470.430000  48.735000 470.600000  53.135000 ;
      RECT 470.430000  56.125000 470.600000  60.525000 ;
      RECT 470.430000  60.845000 470.600000  60.875000 ;
      RECT 470.430000  64.575000 470.600000  64.605000 ;
      RECT 470.430000  64.925000 470.600000  69.325000 ;
      RECT 470.430000  72.085000 470.600000  76.485000 ;
      RECT 470.430000  76.805000 470.600000  76.835000 ;
      RECT 470.430000  80.535000 470.600000  80.565000 ;
      RECT 470.430000  80.885000 470.600000  85.285000 ;
      RECT 470.655000  47.705000 471.325000  47.875000 ;
      RECT 470.655000  61.385000 471.325000  61.555000 ;
      RECT 470.655000  63.895000 471.325000  64.065000 ;
      RECT 470.655000  77.345000 471.325000  77.515000 ;
      RECT 470.655000  79.855000 471.325000  80.025000 ;
      RECT 470.735000  46.665000 471.265000  47.705000 ;
      RECT 470.735000  61.555000 471.265000  62.595000 ;
      RECT 470.735000  62.855000 471.265000  63.895000 ;
      RECT 470.735000  77.515000 471.265000  78.555000 ;
      RECT 470.735000  78.815000 471.265000  79.855000 ;
      RECT 471.210000  48.385000 471.380000  53.135000 ;
      RECT 471.210000  56.125000 471.380000  60.875000 ;
      RECT 471.210000  64.575000 471.380000  69.325000 ;
      RECT 471.210000  72.085000 471.380000  76.835000 ;
      RECT 471.210000  80.535000 471.380000  85.285000 ;
      RECT 471.245000  88.295000 477.515000 253.585000 ;
      RECT 472.255000  45.815000 477.515000  88.295000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 480.000000 253.715000 ;
    LAYER met2 ;
      RECT   0.000000   0.000000  84.980000  30.825000 ;
      RECT   0.000000   0.000000  84.980000  33.515000 ;
      RECT   0.000000   0.000000  85.120000  30.685000 ;
      RECT   0.000000  30.685000  86.105000  33.375000 ;
      RECT   0.000000  30.825000  85.965000  33.515000 ;
      RECT   0.000000  30.825000  85.965000  45.365000 ;
      RECT   0.000000  33.375000 109.675000  36.470000 ;
      RECT   0.000000  33.515000 109.535000  36.525000 ;
      RECT   0.000000  33.515000 109.535000  45.365000 ;
      RECT   0.000000  36.470000 109.695000  36.490000 ;
      RECT   0.000000  36.490000 109.695000  45.420000 ;
      RECT   0.000000  36.525000 109.535000  36.535000 ;
      RECT   0.000000  36.525000 109.535000  36.535000 ;
      RECT   0.000000  36.535000 109.545000  36.545000 ;
      RECT   0.000000  36.535000 109.545000  36.545000 ;
      RECT   0.000000  36.545000 109.555000  45.365000 ;
      RECT   0.000000  45.365000 109.485000  45.435000 ;
      RECT   0.000000  45.365000 109.485000  45.435000 ;
      RECT   0.000000  45.420000 109.325000  45.790000 ;
      RECT   0.000000  45.435000 109.415000  45.505000 ;
      RECT   0.000000  45.435000 109.415000  45.505000 ;
      RECT   0.000000  45.505000 109.345000  45.575000 ;
      RECT   0.000000  45.505000 109.345000  45.575000 ;
      RECT   0.000000  45.575000 109.275000  45.645000 ;
      RECT   0.000000  45.575000 109.275000  45.645000 ;
      RECT   0.000000  45.645000 109.205000  45.715000 ;
      RECT   0.000000  45.645000 109.205000  45.715000 ;
      RECT   0.000000  45.715000 109.185000  45.735000 ;
      RECT   0.000000  45.715000 109.185000  45.735000 ;
      RECT   0.000000  45.735000 109.185000  46.450000 ;
      RECT   0.000000  45.790000 109.325000  46.505000 ;
      RECT   0.000000  46.450000 109.115000  46.520000 ;
      RECT   0.000000  46.450000 109.115000  46.520000 ;
      RECT   0.000000  46.505000 108.430000  47.400000 ;
      RECT   0.000000  46.520000 109.045000  46.590000 ;
      RECT   0.000000  46.520000 109.045000  46.590000 ;
      RECT   0.000000  46.590000 108.975000  46.660000 ;
      RECT   0.000000  46.590000 108.975000  46.660000 ;
      RECT   0.000000  46.660000 108.905000  46.730000 ;
      RECT   0.000000  46.660000 108.905000  46.730000 ;
      RECT   0.000000  46.730000 108.835000  46.800000 ;
      RECT   0.000000  46.730000 108.835000  46.800000 ;
      RECT   0.000000  46.800000 108.765000  46.870000 ;
      RECT   0.000000  46.800000 108.765000  46.870000 ;
      RECT   0.000000  46.870000 108.695000  46.940000 ;
      RECT   0.000000  46.870000 108.695000  46.940000 ;
      RECT   0.000000  46.940000 108.625000  47.010000 ;
      RECT   0.000000  46.940000 108.625000  47.010000 ;
      RECT   0.000000  47.010000 108.555000  47.080000 ;
      RECT   0.000000  47.010000 108.555000  47.080000 ;
      RECT   0.000000  47.080000 108.485000  47.150000 ;
      RECT   0.000000  47.080000 108.485000  47.150000 ;
      RECT   0.000000  47.150000 108.415000  47.220000 ;
      RECT   0.000000  47.150000 108.415000  47.220000 ;
      RECT   0.000000  47.220000 108.345000  47.290000 ;
      RECT   0.000000  47.220000 108.345000  47.290000 ;
      RECT   0.000000  47.290000 108.290000  47.345000 ;
      RECT   0.000000  47.290000 108.290000  47.345000 ;
      RECT   0.000000  47.345000 108.290000  74.765000 ;
      RECT   0.000000  47.400000 108.430000  56.625000 ;
      RECT   0.000000  56.625000 109.240000  57.435000 ;
      RECT   0.000000  56.680000 108.290000  56.750000 ;
      RECT   0.000000  56.680000 108.290000  56.750000 ;
      RECT   0.000000  56.750000 108.360000  56.820000 ;
      RECT   0.000000  56.750000 108.360000  56.820000 ;
      RECT   0.000000  56.820000 108.430000  56.890000 ;
      RECT   0.000000  56.820000 108.430000  56.890000 ;
      RECT   0.000000  56.890000 108.500000  56.960000 ;
      RECT   0.000000  56.890000 108.500000  56.960000 ;
      RECT   0.000000  56.960000 108.570000  57.030000 ;
      RECT   0.000000  56.960000 108.570000  57.030000 ;
      RECT   0.000000  57.030000 108.640000  57.100000 ;
      RECT   0.000000  57.030000 108.640000  57.100000 ;
      RECT   0.000000  57.100000 108.710000  57.170000 ;
      RECT   0.000000  57.100000 108.710000  57.170000 ;
      RECT   0.000000  57.170000 108.780000  57.240000 ;
      RECT   0.000000  57.170000 108.780000  57.240000 ;
      RECT   0.000000  57.240000 108.850000  57.310000 ;
      RECT   0.000000  57.240000 108.850000  57.310000 ;
      RECT   0.000000  57.310000 108.920000  57.380000 ;
      RECT   0.000000  57.310000 108.920000  57.380000 ;
      RECT   0.000000  57.380000 108.990000  57.450000 ;
      RECT   0.000000  57.380000 108.990000  57.450000 ;
      RECT   0.000000  57.435000 109.240000  74.820000 ;
      RECT   0.000000  57.450000 109.060000  57.490000 ;
      RECT   0.000000  57.450000 109.060000  57.490000 ;
      RECT   0.000000  57.490000 109.100000  74.765000 ;
      RECT   0.000000  74.765000 109.030000  74.835000 ;
      RECT   0.000000  74.765000 109.030000  74.835000 ;
      RECT   0.000000  74.820000 107.610000  76.450000 ;
      RECT   0.000000  74.835000 108.960000  74.905000 ;
      RECT   0.000000  74.835000 108.960000  74.905000 ;
      RECT   0.000000  74.905000 108.890000  74.975000 ;
      RECT   0.000000  74.905000 108.890000  74.975000 ;
      RECT   0.000000  74.975000 108.820000  75.045000 ;
      RECT   0.000000  74.975000 108.820000  75.045000 ;
      RECT   0.000000  75.045000 108.750000  75.115000 ;
      RECT   0.000000  75.045000 108.750000  75.115000 ;
      RECT   0.000000  75.115000 108.680000  75.185000 ;
      RECT   0.000000  75.115000 108.680000  75.185000 ;
      RECT   0.000000  75.185000 108.610000  75.255000 ;
      RECT   0.000000  75.185000 108.610000  75.255000 ;
      RECT   0.000000  75.255000 108.540000  75.325000 ;
      RECT   0.000000  75.255000 108.540000  75.325000 ;
      RECT   0.000000  75.325000 108.470000  75.395000 ;
      RECT   0.000000  75.325000 108.470000  75.395000 ;
      RECT   0.000000  75.395000 108.400000  75.465000 ;
      RECT   0.000000  75.395000 108.400000  75.465000 ;
      RECT   0.000000  75.465000 108.330000  75.535000 ;
      RECT   0.000000  75.465000 108.330000  75.535000 ;
      RECT   0.000000  75.535000 108.260000  75.605000 ;
      RECT   0.000000  75.535000 108.260000  75.605000 ;
      RECT   0.000000  75.605000 108.190000  75.675000 ;
      RECT   0.000000  75.605000 108.190000  75.675000 ;
      RECT   0.000000  75.675000 108.120000  75.745000 ;
      RECT   0.000000  75.675000 108.120000  75.745000 ;
      RECT   0.000000  75.745000 108.050000  75.815000 ;
      RECT   0.000000  75.745000 108.050000  75.815000 ;
      RECT   0.000000  75.815000 107.980000  75.885000 ;
      RECT   0.000000  75.815000 107.980000  75.885000 ;
      RECT   0.000000  75.885000 107.910000  75.955000 ;
      RECT   0.000000  75.885000 107.910000  75.955000 ;
      RECT   0.000000  75.955000 107.840000  76.025000 ;
      RECT   0.000000  75.955000 107.840000  76.025000 ;
      RECT   0.000000  76.025000 107.770000  76.095000 ;
      RECT   0.000000  76.025000 107.770000  76.095000 ;
      RECT   0.000000  76.095000 107.700000  76.165000 ;
      RECT   0.000000  76.095000 107.700000  76.165000 ;
      RECT   0.000000  76.165000 107.630000  76.235000 ;
      RECT   0.000000  76.165000 107.630000  76.235000 ;
      RECT   0.000000  76.235000 107.560000  76.305000 ;
      RECT   0.000000  76.235000 107.560000  76.305000 ;
      RECT   0.000000  76.305000 107.490000  76.375000 ;
      RECT   0.000000  76.305000 107.490000  76.375000 ;
      RECT   0.000000  76.375000 107.470000  76.395000 ;
      RECT   0.000000  76.375000 107.470000  76.395000 ;
      RECT   0.000000  76.395000 107.470000  87.425000 ;
      RECT   0.000000  76.450000 107.610000  87.480000 ;
      RECT   0.000000  87.425000 107.400000  87.495000 ;
      RECT   0.000000  87.425000 107.400000  87.495000 ;
      RECT   0.000000  87.480000 105.670000  89.420000 ;
      RECT   0.000000  87.495000 107.330000  87.565000 ;
      RECT   0.000000  87.495000 107.330000  87.565000 ;
      RECT   0.000000  87.565000 107.260000  87.635000 ;
      RECT   0.000000  87.565000 107.260000  87.635000 ;
      RECT   0.000000  87.635000 107.190000  87.705000 ;
      RECT   0.000000  87.635000 107.190000  87.705000 ;
      RECT   0.000000  87.705000 107.120000  87.775000 ;
      RECT   0.000000  87.705000 107.120000  87.775000 ;
      RECT   0.000000  87.775000 107.050000  87.845000 ;
      RECT   0.000000  87.775000 107.050000  87.845000 ;
      RECT   0.000000  87.845000 106.980000  87.915000 ;
      RECT   0.000000  87.845000 106.980000  87.915000 ;
      RECT   0.000000  87.915000 106.910000  87.985000 ;
      RECT   0.000000  87.915000 106.910000  87.985000 ;
      RECT   0.000000  87.985000 106.840000  88.055000 ;
      RECT   0.000000  87.985000 106.840000  88.055000 ;
      RECT   0.000000  88.055000 106.770000  88.125000 ;
      RECT   0.000000  88.055000 106.770000  88.125000 ;
      RECT   0.000000  88.125000 106.700000  88.195000 ;
      RECT   0.000000  88.125000 106.700000  88.195000 ;
      RECT   0.000000  88.195000 106.630000  88.265000 ;
      RECT   0.000000  88.195000 106.630000  88.265000 ;
      RECT   0.000000  88.265000 106.560000  88.335000 ;
      RECT   0.000000  88.265000 106.560000  88.335000 ;
      RECT   0.000000  88.335000 106.490000  88.405000 ;
      RECT   0.000000  88.335000 106.490000  88.405000 ;
      RECT   0.000000  88.405000 106.420000  88.475000 ;
      RECT   0.000000  88.405000 106.420000  88.475000 ;
      RECT   0.000000  88.475000 106.350000  88.545000 ;
      RECT   0.000000  88.475000 106.350000  88.545000 ;
      RECT   0.000000  88.545000 106.280000  88.615000 ;
      RECT   0.000000  88.545000 106.280000  88.615000 ;
      RECT   0.000000  88.615000 106.210000  88.685000 ;
      RECT   0.000000  88.615000 106.210000  88.685000 ;
      RECT   0.000000  88.685000 106.140000  88.755000 ;
      RECT   0.000000  88.685000 106.140000  88.755000 ;
      RECT   0.000000  88.755000 106.070000  88.825000 ;
      RECT   0.000000  88.755000 106.070000  88.825000 ;
      RECT   0.000000  88.825000 106.000000  88.895000 ;
      RECT   0.000000  88.825000 106.000000  88.895000 ;
      RECT   0.000000  88.895000 105.930000  88.965000 ;
      RECT   0.000000  88.895000 105.930000  88.965000 ;
      RECT   0.000000  88.965000 105.860000  89.035000 ;
      RECT   0.000000  88.965000 105.860000  89.035000 ;
      RECT   0.000000  89.035000 105.790000  89.105000 ;
      RECT   0.000000  89.035000 105.790000  89.105000 ;
      RECT   0.000000  89.105000 105.720000  89.175000 ;
      RECT   0.000000  89.105000 105.720000  89.175000 ;
      RECT   0.000000  89.175000 105.650000  89.245000 ;
      RECT   0.000000  89.175000 105.650000  89.245000 ;
      RECT   0.000000  89.245000 105.580000  89.315000 ;
      RECT   0.000000  89.245000 105.580000  89.315000 ;
      RECT   0.000000  89.315000 105.530000  89.365000 ;
      RECT   0.000000  89.315000 105.530000  89.365000 ;
      RECT   0.000000  89.365000 105.530000  94.050000 ;
      RECT   0.000000  89.420000 105.670000  94.105000 ;
      RECT   0.000000  94.050000 105.460000  94.120000 ;
      RECT   0.000000  94.050000 105.460000  94.120000 ;
      RECT   0.000000  94.105000 105.215000  94.560000 ;
      RECT   0.000000  94.120000 105.390000  94.190000 ;
      RECT   0.000000  94.120000 105.390000  94.190000 ;
      RECT   0.000000  94.190000 105.320000  94.260000 ;
      RECT   0.000000  94.190000 105.320000  94.260000 ;
      RECT   0.000000  94.260000 105.250000  94.330000 ;
      RECT   0.000000  94.260000 105.250000  94.330000 ;
      RECT   0.000000  94.330000 105.180000  94.400000 ;
      RECT   0.000000  94.330000 105.180000  94.400000 ;
      RECT   0.000000  94.400000 105.160000  94.420000 ;
      RECT   0.000000  94.400000 105.160000  94.420000 ;
      RECT   0.000000  94.420000 100.405000  94.490000 ;
      RECT   0.000000  94.420000 100.405000  94.490000 ;
      RECT   0.000000  94.490000 100.335000  94.560000 ;
      RECT   0.000000  94.490000 100.335000  94.560000 ;
      RECT   0.000000  94.560000  92.165000 102.925000 ;
      RECT   0.000000  94.560000 100.265000  94.630000 ;
      RECT   0.000000  94.560000 100.265000  94.630000 ;
      RECT   0.000000  94.630000 100.195000  94.700000 ;
      RECT   0.000000  94.630000 100.195000  94.700000 ;
      RECT   0.000000  94.700000 100.125000  94.770000 ;
      RECT   0.000000  94.700000 100.125000  94.770000 ;
      RECT   0.000000  94.770000 100.055000  94.840000 ;
      RECT   0.000000  94.770000 100.055000  94.840000 ;
      RECT   0.000000  94.840000  99.985000  94.910000 ;
      RECT   0.000000  94.840000  99.985000  94.910000 ;
      RECT   0.000000  94.910000  99.915000  94.980000 ;
      RECT   0.000000  94.910000  99.915000  94.980000 ;
      RECT   0.000000  94.980000  99.845000  95.050000 ;
      RECT   0.000000  94.980000  99.845000  95.050000 ;
      RECT   0.000000  95.050000  99.775000  95.120000 ;
      RECT   0.000000  95.050000  99.775000  95.120000 ;
      RECT   0.000000  95.120000  99.705000  95.190000 ;
      RECT   0.000000  95.120000  99.705000  95.190000 ;
      RECT   0.000000  95.190000  99.635000  95.260000 ;
      RECT   0.000000  95.190000  99.635000  95.260000 ;
      RECT   0.000000  95.260000  99.565000  95.330000 ;
      RECT   0.000000  95.260000  99.565000  95.330000 ;
      RECT   0.000000  95.330000  99.495000  95.400000 ;
      RECT   0.000000  95.330000  99.495000  95.400000 ;
      RECT   0.000000  95.400000  99.425000  95.470000 ;
      RECT   0.000000  95.400000  99.425000  95.470000 ;
      RECT   0.000000  95.470000  99.355000  95.540000 ;
      RECT   0.000000  95.470000  99.355000  95.540000 ;
      RECT   0.000000  95.540000  99.285000  95.610000 ;
      RECT   0.000000  95.540000  99.285000  95.610000 ;
      RECT   0.000000  95.610000  99.215000  95.680000 ;
      RECT   0.000000  95.610000  99.215000  95.680000 ;
      RECT   0.000000  95.680000  99.145000  95.750000 ;
      RECT   0.000000  95.680000  99.145000  95.750000 ;
      RECT   0.000000  95.750000  99.075000  95.820000 ;
      RECT   0.000000  95.750000  99.075000  95.820000 ;
      RECT   0.000000  95.820000  99.005000  95.890000 ;
      RECT   0.000000  95.820000  99.005000  95.890000 ;
      RECT   0.000000  95.890000  98.935000  95.960000 ;
      RECT   0.000000  95.890000  98.935000  95.960000 ;
      RECT   0.000000  95.960000  98.865000  96.030000 ;
      RECT   0.000000  95.960000  98.865000  96.030000 ;
      RECT   0.000000  96.030000  98.795000  96.100000 ;
      RECT   0.000000  96.030000  98.795000  96.100000 ;
      RECT   0.000000  96.100000  98.725000  96.170000 ;
      RECT   0.000000  96.100000  98.725000  96.170000 ;
      RECT   0.000000  96.170000  98.655000  96.240000 ;
      RECT   0.000000  96.170000  98.655000  96.240000 ;
      RECT   0.000000  96.240000  98.585000  96.310000 ;
      RECT   0.000000  96.240000  98.585000  96.310000 ;
      RECT   0.000000  96.310000  98.515000  96.380000 ;
      RECT   0.000000  96.310000  98.515000  96.380000 ;
      RECT   0.000000  96.380000  98.445000  96.450000 ;
      RECT   0.000000  96.380000  98.445000  96.450000 ;
      RECT   0.000000  96.450000  98.375000  96.520000 ;
      RECT   0.000000  96.450000  98.375000  96.520000 ;
      RECT   0.000000  96.520000  98.305000  96.590000 ;
      RECT   0.000000  96.520000  98.305000  96.590000 ;
      RECT   0.000000  96.590000  98.235000  96.660000 ;
      RECT   0.000000  96.590000  98.235000  96.660000 ;
      RECT   0.000000  96.660000  98.165000  96.730000 ;
      RECT   0.000000  96.660000  98.165000  96.730000 ;
      RECT   0.000000  96.730000  98.095000  96.800000 ;
      RECT   0.000000  96.730000  98.095000  96.800000 ;
      RECT   0.000000  96.800000  98.025000  96.870000 ;
      RECT   0.000000  96.800000  98.025000  96.870000 ;
      RECT   0.000000  96.870000  97.955000  96.940000 ;
      RECT   0.000000  96.870000  97.955000  96.940000 ;
      RECT   0.000000  96.940000  97.885000  97.010000 ;
      RECT   0.000000  96.940000  97.885000  97.010000 ;
      RECT   0.000000  97.010000  97.815000  97.080000 ;
      RECT   0.000000  97.010000  97.815000  97.080000 ;
      RECT   0.000000  97.080000  97.745000  97.150000 ;
      RECT   0.000000  97.080000  97.745000  97.150000 ;
      RECT   0.000000  97.150000  97.675000  97.220000 ;
      RECT   0.000000  97.150000  97.675000  97.220000 ;
      RECT   0.000000  97.220000  97.605000  97.290000 ;
      RECT   0.000000  97.220000  97.605000  97.290000 ;
      RECT   0.000000  97.290000  97.535000  97.360000 ;
      RECT   0.000000  97.290000  97.535000  97.360000 ;
      RECT   0.000000  97.360000  97.465000  97.430000 ;
      RECT   0.000000  97.360000  97.465000  97.430000 ;
      RECT   0.000000  97.430000  97.395000  97.500000 ;
      RECT   0.000000  97.430000  97.395000  97.500000 ;
      RECT   0.000000  97.500000  97.325000  97.570000 ;
      RECT   0.000000  97.500000  97.325000  97.570000 ;
      RECT   0.000000  97.570000  97.255000  97.640000 ;
      RECT   0.000000  97.570000  97.255000  97.640000 ;
      RECT   0.000000  97.640000  97.185000  97.710000 ;
      RECT   0.000000  97.640000  97.185000  97.710000 ;
      RECT   0.000000  97.710000  97.115000  97.780000 ;
      RECT   0.000000  97.710000  97.115000  97.780000 ;
      RECT   0.000000  97.780000  97.045000  97.850000 ;
      RECT   0.000000  97.780000  97.045000  97.850000 ;
      RECT   0.000000  97.850000  96.975000  97.920000 ;
      RECT   0.000000  97.850000  96.975000  97.920000 ;
      RECT   0.000000  97.920000  96.905000  97.990000 ;
      RECT   0.000000  97.920000  96.905000  97.990000 ;
      RECT   0.000000  97.990000  96.835000  98.060000 ;
      RECT   0.000000  97.990000  96.835000  98.060000 ;
      RECT   0.000000  98.060000  96.765000  98.130000 ;
      RECT   0.000000  98.060000  96.765000  98.130000 ;
      RECT   0.000000  98.130000  96.695000  98.200000 ;
      RECT   0.000000  98.130000  96.695000  98.200000 ;
      RECT   0.000000  98.200000  96.625000  98.270000 ;
      RECT   0.000000  98.200000  96.625000  98.270000 ;
      RECT   0.000000  98.270000  96.555000  98.340000 ;
      RECT   0.000000  98.270000  96.555000  98.340000 ;
      RECT   0.000000  98.340000  96.485000  98.410000 ;
      RECT   0.000000  98.340000  96.485000  98.410000 ;
      RECT   0.000000  98.410000  96.415000  98.480000 ;
      RECT   0.000000  98.410000  96.415000  98.480000 ;
      RECT   0.000000  98.480000  96.345000  98.550000 ;
      RECT   0.000000  98.480000  96.345000  98.550000 ;
      RECT   0.000000  98.550000  96.275000  98.620000 ;
      RECT   0.000000  98.550000  96.275000  98.620000 ;
      RECT   0.000000  98.620000  96.205000  98.690000 ;
      RECT   0.000000  98.620000  96.205000  98.690000 ;
      RECT   0.000000  98.690000  96.135000  98.760000 ;
      RECT   0.000000  98.690000  96.135000  98.760000 ;
      RECT   0.000000  98.760000  96.065000  98.830000 ;
      RECT   0.000000  98.760000  96.065000  98.830000 ;
      RECT   0.000000  98.830000  95.995000  98.900000 ;
      RECT   0.000000  98.830000  95.995000  98.900000 ;
      RECT   0.000000  98.900000  95.925000  98.970000 ;
      RECT   0.000000  98.900000  95.925000  98.970000 ;
      RECT   0.000000  98.970000  95.855000  99.040000 ;
      RECT   0.000000  98.970000  95.855000  99.040000 ;
      RECT   0.000000  99.040000  95.785000  99.110000 ;
      RECT   0.000000  99.040000  95.785000  99.110000 ;
      RECT   0.000000  99.110000  95.715000  99.180000 ;
      RECT   0.000000  99.110000  95.715000  99.180000 ;
      RECT   0.000000  99.180000  95.645000  99.250000 ;
      RECT   0.000000  99.180000  95.645000  99.250000 ;
      RECT   0.000000  99.250000  95.575000  99.320000 ;
      RECT   0.000000  99.250000  95.575000  99.320000 ;
      RECT   0.000000  99.320000  95.505000  99.390000 ;
      RECT   0.000000  99.320000  95.505000  99.390000 ;
      RECT   0.000000  99.390000  95.435000  99.460000 ;
      RECT   0.000000  99.390000  95.435000  99.460000 ;
      RECT   0.000000  99.460000  95.365000  99.530000 ;
      RECT   0.000000  99.460000  95.365000  99.530000 ;
      RECT   0.000000  99.530000  95.295000  99.600000 ;
      RECT   0.000000  99.530000  95.295000  99.600000 ;
      RECT   0.000000  99.600000  95.225000  99.670000 ;
      RECT   0.000000  99.600000  95.225000  99.670000 ;
      RECT   0.000000  99.670000  95.155000  99.740000 ;
      RECT   0.000000  99.670000  95.155000  99.740000 ;
      RECT   0.000000  99.740000  95.085000  99.810000 ;
      RECT   0.000000  99.740000  95.085000  99.810000 ;
      RECT   0.000000  99.810000  95.015000  99.880000 ;
      RECT   0.000000  99.810000  95.015000  99.880000 ;
      RECT   0.000000  99.880000  94.945000  99.950000 ;
      RECT   0.000000  99.880000  94.945000  99.950000 ;
      RECT   0.000000  99.950000  94.875000 100.020000 ;
      RECT   0.000000  99.950000  94.875000 100.020000 ;
      RECT   0.000000 100.020000  94.805000 100.090000 ;
      RECT   0.000000 100.020000  94.805000 100.090000 ;
      RECT   0.000000 100.090000  94.735000 100.160000 ;
      RECT   0.000000 100.090000  94.735000 100.160000 ;
      RECT   0.000000 100.160000  94.665000 100.230000 ;
      RECT   0.000000 100.160000  94.665000 100.230000 ;
      RECT   0.000000 100.230000  94.595000 100.300000 ;
      RECT   0.000000 100.230000  94.595000 100.300000 ;
      RECT   0.000000 100.300000  94.525000 100.370000 ;
      RECT   0.000000 100.300000  94.525000 100.370000 ;
      RECT   0.000000 100.370000  94.455000 100.440000 ;
      RECT   0.000000 100.370000  94.455000 100.440000 ;
      RECT   0.000000 100.440000  94.385000 100.510000 ;
      RECT   0.000000 100.440000  94.385000 100.510000 ;
      RECT   0.000000 100.510000  94.315000 100.580000 ;
      RECT   0.000000 100.510000  94.315000 100.580000 ;
      RECT   0.000000 100.580000  94.245000 100.650000 ;
      RECT   0.000000 100.580000  94.245000 100.650000 ;
      RECT   0.000000 100.650000  94.175000 100.720000 ;
      RECT   0.000000 100.650000  94.175000 100.720000 ;
      RECT   0.000000 100.720000  94.105000 100.790000 ;
      RECT   0.000000 100.720000  94.105000 100.790000 ;
      RECT   0.000000 100.790000  94.035000 100.860000 ;
      RECT   0.000000 100.790000  94.035000 100.860000 ;
      RECT   0.000000 100.860000  93.965000 100.930000 ;
      RECT   0.000000 100.860000  93.965000 100.930000 ;
      RECT   0.000000 100.930000  93.895000 101.000000 ;
      RECT   0.000000 100.930000  93.895000 101.000000 ;
      RECT   0.000000 101.000000  93.825000 101.070000 ;
      RECT   0.000000 101.000000  93.825000 101.070000 ;
      RECT   0.000000 101.070000  93.755000 101.140000 ;
      RECT   0.000000 101.070000  93.755000 101.140000 ;
      RECT   0.000000 101.140000  93.685000 101.210000 ;
      RECT   0.000000 101.140000  93.685000 101.210000 ;
      RECT   0.000000 101.210000  93.615000 101.280000 ;
      RECT   0.000000 101.210000  93.615000 101.280000 ;
      RECT   0.000000 101.280000  93.545000 101.350000 ;
      RECT   0.000000 101.280000  93.545000 101.350000 ;
      RECT   0.000000 101.350000  93.475000 101.420000 ;
      RECT   0.000000 101.350000  93.475000 101.420000 ;
      RECT   0.000000 101.420000  93.405000 101.490000 ;
      RECT   0.000000 101.420000  93.405000 101.490000 ;
      RECT   0.000000 101.490000  93.335000 101.560000 ;
      RECT   0.000000 101.490000  93.335000 101.560000 ;
      RECT   0.000000 101.560000  93.265000 101.630000 ;
      RECT   0.000000 101.560000  93.265000 101.630000 ;
      RECT   0.000000 101.630000  93.195000 101.700000 ;
      RECT   0.000000 101.630000  93.195000 101.700000 ;
      RECT   0.000000 101.700000  93.125000 101.770000 ;
      RECT   0.000000 101.700000  93.125000 101.770000 ;
      RECT   0.000000 101.770000  93.055000 101.840000 ;
      RECT   0.000000 101.770000  93.055000 101.840000 ;
      RECT   0.000000 101.840000  92.985000 101.910000 ;
      RECT   0.000000 101.840000  92.985000 101.910000 ;
      RECT   0.000000 101.910000  92.915000 101.980000 ;
      RECT   0.000000 101.910000  92.915000 101.980000 ;
      RECT   0.000000 101.980000  92.845000 102.050000 ;
      RECT   0.000000 101.980000  92.845000 102.050000 ;
      RECT   0.000000 102.050000  92.775000 102.120000 ;
      RECT   0.000000 102.050000  92.775000 102.120000 ;
      RECT   0.000000 102.120000  92.705000 102.190000 ;
      RECT   0.000000 102.120000  92.705000 102.190000 ;
      RECT   0.000000 102.190000  92.635000 102.260000 ;
      RECT   0.000000 102.190000  92.635000 102.260000 ;
      RECT   0.000000 102.260000  92.565000 102.330000 ;
      RECT   0.000000 102.260000  92.565000 102.330000 ;
      RECT   0.000000 102.330000  92.495000 102.400000 ;
      RECT   0.000000 102.330000  92.495000 102.400000 ;
      RECT   0.000000 102.400000  92.425000 102.470000 ;
      RECT   0.000000 102.400000  92.425000 102.470000 ;
      RECT   0.000000 102.470000  92.355000 102.540000 ;
      RECT   0.000000 102.470000  92.355000 102.540000 ;
      RECT   0.000000 102.540000  92.285000 102.610000 ;
      RECT   0.000000 102.540000  92.285000 102.610000 ;
      RECT   0.000000 102.610000  92.215000 102.680000 ;
      RECT   0.000000 102.610000  92.215000 102.680000 ;
      RECT   0.000000 102.680000  92.145000 102.750000 ;
      RECT   0.000000 102.680000  92.145000 102.750000 ;
      RECT   0.000000 102.750000  92.075000 102.820000 ;
      RECT   0.000000 102.750000  92.075000 102.820000 ;
      RECT   0.000000 102.820000  92.025000 102.870000 ;
      RECT   0.000000 102.820000  92.025000 102.870000 ;
      RECT   0.000000 102.870000  92.025000 112.420000 ;
      RECT   0.000000 102.925000  92.165000 111.660000 ;
      RECT   0.000000 111.660000  92.405000 111.900000 ;
      RECT   0.000000 111.715000  92.025000 111.785000 ;
      RECT   0.000000 111.715000  92.025000 111.785000 ;
      RECT   0.000000 111.785000  92.095000 111.855000 ;
      RECT   0.000000 111.785000  92.095000 111.855000 ;
      RECT   0.000000 111.855000  92.165000 111.925000 ;
      RECT   0.000000 111.855000  92.165000 111.925000 ;
      RECT   0.000000 111.900000  92.945000 111.960000 ;
      RECT   0.000000 111.925000  92.235000 111.995000 ;
      RECT   0.000000 111.925000  92.235000 111.995000 ;
      RECT   0.000000 111.960000  92.945000 112.280000 ;
      RECT   0.000000 111.995000  92.305000 112.040000 ;
      RECT   0.000000 111.995000  92.305000 112.040000 ;
      RECT   0.000000 112.280000 446.945000 244.130000 ;
      RECT   0.000000 112.420000 446.640000 253.715000 ;
      RECT   0.000000 112.420000 446.805000 244.075000 ;
      RECT   0.000000 244.075000 446.640000 253.715000 ;
      RECT   0.000000 244.075000 446.640000 253.715000 ;
      RECT   0.000000 244.075000 446.640000 253.715000 ;
      RECT   0.000000 244.075000 446.735000 244.145000 ;
      RECT   0.000000 244.075000 446.735000 244.145000 ;
      RECT   0.000000 244.130000 446.780000 244.295000 ;
      RECT   0.000000 244.145000 446.665000 244.215000 ;
      RECT   0.000000 244.145000 446.665000 244.215000 ;
      RECT   0.000000 244.215000 446.640000 244.240000 ;
      RECT   0.000000 244.215000 446.640000 244.240000 ;
      RECT   0.000000 244.240000 446.640000 244.895000 ;
      RECT   0.000000 244.295000 446.780000 244.755000 ;
      RECT   0.000000 244.755000 447.605000 245.155000 ;
      RECT   0.000000 244.895000 447.465000 245.295000 ;
      RECT   0.000000 244.895000 447.465000 253.715000 ;
      RECT   0.000000 244.895000 447.465000 253.715000 ;
      RECT   0.000000 244.895000 447.465000 253.715000 ;
      RECT   0.000000 244.895000 447.465000 253.715000 ;
      RECT   0.000000 245.155000 448.355000 245.555000 ;
      RECT   0.000000 245.295000 448.215000 245.695000 ;
      RECT   0.000000 245.295000 448.215000 253.715000 ;
      RECT   0.000000 245.295000 448.215000 253.715000 ;
      RECT   0.000000 245.295000 448.215000 253.715000 ;
      RECT   0.000000 245.295000 448.215000 253.715000 ;
      RECT   0.000000 245.555000 449.105000 245.955000 ;
      RECT   0.000000 245.695000 448.965000 246.095000 ;
      RECT   0.000000 245.695000 448.965000 253.715000 ;
      RECT   0.000000 245.695000 448.965000 253.715000 ;
      RECT   0.000000 245.695000 448.965000 253.715000 ;
      RECT   0.000000 245.695000 448.965000 253.715000 ;
      RECT   0.000000 245.955000 480.000000 253.715000 ;
      RECT   0.000000 246.095000 480.000000 253.715000 ;
      RECT  87.235000   0.000000 106.570000   1.410000 ;
      RECT  87.235000   1.410000 107.285000   2.125000 ;
      RECT  87.235000   2.125000 107.285000  18.295000 ;
      RECT  87.235000  18.295000 109.675000  33.375000 ;
      RECT  87.375000   0.000000 106.430000   1.465000 ;
      RECT  87.375000   1.465000 106.430000   1.535000 ;
      RECT  87.375000   1.465000 106.430000   1.535000 ;
      RECT  87.375000   1.535000 106.500000   1.605000 ;
      RECT  87.375000   1.535000 106.500000   1.605000 ;
      RECT  87.375000   1.605000 106.570000   1.675000 ;
      RECT  87.375000   1.605000 106.570000   1.675000 ;
      RECT  87.375000   1.675000 106.640000   1.745000 ;
      RECT  87.375000   1.675000 106.640000   1.745000 ;
      RECT  87.375000   1.745000 106.710000   1.815000 ;
      RECT  87.375000   1.745000 106.710000   1.815000 ;
      RECT  87.375000   1.815000 106.780000   1.885000 ;
      RECT  87.375000   1.815000 106.780000   1.885000 ;
      RECT  87.375000   1.885000 106.850000   1.955000 ;
      RECT  87.375000   1.885000 106.850000   1.955000 ;
      RECT  87.375000   1.955000 106.920000   2.025000 ;
      RECT  87.375000   1.955000 106.920000   2.025000 ;
      RECT  87.375000   2.025000 106.990000   2.095000 ;
      RECT  87.375000   2.025000 106.990000   2.095000 ;
      RECT  87.375000   2.095000 107.060000   2.165000 ;
      RECT  87.375000   2.095000 107.060000   2.165000 ;
      RECT  87.375000   2.165000 107.130000   2.180000 ;
      RECT  87.375000   2.165000 107.130000   2.180000 ;
      RECT  87.375000   2.180000 107.145000   2.280000 ;
      RECT  87.375000   2.280000 107.200000  18.435000 ;
      RECT  87.375000  18.435000 109.535000  33.515000 ;
      RECT  87.375000  18.435000 109.535000  45.365000 ;
      RECT  89.800000 112.040000  92.805000 112.420000 ;
      RECT  92.735000 103.125000 297.270000 111.315000 ;
      RECT  92.735000 111.315000 297.225000 111.360000 ;
      RECT  92.875000 103.180000 297.130000 111.220000 ;
      RECT  92.905000 103.150000 297.100000 103.180000 ;
      RECT  92.905000 103.150000 297.100000 103.180000 ;
      RECT  92.975000 103.080000 297.030000 103.150000 ;
      RECT  92.975000 103.080000 297.030000 103.150000 ;
      RECT  93.045000 103.010000 296.960000 103.080000 ;
      RECT  93.045000 103.010000 296.960000 103.080000 ;
      RECT  93.115000 102.940000 296.890000 103.010000 ;
      RECT  93.115000 102.940000 296.890000 103.010000 ;
      RECT  93.185000 102.870000 296.820000 102.940000 ;
      RECT  93.185000 102.870000 296.820000 102.940000 ;
      RECT  93.255000 102.800000 296.750000 102.870000 ;
      RECT  93.255000 102.800000 296.750000 102.870000 ;
      RECT  93.325000 102.730000 296.680000 102.800000 ;
      RECT  93.325000 102.730000 296.680000 102.800000 ;
      RECT  93.395000 102.660000 296.610000 102.730000 ;
      RECT  93.395000 102.660000 296.610000 102.730000 ;
      RECT  93.465000 102.590000 296.540000 102.660000 ;
      RECT  93.465000 102.590000 296.540000 102.660000 ;
      RECT  93.485000 111.360000 296.520000 112.280000 ;
      RECT  93.535000 102.520000 296.470000 102.590000 ;
      RECT  93.535000 102.520000 296.470000 102.590000 ;
      RECT  93.605000 102.450000 296.400000 102.520000 ;
      RECT  93.605000 102.450000 296.400000 102.520000 ;
      RECT  93.625000 111.220000 296.380000 112.420000 ;
      RECT  93.675000 102.380000 296.330000 102.450000 ;
      RECT  93.675000 102.380000 296.330000 102.450000 ;
      RECT  93.745000 102.310000 296.260000 102.380000 ;
      RECT  93.745000 102.310000 296.260000 102.380000 ;
      RECT  93.815000 102.240000 296.190000 102.310000 ;
      RECT  93.815000 102.240000 296.190000 102.310000 ;
      RECT  93.885000 102.170000 296.120000 102.240000 ;
      RECT  93.885000 102.170000 296.120000 102.240000 ;
      RECT  93.955000 102.100000 296.050000 102.170000 ;
      RECT  93.955000 102.100000 296.050000 102.170000 ;
      RECT  94.025000 102.030000 295.980000 102.100000 ;
      RECT  94.025000 102.030000 295.980000 102.100000 ;
      RECT  94.095000 101.960000 295.910000 102.030000 ;
      RECT  94.095000 101.960000 295.910000 102.030000 ;
      RECT  94.165000 101.890000 295.840000 101.960000 ;
      RECT  94.165000 101.890000 295.840000 101.960000 ;
      RECT  94.235000 101.820000 295.770000 101.890000 ;
      RECT  94.235000 101.820000 295.770000 101.890000 ;
      RECT  94.305000 101.750000 295.700000 101.820000 ;
      RECT  94.305000 101.750000 295.700000 101.820000 ;
      RECT  94.375000 101.680000 295.630000 101.750000 ;
      RECT  94.375000 101.680000 295.630000 101.750000 ;
      RECT  94.445000 101.610000 295.560000 101.680000 ;
      RECT  94.445000 101.610000 295.560000 101.680000 ;
      RECT  94.515000 101.540000 295.490000 101.610000 ;
      RECT  94.515000 101.540000 295.490000 101.610000 ;
      RECT  94.585000 101.470000 295.420000 101.540000 ;
      RECT  94.585000 101.470000 295.420000 101.540000 ;
      RECT  94.655000 101.400000 295.350000 101.470000 ;
      RECT  94.655000 101.400000 295.350000 101.470000 ;
      RECT  94.725000 101.330000 295.280000 101.400000 ;
      RECT  94.725000 101.330000 295.280000 101.400000 ;
      RECT  94.795000 101.260000 295.210000 101.330000 ;
      RECT  94.795000 101.260000 295.210000 101.330000 ;
      RECT  94.865000 101.190000 295.140000 101.260000 ;
      RECT  94.865000 101.190000 295.140000 101.260000 ;
      RECT  94.935000 101.120000 295.070000 101.190000 ;
      RECT  94.935000 101.120000 295.070000 101.190000 ;
      RECT  95.005000 101.050000 295.000000 101.120000 ;
      RECT  95.005000 101.050000 295.000000 101.120000 ;
      RECT  95.075000 100.980000 294.930000 101.050000 ;
      RECT  95.075000 100.980000 294.930000 101.050000 ;
      RECT  95.145000 100.910000 294.860000 100.980000 ;
      RECT  95.145000 100.910000 294.860000 100.980000 ;
      RECT  95.215000 100.840000 294.790000 100.910000 ;
      RECT  95.215000 100.840000 294.790000 100.910000 ;
      RECT  95.285000 100.770000 294.720000 100.840000 ;
      RECT  95.285000 100.770000 294.720000 100.840000 ;
      RECT  95.355000 100.700000 294.650000 100.770000 ;
      RECT  95.355000 100.700000 294.650000 100.770000 ;
      RECT  95.425000 100.630000 294.580000 100.700000 ;
      RECT  95.425000 100.630000 294.580000 100.700000 ;
      RECT  95.495000 100.560000 294.510000 100.630000 ;
      RECT  95.495000 100.560000 294.510000 100.630000 ;
      RECT  95.565000 100.490000 294.440000 100.560000 ;
      RECT  95.565000 100.490000 294.440000 100.560000 ;
      RECT  95.635000 100.420000 294.370000 100.490000 ;
      RECT  95.635000 100.420000 294.370000 100.490000 ;
      RECT  95.705000 100.350000 294.300000 100.420000 ;
      RECT  95.705000 100.350000 294.300000 100.420000 ;
      RECT  95.775000 100.280000 294.230000 100.350000 ;
      RECT  95.775000 100.280000 294.230000 100.350000 ;
      RECT  95.845000 100.210000 294.160000 100.280000 ;
      RECT  95.845000 100.210000 294.160000 100.280000 ;
      RECT  95.915000 100.140000 294.090000 100.210000 ;
      RECT  95.915000 100.140000 294.090000 100.210000 ;
      RECT  95.985000 100.070000 294.020000 100.140000 ;
      RECT  95.985000 100.070000 294.020000 100.140000 ;
      RECT  96.055000 100.000000 293.950000 100.070000 ;
      RECT  96.055000 100.000000 293.950000 100.070000 ;
      RECT  96.125000  99.930000 293.880000 100.000000 ;
      RECT  96.125000  99.930000 293.880000 100.000000 ;
      RECT  96.195000  99.860000 293.810000  99.930000 ;
      RECT  96.195000  99.860000 293.810000  99.930000 ;
      RECT  96.265000  99.790000 293.740000  99.860000 ;
      RECT  96.265000  99.790000 293.740000  99.860000 ;
      RECT  96.335000  99.720000 293.670000  99.790000 ;
      RECT  96.335000  99.720000 293.670000  99.790000 ;
      RECT  96.405000  99.650000 293.600000  99.720000 ;
      RECT  96.405000  99.650000 293.600000  99.720000 ;
      RECT  96.475000  99.580000 293.530000  99.650000 ;
      RECT  96.475000  99.580000 293.530000  99.650000 ;
      RECT  96.545000  99.510000 293.460000  99.580000 ;
      RECT  96.545000  99.510000 293.460000  99.580000 ;
      RECT  96.615000  99.440000 293.390000  99.510000 ;
      RECT  96.615000  99.440000 293.390000  99.510000 ;
      RECT  96.685000  99.370000 293.320000  99.440000 ;
      RECT  96.685000  99.370000 293.320000  99.440000 ;
      RECT  96.755000  99.300000 293.250000  99.370000 ;
      RECT  96.755000  99.300000 293.250000  99.370000 ;
      RECT  96.825000  99.230000 293.180000  99.300000 ;
      RECT  96.825000  99.230000 293.180000  99.300000 ;
      RECT  96.895000  99.160000 293.110000  99.230000 ;
      RECT  96.895000  99.160000 293.110000  99.230000 ;
      RECT  96.965000  99.090000 293.040000  99.160000 ;
      RECT  96.965000  99.090000 293.040000  99.160000 ;
      RECT  97.035000  99.020000 292.970000  99.090000 ;
      RECT  97.035000  99.020000 292.970000  99.090000 ;
      RECT  97.105000  98.950000 292.900000  99.020000 ;
      RECT  97.105000  98.950000 292.900000  99.020000 ;
      RECT  97.175000  98.880000 292.830000  98.950000 ;
      RECT  97.175000  98.880000 292.830000  98.950000 ;
      RECT  97.245000  98.810000 292.760000  98.880000 ;
      RECT  97.245000  98.810000 292.760000  98.880000 ;
      RECT  97.315000  98.740000 292.690000  98.810000 ;
      RECT  97.315000  98.740000 292.690000  98.810000 ;
      RECT  97.385000  98.670000 292.620000  98.740000 ;
      RECT  97.385000  98.670000 292.620000  98.740000 ;
      RECT  97.455000  98.600000 292.550000  98.670000 ;
      RECT  97.455000  98.600000 292.550000  98.670000 ;
      RECT  97.525000  98.530000 292.480000  98.600000 ;
      RECT  97.525000  98.530000 292.480000  98.600000 ;
      RECT  97.595000  98.460000 292.410000  98.530000 ;
      RECT  97.595000  98.460000 292.410000  98.530000 ;
      RECT  97.665000  98.390000 292.340000  98.460000 ;
      RECT  97.665000  98.390000 292.340000  98.460000 ;
      RECT  97.735000  98.320000 292.270000  98.390000 ;
      RECT  97.735000  98.320000 292.270000  98.390000 ;
      RECT  97.805000  98.250000 292.200000  98.320000 ;
      RECT  97.805000  98.250000 292.200000  98.320000 ;
      RECT  97.875000  98.180000 292.130000  98.250000 ;
      RECT  97.875000  98.180000 292.130000  98.250000 ;
      RECT  97.945000  98.110000 292.060000  98.180000 ;
      RECT  97.945000  98.110000 292.060000  98.180000 ;
      RECT  98.015000  98.040000 291.990000  98.110000 ;
      RECT  98.015000  98.040000 291.990000  98.110000 ;
      RECT  98.085000  97.970000 291.920000  98.040000 ;
      RECT  98.085000  97.970000 291.920000  98.040000 ;
      RECT  98.155000  97.900000 291.850000  97.970000 ;
      RECT  98.155000  97.900000 291.850000  97.970000 ;
      RECT  98.225000  97.830000 291.780000  97.900000 ;
      RECT  98.225000  97.830000 291.780000  97.900000 ;
      RECT  98.295000  97.760000 291.710000  97.830000 ;
      RECT  98.295000  97.760000 291.710000  97.830000 ;
      RECT  98.365000  97.690000 291.640000  97.760000 ;
      RECT  98.365000  97.690000 291.640000  97.760000 ;
      RECT  98.435000  97.620000 291.570000  97.690000 ;
      RECT  98.435000  97.620000 291.570000  97.690000 ;
      RECT  98.505000  97.550000 291.500000  97.620000 ;
      RECT  98.505000  97.550000 291.500000  97.620000 ;
      RECT  98.575000  97.480000 291.430000  97.550000 ;
      RECT  98.575000  97.480000 291.430000  97.550000 ;
      RECT  98.645000  97.410000 291.360000  97.480000 ;
      RECT  98.645000  97.410000 291.360000  97.480000 ;
      RECT  98.715000  97.340000 291.290000  97.410000 ;
      RECT  98.715000  97.340000 291.290000  97.410000 ;
      RECT  98.785000  97.270000 291.220000  97.340000 ;
      RECT  98.785000  97.270000 291.220000  97.340000 ;
      RECT  98.855000  97.200000 291.150000  97.270000 ;
      RECT  98.855000  97.200000 291.150000  97.270000 ;
      RECT  98.925000  97.130000 291.080000  97.200000 ;
      RECT  98.925000  97.130000 291.080000  97.200000 ;
      RECT  98.995000  97.060000 291.010000  97.130000 ;
      RECT  98.995000  97.060000 291.010000  97.130000 ;
      RECT  99.065000  96.990000 290.940000  97.060000 ;
      RECT  99.065000  96.990000 290.940000  97.060000 ;
      RECT  99.135000  96.920000 290.870000  96.990000 ;
      RECT  99.135000  96.920000 290.870000  96.990000 ;
      RECT  99.205000  96.850000 290.800000  96.920000 ;
      RECT  99.205000  96.850000 290.800000  96.920000 ;
      RECT  99.275000  96.780000 290.730000  96.850000 ;
      RECT  99.275000  96.780000 290.730000  96.850000 ;
      RECT  99.345000  96.710000 290.660000  96.780000 ;
      RECT  99.345000  96.710000 290.660000  96.780000 ;
      RECT  99.415000  96.640000 290.590000  96.710000 ;
      RECT  99.415000  96.640000 290.590000  96.710000 ;
      RECT  99.485000  96.570000 290.520000  96.640000 ;
      RECT  99.485000  96.570000 290.520000  96.640000 ;
      RECT  99.555000  96.500000 290.450000  96.570000 ;
      RECT  99.555000  96.500000 290.450000  96.570000 ;
      RECT  99.625000  96.430000 290.380000  96.500000 ;
      RECT  99.625000  96.430000 290.380000  96.500000 ;
      RECT  99.695000  96.360000 290.310000  96.430000 ;
      RECT  99.695000  96.360000 290.310000  96.430000 ;
      RECT  99.765000  96.290000 290.240000  96.360000 ;
      RECT  99.765000  96.290000 290.240000  96.360000 ;
      RECT  99.835000  96.220000 290.170000  96.290000 ;
      RECT  99.835000  96.220000 290.170000  96.290000 ;
      RECT  99.905000  96.150000 290.100000  96.220000 ;
      RECT  99.905000  96.150000 290.100000  96.220000 ;
      RECT  99.975000  96.080000 290.030000  96.150000 ;
      RECT  99.975000  96.080000 290.030000  96.150000 ;
      RECT 100.045000  96.010000 289.960000  96.080000 ;
      RECT 100.045000  96.010000 289.960000  96.080000 ;
      RECT 100.115000  95.940000 289.890000  96.010000 ;
      RECT 100.115000  95.940000 289.890000  96.010000 ;
      RECT 100.185000  95.870000 289.820000  95.940000 ;
      RECT 100.185000  95.870000 289.820000  95.940000 ;
      RECT 100.255000  95.800000 289.750000  95.870000 ;
      RECT 100.255000  95.800000 289.750000  95.870000 ;
      RECT 100.325000  95.730000 289.680000  95.800000 ;
      RECT 100.325000  95.730000 289.680000  95.800000 ;
      RECT 100.395000  95.660000 289.610000  95.730000 ;
      RECT 100.395000  95.660000 289.610000  95.730000 ;
      RECT 100.465000  95.590000 289.540000  95.660000 ;
      RECT 100.465000  95.590000 289.540000  95.660000 ;
      RECT 100.535000  95.520000 289.470000  95.590000 ;
      RECT 100.535000  95.520000 289.470000  95.590000 ;
      RECT 100.605000  95.450000 289.400000  95.520000 ;
      RECT 100.605000  95.450000 289.400000  95.520000 ;
      RECT 100.675000  95.380000 289.330000  95.450000 ;
      RECT 100.675000  95.380000 289.330000  95.450000 ;
      RECT 100.745000  95.310000 289.260000  95.380000 ;
      RECT 100.745000  95.310000 289.260000  95.380000 ;
      RECT 100.755000  95.100000 297.270000 103.125000 ;
      RECT 100.815000  95.240000 289.190000  95.310000 ;
      RECT 100.815000  95.240000 289.190000  95.310000 ;
      RECT 105.535000  95.205000 284.470000  95.240000 ;
      RECT 105.535000  95.205000 284.470000  95.240000 ;
      RECT 105.605000  95.135000 284.400000  95.205000 ;
      RECT 105.605000  95.135000 284.400000  95.205000 ;
      RECT 105.675000  95.065000 284.330000  95.135000 ;
      RECT 105.675000  95.065000 284.330000  95.135000 ;
      RECT 105.745000  94.995000 284.260000  95.065000 ;
      RECT 105.745000  94.995000 284.260000  95.065000 ;
      RECT 105.815000  94.925000 284.190000  94.995000 ;
      RECT 105.815000  94.925000 284.190000  94.995000 ;
      RECT 105.885000  94.855000 284.120000  94.925000 ;
      RECT 105.885000  94.855000 284.120000  94.925000 ;
      RECT 105.955000  94.785000 284.050000  94.855000 ;
      RECT 105.955000  94.785000 284.050000  94.855000 ;
      RECT 106.025000  94.715000 283.980000  94.785000 ;
      RECT 106.025000  94.715000 283.980000  94.785000 ;
      RECT 106.095000  94.645000 283.910000  94.715000 ;
      RECT 106.095000  94.645000 283.910000  94.715000 ;
      RECT 106.165000  94.575000 283.840000  94.645000 ;
      RECT 106.165000  94.575000 283.840000  94.645000 ;
      RECT 106.235000  89.625000 283.770000  94.310000 ;
      RECT 106.235000  94.310000 284.560000  95.100000 ;
      RECT 106.235000  94.505000 283.770000  94.575000 ;
      RECT 106.235000  94.505000 283.770000  94.575000 ;
      RECT 106.305000  94.435000 283.700000  94.505000 ;
      RECT 106.305000  94.435000 283.700000  94.505000 ;
      RECT 106.375000  89.680000 283.630000  94.365000 ;
      RECT 106.375000  94.365000 283.630000  94.435000 ;
      RECT 106.375000  94.365000 283.630000  94.435000 ;
      RECT 106.400000  89.655000 283.605000  89.680000 ;
      RECT 106.400000  89.655000 283.605000  89.680000 ;
      RECT 106.470000  89.585000 283.535000  89.655000 ;
      RECT 106.470000  89.585000 283.535000  89.655000 ;
      RECT 106.540000  89.515000 283.465000  89.585000 ;
      RECT 106.540000  89.515000 283.465000  89.585000 ;
      RECT 106.610000  89.445000 283.395000  89.515000 ;
      RECT 106.610000  89.445000 283.395000  89.515000 ;
      RECT 106.680000  89.375000 283.325000  89.445000 ;
      RECT 106.680000  89.375000 283.325000  89.445000 ;
      RECT 106.750000  89.305000 283.255000  89.375000 ;
      RECT 106.750000  89.305000 283.255000  89.375000 ;
      RECT 106.820000  89.235000 283.185000  89.305000 ;
      RECT 106.820000  89.235000 283.185000  89.305000 ;
      RECT 106.890000  89.165000 283.115000  89.235000 ;
      RECT 106.890000  89.165000 283.115000  89.235000 ;
      RECT 106.960000  89.095000 283.045000  89.165000 ;
      RECT 106.960000  89.095000 283.045000  89.165000 ;
      RECT 107.030000  89.025000 282.975000  89.095000 ;
      RECT 107.030000  89.025000 282.975000  89.095000 ;
      RECT 107.100000  88.955000 282.905000  89.025000 ;
      RECT 107.100000  88.955000 282.905000  89.025000 ;
      RECT 107.110000   0.000000 109.950000   1.180000 ;
      RECT 107.110000   1.180000 109.950000   1.895000 ;
      RECT 107.170000  88.885000 282.835000  88.955000 ;
      RECT 107.170000  88.885000 282.835000  88.955000 ;
      RECT 107.240000  88.815000 282.765000  88.885000 ;
      RECT 107.240000  88.815000 282.765000  88.885000 ;
      RECT 107.250000   0.000000 109.810000   1.125000 ;
      RECT 107.310000  88.745000 282.695000  88.815000 ;
      RECT 107.310000  88.745000 282.695000  88.815000 ;
      RECT 107.320000   1.125000 109.810000   1.195000 ;
      RECT 107.380000  88.675000 282.625000  88.745000 ;
      RECT 107.380000  88.675000 282.625000  88.745000 ;
      RECT 107.390000   1.195000 109.810000   1.265000 ;
      RECT 107.450000  88.605000 282.555000  88.675000 ;
      RECT 107.450000  88.605000 282.555000  88.675000 ;
      RECT 107.460000   1.265000 109.810000   1.335000 ;
      RECT 107.520000  88.535000 282.485000  88.605000 ;
      RECT 107.520000  88.535000 282.485000  88.605000 ;
      RECT 107.530000   1.335000 109.810000   1.405000 ;
      RECT 107.590000  88.465000 282.415000  88.535000 ;
      RECT 107.590000  88.465000 282.415000  88.535000 ;
      RECT 107.600000   1.405000 109.810000   1.475000 ;
      RECT 107.660000  88.395000 282.345000  88.465000 ;
      RECT 107.660000  88.395000 282.345000  88.465000 ;
      RECT 107.670000   1.475000 109.810000   1.545000 ;
      RECT 107.730000  88.325000 282.275000  88.395000 ;
      RECT 107.730000  88.325000 282.275000  88.395000 ;
      RECT 107.740000   1.545000 109.810000   1.615000 ;
      RECT 107.800000  88.255000 282.205000  88.325000 ;
      RECT 107.800000  88.255000 282.205000  88.325000 ;
      RECT 107.810000   1.615000 109.810000   1.685000 ;
      RECT 107.825000   1.895000 109.950000  17.295000 ;
      RECT 107.825000  17.295000 109.675000  17.570000 ;
      RECT 107.825000  17.570000 109.675000  18.295000 ;
      RECT 107.870000  88.185000 282.135000  88.255000 ;
      RECT 107.870000  88.185000 282.135000  88.255000 ;
      RECT 107.880000   1.685000 109.810000   1.755000 ;
      RECT 107.935000   2.680000 109.810000   7.155000 ;
      RECT 107.940000  88.115000 282.065000  88.185000 ;
      RECT 107.940000  88.115000 282.065000  88.185000 ;
      RECT 107.950000   1.755000 109.810000   1.825000 ;
      RECT 107.965000   1.825000 109.810000   1.840000 ;
      RECT 107.965000   1.840000 109.810000   2.680000 ;
      RECT 107.965000   7.155000 109.810000  17.240000 ;
      RECT 107.965000  17.240000 109.740000  17.310000 ;
      RECT 107.965000  17.310000 109.670000  17.380000 ;
      RECT 107.965000  17.380000 109.600000  17.450000 ;
      RECT 107.965000  17.450000 109.535000  17.515000 ;
      RECT 107.965000  17.515000 109.535000  18.435000 ;
      RECT 108.010000  88.045000 281.995000  88.115000 ;
      RECT 108.010000  88.045000 281.995000  88.115000 ;
      RECT 108.080000  87.975000 281.925000  88.045000 ;
      RECT 108.080000  87.975000 281.925000  88.045000 ;
      RECT 108.150000  76.675000 281.855000  87.710000 ;
      RECT 108.150000  87.710000 283.770000  89.625000 ;
      RECT 108.150000  87.905000 281.855000  87.975000 ;
      RECT 108.150000  87.905000 281.855000  87.975000 ;
      RECT 108.220000  87.835000 281.785000  87.905000 ;
      RECT 108.220000  87.835000 281.785000  87.905000 ;
      RECT 108.290000  76.735000 281.715000  87.765000 ;
      RECT 108.290000  76.735000 281.715000  89.680000 ;
      RECT 108.290000  76.735000 281.715000  94.365000 ;
      RECT 108.290000  87.765000 281.715000  87.835000 ;
      RECT 108.290000  87.765000 281.715000  87.835000 ;
      RECT 108.310000  76.715000 281.695000  76.735000 ;
      RECT 108.310000  76.715000 281.695000  76.735000 ;
      RECT 108.380000  76.645000 281.625000  76.715000 ;
      RECT 108.380000  76.645000 281.625000  76.715000 ;
      RECT 108.450000  76.575000 281.555000  76.645000 ;
      RECT 108.450000  76.575000 281.555000  76.645000 ;
      RECT 108.520000  76.505000 281.485000  76.575000 ;
      RECT 108.520000  76.505000 281.485000  76.575000 ;
      RECT 108.590000  76.435000 281.415000  76.505000 ;
      RECT 108.590000  76.435000 281.415000  76.505000 ;
      RECT 108.660000  76.365000 281.345000  76.435000 ;
      RECT 108.660000  76.365000 281.345000  76.435000 ;
      RECT 108.730000  76.295000 281.275000  76.365000 ;
      RECT 108.730000  76.295000 281.275000  76.365000 ;
      RECT 108.800000  76.225000 281.205000  76.295000 ;
      RECT 108.800000  76.225000 281.205000  76.295000 ;
      RECT 108.870000  76.155000 281.135000  76.225000 ;
      RECT 108.870000  76.155000 281.135000  76.225000 ;
      RECT 108.940000  76.085000 281.065000  76.155000 ;
      RECT 108.940000  76.085000 281.065000  76.155000 ;
      RECT 108.970000  47.630000 125.515000  48.605000 ;
      RECT 108.970000  48.605000 125.210000  48.910000 ;
      RECT 108.970000  48.910000 125.210000  51.985000 ;
      RECT 108.970000  51.985000 149.665000  56.395000 ;
      RECT 108.970000  56.395000 149.665000  57.205000 ;
      RECT 109.010000  76.015000 280.995000  76.085000 ;
      RECT 109.010000  76.015000 280.995000  76.085000 ;
      RECT 109.070000  47.530000 125.515000  47.630000 ;
      RECT 109.080000  75.945000 280.925000  76.015000 ;
      RECT 109.080000  75.945000 280.925000  76.015000 ;
      RECT 109.110000  47.685000 125.375000  48.070000 ;
      RECT 109.110000  48.070000 125.375000  48.550000 ;
      RECT 109.110000  48.550000 125.070000  52.125000 ;
      RECT 109.110000  48.550000 125.070000  52.125000 ;
      RECT 109.110000  48.550000 125.070000  52.125000 ;
      RECT 109.110000  48.550000 125.070000  52.125000 ;
      RECT 109.110000  48.550000 125.305000  48.620000 ;
      RECT 109.110000  48.550000 125.305000  48.620000 ;
      RECT 109.110000  48.620000 125.235000  48.690000 ;
      RECT 109.110000  48.620000 125.235000  48.690000 ;
      RECT 109.110000  48.690000 125.165000  48.760000 ;
      RECT 109.110000  48.690000 125.165000  48.760000 ;
      RECT 109.110000  48.760000 125.095000  48.830000 ;
      RECT 109.110000  48.760000 125.095000  48.830000 ;
      RECT 109.110000  48.830000 125.070000  48.855000 ;
      RECT 109.110000  48.830000 125.070000  48.855000 ;
      RECT 109.110000  48.855000 125.070000  48.855000 ;
      RECT 109.110000  48.855000 125.070000  52.125000 ;
      RECT 109.110000  52.125000 149.525000  56.340000 ;
      RECT 109.150000  75.875000 280.855000  75.945000 ;
      RECT 109.150000  75.875000 280.855000  75.945000 ;
      RECT 109.160000  47.635000 125.375000  47.685000 ;
      RECT 109.160000  47.635000 125.375000  47.685000 ;
      RECT 109.180000  56.340000 149.525000  56.410000 ;
      RECT 109.180000  56.340000 149.525000  56.410000 ;
      RECT 109.210000  47.585000 125.375000  47.635000 ;
      RECT 109.210000  47.585000 125.375000  47.635000 ;
      RECT 109.220000  75.805000 280.785000  75.875000 ;
      RECT 109.220000  75.805000 280.785000  75.875000 ;
      RECT 109.235000  47.560000 125.350000  47.585000 ;
      RECT 109.235000  47.560000 125.350000  47.585000 ;
      RECT 109.250000  56.410000 149.525000  56.480000 ;
      RECT 109.250000  56.410000 149.525000  56.480000 ;
      RECT 109.290000  75.735000 280.715000  75.805000 ;
      RECT 109.290000  75.735000 280.715000  75.805000 ;
      RECT 109.305000  47.490000 125.280000  47.560000 ;
      RECT 109.305000  47.490000 125.280000  47.560000 ;
      RECT 109.320000  56.480000 149.525000  56.550000 ;
      RECT 109.320000  56.480000 149.525000  56.550000 ;
      RECT 109.360000  75.665000 280.645000  75.735000 ;
      RECT 109.360000  75.665000 280.645000  75.735000 ;
      RECT 109.375000  47.420000 125.210000  47.490000 ;
      RECT 109.375000  47.420000 125.210000  47.490000 ;
      RECT 109.390000  56.550000 149.525000  56.620000 ;
      RECT 109.390000  56.550000 149.525000  56.620000 ;
      RECT 109.430000  75.595000 280.575000  75.665000 ;
      RECT 109.430000  75.595000 280.575000  75.665000 ;
      RECT 109.445000  47.350000 125.140000  47.420000 ;
      RECT 109.445000  47.350000 125.140000  47.420000 ;
      RECT 109.460000  56.620000 149.525000  56.690000 ;
      RECT 109.460000  56.620000 149.525000  56.690000 ;
      RECT 109.500000  75.525000 280.505000  75.595000 ;
      RECT 109.500000  75.525000 280.505000  75.595000 ;
      RECT 109.515000  47.280000 125.070000  47.350000 ;
      RECT 109.515000  47.280000 125.070000  47.350000 ;
      RECT 109.530000  56.690000 149.525000  56.760000 ;
      RECT 109.530000  56.690000 149.525000  56.760000 ;
      RECT 109.570000  75.455000 280.435000  75.525000 ;
      RECT 109.570000  75.455000 280.435000  75.525000 ;
      RECT 109.585000  47.210000 125.000000  47.280000 ;
      RECT 109.585000  47.210000 125.000000  47.280000 ;
      RECT 109.600000  56.760000 149.525000  56.830000 ;
      RECT 109.600000  56.760000 149.525000  56.830000 ;
      RECT 109.640000  75.385000 280.365000  75.455000 ;
      RECT 109.640000  75.385000 280.365000  75.455000 ;
      RECT 109.655000  47.140000 124.930000  47.210000 ;
      RECT 109.655000  47.140000 124.930000  47.210000 ;
      RECT 109.670000  56.830000 149.525000  56.900000 ;
      RECT 109.670000  56.830000 149.525000  56.900000 ;
      RECT 109.710000  75.315000 280.295000  75.385000 ;
      RECT 109.710000  75.315000 280.295000  75.385000 ;
      RECT 109.725000  47.070000 124.860000  47.140000 ;
      RECT 109.725000  47.070000 124.860000  47.140000 ;
      RECT 109.740000  56.900000 149.525000  56.970000 ;
      RECT 109.740000  56.900000 149.525000  56.970000 ;
      RECT 109.780000  57.205000 149.665000  58.665000 ;
      RECT 109.780000  58.665000 280.225000  75.050000 ;
      RECT 109.780000  75.050000 281.855000  76.675000 ;
      RECT 109.780000  75.245000 280.225000  75.315000 ;
      RECT 109.780000  75.245000 280.225000  75.315000 ;
      RECT 109.795000  47.000000 124.790000  47.070000 ;
      RECT 109.795000  47.000000 124.790000  47.070000 ;
      RECT 109.810000  56.970000 149.525000  57.040000 ;
      RECT 109.810000  56.970000 149.525000  57.040000 ;
      RECT 109.850000  75.175000 280.155000  75.245000 ;
      RECT 109.850000  75.175000 280.155000  75.245000 ;
      RECT 109.865000  46.020000 121.315000  46.420000 ;
      RECT 109.865000  46.420000 124.720000  46.735000 ;
      RECT 109.865000  46.735000 125.515000  47.530000 ;
      RECT 109.865000  46.930000 124.720000  47.000000 ;
      RECT 109.865000  46.930000 124.720000  47.000000 ;
      RECT 109.880000  57.040000 149.525000  57.110000 ;
      RECT 109.880000  57.040000 149.525000  57.110000 ;
      RECT 109.920000  52.125000 149.525000  75.105000 ;
      RECT 109.920000  52.125000 149.525000  75.105000 ;
      RECT 109.920000  57.110000 149.525000  57.150000 ;
      RECT 109.920000  57.110000 149.525000  57.150000 ;
      RECT 109.920000  57.150000 149.525000  58.805000 ;
      RECT 109.920000  58.805000 280.085000  75.105000 ;
      RECT 109.920000  75.105000 280.085000  75.175000 ;
      RECT 109.920000  75.105000 280.085000  75.175000 ;
      RECT 109.935000  46.860000 124.650000  46.930000 ;
      RECT 109.935000  46.860000 124.650000  46.930000 ;
      RECT 110.005000  46.075000 121.175000  46.560000 ;
      RECT 110.005000  46.560000 124.350000  46.630000 ;
      RECT 110.005000  46.560000 124.350000  46.630000 ;
      RECT 110.005000  46.630000 124.420000  46.700000 ;
      RECT 110.005000  46.630000 124.420000  46.700000 ;
      RECT 110.005000  46.700000 124.490000  46.770000 ;
      RECT 110.005000  46.700000 124.490000  46.770000 ;
      RECT 110.005000  46.770000 124.560000  46.790000 ;
      RECT 110.005000  46.770000 124.560000  46.790000 ;
      RECT 110.005000  46.790000 124.580000  46.860000 ;
      RECT 110.005000  46.790000 124.580000  46.860000 ;
      RECT 110.025000  46.055000 121.175000  46.075000 ;
      RECT 110.025000  46.055000 121.175000  46.075000 ;
      RECT 110.095000  45.985000 121.175000  46.055000 ;
      RECT 110.095000  45.985000 121.175000  46.055000 ;
      RECT 110.165000  45.915000 121.175000  45.985000 ;
      RECT 110.165000  45.915000 121.175000  45.985000 ;
      RECT 110.215000  17.795000 121.315000  36.240000 ;
      RECT 110.215000  36.240000 121.315000  36.260000 ;
      RECT 110.235000  36.260000 121.315000  45.650000 ;
      RECT 110.235000  45.650000 121.315000  46.020000 ;
      RECT 110.235000  45.845000 121.175000  45.915000 ;
      RECT 110.235000  45.845000 121.175000  45.915000 ;
      RECT 110.305000  45.775000 121.175000  45.845000 ;
      RECT 110.305000  45.775000 121.175000  45.845000 ;
      RECT 110.355000  17.855000 121.175000  36.185000 ;
      RECT 110.365000  36.185000 121.175000  36.195000 ;
      RECT 110.365000  36.185000 121.175000  36.195000 ;
      RECT 110.375000  36.195000 121.175000  36.205000 ;
      RECT 110.375000  36.195000 121.175000  36.205000 ;
      RECT 110.375000  36.205000 121.175000  46.790000 ;
      RECT 110.375000  45.705000 121.175000  45.775000 ;
      RECT 110.375000  45.705000 121.175000  45.775000 ;
      RECT 110.420000  17.790000 121.175000  17.855000 ;
      RECT 110.420000  17.790000 121.175000  17.855000 ;
      RECT 110.490000   0.000000 121.315000  17.525000 ;
      RECT 110.490000  17.525000 121.315000  17.795000 ;
      RECT 110.490000  17.720000 121.175000  17.790000 ;
      RECT 110.490000  17.720000 121.175000  17.790000 ;
      RECT 110.560000  17.650000 121.175000  17.720000 ;
      RECT 110.560000  17.650000 121.175000  17.720000 ;
      RECT 110.630000   0.000000 121.175000  17.580000 ;
      RECT 110.630000  17.580000 121.175000  17.650000 ;
      RECT 110.630000  17.580000 121.175000  17.650000 ;
      RECT 121.855000   0.000000 127.985000  10.005000 ;
      RECT 121.855000  10.005000 127.120000  10.870000 ;
      RECT 121.855000  10.870000 127.120000  23.830000 ;
      RECT 121.855000  23.830000 127.720000  24.435000 ;
      RECT 121.855000  24.435000 127.720000  43.050000 ;
      RECT 121.855000  43.050000 145.495000  45.780000 ;
      RECT 121.855000  45.780000 145.495000  45.880000 ;
      RECT 121.995000   0.000000 127.845000   2.610000 ;
      RECT 121.995000   0.000000 127.845000   7.810000 ;
      RECT 121.995000   0.000000 127.845000   7.810000 ;
      RECT 121.995000   2.610000 127.980000   7.810000 ;
      RECT 121.995000   7.810000 127.845000   9.950000 ;
      RECT 121.995000   9.950000 126.980000  23.890000 ;
      RECT 121.995000   9.950000 126.980000  23.890000 ;
      RECT 121.995000   9.950000 127.775000  10.020000 ;
      RECT 121.995000   9.950000 127.775000  10.020000 ;
      RECT 121.995000  10.020000 127.705000  10.090000 ;
      RECT 121.995000  10.020000 127.705000  10.090000 ;
      RECT 121.995000  10.090000 127.635000  10.160000 ;
      RECT 121.995000  10.090000 127.635000  10.160000 ;
      RECT 121.995000  10.160000 127.565000  10.230000 ;
      RECT 121.995000  10.160000 127.565000  10.230000 ;
      RECT 121.995000  10.230000 127.495000  10.300000 ;
      RECT 121.995000  10.230000 127.495000  10.300000 ;
      RECT 121.995000  10.300000 127.425000  10.370000 ;
      RECT 121.995000  10.300000 127.425000  10.370000 ;
      RECT 121.995000  10.370000 127.355000  10.440000 ;
      RECT 121.995000  10.370000 127.355000  10.440000 ;
      RECT 121.995000  10.440000 127.285000  10.510000 ;
      RECT 121.995000  10.440000 127.285000  10.510000 ;
      RECT 121.995000  10.510000 127.215000  10.580000 ;
      RECT 121.995000  10.510000 127.215000  10.580000 ;
      RECT 121.995000  10.580000 127.145000  10.650000 ;
      RECT 121.995000  10.580000 127.145000  10.650000 ;
      RECT 121.995000  10.650000 127.075000  10.720000 ;
      RECT 121.995000  10.650000 127.075000  10.720000 ;
      RECT 121.995000  10.720000 127.005000  10.790000 ;
      RECT 121.995000  10.720000 127.005000  10.790000 ;
      RECT 121.995000  10.790000 126.980000  10.815000 ;
      RECT 121.995000  10.790000 126.980000  10.815000 ;
      RECT 121.995000  10.815000 126.980000  23.890000 ;
      RECT 121.995000  23.890000 126.980000  23.960000 ;
      RECT 121.995000  23.890000 126.980000  23.960000 ;
      RECT 121.995000  23.960000 127.050000  24.030000 ;
      RECT 121.995000  23.960000 127.050000  24.030000 ;
      RECT 121.995000  24.030000 127.120000  24.100000 ;
      RECT 121.995000  24.030000 127.120000  24.100000 ;
      RECT 121.995000  24.100000 127.190000  24.170000 ;
      RECT 121.995000  24.100000 127.190000  24.170000 ;
      RECT 121.995000  24.170000 127.260000  24.240000 ;
      RECT 121.995000  24.170000 127.260000  24.240000 ;
      RECT 121.995000  24.240000 127.330000  24.310000 ;
      RECT 121.995000  24.240000 127.330000  24.310000 ;
      RECT 121.995000  24.310000 127.400000  24.380000 ;
      RECT 121.995000  24.310000 127.400000  24.380000 ;
      RECT 121.995000  24.380000 127.470000  24.450000 ;
      RECT 121.995000  24.380000 127.470000  24.450000 ;
      RECT 121.995000  24.450000 127.540000  24.490000 ;
      RECT 121.995000  24.450000 127.540000  24.490000 ;
      RECT 121.995000  24.490000 127.580000  43.190000 ;
      RECT 121.995000  24.490000 127.580000  45.740000 ;
      RECT 121.995000  24.490000 127.580000  45.740000 ;
      RECT 121.995000  24.490000 127.580000  45.740000 ;
      RECT 121.995000  24.490000 127.580000  45.740000 ;
      RECT 121.995000  43.190000 145.355000  45.740000 ;
      RECT 124.630000  45.880000 145.495000  47.300000 ;
      RECT 124.760000  45.740000 145.355000  45.810000 ;
      RECT 124.760000  45.740000 145.355000  45.810000 ;
      RECT 124.830000  45.810000 145.355000  45.880000 ;
      RECT 124.830000  45.810000 145.355000  45.880000 ;
      RECT 124.900000  45.880000 145.355000  45.950000 ;
      RECT 124.900000  45.880000 145.355000  45.950000 ;
      RECT 124.970000  45.950000 145.355000  46.020000 ;
      RECT 124.970000  45.950000 145.355000  46.020000 ;
      RECT 125.040000  46.020000 145.355000  46.090000 ;
      RECT 125.040000  46.020000 145.355000  46.090000 ;
      RECT 125.110000  46.090000 145.355000  46.160000 ;
      RECT 125.110000  46.090000 145.355000  46.160000 ;
      RECT 125.180000  46.160000 145.355000  46.230000 ;
      RECT 125.180000  46.160000 145.355000  46.230000 ;
      RECT 125.250000  46.230000 145.355000  46.300000 ;
      RECT 125.250000  46.230000 145.355000  46.300000 ;
      RECT 125.320000  46.300000 145.355000  46.370000 ;
      RECT 125.320000  46.300000 145.355000  46.370000 ;
      RECT 125.390000  46.370000 145.355000  46.440000 ;
      RECT 125.390000  46.370000 145.355000  46.440000 ;
      RECT 125.460000  46.440000 145.355000  46.510000 ;
      RECT 125.460000  46.440000 145.355000  46.510000 ;
      RECT 125.530000  46.510000 145.355000  46.580000 ;
      RECT 125.530000  46.510000 145.355000  46.580000 ;
      RECT 125.600000  46.580000 145.355000  46.650000 ;
      RECT 125.600000  46.580000 145.355000  46.650000 ;
      RECT 125.670000  46.650000 145.355000  46.720000 ;
      RECT 125.670000  46.650000 145.355000  46.720000 ;
      RECT 125.740000  46.720000 145.355000  46.790000 ;
      RECT 125.740000  46.720000 145.355000  46.790000 ;
      RECT 125.810000  46.790000 145.355000  46.860000 ;
      RECT 125.810000  46.790000 145.355000  46.860000 ;
      RECT 125.880000  46.860000 145.355000  46.930000 ;
      RECT 125.880000  46.860000 145.355000  46.930000 ;
      RECT 125.950000  46.930000 145.355000  47.000000 ;
      RECT 125.950000  46.930000 145.355000  47.000000 ;
      RECT 126.020000  47.000000 145.355000  47.070000 ;
      RECT 126.020000  47.000000 145.355000  47.070000 ;
      RECT 126.055000  47.300000 145.495000  48.770000 ;
      RECT 126.055000  48.770000 145.495000  48.910000 ;
      RECT 126.090000  47.070000 145.355000  47.140000 ;
      RECT 126.090000  47.070000 145.355000  47.140000 ;
      RECT 126.160000  47.140000 145.355000  47.210000 ;
      RECT 126.160000  47.140000 145.355000  47.210000 ;
      RECT 126.195000  47.210000 145.355000  47.245000 ;
      RECT 126.195000  47.210000 145.355000  47.245000 ;
      RECT 126.195000  47.245000 145.355000  48.715000 ;
      RECT 126.195000  48.910000 145.495000  49.170000 ;
      RECT 126.195000  49.170000 145.450000  49.215000 ;
      RECT 126.195000  49.215000 145.115000  49.755000 ;
      RECT 126.195000  49.755000 149.665000  51.985000 ;
      RECT 126.265000  48.715000 145.355000  48.785000 ;
      RECT 126.265000  48.715000 145.355000  48.785000 ;
      RECT 126.335000  48.715000 144.975000  56.340000 ;
      RECT 126.335000  48.715000 144.975000  56.340000 ;
      RECT 126.335000  48.715000 144.975000  56.340000 ;
      RECT 126.335000  48.785000 145.355000  48.855000 ;
      RECT 126.335000  48.785000 145.355000  48.855000 ;
      RECT 126.335000  48.855000 145.355000  49.075000 ;
      RECT 126.335000  49.895000 149.525000  52.125000 ;
      RECT 126.335000  49.895000 149.525000  56.340000 ;
      RECT 126.335000  49.895000 149.525000  56.340000 ;
      RECT 126.335000  49.895000 149.525000  56.340000 ;
      RECT 127.660000  11.100000 135.035000  23.605000 ;
      RECT 127.660000  23.605000 135.035000  24.205000 ;
      RECT 127.800000  11.155000 134.895000  23.550000 ;
      RECT 127.825000  11.130000 134.895000  11.155000 ;
      RECT 127.825000  11.130000 134.895000  11.155000 ;
      RECT 127.870000  23.550000 134.895000  23.620000 ;
      RECT 127.870000  23.550000 134.895000  23.620000 ;
      RECT 127.895000  11.060000 134.895000  11.130000 ;
      RECT 127.895000  11.060000 134.895000  11.130000 ;
      RECT 127.940000  23.620000 134.895000  23.690000 ;
      RECT 127.940000  23.620000 134.895000  23.690000 ;
      RECT 127.965000  10.990000 134.895000  11.060000 ;
      RECT 127.965000  10.990000 134.895000  11.060000 ;
      RECT 128.010000  23.690000 134.895000  23.760000 ;
      RECT 128.010000  23.690000 134.895000  23.760000 ;
      RECT 128.035000  10.920000 134.895000  10.990000 ;
      RECT 128.035000  10.920000 134.895000  10.990000 ;
      RECT 128.080000  23.760000 134.895000  23.830000 ;
      RECT 128.080000  23.760000 134.895000  23.830000 ;
      RECT 128.105000  10.850000 134.895000  10.920000 ;
      RECT 128.105000  10.850000 134.895000  10.920000 ;
      RECT 128.150000  23.830000 134.895000  23.900000 ;
      RECT 128.150000  23.830000 134.895000  23.900000 ;
      RECT 128.175000  10.780000 134.895000  10.850000 ;
      RECT 128.175000  10.780000 134.895000  10.850000 ;
      RECT 128.220000  23.900000 134.895000  23.970000 ;
      RECT 128.220000  23.900000 134.895000  23.970000 ;
      RECT 128.245000  10.710000 134.895000  10.780000 ;
      RECT 128.245000  10.710000 134.895000  10.780000 ;
      RECT 128.260000  24.205000 135.035000  28.780000 ;
      RECT 128.260000  28.780000 134.505000  29.310000 ;
      RECT 128.260000  29.310000 134.505000  29.800000 ;
      RECT 128.260000  29.800000 134.460000  29.845000 ;
      RECT 128.260000  29.845000 133.615000  30.385000 ;
      RECT 128.260000  30.385000 133.995000  30.430000 ;
      RECT 128.260000  30.430000 133.995000  42.465000 ;
      RECT 128.260000  42.465000 133.995000  42.510000 ;
      RECT 128.290000  23.970000 134.895000  24.040000 ;
      RECT 128.290000  23.970000 134.895000  24.040000 ;
      RECT 128.315000  10.640000 134.895000  10.710000 ;
      RECT 128.315000  10.640000 134.895000  10.710000 ;
      RECT 128.360000  24.040000 134.895000  24.110000 ;
      RECT 128.360000  24.040000 134.895000  24.110000 ;
      RECT 128.385000  10.570000 134.895000  10.640000 ;
      RECT 128.385000  10.570000 134.895000  10.640000 ;
      RECT 128.400000  24.110000 134.895000  24.150000 ;
      RECT 128.400000  24.110000 134.895000  24.150000 ;
      RECT 128.400000  24.150000 134.895000  28.725000 ;
      RECT 128.400000  28.725000 133.475000  42.370000 ;
      RECT 128.400000  28.725000 134.825000  28.795000 ;
      RECT 128.400000  28.725000 134.825000  28.795000 ;
      RECT 128.400000  28.795000 134.755000  28.865000 ;
      RECT 128.400000  28.795000 134.755000  28.865000 ;
      RECT 128.400000  28.865000 134.685000  28.935000 ;
      RECT 128.400000  28.865000 134.685000  28.935000 ;
      RECT 128.400000  28.935000 134.615000  29.005000 ;
      RECT 128.400000  28.935000 134.615000  29.005000 ;
      RECT 128.400000  29.005000 134.545000  29.075000 ;
      RECT 128.400000  29.005000 134.545000  29.075000 ;
      RECT 128.400000  29.075000 134.475000  29.145000 ;
      RECT 128.400000  29.075000 134.475000  29.145000 ;
      RECT 128.400000  29.145000 134.405000  29.215000 ;
      RECT 128.400000  29.145000 134.405000  29.215000 ;
      RECT 128.400000  29.215000 134.365000  29.255000 ;
      RECT 128.400000  29.215000 134.365000  29.255000 ;
      RECT 128.400000  29.255000 134.295000  29.325000 ;
      RECT 128.400000  29.255000 134.295000  29.325000 ;
      RECT 128.400000  29.325000 134.225000  29.395000 ;
      RECT 128.400000  29.325000 134.225000  29.395000 ;
      RECT 128.400000  29.395000 134.155000  29.465000 ;
      RECT 128.400000  29.395000 134.155000  29.465000 ;
      RECT 128.400000  29.465000 134.085000  29.535000 ;
      RECT 128.400000  29.465000 134.085000  29.535000 ;
      RECT 128.400000  29.535000 134.015000  29.605000 ;
      RECT 128.400000  29.535000 134.015000  29.605000 ;
      RECT 128.400000  29.605000 133.945000  29.675000 ;
      RECT 128.400000  29.605000 133.945000  29.675000 ;
      RECT 128.400000  29.675000 133.915000  29.705000 ;
      RECT 128.400000  29.675000 133.915000  29.705000 ;
      RECT 128.400000  29.705000 133.475000  30.525000 ;
      RECT 128.400000  30.525000 133.855000  42.370000 ;
      RECT 128.455000  10.500000 134.895000  10.570000 ;
      RECT 128.455000  10.500000 134.895000  10.570000 ;
      RECT 128.525000   0.000000 135.035000  10.235000 ;
      RECT 128.525000  10.235000 135.035000  11.100000 ;
      RECT 128.525000  10.430000 134.895000  10.500000 ;
      RECT 128.525000  10.430000 134.895000  10.500000 ;
      RECT 128.595000  10.360000 134.895000  10.430000 ;
      RECT 128.595000  10.360000 134.895000  10.430000 ;
      RECT 128.665000   0.000000 134.895000   3.005000 ;
      RECT 128.665000   2.610000 134.895000  11.155000 ;
      RECT 128.665000   2.610000 134.895000  11.155000 ;
      RECT 128.665000   2.610000 134.895000  11.155000 ;
      RECT 128.665000   2.610000 135.035000   7.810000 ;
      RECT 128.665000   7.810000 134.895000  10.290000 ;
      RECT 128.665000  10.290000 134.895000  10.360000 ;
      RECT 128.665000  10.290000 134.895000  10.360000 ;
      RECT 129.020000  42.510000 133.995000  42.880000 ;
      RECT 129.020000  42.880000 145.495000  43.050000 ;
      RECT 129.160000  30.525000 133.855000  43.190000 ;
      RECT 129.160000  30.525000 133.855000  43.190000 ;
      RECT 129.160000  30.525000 133.855000  43.190000 ;
      RECT 129.160000  42.370000 133.855000  43.020000 ;
      RECT 129.160000  43.020000 145.355000  43.190000 ;
      RECT 134.535000  30.430000 135.435000  36.505000 ;
      RECT 134.535000  36.505000 135.390000  36.550000 ;
      RECT 134.535000  36.550000 135.055000  37.090000 ;
      RECT 134.535000  37.090000 145.495000  42.880000 ;
      RECT 134.580000  30.385000 135.435000  30.430000 ;
      RECT 134.675000  30.525000 135.295000  36.410000 ;
      RECT 134.675000  36.410000 134.915000  37.230000 ;
      RECT 134.675000  37.230000 145.355000  43.020000 ;
      RECT 134.675000  37.230000 145.355000  43.190000 ;
      RECT 134.675000  37.230000 145.355000  43.190000 ;
      RECT 134.675000  37.230000 145.355000  43.190000 ;
      RECT 134.805000  30.465000 135.295000  30.525000 ;
      RECT 134.875000  30.395000 135.295000  30.465000 ;
      RECT 134.945000  30.325000 135.295000  30.395000 ;
      RECT 135.015000  30.255000 135.295000  30.325000 ;
      RECT 135.045000  29.540000 135.435000  30.025000 ;
      RECT 135.045000  30.025000 135.435000  30.385000 ;
      RECT 135.085000  30.185000 135.295000  30.255000 ;
      RECT 135.155000  30.115000 135.295000  30.185000 ;
      RECT 135.225000  30.045000 135.295000  30.115000 ;
      RECT 135.975000   0.000000 141.060000   1.820000 ;
      RECT 135.975000   1.570000 140.715000   1.765000 ;
      RECT 135.975000   1.765000 140.715000   4.770000 ;
      RECT 135.975000   1.765000 140.850000   1.835000 ;
      RECT 135.975000   1.820000 140.855000   2.025000 ;
      RECT 135.975000   1.835000 140.780000   1.905000 ;
      RECT 135.975000   1.905000 140.715000   1.970000 ;
      RECT 135.975000   2.025000 140.855000   2.485000 ;
      RECT 135.975000   2.485000 141.865000   7.720000 ;
      RECT 135.975000   2.625000 141.725000   6.100000 ;
      RECT 135.975000   7.720000 142.265000  10.730000 ;
      RECT 135.975000  10.730000 147.075000  26.750000 ;
      RECT 135.975000  26.750000 145.495000  28.330000 ;
      RECT 135.975000  28.330000 145.495000  37.090000 ;
      RECT 136.115000   0.000000 140.715000   1.570000 ;
      RECT 136.115000   2.625000 141.725000  10.870000 ;
      RECT 136.115000   2.625000 141.725000  10.870000 ;
      RECT 136.115000   6.100000 141.725000   7.860000 ;
      RECT 136.115000   7.860000 142.125000  10.870000 ;
      RECT 136.115000   7.860000 142.125000  26.695000 ;
      RECT 136.115000   7.860000 142.125000  26.695000 ;
      RECT 136.115000  10.870000 146.935000  26.695000 ;
      RECT 136.115000  26.695000 145.355000  37.230000 ;
      RECT 136.115000  26.695000 146.865000  26.765000 ;
      RECT 136.115000  26.695000 146.865000  26.765000 ;
      RECT 136.115000  26.765000 146.795000  26.835000 ;
      RECT 136.115000  26.765000 146.795000  26.835000 ;
      RECT 136.115000  26.835000 146.725000  26.905000 ;
      RECT 136.115000  26.835000 146.725000  26.905000 ;
      RECT 136.115000  26.905000 146.655000  26.975000 ;
      RECT 136.115000  26.905000 146.655000  26.975000 ;
      RECT 136.115000  26.975000 146.585000  27.045000 ;
      RECT 136.115000  26.975000 146.585000  27.045000 ;
      RECT 136.115000  27.045000 146.515000  27.115000 ;
      RECT 136.115000  27.045000 146.515000  27.115000 ;
      RECT 136.115000  27.115000 146.445000  27.185000 ;
      RECT 136.115000  27.115000 146.445000  27.185000 ;
      RECT 136.115000  27.185000 146.375000  27.255000 ;
      RECT 136.115000  27.185000 146.375000  27.255000 ;
      RECT 136.115000  27.255000 146.305000  27.325000 ;
      RECT 136.115000  27.255000 146.305000  27.325000 ;
      RECT 136.115000  27.325000 146.235000  27.395000 ;
      RECT 136.115000  27.325000 146.235000  27.395000 ;
      RECT 136.115000  27.395000 146.165000  27.465000 ;
      RECT 136.115000  27.395000 146.165000  27.465000 ;
      RECT 136.115000  27.465000 146.095000  27.535000 ;
      RECT 136.115000  27.465000 146.095000  27.535000 ;
      RECT 136.115000  27.535000 146.025000  27.605000 ;
      RECT 136.115000  27.535000 146.025000  27.605000 ;
      RECT 136.115000  27.605000 145.955000  27.675000 ;
      RECT 136.115000  27.605000 145.955000  27.675000 ;
      RECT 136.115000  27.675000 145.885000  27.745000 ;
      RECT 136.115000  27.675000 145.885000  27.745000 ;
      RECT 136.115000  27.745000 145.815000  27.815000 ;
      RECT 136.115000  27.745000 145.815000  27.815000 ;
      RECT 136.115000  27.815000 145.745000  27.885000 ;
      RECT 136.115000  27.815000 145.745000  27.885000 ;
      RECT 136.115000  27.885000 145.675000  27.955000 ;
      RECT 136.115000  27.885000 145.675000  27.955000 ;
      RECT 136.115000  27.955000 145.605000  28.025000 ;
      RECT 136.115000  27.955000 145.605000  28.025000 ;
      RECT 136.115000  28.025000 145.535000  28.095000 ;
      RECT 136.115000  28.025000 145.535000  28.095000 ;
      RECT 136.115000  28.095000 145.465000  28.165000 ;
      RECT 136.115000  28.095000 145.465000  28.165000 ;
      RECT 136.115000  28.165000 145.395000  28.235000 ;
      RECT 136.115000  28.165000 145.395000  28.235000 ;
      RECT 136.115000  28.235000 145.355000  28.275000 ;
      RECT 136.115000  28.235000 145.355000  28.275000 ;
      RECT 136.115000  28.275000 145.355000  37.230000 ;
      RECT 140.715000   0.000000 140.920000   1.765000 ;
      RECT 141.685000   0.000000 141.865000   1.935000 ;
      RECT 141.685000   1.935000 141.865000   2.025000 ;
      RECT 141.775000   2.025000 141.865000   2.485000 ;
      RECT 142.805000   0.000000 147.075000  10.730000 ;
      RECT 142.945000   0.000000 146.935000  10.870000 ;
      RECT 142.945000   0.000000 146.935000  26.695000 ;
      RECT 146.035000  28.560000 147.475000  46.275000 ;
      RECT 146.035000  46.275000 149.665000  49.755000 ;
      RECT 146.175000  28.615000 147.335000  46.415000 ;
      RECT 146.175000  46.415000 149.525000  49.895000 ;
      RECT 146.175000  46.415000 149.525000  52.125000 ;
      RECT 146.175000  46.415000 149.525000  56.340000 ;
      RECT 146.175000  46.415000 149.525000  56.340000 ;
      RECT 146.175000  46.415000 149.525000  56.340000 ;
      RECT 146.215000  28.575000 147.335000  28.615000 ;
      RECT 146.285000  28.505000 147.335000  28.575000 ;
      RECT 146.355000  28.435000 147.335000  28.505000 ;
      RECT 146.425000  28.365000 147.335000  28.435000 ;
      RECT 146.495000  28.295000 147.335000  28.365000 ;
      RECT 146.565000  28.225000 147.335000  28.295000 ;
      RECT 146.635000  28.155000 147.335000  28.225000 ;
      RECT 146.705000  28.085000 147.335000  28.155000 ;
      RECT 146.775000  28.015000 147.335000  28.085000 ;
      RECT 146.845000  27.945000 147.335000  28.015000 ;
      RECT 146.915000  27.875000 147.335000  27.945000 ;
      RECT 146.985000  27.805000 147.335000  27.875000 ;
      RECT 147.055000  27.735000 147.335000  27.805000 ;
      RECT 147.125000  27.665000 147.335000  27.735000 ;
      RECT 147.195000  27.595000 147.335000  27.665000 ;
      RECT 147.265000  27.525000 147.335000  27.595000 ;
      RECT 148.015000   0.000000 149.665000  28.310000 ;
      RECT 148.015000  28.310000 150.205000  28.845000 ;
      RECT 148.015000  28.845000 150.205000  30.665000 ;
      RECT 148.015000  30.665000 149.665000  31.205000 ;
      RECT 148.015000  31.205000 149.665000  46.275000 ;
      RECT 148.155000   0.000000 149.525000  28.365000 ;
      RECT 148.155000  28.365000 149.525000  28.435000 ;
      RECT 148.155000  28.435000 149.595000  28.505000 ;
      RECT 148.155000  28.505000 149.665000  28.575000 ;
      RECT 148.155000  28.575000 149.735000  28.645000 ;
      RECT 148.155000  28.645000 149.805000  28.715000 ;
      RECT 148.155000  28.715000 149.875000  28.785000 ;
      RECT 148.155000  28.785000 149.945000  28.855000 ;
      RECT 148.155000  28.855000 150.015000  28.905000 ;
      RECT 148.155000  28.905000 150.065000  30.610000 ;
      RECT 148.155000  30.610000 149.995000  30.680000 ;
      RECT 148.155000  30.680000 149.925000  30.750000 ;
      RECT 148.155000  30.750000 149.855000  30.820000 ;
      RECT 148.155000  30.820000 149.785000  30.890000 ;
      RECT 148.155000  30.890000 149.715000  30.960000 ;
      RECT 148.155000  30.960000 149.645000  31.030000 ;
      RECT 148.155000  31.030000 149.575000  31.100000 ;
      RECT 148.155000  31.100000 149.525000  31.150000 ;
      RECT 148.155000  31.150000 149.525000  46.415000 ;
      RECT 150.205000   0.000000 153.270000   2.155000 ;
      RECT 150.205000   2.155000 153.250000   2.175000 ;
      RECT 150.205000   2.175000 153.250000   3.065000 ;
      RECT 150.205000   3.065000 153.270000   3.085000 ;
      RECT 150.205000   3.085000 153.270000  27.815000 ;
      RECT 150.205000  27.815000 153.270000  28.355000 ;
      RECT 150.205000  31.700000 153.270000  35.085000 ;
      RECT 150.205000  35.085000 153.670000  42.155000 ;
      RECT 150.205000  42.155000 153.680000  42.165000 ;
      RECT 150.205000  42.165000 153.680000  43.050000 ;
      RECT 150.205000  43.050000 239.800000  58.080000 ;
      RECT 150.205000  58.080000 239.755000  58.125000 ;
      RECT 150.345000   0.000000 153.130000   2.100000 ;
      RECT 150.345000   2.100000 153.120000   2.110000 ;
      RECT 150.345000   2.110000 153.110000   2.120000 ;
      RECT 150.345000   2.120000 153.110000   3.120000 ;
      RECT 150.345000   3.120000 153.110000   3.130000 ;
      RECT 150.345000   3.130000 153.120000   3.140000 ;
      RECT 150.345000   3.140000 153.130000  27.760000 ;
      RECT 150.345000  31.755000 153.130000  35.225000 ;
      RECT 150.345000  35.225000 153.530000  42.210000 ;
      RECT 150.345000  35.225000 153.530000  57.985000 ;
      RECT 150.345000  35.225000 153.530000  57.985000 ;
      RECT 150.345000  42.210000 153.530000  42.215000 ;
      RECT 150.345000  42.210000 153.530000  42.215000 ;
      RECT 150.345000  42.215000 153.535000  42.220000 ;
      RECT 150.345000  42.215000 153.535000  42.220000 ;
      RECT 150.345000  42.220000 153.540000  43.190000 ;
      RECT 150.345000  43.190000 239.660000  57.985000 ;
      RECT 150.395000  31.705000 153.130000  31.755000 ;
      RECT 150.415000  27.760000 153.130000  27.830000 ;
      RECT 150.465000  31.635000 153.130000  31.705000 ;
      RECT 150.485000  27.830000 153.130000  27.900000 ;
      RECT 150.535000  31.565000 153.130000  31.635000 ;
      RECT 150.555000  27.900000 153.130000  27.970000 ;
      RECT 150.585000  58.125000 239.420000  58.665000 ;
      RECT 150.605000  31.495000 153.130000  31.565000 ;
      RECT 150.625000  27.970000 153.130000  28.040000 ;
      RECT 150.675000  31.425000 153.130000  31.495000 ;
      RECT 150.695000  28.040000 153.130000  28.110000 ;
      RECT 150.725000  43.190000 239.280000  58.805000 ;
      RECT 150.725000  43.190000 239.280000  58.805000 ;
      RECT 150.725000  43.190000 239.280000  58.805000 ;
      RECT 150.725000  57.985000 239.280000  58.805000 ;
      RECT 150.745000  28.355000 153.270000  31.160000 ;
      RECT 150.745000  31.160000 153.270000  31.700000 ;
      RECT 150.745000  31.355000 153.130000  31.425000 ;
      RECT 150.765000  28.110000 153.130000  28.180000 ;
      RECT 150.815000  31.285000 153.130000  31.355000 ;
      RECT 150.835000  28.180000 153.130000  28.250000 ;
      RECT 150.885000  28.250000 153.130000  28.300000 ;
      RECT 150.885000  28.300000 153.130000  31.215000 ;
      RECT 150.885000  31.215000 153.130000  31.285000 ;
      RECT 154.210000   0.000000 155.840000  33.975000 ;
      RECT 154.210000  33.975000 235.795000  41.925000 ;
      RECT 154.210000  41.925000 235.785000  41.935000 ;
      RECT 154.220000  41.935000 235.785000  43.050000 ;
      RECT 154.350000   0.000000 155.700000  34.115000 ;
      RECT 154.350000  34.115000 235.655000  41.870000 ;
      RECT 154.355000  41.870000 235.650000  41.875000 ;
      RECT 154.355000  41.870000 235.650000  41.875000 ;
      RECT 154.360000  41.870000 235.645000  57.985000 ;
      RECT 154.360000  41.870000 235.645000  57.985000 ;
      RECT 154.360000  41.875000 235.645000  41.880000 ;
      RECT 154.360000  41.875000 235.645000  41.880000 ;
      RECT 154.360000  41.880000 235.645000  43.190000 ;
      RECT 156.380000  33.235000 233.625000  33.975000 ;
      RECT 156.520000  33.375000 233.485000  34.115000 ;
      RECT 156.520000  33.375000 233.485000  41.870000 ;
      RECT 156.780000   0.000000 176.850000  24.370000 ;
      RECT 156.780000  24.370000 233.225000  33.235000 ;
      RECT 156.920000   0.000000 176.710000  24.510000 ;
      RECT 156.920000  24.510000 233.085000  33.375000 ;
      RECT 156.920000  24.510000 233.085000  41.870000 ;
      RECT 179.130000   0.000000 210.875000  24.370000 ;
      RECT 179.270000   0.000000 210.735000  24.510000 ;
      RECT 213.155000   0.000000 233.225000  24.370000 ;
      RECT 213.295000   0.000000 233.085000  24.510000 ;
      RECT 234.165000   0.000000 235.795000  33.975000 ;
      RECT 234.305000   0.000000 235.655000  34.115000 ;
      RECT 236.325000  42.165000 239.800000  43.050000 ;
      RECT 236.335000  35.085000 239.800000  42.155000 ;
      RECT 236.335000  42.155000 239.800000  42.165000 ;
      RECT 236.465000  42.220000 239.660000  43.190000 ;
      RECT 236.465000  42.220000 239.660000  57.985000 ;
      RECT 236.465000  42.220000 239.660000  57.985000 ;
      RECT 236.470000  42.215000 239.660000  42.220000 ;
      RECT 236.470000  42.215000 239.660000  42.220000 ;
      RECT 236.475000  35.225000 239.660000  42.210000 ;
      RECT 236.475000  35.225000 239.660000  42.220000 ;
      RECT 236.475000  35.225000 239.660000  42.220000 ;
      RECT 236.475000  42.210000 239.660000  42.215000 ;
      RECT 236.475000  42.210000 239.660000  42.215000 ;
      RECT 236.735000   0.000000 239.800000   2.130000 ;
      RECT 236.735000   2.130000 239.800000   2.175000 ;
      RECT 236.735000   3.110000 239.800000  27.815000 ;
      RECT 236.735000  27.815000 239.260000  28.355000 ;
      RECT 236.735000  28.355000 239.260000  31.160000 ;
      RECT 236.735000  31.160000 239.800000  31.700000 ;
      RECT 236.735000  31.700000 239.800000  35.085000 ;
      RECT 236.780000   2.175000 239.800000   3.065000 ;
      RECT 236.780000   3.065000 239.800000   3.110000 ;
      RECT 236.875000   0.000000 239.660000   2.075000 ;
      RECT 236.875000   3.165000 239.660000  27.760000 ;
      RECT 236.875000  27.760000 239.590000  27.830000 ;
      RECT 236.875000  27.830000 239.520000  27.900000 ;
      RECT 236.875000  27.900000 239.450000  27.970000 ;
      RECT 236.875000  27.970000 239.380000  28.040000 ;
      RECT 236.875000  28.040000 239.310000  28.110000 ;
      RECT 236.875000  28.110000 239.240000  28.180000 ;
      RECT 236.875000  28.180000 239.170000  28.250000 ;
      RECT 236.875000  28.250000 239.120000  28.300000 ;
      RECT 236.875000  28.300000 239.120000  31.215000 ;
      RECT 236.875000  31.215000 239.120000  31.285000 ;
      RECT 236.875000  31.285000 239.190000  31.355000 ;
      RECT 236.875000  31.355000 239.260000  31.425000 ;
      RECT 236.875000  31.425000 239.330000  31.495000 ;
      RECT 236.875000  31.495000 239.400000  31.565000 ;
      RECT 236.875000  31.565000 239.470000  31.635000 ;
      RECT 236.875000  31.635000 239.540000  31.705000 ;
      RECT 236.875000  31.705000 239.610000  31.755000 ;
      RECT 236.875000  31.755000 239.660000  35.225000 ;
      RECT 236.895000   2.075000 239.660000   2.095000 ;
      RECT 236.895000   3.145000 239.660000   3.165000 ;
      RECT 236.915000   2.095000 239.660000   2.115000 ;
      RECT 236.920000   2.115000 239.660000   2.120000 ;
      RECT 236.920000   2.120000 239.660000   3.120000 ;
      RECT 236.920000   3.120000 239.660000   3.145000 ;
      RECT 239.800000  28.845000 241.990000  30.665000 ;
      RECT 239.800000  30.665000 241.990000  31.205000 ;
      RECT 239.940000  28.905000 241.850000  30.610000 ;
      RECT 239.990000  28.855000 241.850000  28.905000 ;
      RECT 240.010000  30.610000 241.850000  30.680000 ;
      RECT 240.060000  28.785000 241.850000  28.855000 ;
      RECT 240.080000  30.680000 241.850000  30.750000 ;
      RECT 240.130000  28.715000 241.850000  28.785000 ;
      RECT 240.150000  30.750000 241.850000  30.820000 ;
      RECT 240.200000  28.645000 241.850000  28.715000 ;
      RECT 240.220000  30.820000 241.850000  30.890000 ;
      RECT 240.270000  28.575000 241.850000  28.645000 ;
      RECT 240.290000  30.890000 241.850000  30.960000 ;
      RECT 240.340000   0.000000 241.990000  28.310000 ;
      RECT 240.340000  28.310000 241.990000  28.845000 ;
      RECT 240.340000  28.505000 241.850000  28.575000 ;
      RECT 240.340000  31.205000 241.990000  46.275000 ;
      RECT 240.340000  46.275000 243.970000  49.755000 ;
      RECT 240.340000  49.755000 263.810000  51.985000 ;
      RECT 240.340000  51.985000 281.035000  56.395000 ;
      RECT 240.340000  56.395000 280.225000  57.205000 ;
      RECT 240.340000  57.205000 280.225000  58.665000 ;
      RECT 240.360000  30.960000 241.850000  31.030000 ;
      RECT 240.410000  28.435000 241.850000  28.505000 ;
      RECT 240.430000  31.030000 241.850000  31.100000 ;
      RECT 240.480000   0.000000 241.850000  28.365000 ;
      RECT 240.480000  28.365000 241.850000  28.435000 ;
      RECT 240.480000  31.100000 241.850000  31.150000 ;
      RECT 240.480000  31.150000 241.850000  46.415000 ;
      RECT 240.480000  46.415000 243.830000  49.895000 ;
      RECT 240.480000  46.415000 243.830000  52.125000 ;
      RECT 240.480000  46.415000 243.830000  56.340000 ;
      RECT 240.480000  46.415000 243.830000  56.340000 ;
      RECT 240.480000  46.415000 243.830000  56.340000 ;
      RECT 240.480000  49.895000 263.670000  52.125000 ;
      RECT 240.480000  49.895000 263.670000  56.340000 ;
      RECT 240.480000  49.895000 263.670000  56.340000 ;
      RECT 240.480000  49.895000 263.670000  56.340000 ;
      RECT 240.480000  52.125000 280.085000  75.105000 ;
      RECT 240.480000  52.125000 280.085000  75.105000 ;
      RECT 240.480000  52.125000 280.895000  56.340000 ;
      RECT 240.480000  56.340000 280.825000  56.410000 ;
      RECT 240.480000  56.340000 280.825000  56.410000 ;
      RECT 240.480000  56.410000 280.755000  56.480000 ;
      RECT 240.480000  56.410000 280.755000  56.480000 ;
      RECT 240.480000  56.480000 280.685000  56.550000 ;
      RECT 240.480000  56.480000 280.685000  56.550000 ;
      RECT 240.480000  56.550000 280.615000  56.620000 ;
      RECT 240.480000  56.550000 280.615000  56.620000 ;
      RECT 240.480000  56.620000 280.545000  56.690000 ;
      RECT 240.480000  56.620000 280.545000  56.690000 ;
      RECT 240.480000  56.690000 280.475000  56.760000 ;
      RECT 240.480000  56.690000 280.475000  56.760000 ;
      RECT 240.480000  56.760000 280.405000  56.830000 ;
      RECT 240.480000  56.760000 280.405000  56.830000 ;
      RECT 240.480000  56.830000 280.335000  56.900000 ;
      RECT 240.480000  56.830000 280.335000  56.900000 ;
      RECT 240.480000  56.900000 280.265000  56.970000 ;
      RECT 240.480000  56.900000 280.265000  56.970000 ;
      RECT 240.480000  56.970000 280.195000  57.040000 ;
      RECT 240.480000  56.970000 280.195000  57.040000 ;
      RECT 240.480000  57.040000 280.125000  57.110000 ;
      RECT 240.480000  57.040000 280.125000  57.110000 ;
      RECT 240.480000  57.110000 280.085000  57.150000 ;
      RECT 240.480000  57.110000 280.085000  57.150000 ;
      RECT 240.480000  57.150000 280.085000  58.805000 ;
      RECT 242.530000  27.115000 243.970000  28.560000 ;
      RECT 242.530000  28.560000 243.970000  46.275000 ;
      RECT 242.670000  27.525000 242.740000  27.595000 ;
      RECT 242.670000  27.595000 242.810000  27.665000 ;
      RECT 242.670000  27.665000 242.880000  27.735000 ;
      RECT 242.670000  27.735000 242.950000  27.805000 ;
      RECT 242.670000  27.805000 243.020000  27.875000 ;
      RECT 242.670000  27.875000 243.090000  27.945000 ;
      RECT 242.670000  27.945000 243.160000  28.015000 ;
      RECT 242.670000  28.015000 243.230000  28.085000 ;
      RECT 242.670000  28.085000 243.300000  28.155000 ;
      RECT 242.670000  28.155000 243.370000  28.225000 ;
      RECT 242.670000  28.225000 243.440000  28.295000 ;
      RECT 242.670000  28.295000 243.510000  28.365000 ;
      RECT 242.670000  28.365000 243.580000  28.435000 ;
      RECT 242.670000  28.435000 243.650000  28.505000 ;
      RECT 242.670000  28.505000 243.720000  28.575000 ;
      RECT 242.670000  28.575000 243.790000  28.615000 ;
      RECT 242.670000  28.615000 243.830000  46.415000 ;
      RECT 242.930000   0.000000 247.200000  10.730000 ;
      RECT 242.930000  10.730000 254.030000  26.750000 ;
      RECT 242.930000  26.750000 254.030000  28.330000 ;
      RECT 243.070000   0.000000 247.060000  10.870000 ;
      RECT 243.070000   0.000000 247.060000  26.695000 ;
      RECT 243.070000  10.870000 253.890000  26.695000 ;
      RECT 243.140000  26.695000 253.890000  26.765000 ;
      RECT 243.140000  26.695000 253.890000  26.765000 ;
      RECT 243.210000  26.765000 253.890000  26.835000 ;
      RECT 243.210000  26.765000 253.890000  26.835000 ;
      RECT 243.280000  26.835000 253.890000  26.905000 ;
      RECT 243.280000  26.835000 253.890000  26.905000 ;
      RECT 243.350000  26.905000 253.890000  26.975000 ;
      RECT 243.350000  26.905000 253.890000  26.975000 ;
      RECT 243.420000  26.975000 253.890000  27.045000 ;
      RECT 243.420000  26.975000 253.890000  27.045000 ;
      RECT 243.490000  27.045000 253.890000  27.115000 ;
      RECT 243.490000  27.045000 253.890000  27.115000 ;
      RECT 243.560000  27.115000 253.890000  27.185000 ;
      RECT 243.560000  27.115000 253.890000  27.185000 ;
      RECT 243.630000  27.185000 253.890000  27.255000 ;
      RECT 243.630000  27.185000 253.890000  27.255000 ;
      RECT 243.700000  27.255000 253.890000  27.325000 ;
      RECT 243.700000  27.255000 253.890000  27.325000 ;
      RECT 243.770000  27.325000 253.890000  27.395000 ;
      RECT 243.770000  27.325000 253.890000  27.395000 ;
      RECT 243.840000  27.395000 253.890000  27.465000 ;
      RECT 243.840000  27.395000 253.890000  27.465000 ;
      RECT 243.910000  27.465000 253.890000  27.535000 ;
      RECT 243.910000  27.465000 253.890000  27.535000 ;
      RECT 243.980000  27.535000 253.890000  27.605000 ;
      RECT 243.980000  27.535000 253.890000  27.605000 ;
      RECT 244.050000  27.605000 253.890000  27.675000 ;
      RECT 244.050000  27.605000 253.890000  27.675000 ;
      RECT 244.120000  27.675000 253.890000  27.745000 ;
      RECT 244.120000  27.675000 253.890000  27.745000 ;
      RECT 244.190000  27.745000 253.890000  27.815000 ;
      RECT 244.190000  27.745000 253.890000  27.815000 ;
      RECT 244.260000  27.815000 253.890000  27.885000 ;
      RECT 244.260000  27.815000 253.890000  27.885000 ;
      RECT 244.330000  27.885000 253.890000  27.955000 ;
      RECT 244.330000  27.885000 253.890000  27.955000 ;
      RECT 244.400000  27.955000 253.890000  28.025000 ;
      RECT 244.400000  27.955000 253.890000  28.025000 ;
      RECT 244.470000  28.025000 253.890000  28.095000 ;
      RECT 244.470000  28.025000 253.890000  28.095000 ;
      RECT 244.510000  28.330000 254.030000  37.090000 ;
      RECT 244.510000  37.090000 255.470000  42.880000 ;
      RECT 244.510000  42.880000 260.985000  43.050000 ;
      RECT 244.510000  43.050000 268.150000  45.780000 ;
      RECT 244.510000  45.780000 268.050000  45.880000 ;
      RECT 244.510000  45.880000 263.950000  47.300000 ;
      RECT 244.510000  47.300000 263.950000  48.770000 ;
      RECT 244.510000  48.770000 263.810000  48.910000 ;
      RECT 244.510000  48.910000 263.810000  49.170000 ;
      RECT 244.510000  49.170000 263.810000  49.215000 ;
      RECT 244.540000  28.095000 253.890000  28.165000 ;
      RECT 244.540000  28.095000 253.890000  28.165000 ;
      RECT 244.610000  28.165000 253.890000  28.235000 ;
      RECT 244.610000  28.165000 253.890000  28.235000 ;
      RECT 244.650000  10.870000 253.890000  37.230000 ;
      RECT 244.650000  28.235000 253.890000  28.275000 ;
      RECT 244.650000  28.235000 253.890000  28.275000 ;
      RECT 244.650000  28.275000 253.890000  37.230000 ;
      RECT 244.650000  37.230000 255.330000  43.020000 ;
      RECT 244.650000  37.230000 255.330000  43.190000 ;
      RECT 244.650000  37.230000 255.330000  43.190000 ;
      RECT 244.650000  37.230000 255.330000  43.190000 ;
      RECT 244.650000  43.020000 260.845000  43.190000 ;
      RECT 244.650000  43.190000 268.010000  45.740000 ;
      RECT 244.650000  45.740000 265.245000  45.810000 ;
      RECT 244.650000  45.740000 265.245000  45.810000 ;
      RECT 244.650000  45.810000 265.175000  45.880000 ;
      RECT 244.650000  45.810000 265.175000  45.880000 ;
      RECT 244.650000  45.880000 265.105000  45.950000 ;
      RECT 244.650000  45.880000 265.105000  45.950000 ;
      RECT 244.650000  45.950000 265.035000  46.020000 ;
      RECT 244.650000  45.950000 265.035000  46.020000 ;
      RECT 244.650000  46.020000 264.965000  46.090000 ;
      RECT 244.650000  46.020000 264.965000  46.090000 ;
      RECT 244.650000  46.090000 264.895000  46.160000 ;
      RECT 244.650000  46.090000 264.895000  46.160000 ;
      RECT 244.650000  46.160000 264.825000  46.230000 ;
      RECT 244.650000  46.160000 264.825000  46.230000 ;
      RECT 244.650000  46.230000 264.755000  46.300000 ;
      RECT 244.650000  46.230000 264.755000  46.300000 ;
      RECT 244.650000  46.300000 264.685000  46.370000 ;
      RECT 244.650000  46.300000 264.685000  46.370000 ;
      RECT 244.650000  46.370000 264.615000  46.440000 ;
      RECT 244.650000  46.370000 264.615000  46.440000 ;
      RECT 244.650000  46.440000 264.545000  46.510000 ;
      RECT 244.650000  46.440000 264.545000  46.510000 ;
      RECT 244.650000  46.510000 264.475000  46.580000 ;
      RECT 244.650000  46.510000 264.475000  46.580000 ;
      RECT 244.650000  46.580000 264.405000  46.650000 ;
      RECT 244.650000  46.580000 264.405000  46.650000 ;
      RECT 244.650000  46.650000 264.335000  46.720000 ;
      RECT 244.650000  46.650000 264.335000  46.720000 ;
      RECT 244.650000  46.720000 264.265000  46.790000 ;
      RECT 244.650000  46.720000 264.265000  46.790000 ;
      RECT 244.650000  46.790000 264.195000  46.860000 ;
      RECT 244.650000  46.790000 264.195000  46.860000 ;
      RECT 244.650000  46.860000 264.125000  46.930000 ;
      RECT 244.650000  46.860000 264.125000  46.930000 ;
      RECT 244.650000  46.930000 264.055000  47.000000 ;
      RECT 244.650000  46.930000 264.055000  47.000000 ;
      RECT 244.650000  47.000000 263.985000  47.070000 ;
      RECT 244.650000  47.000000 263.985000  47.070000 ;
      RECT 244.650000  47.070000 263.915000  47.140000 ;
      RECT 244.650000  47.070000 263.915000  47.140000 ;
      RECT 244.650000  47.140000 263.845000  47.210000 ;
      RECT 244.650000  47.140000 263.845000  47.210000 ;
      RECT 244.650000  47.210000 263.810000  47.245000 ;
      RECT 244.650000  47.210000 263.810000  47.245000 ;
      RECT 244.650000  47.245000 263.810000  48.715000 ;
      RECT 244.650000  48.715000 263.740000  48.785000 ;
      RECT 244.650000  48.715000 263.740000  48.785000 ;
      RECT 244.650000  48.785000 263.670000  48.855000 ;
      RECT 244.650000  48.785000 263.670000  48.855000 ;
      RECT 244.650000  48.855000 247.655000  49.075000 ;
      RECT 244.890000  49.215000 263.810000  49.755000 ;
      RECT 245.030000  48.715000 263.670000  56.340000 ;
      RECT 245.030000  48.715000 263.670000  56.340000 ;
      RECT 245.030000  48.715000 263.670000  56.340000 ;
      RECT 247.740000   7.720000 254.030000  10.730000 ;
      RECT 247.880000   7.860000 253.890000  10.870000 ;
      RECT 247.880000   7.860000 253.890000  26.695000 ;
      RECT 247.880000   7.860000 253.890000  26.695000 ;
      RECT 248.140000   0.000000 248.320000   1.935000 ;
      RECT 248.140000   1.935000 248.230000   2.025000 ;
      RECT 248.140000   2.025000 248.230000   2.485000 ;
      RECT 248.140000   2.485000 254.030000   7.720000 ;
      RECT 248.280000   2.625000 253.890000  10.870000 ;
      RECT 248.280000   2.625000 253.890000  10.870000 ;
      RECT 248.280000   2.625000 254.030000   6.100000 ;
      RECT 248.280000   6.100000 253.890000   7.860000 ;
      RECT 248.945000   0.000000 254.030000   1.820000 ;
      RECT 248.945000   1.820000 254.030000   2.025000 ;
      RECT 249.085000   0.000000 249.290000   1.765000 ;
      RECT 249.150000   2.025000 254.030000   2.485000 ;
      RECT 249.155000   1.765000 254.030000   1.835000 ;
      RECT 249.225000   1.835000 254.030000   1.905000 ;
      RECT 249.290000   0.000000 253.890000   1.570000 ;
      RECT 249.290000   1.570000 254.030000   1.765000 ;
      RECT 249.290000   1.765000 254.030000   1.970000 ;
      RECT 249.290000   1.905000 254.030000   1.970000 ;
      RECT 249.290000   1.970000 254.030000   2.625000 ;
      RECT 254.570000  29.150000 254.960000  29.540000 ;
      RECT 254.570000  29.540000 254.960000  30.025000 ;
      RECT 254.570000  30.025000 255.315000  30.385000 ;
      RECT 254.570000  30.385000 255.470000  30.430000 ;
      RECT 254.570000  30.430000 255.470000  36.505000 ;
      RECT 254.570000  36.505000 255.470000  36.550000 ;
      RECT 254.710000  30.045000 254.780000  30.115000 ;
      RECT 254.710000  30.115000 254.850000  30.185000 ;
      RECT 254.710000  30.185000 254.920000  30.255000 ;
      RECT 254.710000  30.255000 254.990000  30.325000 ;
      RECT 254.710000  30.325000 255.060000  30.395000 ;
      RECT 254.710000  30.395000 255.130000  30.465000 ;
      RECT 254.710000  30.465000 255.200000  30.525000 ;
      RECT 254.710000  30.525000 255.330000  36.410000 ;
      RECT 254.950000  36.550000 255.470000  37.090000 ;
      RECT 254.970000   0.000000 261.480000  10.235000 ;
      RECT 254.970000   2.610000 261.340000   7.810000 ;
      RECT 254.970000  10.235000 262.345000  11.100000 ;
      RECT 254.970000  11.100000 262.345000  23.605000 ;
      RECT 254.970000  23.605000 261.745000  24.205000 ;
      RECT 254.970000  24.205000 261.745000  28.780000 ;
      RECT 254.970000  28.780000 261.745000  29.310000 ;
      RECT 255.090000  36.410000 255.330000  37.230000 ;
      RECT 255.110000   0.000000 261.340000   3.005000 ;
      RECT 255.110000   2.610000 261.340000  11.155000 ;
      RECT 255.110000   2.610000 261.340000  11.155000 ;
      RECT 255.110000   2.610000 261.340000  11.155000 ;
      RECT 255.110000   7.810000 261.340000  10.290000 ;
      RECT 255.110000  10.290000 261.340000  10.360000 ;
      RECT 255.110000  10.290000 261.340000  10.360000 ;
      RECT 255.110000  10.360000 261.410000  10.430000 ;
      RECT 255.110000  10.360000 261.410000  10.430000 ;
      RECT 255.110000  10.430000 261.480000  10.500000 ;
      RECT 255.110000  10.430000 261.480000  10.500000 ;
      RECT 255.110000  10.500000 261.550000  10.570000 ;
      RECT 255.110000  10.500000 261.550000  10.570000 ;
      RECT 255.110000  10.570000 261.620000  10.640000 ;
      RECT 255.110000  10.570000 261.620000  10.640000 ;
      RECT 255.110000  10.640000 261.690000  10.710000 ;
      RECT 255.110000  10.640000 261.690000  10.710000 ;
      RECT 255.110000  10.710000 261.760000  10.780000 ;
      RECT 255.110000  10.710000 261.760000  10.780000 ;
      RECT 255.110000  10.780000 261.830000  10.850000 ;
      RECT 255.110000  10.780000 261.830000  10.850000 ;
      RECT 255.110000  10.850000 261.900000  10.920000 ;
      RECT 255.110000  10.850000 261.900000  10.920000 ;
      RECT 255.110000  10.920000 261.970000  10.990000 ;
      RECT 255.110000  10.920000 261.970000  10.990000 ;
      RECT 255.110000  10.990000 262.040000  11.060000 ;
      RECT 255.110000  10.990000 262.040000  11.060000 ;
      RECT 255.110000  11.060000 262.110000  11.130000 ;
      RECT 255.110000  11.060000 262.110000  11.130000 ;
      RECT 255.110000  11.130000 262.180000  11.155000 ;
      RECT 255.110000  11.130000 262.180000  11.155000 ;
      RECT 255.110000  11.155000 262.205000  23.550000 ;
      RECT 255.110000  23.550000 262.135000  23.620000 ;
      RECT 255.110000  23.550000 262.135000  23.620000 ;
      RECT 255.110000  23.620000 262.065000  23.690000 ;
      RECT 255.110000  23.620000 262.065000  23.690000 ;
      RECT 255.110000  23.690000 261.995000  23.760000 ;
      RECT 255.110000  23.690000 261.995000  23.760000 ;
      RECT 255.110000  23.760000 261.925000  23.830000 ;
      RECT 255.110000  23.760000 261.925000  23.830000 ;
      RECT 255.110000  23.830000 261.855000  23.900000 ;
      RECT 255.110000  23.830000 261.855000  23.900000 ;
      RECT 255.110000  23.900000 261.785000  23.970000 ;
      RECT 255.110000  23.900000 261.785000  23.970000 ;
      RECT 255.110000  23.970000 261.715000  24.040000 ;
      RECT 255.110000  23.970000 261.715000  24.040000 ;
      RECT 255.110000  24.040000 261.645000  24.110000 ;
      RECT 255.110000  24.040000 261.645000  24.110000 ;
      RECT 255.110000  24.110000 261.605000  24.150000 ;
      RECT 255.110000  24.110000 261.605000  24.150000 ;
      RECT 255.110000  24.150000 261.605000  28.725000 ;
      RECT 255.180000  28.725000 261.605000  28.795000 ;
      RECT 255.180000  28.725000 261.605000  28.795000 ;
      RECT 255.250000  28.795000 261.605000  28.865000 ;
      RECT 255.250000  28.795000 261.605000  28.865000 ;
      RECT 255.320000  28.865000 261.605000  28.935000 ;
      RECT 255.320000  28.865000 261.605000  28.935000 ;
      RECT 255.390000  28.935000 261.605000  29.005000 ;
      RECT 255.390000  28.935000 261.605000  29.005000 ;
      RECT 255.460000  29.005000 261.605000  29.075000 ;
      RECT 255.460000  29.005000 261.605000  29.075000 ;
      RECT 255.500000  29.310000 261.745000  29.800000 ;
      RECT 255.500000  29.800000 261.745000  29.845000 ;
      RECT 255.530000  29.075000 261.605000  29.145000 ;
      RECT 255.530000  29.075000 261.605000  29.145000 ;
      RECT 255.600000  29.145000 261.605000  29.215000 ;
      RECT 255.600000  29.145000 261.605000  29.215000 ;
      RECT 255.640000  24.150000 261.605000  29.705000 ;
      RECT 255.640000  29.215000 261.605000  29.255000 ;
      RECT 255.640000  29.215000 261.605000  29.255000 ;
      RECT 255.710000  29.255000 261.605000  29.325000 ;
      RECT 255.710000  29.255000 261.605000  29.325000 ;
      RECT 255.780000  29.325000 261.605000  29.395000 ;
      RECT 255.780000  29.325000 261.605000  29.395000 ;
      RECT 255.850000  29.395000 261.605000  29.465000 ;
      RECT 255.850000  29.395000 261.605000  29.465000 ;
      RECT 255.920000  29.465000 261.605000  29.535000 ;
      RECT 255.920000  29.465000 261.605000  29.535000 ;
      RECT 255.990000  29.535000 261.605000  29.605000 ;
      RECT 255.990000  29.535000 261.605000  29.605000 ;
      RECT 256.010000  30.430000 261.745000  42.465000 ;
      RECT 256.010000  42.465000 261.700000  42.510000 ;
      RECT 256.010000  42.510000 260.985000  42.880000 ;
      RECT 256.055000  30.385000 261.745000  30.430000 ;
      RECT 256.060000  29.605000 261.605000  29.675000 ;
      RECT 256.060000  29.605000 261.605000  29.675000 ;
      RECT 256.090000  29.675000 261.605000  29.705000 ;
      RECT 256.090000  29.675000 261.605000  29.705000 ;
      RECT 256.150000  30.525000 261.605000  42.370000 ;
      RECT 256.150000  42.370000 260.845000  43.020000 ;
      RECT 256.390000  29.845000 261.745000  30.385000 ;
      RECT 256.530000  24.150000 261.605000  42.370000 ;
      RECT 256.530000  29.705000 261.605000  30.525000 ;
      RECT 262.020000   0.000000 268.150000  10.005000 ;
      RECT 262.020000  10.005000 268.150000  10.870000 ;
      RECT 262.025000   2.610000 268.010000   7.810000 ;
      RECT 262.160000   0.000000 268.010000   2.610000 ;
      RECT 262.160000   0.000000 268.010000   7.810000 ;
      RECT 262.160000   0.000000 268.010000   7.810000 ;
      RECT 262.160000   7.810000 268.010000   9.950000 ;
      RECT 262.230000   9.950000 268.010000  10.020000 ;
      RECT 262.230000   9.950000 268.010000  10.020000 ;
      RECT 262.285000  24.435000 268.150000  43.050000 ;
      RECT 262.300000  10.020000 268.010000  10.090000 ;
      RECT 262.300000  10.020000 268.010000  10.090000 ;
      RECT 262.370000  10.090000 268.010000  10.160000 ;
      RECT 262.370000  10.090000 268.010000  10.160000 ;
      RECT 262.425000  24.490000 268.010000  43.190000 ;
      RECT 262.425000  24.490000 268.010000  45.740000 ;
      RECT 262.425000  24.490000 268.010000  45.740000 ;
      RECT 262.425000  24.490000 268.010000  45.740000 ;
      RECT 262.425000  24.490000 268.010000  45.740000 ;
      RECT 262.440000  10.160000 268.010000  10.230000 ;
      RECT 262.440000  10.160000 268.010000  10.230000 ;
      RECT 262.465000  24.450000 268.010000  24.490000 ;
      RECT 262.465000  24.450000 268.010000  24.490000 ;
      RECT 262.510000  10.230000 268.010000  10.300000 ;
      RECT 262.510000  10.230000 268.010000  10.300000 ;
      RECT 262.535000  24.380000 268.010000  24.450000 ;
      RECT 262.535000  24.380000 268.010000  24.450000 ;
      RECT 262.580000  10.300000 268.010000  10.370000 ;
      RECT 262.580000  10.300000 268.010000  10.370000 ;
      RECT 262.605000  24.310000 268.010000  24.380000 ;
      RECT 262.605000  24.310000 268.010000  24.380000 ;
      RECT 262.650000  10.370000 268.010000  10.440000 ;
      RECT 262.650000  10.370000 268.010000  10.440000 ;
      RECT 262.675000  24.240000 268.010000  24.310000 ;
      RECT 262.675000  24.240000 268.010000  24.310000 ;
      RECT 262.720000  10.440000 268.010000  10.510000 ;
      RECT 262.720000  10.440000 268.010000  10.510000 ;
      RECT 262.745000  24.170000 268.010000  24.240000 ;
      RECT 262.745000  24.170000 268.010000  24.240000 ;
      RECT 262.790000  10.510000 268.010000  10.580000 ;
      RECT 262.790000  10.510000 268.010000  10.580000 ;
      RECT 262.815000  24.100000 268.010000  24.170000 ;
      RECT 262.815000  24.100000 268.010000  24.170000 ;
      RECT 262.860000  10.580000 268.010000  10.650000 ;
      RECT 262.860000  10.580000 268.010000  10.650000 ;
      RECT 262.885000  10.870000 268.150000  23.830000 ;
      RECT 262.885000  23.830000 268.150000  24.435000 ;
      RECT 262.885000  24.030000 268.010000  24.100000 ;
      RECT 262.885000  24.030000 268.010000  24.100000 ;
      RECT 262.930000  10.650000 268.010000  10.720000 ;
      RECT 262.930000  10.650000 268.010000  10.720000 ;
      RECT 262.955000  23.960000 268.010000  24.030000 ;
      RECT 262.955000  23.960000 268.010000  24.030000 ;
      RECT 263.000000  10.720000 268.010000  10.790000 ;
      RECT 263.000000  10.720000 268.010000  10.790000 ;
      RECT 263.025000   9.950000 268.010000  23.890000 ;
      RECT 263.025000   9.950000 268.010000  23.890000 ;
      RECT 263.025000  10.790000 268.010000  10.815000 ;
      RECT 263.025000  10.790000 268.010000  10.815000 ;
      RECT 263.025000  10.815000 268.010000  23.890000 ;
      RECT 263.025000  23.890000 268.010000  23.960000 ;
      RECT 263.025000  23.890000 268.010000  23.960000 ;
      RECT 264.490000  47.530000 281.035000  47.630000 ;
      RECT 264.490000  47.630000 281.035000  48.605000 ;
      RECT 264.490000  48.605000 281.035000  48.910000 ;
      RECT 264.630000  47.585000 280.795000  47.635000 ;
      RECT 264.630000  47.635000 280.845000  47.685000 ;
      RECT 264.630000  47.680000 280.885000  47.685000 ;
      RECT 264.630000  47.680000 280.885000  47.685000 ;
      RECT 264.630000  47.685000 280.895000  48.145000 ;
      RECT 264.630000  48.145000 280.895000  48.550000 ;
      RECT 264.635000  47.675000 280.885000  47.680000 ;
      RECT 264.635000  47.675000 280.885000  47.680000 ;
      RECT 264.655000  47.560000 280.770000  47.585000 ;
      RECT 264.670000  47.630000 280.840000  47.675000 ;
      RECT 264.670000  47.630000 280.840000  47.675000 ;
      RECT 264.700000  48.550000 280.895000  48.620000 ;
      RECT 264.700000  48.550000 280.895000  48.620000 ;
      RECT 264.710000  47.585000 280.795000  47.630000 ;
      RECT 264.710000  47.585000 280.795000  47.630000 ;
      RECT 264.725000  47.490000 280.700000  47.560000 ;
      RECT 264.760000  47.525000 280.735000  47.585000 ;
      RECT 264.760000  47.525000 280.735000  47.585000 ;
      RECT 264.770000  48.620000 280.895000  48.690000 ;
      RECT 264.770000  48.620000 280.895000  48.690000 ;
      RECT 264.795000  47.420000 280.630000  47.490000 ;
      RECT 264.795000  48.910000 281.035000  51.985000 ;
      RECT 264.820000  47.455000 280.665000  47.525000 ;
      RECT 264.820000  47.455000 280.665000  47.525000 ;
      RECT 264.840000  48.690000 280.895000  48.760000 ;
      RECT 264.840000  48.690000 280.895000  48.760000 ;
      RECT 264.865000  47.350000 280.560000  47.420000 ;
      RECT 264.880000  47.385000 280.595000  47.455000 ;
      RECT 264.880000  47.385000 280.595000  47.455000 ;
      RECT 264.910000  48.760000 280.895000  48.830000 ;
      RECT 264.910000  48.760000 280.895000  48.830000 ;
      RECT 264.935000  47.280000 280.490000  47.350000 ;
      RECT 264.935000  47.685000 280.895000  56.340000 ;
      RECT 264.935000  47.685000 280.895000  56.340000 ;
      RECT 264.935000  47.685000 280.895000  56.340000 ;
      RECT 264.935000  48.830000 280.895000  48.855000 ;
      RECT 264.935000  48.830000 280.895000  48.855000 ;
      RECT 264.940000  47.315000 280.525000  47.385000 ;
      RECT 264.940000  47.315000 280.525000  47.385000 ;
      RECT 265.000000  47.245000 280.455000  47.315000 ;
      RECT 265.000000  47.245000 280.455000  47.315000 ;
      RECT 265.005000  47.210000 280.420000  47.280000 ;
      RECT 265.060000  47.175000 280.385000  47.245000 ;
      RECT 265.060000  47.175000 280.385000  47.245000 ;
      RECT 265.075000  47.140000 280.350000  47.210000 ;
      RECT 265.120000  47.105000 280.315000  47.175000 ;
      RECT 265.120000  47.105000 280.315000  47.175000 ;
      RECT 265.145000  47.070000 280.280000  47.140000 ;
      RECT 265.180000  47.035000 280.245000  47.105000 ;
      RECT 265.180000  47.035000 280.245000  47.105000 ;
      RECT 265.215000  47.000000 280.210000  47.035000 ;
      RECT 265.215000  47.000000 280.210000  47.035000 ;
      RECT 265.215000  47.000000 280.210000  47.070000 ;
      RECT 265.285000  46.735000 280.935000  47.530000 ;
      RECT 265.285000  46.930000 280.140000  47.000000 ;
      RECT 265.285000  46.930000 280.140000  47.000000 ;
      RECT 265.285000  46.930000 280.140000  47.000000 ;
      RECT 265.355000  46.860000 280.070000  46.930000 ;
      RECT 265.355000  46.860000 280.070000  46.930000 ;
      RECT 265.355000  46.860000 280.070000  46.930000 ;
      RECT 265.425000  46.790000 280.000000  46.860000 ;
      RECT 265.425000  46.790000 280.000000  46.860000 ;
      RECT 265.425000  46.790000 280.000000  46.860000 ;
      RECT 265.445000  46.770000 280.000000  46.790000 ;
      RECT 265.445000  46.770000 280.000000  46.790000 ;
      RECT 265.515000  46.700000 280.000000  46.770000 ;
      RECT 265.515000  46.700000 280.000000  46.770000 ;
      RECT 265.585000  46.630000 280.000000  46.700000 ;
      RECT 265.585000  46.630000 280.000000  46.700000 ;
      RECT 265.600000  46.420000 280.140000  46.735000 ;
      RECT 265.655000  46.560000 280.000000  46.630000 ;
      RECT 265.655000  46.560000 280.000000  46.630000 ;
      RECT 268.690000   0.000000 279.515000  17.525000 ;
      RECT 268.690000  17.525000 279.790000  17.795000 ;
      RECT 268.690000  17.795000 279.790000  36.240000 ;
      RECT 268.690000  36.240000 279.770000  36.260000 ;
      RECT 268.690000  36.260000 279.770000  45.650000 ;
      RECT 268.690000  45.650000 280.140000  46.020000 ;
      RECT 268.690000  46.020000 280.140000  46.420000 ;
      RECT 268.830000   0.000000 279.375000  17.580000 ;
      RECT 268.830000  17.580000 279.375000  17.650000 ;
      RECT 268.830000  17.580000 279.375000  17.650000 ;
      RECT 268.830000  17.650000 279.445000  17.720000 ;
      RECT 268.830000  17.650000 279.445000  17.720000 ;
      RECT 268.830000  17.720000 279.515000  17.790000 ;
      RECT 268.830000  17.720000 279.515000  17.790000 ;
      RECT 268.830000  17.790000 279.585000  17.855000 ;
      RECT 268.830000  17.790000 279.585000  17.855000 ;
      RECT 268.830000  17.855000 279.650000  36.185000 ;
      RECT 268.830000  36.185000 279.640000  36.195000 ;
      RECT 268.830000  36.185000 279.640000  36.195000 ;
      RECT 268.830000  36.195000 279.630000  36.205000 ;
      RECT 268.830000  36.195000 279.630000  36.205000 ;
      RECT 268.830000  36.205000 279.630000  46.790000 ;
      RECT 268.830000  36.205000 279.630000  46.790000 ;
      RECT 268.830000  45.705000 279.630000  45.775000 ;
      RECT 268.830000  45.705000 279.630000  45.775000 ;
      RECT 268.830000  45.775000 279.700000  45.845000 ;
      RECT 268.830000  45.775000 279.700000  45.845000 ;
      RECT 268.830000  45.845000 279.770000  45.915000 ;
      RECT 268.830000  45.845000 279.770000  45.915000 ;
      RECT 268.830000  45.915000 279.840000  45.985000 ;
      RECT 268.830000  45.915000 279.840000  45.985000 ;
      RECT 268.830000  45.985000 279.910000  46.055000 ;
      RECT 268.830000  45.985000 279.910000  46.055000 ;
      RECT 268.830000  46.055000 279.980000  46.075000 ;
      RECT 268.830000  46.055000 279.980000  46.075000 ;
      RECT 268.830000  46.075000 280.000000  46.560000 ;
      RECT 280.055000   0.000000 282.895000   1.180000 ;
      RECT 280.055000   1.180000 282.180000   1.895000 ;
      RECT 280.055000   1.895000 282.180000  17.295000 ;
      RECT 280.055000  17.295000 282.180000  17.570000 ;
      RECT 280.195000   0.000000 282.755000   1.125000 ;
      RECT 280.195000   1.125000 282.685000   1.195000 ;
      RECT 280.195000   1.195000 282.615000   1.265000 ;
      RECT 280.195000   1.265000 282.545000   1.335000 ;
      RECT 280.195000   1.335000 282.475000   1.405000 ;
      RECT 280.195000   1.405000 282.405000   1.475000 ;
      RECT 280.195000   1.475000 282.335000   1.545000 ;
      RECT 280.195000   1.545000 282.265000   1.615000 ;
      RECT 280.195000   1.615000 282.195000   1.685000 ;
      RECT 280.195000   1.685000 282.125000   1.755000 ;
      RECT 280.195000   1.755000 282.055000   1.825000 ;
      RECT 280.195000   1.825000 282.040000   1.840000 ;
      RECT 280.195000   1.840000 282.040000   2.680000 ;
      RECT 280.195000   2.680000 282.070000   7.155000 ;
      RECT 280.195000   7.155000 282.040000  17.240000 ;
      RECT 280.265000  17.240000 282.040000  17.310000 ;
      RECT 280.310000  36.490000 447.765000  45.420000 ;
      RECT 280.310000  45.420000 447.765000  45.790000 ;
      RECT 280.330000  17.570000 282.180000  18.295000 ;
      RECT 280.330000  18.295000 302.770000  33.375000 ;
      RECT 280.330000  33.375000 447.765000  36.470000 ;
      RECT 280.330000  36.470000 447.765000  36.490000 ;
      RECT 280.335000  17.310000 282.040000  17.380000 ;
      RECT 280.405000  17.380000 282.040000  17.450000 ;
      RECT 280.450000  36.545000 447.625000  45.365000 ;
      RECT 280.460000  36.535000 447.625000  36.545000 ;
      RECT 280.460000  36.535000 447.625000  36.545000 ;
      RECT 280.470000  17.450000 282.040000  17.515000 ;
      RECT 280.470000  17.515000 282.040000  18.435000 ;
      RECT 280.470000  18.435000 302.630000  33.515000 ;
      RECT 280.470000  18.435000 302.630000  36.525000 ;
      RECT 280.470000  33.515000 447.625000  36.525000 ;
      RECT 280.470000  33.515000 447.625000  45.365000 ;
      RECT 280.470000  36.525000 447.625000  36.535000 ;
      RECT 280.470000  36.525000 447.625000  36.535000 ;
      RECT 280.520000  45.365000 447.625000  45.435000 ;
      RECT 280.520000  45.365000 447.625000  45.435000 ;
      RECT 280.590000  45.435000 447.625000  45.505000 ;
      RECT 280.590000  45.435000 447.625000  45.505000 ;
      RECT 280.660000  45.505000 447.625000  45.575000 ;
      RECT 280.660000  45.505000 447.625000  45.575000 ;
      RECT 280.680000  45.790000 447.765000  46.505000 ;
      RECT 280.680000  46.505000 447.765000  47.400000 ;
      RECT 280.730000  45.575000 447.625000  45.645000 ;
      RECT 280.730000  45.575000 447.625000  45.645000 ;
      RECT 280.765000  57.435000 447.765000  74.820000 ;
      RECT 280.765000  74.820000 447.765000  76.450000 ;
      RECT 280.800000  45.645000 447.625000  45.715000 ;
      RECT 280.800000  45.645000 447.625000  45.715000 ;
      RECT 280.820000  45.715000 447.625000  45.735000 ;
      RECT 280.820000  45.715000 447.625000  45.735000 ;
      RECT 280.820000  45.735000 447.625000  46.450000 ;
      RECT 280.890000  46.450000 447.625000  46.520000 ;
      RECT 280.890000  46.450000 447.625000  46.520000 ;
      RECT 280.905000  57.490000 447.625000  74.765000 ;
      RECT 280.945000  57.450000 447.625000  57.490000 ;
      RECT 280.945000  57.450000 447.625000  57.490000 ;
      RECT 280.960000  46.520000 447.625000  46.590000 ;
      RECT 280.960000  46.520000 447.625000  46.590000 ;
      RECT 280.975000  74.765000 447.625000  74.835000 ;
      RECT 280.975000  74.765000 447.625000  74.835000 ;
      RECT 281.015000  57.380000 447.625000  57.450000 ;
      RECT 281.015000  57.380000 447.625000  57.450000 ;
      RECT 281.030000  46.590000 447.625000  46.660000 ;
      RECT 281.030000  46.590000 447.625000  46.660000 ;
      RECT 281.045000  74.835000 447.625000  74.905000 ;
      RECT 281.045000  74.835000 447.625000  74.905000 ;
      RECT 281.085000  57.310000 447.625000  57.380000 ;
      RECT 281.085000  57.310000 447.625000  57.380000 ;
      RECT 281.100000  46.660000 447.625000  46.730000 ;
      RECT 281.100000  46.660000 447.625000  46.730000 ;
      RECT 281.115000  74.905000 447.625000  74.975000 ;
      RECT 281.115000  74.905000 447.625000  74.975000 ;
      RECT 281.155000  57.240000 447.625000  57.310000 ;
      RECT 281.155000  57.240000 447.625000  57.310000 ;
      RECT 281.170000  46.730000 447.625000  46.800000 ;
      RECT 281.170000  46.730000 447.625000  46.800000 ;
      RECT 281.185000  74.975000 447.625000  75.045000 ;
      RECT 281.185000  74.975000 447.625000  75.045000 ;
      RECT 281.225000  57.170000 447.625000  57.240000 ;
      RECT 281.225000  57.170000 447.625000  57.240000 ;
      RECT 281.240000  46.800000 447.625000  46.870000 ;
      RECT 281.240000  46.800000 447.625000  46.870000 ;
      RECT 281.255000  75.045000 447.625000  75.115000 ;
      RECT 281.255000  75.045000 447.625000  75.115000 ;
      RECT 281.295000  57.100000 447.625000  57.170000 ;
      RECT 281.295000  57.100000 447.625000  57.170000 ;
      RECT 281.310000  46.870000 447.625000  46.940000 ;
      RECT 281.310000  46.870000 447.625000  46.940000 ;
      RECT 281.325000  75.115000 447.625000  75.185000 ;
      RECT 281.325000  75.115000 447.625000  75.185000 ;
      RECT 281.365000  57.030000 447.625000  57.100000 ;
      RECT 281.365000  57.030000 447.625000  57.100000 ;
      RECT 281.380000  46.940000 447.625000  47.010000 ;
      RECT 281.380000  46.940000 447.625000  47.010000 ;
      RECT 281.395000  75.185000 447.625000  75.255000 ;
      RECT 281.395000  75.185000 447.625000  75.255000 ;
      RECT 281.435000  56.960000 447.625000  57.030000 ;
      RECT 281.435000  56.960000 447.625000  57.030000 ;
      RECT 281.450000  47.010000 447.625000  47.080000 ;
      RECT 281.450000  47.010000 447.625000  47.080000 ;
      RECT 281.465000  75.255000 447.625000  75.325000 ;
      RECT 281.465000  75.255000 447.625000  75.325000 ;
      RECT 281.505000  56.890000 447.625000  56.960000 ;
      RECT 281.505000  56.890000 447.625000  56.960000 ;
      RECT 281.520000  47.080000 447.625000  47.150000 ;
      RECT 281.520000  47.080000 447.625000  47.150000 ;
      RECT 281.535000  75.325000 447.625000  75.395000 ;
      RECT 281.535000  75.325000 447.625000  75.395000 ;
      RECT 281.575000  47.400000 447.765000  56.625000 ;
      RECT 281.575000  56.625000 447.765000  57.435000 ;
      RECT 281.575000  56.820000 447.625000  56.890000 ;
      RECT 281.575000  56.820000 447.625000  56.890000 ;
      RECT 281.590000  47.150000 447.625000  47.220000 ;
      RECT 281.590000  47.150000 447.625000  47.220000 ;
      RECT 281.605000  75.395000 447.625000  75.465000 ;
      RECT 281.605000  75.395000 447.625000  75.465000 ;
      RECT 281.645000  56.750000 447.625000  56.820000 ;
      RECT 281.645000  56.750000 447.625000  56.820000 ;
      RECT 281.660000  47.220000 447.625000  47.290000 ;
      RECT 281.660000  47.220000 447.625000  47.290000 ;
      RECT 281.675000  75.465000 447.625000  75.535000 ;
      RECT 281.675000  75.465000 447.625000  75.535000 ;
      RECT 281.715000  47.290000 447.625000  47.345000 ;
      RECT 281.715000  47.290000 447.625000  47.345000 ;
      RECT 281.715000  47.345000 447.625000  74.765000 ;
      RECT 281.715000  56.680000 447.625000  56.750000 ;
      RECT 281.715000  56.680000 447.625000  56.750000 ;
      RECT 281.745000  75.535000 447.625000  75.605000 ;
      RECT 281.745000  75.535000 447.625000  75.605000 ;
      RECT 281.815000  75.605000 447.625000  75.675000 ;
      RECT 281.815000  75.605000 447.625000  75.675000 ;
      RECT 281.885000  75.675000 447.625000  75.745000 ;
      RECT 281.885000  75.675000 447.625000  75.745000 ;
      RECT 281.955000  75.745000 447.625000  75.815000 ;
      RECT 281.955000  75.745000 447.625000  75.815000 ;
      RECT 282.025000  75.815000 447.625000  75.885000 ;
      RECT 282.025000  75.815000 447.625000  75.885000 ;
      RECT 282.095000  75.885000 447.625000  75.955000 ;
      RECT 282.095000  75.885000 447.625000  75.955000 ;
      RECT 282.165000  75.955000 447.625000  76.025000 ;
      RECT 282.165000  75.955000 447.625000  76.025000 ;
      RECT 282.235000  76.025000 447.625000  76.095000 ;
      RECT 282.235000  76.025000 447.625000  76.095000 ;
      RECT 282.305000  76.095000 447.625000  76.165000 ;
      RECT 282.305000  76.095000 447.625000  76.165000 ;
      RECT 282.375000  76.165000 447.625000  76.235000 ;
      RECT 282.375000  76.165000 447.625000  76.235000 ;
      RECT 282.395000  76.450000 447.765000  83.500000 ;
      RECT 282.395000  83.500000 446.945000  85.775000 ;
      RECT 282.395000  85.775000 446.945000  87.480000 ;
      RECT 282.395000  87.480000 446.945000  89.420000 ;
      RECT 282.445000  76.235000 447.625000  76.305000 ;
      RECT 282.445000  76.235000 447.625000  76.305000 ;
      RECT 282.515000  76.305000 447.625000  76.375000 ;
      RECT 282.515000  76.305000 447.625000  76.375000 ;
      RECT 282.535000  76.375000 447.625000  76.395000 ;
      RECT 282.535000  76.375000 447.625000  76.395000 ;
      RECT 282.535000  76.395000 447.625000  83.640000 ;
      RECT 282.535000  83.640000 447.625000  84.900000 ;
      RECT 282.535000  83.640000 448.815000  83.710000 ;
      RECT 282.535000  83.710000 448.745000  83.780000 ;
      RECT 282.535000  83.780000 448.675000  83.850000 ;
      RECT 282.535000  83.850000 448.605000  83.920000 ;
      RECT 282.535000  83.920000 448.535000  83.990000 ;
      RECT 282.535000  83.990000 448.465000  84.060000 ;
      RECT 282.535000  84.060000 448.395000  84.130000 ;
      RECT 282.535000  84.130000 448.325000  84.200000 ;
      RECT 282.535000  84.200000 448.255000  84.270000 ;
      RECT 282.535000  84.270000 448.185000  84.340000 ;
      RECT 282.535000  84.340000 448.115000  84.410000 ;
      RECT 282.535000  84.410000 448.045000  84.480000 ;
      RECT 282.535000  84.480000 447.975000  84.550000 ;
      RECT 282.535000  84.550000 447.905000  84.620000 ;
      RECT 282.535000  84.620000 447.835000  84.690000 ;
      RECT 282.535000  84.690000 447.765000  84.760000 ;
      RECT 282.535000  84.760000 447.695000  84.830000 ;
      RECT 282.535000  84.830000 447.625000  84.900000 ;
      RECT 282.535000  84.900000 447.555000  84.970000 ;
      RECT 282.535000  84.900000 447.555000  84.970000 ;
      RECT 282.535000  84.900000 447.555000  84.970000 ;
      RECT 282.535000  84.970000 447.485000  85.040000 ;
      RECT 282.535000  84.970000 447.485000  85.040000 ;
      RECT 282.535000  84.970000 447.485000  85.040000 ;
      RECT 282.535000  85.040000 447.415000  85.110000 ;
      RECT 282.535000  85.040000 447.415000  85.110000 ;
      RECT 282.535000  85.040000 447.415000  85.110000 ;
      RECT 282.535000  85.110000 447.345000  85.180000 ;
      RECT 282.535000  85.110000 447.345000  85.180000 ;
      RECT 282.535000  85.110000 447.345000  85.180000 ;
      RECT 282.535000  85.180000 447.275000  85.250000 ;
      RECT 282.535000  85.180000 447.275000  85.250000 ;
      RECT 282.535000  85.180000 447.275000  85.250000 ;
      RECT 282.535000  85.250000 447.205000  85.320000 ;
      RECT 282.535000  85.250000 447.205000  85.320000 ;
      RECT 282.535000  85.250000 447.205000  85.320000 ;
      RECT 282.535000  85.320000 447.135000  85.390000 ;
      RECT 282.535000  85.320000 447.135000  85.390000 ;
      RECT 282.535000  85.320000 447.135000  85.390000 ;
      RECT 282.535000  85.390000 447.065000  85.460000 ;
      RECT 282.535000  85.390000 447.065000  85.460000 ;
      RECT 282.535000  85.390000 447.065000  85.460000 ;
      RECT 282.535000  85.460000 446.995000  85.530000 ;
      RECT 282.535000  85.460000 446.995000  85.530000 ;
      RECT 282.535000  85.460000 446.995000  85.530000 ;
      RECT 282.535000  85.530000 446.925000  85.600000 ;
      RECT 282.535000  85.530000 446.925000  85.600000 ;
      RECT 282.535000  85.530000 446.925000  85.600000 ;
      RECT 282.535000  85.600000 446.855000  85.670000 ;
      RECT 282.535000  85.600000 446.855000  85.670000 ;
      RECT 282.535000  85.600000 446.855000  85.670000 ;
      RECT 282.535000  85.670000 446.805000  85.720000 ;
      RECT 282.535000  85.670000 446.805000  85.720000 ;
      RECT 282.535000  85.670000 446.805000  85.720000 ;
      RECT 282.535000  85.720000 446.805000  87.425000 ;
      RECT 282.605000  87.425000 446.805000  87.495000 ;
      RECT 282.605000  87.425000 446.805000  87.495000 ;
      RECT 282.675000  87.495000 446.805000  87.565000 ;
      RECT 282.675000  87.495000 446.805000  87.565000 ;
      RECT 282.720000   2.125000 302.770000  18.295000 ;
      RECT 282.745000  87.565000 446.805000  87.635000 ;
      RECT 282.745000  87.565000 446.805000  87.635000 ;
      RECT 282.805000   2.280000 302.630000  18.435000 ;
      RECT 282.815000  87.635000 446.805000  87.705000 ;
      RECT 282.815000  87.635000 446.805000  87.705000 ;
      RECT 282.860000   2.180000 302.630000   2.280000 ;
      RECT 282.875000   2.165000 302.630000   2.180000 ;
      RECT 282.875000   2.165000 302.630000   2.180000 ;
      RECT 282.885000  87.705000 446.805000  87.775000 ;
      RECT 282.885000  87.705000 446.805000  87.775000 ;
      RECT 282.945000   2.095000 302.630000   2.165000 ;
      RECT 282.945000   2.095000 302.630000   2.165000 ;
      RECT 282.955000  87.775000 446.805000  87.845000 ;
      RECT 282.955000  87.775000 446.805000  87.845000 ;
      RECT 283.015000   2.025000 302.630000   2.095000 ;
      RECT 283.015000   2.025000 302.630000   2.095000 ;
      RECT 283.025000  87.845000 446.805000  87.915000 ;
      RECT 283.025000  87.845000 446.805000  87.915000 ;
      RECT 283.085000   1.955000 302.630000   2.025000 ;
      RECT 283.085000   1.955000 302.630000   2.025000 ;
      RECT 283.095000  87.915000 446.805000  87.985000 ;
      RECT 283.095000  87.915000 446.805000  87.985000 ;
      RECT 283.155000   1.885000 302.630000   1.955000 ;
      RECT 283.155000   1.885000 302.630000   1.955000 ;
      RECT 283.165000  87.985000 446.805000  88.055000 ;
      RECT 283.165000  87.985000 446.805000  88.055000 ;
      RECT 283.225000   1.815000 302.630000   1.885000 ;
      RECT 283.225000   1.815000 302.630000   1.885000 ;
      RECT 283.235000  88.055000 446.805000  88.125000 ;
      RECT 283.235000  88.055000 446.805000  88.125000 ;
      RECT 283.295000   1.745000 302.630000   1.815000 ;
      RECT 283.295000   1.745000 302.630000   1.815000 ;
      RECT 283.305000  88.125000 446.805000  88.195000 ;
      RECT 283.305000  88.125000 446.805000  88.195000 ;
      RECT 283.365000   1.675000 302.630000   1.745000 ;
      RECT 283.365000   1.675000 302.630000   1.745000 ;
      RECT 283.375000  88.195000 446.805000  88.265000 ;
      RECT 283.375000  88.195000 446.805000  88.265000 ;
      RECT 283.435000   0.000000 302.770000   1.410000 ;
      RECT 283.435000   1.410000 302.770000   2.125000 ;
      RECT 283.435000   1.605000 302.630000   1.675000 ;
      RECT 283.435000   1.605000 302.630000   1.675000 ;
      RECT 283.445000  88.265000 446.805000  88.335000 ;
      RECT 283.445000  88.265000 446.805000  88.335000 ;
      RECT 283.505000   1.535000 302.630000   1.605000 ;
      RECT 283.505000   1.535000 302.630000   1.605000 ;
      RECT 283.515000  88.335000 446.805000  88.405000 ;
      RECT 283.515000  88.335000 446.805000  88.405000 ;
      RECT 283.575000   0.000000 302.630000   1.465000 ;
      RECT 283.575000   0.000000 302.630000  18.435000 ;
      RECT 283.575000   0.000000 302.630000  18.435000 ;
      RECT 283.575000   1.465000 302.630000   1.535000 ;
      RECT 283.575000   1.465000 302.630000   1.535000 ;
      RECT 283.585000  88.405000 446.805000  88.475000 ;
      RECT 283.585000  88.405000 446.805000  88.475000 ;
      RECT 283.655000  88.475000 446.805000  88.545000 ;
      RECT 283.655000  88.475000 446.805000  88.545000 ;
      RECT 283.725000  88.545000 446.805000  88.615000 ;
      RECT 283.725000  88.545000 446.805000  88.615000 ;
      RECT 283.795000  88.615000 446.805000  88.685000 ;
      RECT 283.795000  88.615000 446.805000  88.685000 ;
      RECT 283.865000  88.685000 446.805000  88.755000 ;
      RECT 283.865000  88.685000 446.805000  88.755000 ;
      RECT 283.935000  88.755000 446.805000  88.825000 ;
      RECT 283.935000  88.755000 446.805000  88.825000 ;
      RECT 284.005000  88.825000 446.805000  88.895000 ;
      RECT 284.005000  88.825000 446.805000  88.895000 ;
      RECT 284.075000  88.895000 446.805000  88.965000 ;
      RECT 284.075000  88.895000 446.805000  88.965000 ;
      RECT 284.145000  88.965000 446.805000  89.035000 ;
      RECT 284.145000  88.965000 446.805000  89.035000 ;
      RECT 284.215000  89.035000 446.805000  89.105000 ;
      RECT 284.215000  89.035000 446.805000  89.105000 ;
      RECT 284.285000  89.105000 446.805000  89.175000 ;
      RECT 284.285000  89.105000 446.805000  89.175000 ;
      RECT 284.335000  89.420000 446.945000  94.105000 ;
      RECT 284.335000  94.105000 446.945000  94.560000 ;
      RECT 284.355000  89.175000 446.805000  89.245000 ;
      RECT 284.355000  89.175000 446.805000  89.245000 ;
      RECT 284.425000  89.245000 446.805000  89.315000 ;
      RECT 284.425000  89.245000 446.805000  89.315000 ;
      RECT 284.475000  76.395000 446.805000  94.050000 ;
      RECT 284.475000  89.315000 446.805000  89.365000 ;
      RECT 284.475000  89.315000 446.805000  89.365000 ;
      RECT 284.475000  89.365000 446.805000  94.050000 ;
      RECT 284.545000  94.050000 446.805000  94.120000 ;
      RECT 284.545000  94.050000 446.805000  94.120000 ;
      RECT 284.615000  94.120000 446.805000  94.190000 ;
      RECT 284.615000  94.120000 446.805000  94.190000 ;
      RECT 284.685000  94.190000 446.805000  94.260000 ;
      RECT 284.685000  94.190000 446.805000  94.260000 ;
      RECT 284.755000  94.260000 446.805000  94.330000 ;
      RECT 284.755000  94.260000 446.805000  94.330000 ;
      RECT 284.825000  94.330000 446.805000  94.400000 ;
      RECT 284.825000  94.330000 446.805000  94.400000 ;
      RECT 284.845000  94.400000 446.805000  94.420000 ;
      RECT 284.845000  94.400000 446.805000  94.420000 ;
      RECT 289.475000  94.560000 446.945000 102.925000 ;
      RECT 289.600000  94.420000 446.805000  94.490000 ;
      RECT 289.600000  94.420000 446.805000  94.490000 ;
      RECT 289.670000  94.490000 446.805000  94.560000 ;
      RECT 289.670000  94.490000 446.805000  94.560000 ;
      RECT 289.740000  94.560000 446.805000  94.630000 ;
      RECT 289.740000  94.560000 446.805000  94.630000 ;
      RECT 289.810000  94.630000 446.805000  94.700000 ;
      RECT 289.810000  94.630000 446.805000  94.700000 ;
      RECT 289.880000  94.700000 446.805000  94.770000 ;
      RECT 289.880000  94.700000 446.805000  94.770000 ;
      RECT 289.950000  94.770000 446.805000  94.840000 ;
      RECT 289.950000  94.770000 446.805000  94.840000 ;
      RECT 290.020000  94.840000 446.805000  94.910000 ;
      RECT 290.020000  94.840000 446.805000  94.910000 ;
      RECT 290.090000  94.910000 446.805000  94.980000 ;
      RECT 290.090000  94.910000 446.805000  94.980000 ;
      RECT 290.160000  94.980000 446.805000  95.050000 ;
      RECT 290.160000  94.980000 446.805000  95.050000 ;
      RECT 290.230000  95.050000 446.805000  95.120000 ;
      RECT 290.230000  95.050000 446.805000  95.120000 ;
      RECT 290.300000  95.120000 446.805000  95.190000 ;
      RECT 290.300000  95.120000 446.805000  95.190000 ;
      RECT 290.370000  95.190000 446.805000  95.260000 ;
      RECT 290.370000  95.190000 446.805000  95.260000 ;
      RECT 290.440000  95.260000 446.805000  95.330000 ;
      RECT 290.440000  95.260000 446.805000  95.330000 ;
      RECT 290.510000  95.330000 446.805000  95.400000 ;
      RECT 290.510000  95.330000 446.805000  95.400000 ;
      RECT 290.580000  95.400000 446.805000  95.470000 ;
      RECT 290.580000  95.400000 446.805000  95.470000 ;
      RECT 290.650000  95.470000 446.805000  95.540000 ;
      RECT 290.650000  95.470000 446.805000  95.540000 ;
      RECT 290.720000  95.540000 446.805000  95.610000 ;
      RECT 290.720000  95.540000 446.805000  95.610000 ;
      RECT 290.790000  95.610000 446.805000  95.680000 ;
      RECT 290.790000  95.610000 446.805000  95.680000 ;
      RECT 290.860000  95.680000 446.805000  95.750000 ;
      RECT 290.860000  95.680000 446.805000  95.750000 ;
      RECT 290.930000  95.750000 446.805000  95.820000 ;
      RECT 290.930000  95.750000 446.805000  95.820000 ;
      RECT 291.000000  95.820000 446.805000  95.890000 ;
      RECT 291.000000  95.820000 446.805000  95.890000 ;
      RECT 291.070000  95.890000 446.805000  95.960000 ;
      RECT 291.070000  95.890000 446.805000  95.960000 ;
      RECT 291.140000  95.960000 446.805000  96.030000 ;
      RECT 291.140000  95.960000 446.805000  96.030000 ;
      RECT 291.210000  96.030000 446.805000  96.100000 ;
      RECT 291.210000  96.030000 446.805000  96.100000 ;
      RECT 291.280000  96.100000 446.805000  96.170000 ;
      RECT 291.280000  96.100000 446.805000  96.170000 ;
      RECT 291.350000  96.170000 446.805000  96.240000 ;
      RECT 291.350000  96.170000 446.805000  96.240000 ;
      RECT 291.420000  96.240000 446.805000  96.310000 ;
      RECT 291.420000  96.240000 446.805000  96.310000 ;
      RECT 291.490000  96.310000 446.805000  96.380000 ;
      RECT 291.490000  96.310000 446.805000  96.380000 ;
      RECT 291.560000  96.380000 446.805000  96.450000 ;
      RECT 291.560000  96.380000 446.805000  96.450000 ;
      RECT 291.630000  96.450000 446.805000  96.520000 ;
      RECT 291.630000  96.450000 446.805000  96.520000 ;
      RECT 291.700000  96.520000 446.805000  96.590000 ;
      RECT 291.700000  96.520000 446.805000  96.590000 ;
      RECT 291.770000  96.590000 446.805000  96.660000 ;
      RECT 291.770000  96.590000 446.805000  96.660000 ;
      RECT 291.840000  96.660000 446.805000  96.730000 ;
      RECT 291.840000  96.660000 446.805000  96.730000 ;
      RECT 291.910000  96.730000 446.805000  96.800000 ;
      RECT 291.910000  96.730000 446.805000  96.800000 ;
      RECT 291.980000  96.800000 446.805000  96.870000 ;
      RECT 291.980000  96.800000 446.805000  96.870000 ;
      RECT 292.050000  96.870000 446.805000  96.940000 ;
      RECT 292.050000  96.870000 446.805000  96.940000 ;
      RECT 292.120000  96.940000 446.805000  97.010000 ;
      RECT 292.120000  96.940000 446.805000  97.010000 ;
      RECT 292.190000  97.010000 446.805000  97.080000 ;
      RECT 292.190000  97.010000 446.805000  97.080000 ;
      RECT 292.260000  97.080000 446.805000  97.150000 ;
      RECT 292.260000  97.080000 446.805000  97.150000 ;
      RECT 292.330000  97.150000 446.805000  97.220000 ;
      RECT 292.330000  97.150000 446.805000  97.220000 ;
      RECT 292.400000  97.220000 446.805000  97.290000 ;
      RECT 292.400000  97.220000 446.805000  97.290000 ;
      RECT 292.470000  97.290000 446.805000  97.360000 ;
      RECT 292.470000  97.290000 446.805000  97.360000 ;
      RECT 292.540000  97.360000 446.805000  97.430000 ;
      RECT 292.540000  97.360000 446.805000  97.430000 ;
      RECT 292.610000  97.430000 446.805000  97.500000 ;
      RECT 292.610000  97.430000 446.805000  97.500000 ;
      RECT 292.680000  97.500000 446.805000  97.570000 ;
      RECT 292.680000  97.500000 446.805000  97.570000 ;
      RECT 292.750000  97.570000 446.805000  97.640000 ;
      RECT 292.750000  97.570000 446.805000  97.640000 ;
      RECT 292.820000  97.640000 446.805000  97.710000 ;
      RECT 292.820000  97.640000 446.805000  97.710000 ;
      RECT 292.890000  97.710000 446.805000  97.780000 ;
      RECT 292.890000  97.710000 446.805000  97.780000 ;
      RECT 292.960000  97.780000 446.805000  97.850000 ;
      RECT 292.960000  97.780000 446.805000  97.850000 ;
      RECT 293.030000  97.850000 446.805000  97.920000 ;
      RECT 293.030000  97.850000 446.805000  97.920000 ;
      RECT 293.100000  97.920000 446.805000  97.990000 ;
      RECT 293.100000  97.920000 446.805000  97.990000 ;
      RECT 293.170000  97.990000 446.805000  98.060000 ;
      RECT 293.170000  97.990000 446.805000  98.060000 ;
      RECT 293.240000  98.060000 446.805000  98.130000 ;
      RECT 293.240000  98.060000 446.805000  98.130000 ;
      RECT 293.310000  98.130000 446.805000  98.200000 ;
      RECT 293.310000  98.130000 446.805000  98.200000 ;
      RECT 293.380000  98.200000 446.805000  98.270000 ;
      RECT 293.380000  98.200000 446.805000  98.270000 ;
      RECT 293.450000  98.270000 446.805000  98.340000 ;
      RECT 293.450000  98.270000 446.805000  98.340000 ;
      RECT 293.520000  98.340000 446.805000  98.410000 ;
      RECT 293.520000  98.340000 446.805000  98.410000 ;
      RECT 293.590000  98.410000 446.805000  98.480000 ;
      RECT 293.590000  98.410000 446.805000  98.480000 ;
      RECT 293.660000  98.480000 446.805000  98.550000 ;
      RECT 293.660000  98.480000 446.805000  98.550000 ;
      RECT 293.730000  98.550000 446.805000  98.620000 ;
      RECT 293.730000  98.550000 446.805000  98.620000 ;
      RECT 293.800000  98.620000 446.805000  98.690000 ;
      RECT 293.800000  98.620000 446.805000  98.690000 ;
      RECT 293.870000  98.690000 446.805000  98.760000 ;
      RECT 293.870000  98.690000 446.805000  98.760000 ;
      RECT 293.940000  98.760000 446.805000  98.830000 ;
      RECT 293.940000  98.760000 446.805000  98.830000 ;
      RECT 294.010000  98.830000 446.805000  98.900000 ;
      RECT 294.010000  98.830000 446.805000  98.900000 ;
      RECT 294.080000  98.900000 446.805000  98.970000 ;
      RECT 294.080000  98.900000 446.805000  98.970000 ;
      RECT 294.150000  98.970000 446.805000  99.040000 ;
      RECT 294.150000  98.970000 446.805000  99.040000 ;
      RECT 294.220000  99.040000 446.805000  99.110000 ;
      RECT 294.220000  99.040000 446.805000  99.110000 ;
      RECT 294.290000  99.110000 446.805000  99.180000 ;
      RECT 294.290000  99.110000 446.805000  99.180000 ;
      RECT 294.360000  99.180000 446.805000  99.250000 ;
      RECT 294.360000  99.180000 446.805000  99.250000 ;
      RECT 294.430000  99.250000 446.805000  99.320000 ;
      RECT 294.430000  99.250000 446.805000  99.320000 ;
      RECT 294.500000  99.320000 446.805000  99.390000 ;
      RECT 294.500000  99.320000 446.805000  99.390000 ;
      RECT 294.570000  99.390000 446.805000  99.460000 ;
      RECT 294.570000  99.390000 446.805000  99.460000 ;
      RECT 294.640000  99.460000 446.805000  99.530000 ;
      RECT 294.640000  99.460000 446.805000  99.530000 ;
      RECT 294.710000  99.530000 446.805000  99.600000 ;
      RECT 294.710000  99.530000 446.805000  99.600000 ;
      RECT 294.780000  99.600000 446.805000  99.670000 ;
      RECT 294.780000  99.600000 446.805000  99.670000 ;
      RECT 294.850000  99.670000 446.805000  99.740000 ;
      RECT 294.850000  99.670000 446.805000  99.740000 ;
      RECT 294.920000  99.740000 446.805000  99.810000 ;
      RECT 294.920000  99.740000 446.805000  99.810000 ;
      RECT 294.990000  99.810000 446.805000  99.880000 ;
      RECT 294.990000  99.810000 446.805000  99.880000 ;
      RECT 295.060000  99.880000 446.805000  99.950000 ;
      RECT 295.060000  99.880000 446.805000  99.950000 ;
      RECT 295.130000  99.950000 446.805000 100.020000 ;
      RECT 295.130000  99.950000 446.805000 100.020000 ;
      RECT 295.200000 100.020000 446.805000 100.090000 ;
      RECT 295.200000 100.020000 446.805000 100.090000 ;
      RECT 295.270000 100.090000 446.805000 100.160000 ;
      RECT 295.270000 100.090000 446.805000 100.160000 ;
      RECT 295.340000 100.160000 446.805000 100.230000 ;
      RECT 295.340000 100.160000 446.805000 100.230000 ;
      RECT 295.410000 100.230000 446.805000 100.300000 ;
      RECT 295.410000 100.230000 446.805000 100.300000 ;
      RECT 295.480000 100.300000 446.805000 100.370000 ;
      RECT 295.480000 100.300000 446.805000 100.370000 ;
      RECT 295.550000 100.370000 446.805000 100.440000 ;
      RECT 295.550000 100.370000 446.805000 100.440000 ;
      RECT 295.620000 100.440000 446.805000 100.510000 ;
      RECT 295.620000 100.440000 446.805000 100.510000 ;
      RECT 295.690000 100.510000 446.805000 100.580000 ;
      RECT 295.690000 100.510000 446.805000 100.580000 ;
      RECT 295.760000 100.580000 446.805000 100.650000 ;
      RECT 295.760000 100.580000 446.805000 100.650000 ;
      RECT 295.830000 100.650000 446.805000 100.720000 ;
      RECT 295.830000 100.650000 446.805000 100.720000 ;
      RECT 295.900000 100.720000 446.805000 100.790000 ;
      RECT 295.900000 100.720000 446.805000 100.790000 ;
      RECT 295.970000 100.790000 446.805000 100.860000 ;
      RECT 295.970000 100.790000 446.805000 100.860000 ;
      RECT 296.040000 100.860000 446.805000 100.930000 ;
      RECT 296.040000 100.860000 446.805000 100.930000 ;
      RECT 296.110000 100.930000 446.805000 101.000000 ;
      RECT 296.110000 100.930000 446.805000 101.000000 ;
      RECT 296.180000 101.000000 446.805000 101.070000 ;
      RECT 296.180000 101.000000 446.805000 101.070000 ;
      RECT 296.250000 101.070000 446.805000 101.140000 ;
      RECT 296.250000 101.070000 446.805000 101.140000 ;
      RECT 296.320000 101.140000 446.805000 101.210000 ;
      RECT 296.320000 101.140000 446.805000 101.210000 ;
      RECT 296.390000 101.210000 446.805000 101.280000 ;
      RECT 296.390000 101.210000 446.805000 101.280000 ;
      RECT 296.460000 101.280000 446.805000 101.350000 ;
      RECT 296.460000 101.280000 446.805000 101.350000 ;
      RECT 296.530000 101.350000 446.805000 101.420000 ;
      RECT 296.530000 101.350000 446.805000 101.420000 ;
      RECT 296.600000 101.420000 446.805000 101.490000 ;
      RECT 296.600000 101.420000 446.805000 101.490000 ;
      RECT 296.670000 101.490000 446.805000 101.560000 ;
      RECT 296.670000 101.490000 446.805000 101.560000 ;
      RECT 296.740000 101.560000 446.805000 101.630000 ;
      RECT 296.740000 101.560000 446.805000 101.630000 ;
      RECT 296.810000 101.630000 446.805000 101.700000 ;
      RECT 296.810000 101.630000 446.805000 101.700000 ;
      RECT 296.880000 101.700000 446.805000 101.770000 ;
      RECT 296.880000 101.700000 446.805000 101.770000 ;
      RECT 296.950000 101.770000 446.805000 101.840000 ;
      RECT 296.950000 101.770000 446.805000 101.840000 ;
      RECT 297.020000 101.840000 446.805000 101.910000 ;
      RECT 297.020000 101.840000 446.805000 101.910000 ;
      RECT 297.060000 111.960000 446.945000 112.280000 ;
      RECT 297.090000 101.910000 446.805000 101.980000 ;
      RECT 297.090000 101.910000 446.805000 101.980000 ;
      RECT 297.120000 111.900000 446.945000 111.960000 ;
      RECT 297.160000 101.980000 446.805000 102.050000 ;
      RECT 297.160000 101.980000 446.805000 102.050000 ;
      RECT 297.200000 112.040000 300.205000 112.420000 ;
      RECT 297.230000 102.050000 446.805000 102.120000 ;
      RECT 297.230000 102.050000 446.805000 102.120000 ;
      RECT 297.300000 102.120000 446.805000 102.190000 ;
      RECT 297.300000 102.120000 446.805000 102.190000 ;
      RECT 297.305000 112.390000 446.805000 112.420000 ;
      RECT 297.305000 112.390000 446.805000 112.420000 ;
      RECT 297.370000 102.190000 446.805000 102.260000 ;
      RECT 297.370000 102.190000 446.805000 102.260000 ;
      RECT 297.375000 112.320000 446.805000 112.390000 ;
      RECT 297.375000 112.320000 446.805000 112.390000 ;
      RECT 297.440000 102.260000 446.805000 102.330000 ;
      RECT 297.440000 102.260000 446.805000 102.330000 ;
      RECT 297.445000 112.250000 446.805000 112.320000 ;
      RECT 297.445000 112.250000 446.805000 112.320000 ;
      RECT 297.510000 102.330000 446.805000 102.400000 ;
      RECT 297.510000 102.330000 446.805000 102.400000 ;
      RECT 297.515000 112.180000 446.805000 112.250000 ;
      RECT 297.515000 112.180000 446.805000 112.250000 ;
      RECT 297.580000 102.400000 446.805000 102.470000 ;
      RECT 297.580000 102.400000 446.805000 102.470000 ;
      RECT 297.585000 112.110000 446.805000 112.180000 ;
      RECT 297.585000 112.110000 446.805000 112.180000 ;
      RECT 297.650000 102.470000 446.805000 102.540000 ;
      RECT 297.650000 102.470000 446.805000 102.540000 ;
      RECT 297.655000 112.040000 446.805000 112.110000 ;
      RECT 297.655000 112.040000 446.805000 112.110000 ;
      RECT 297.700000 111.995000 446.805000 112.040000 ;
      RECT 297.700000 111.995000 446.805000 112.040000 ;
      RECT 297.720000 102.540000 446.805000 102.610000 ;
      RECT 297.720000 102.540000 446.805000 102.610000 ;
      RECT 297.770000 111.925000 446.805000 111.995000 ;
      RECT 297.770000 111.925000 446.805000 111.995000 ;
      RECT 297.790000 102.610000 446.805000 102.680000 ;
      RECT 297.790000 102.610000 446.805000 102.680000 ;
      RECT 297.840000 102.925000 446.945000 111.660000 ;
      RECT 297.840000 111.660000 446.945000 111.900000 ;
      RECT 297.840000 111.855000 446.805000 111.925000 ;
      RECT 297.840000 111.855000 446.805000 111.925000 ;
      RECT 297.860000 102.680000 446.805000 102.750000 ;
      RECT 297.860000 102.680000 446.805000 102.750000 ;
      RECT 297.910000 111.785000 446.805000 111.855000 ;
      RECT 297.910000 111.785000 446.805000 111.855000 ;
      RECT 297.930000 102.750000 446.805000 102.820000 ;
      RECT 297.930000 102.750000 446.805000 102.820000 ;
      RECT 297.980000 102.820000 446.805000 102.870000 ;
      RECT 297.980000 102.820000 446.805000 102.870000 ;
      RECT 297.980000 102.870000 446.805000 111.715000 ;
      RECT 297.980000 111.715000 446.805000 111.785000 ;
      RECT 297.980000 111.715000 446.805000 111.785000 ;
      RECT 303.900000  30.685000 447.765000  33.375000 ;
      RECT 304.040000  30.825000 447.625000  33.515000 ;
      RECT 304.040000  30.825000 447.625000  45.365000 ;
      RECT 304.885000   0.000000 402.700000  23.280000 ;
      RECT 304.885000  23.280000 447.765000  30.685000 ;
      RECT 305.025000   0.000000 402.560000  23.420000 ;
      RECT 305.025000  23.420000 447.625000  30.825000 ;
      RECT 305.025000  23.420000 447.625000  33.515000 ;
      RECT 403.240000   0.000000 404.855000  14.710000 ;
      RECT 403.240000  14.710000 404.815000  14.750000 ;
      RECT 403.240000  14.750000 404.815000  15.210000 ;
      RECT 403.240000  15.210000 422.550000  23.280000 ;
      RECT 403.380000   0.000000 404.715000  14.655000 ;
      RECT 403.380000  14.655000 404.695000  14.675000 ;
      RECT 403.380000  14.675000 404.675000  14.695000 ;
      RECT 403.380000  14.695000 404.675000  15.350000 ;
      RECT 403.380000  15.350000 422.410000  23.420000 ;
      RECT 403.380000  15.350000 422.410000  30.825000 ;
      RECT 405.395000   0.000000 419.305000   5.175000 ;
      RECT 405.395000   5.175000 422.550000  14.625000 ;
      RECT 405.395000  14.625000 422.550000  14.670000 ;
      RECT 405.535000   0.000000 419.165000   5.315000 ;
      RECT 405.535000   5.315000 422.410000  14.530000 ;
      RECT 405.735000  14.670000 422.550000  15.210000 ;
      RECT 405.875000   5.315000 422.410000  15.350000 ;
      RECT 405.875000  14.530000 422.410000  15.350000 ;
      RECT 419.845000   0.000000 422.550000   5.175000 ;
      RECT 419.985000   0.000000 422.410000   5.315000 ;
      RECT 423.090000   0.000000 444.700000  23.155000 ;
      RECT 423.090000  23.155000 447.765000  23.280000 ;
      RECT 423.230000   0.000000 444.560000  23.295000 ;
      RECT 423.230000   0.000000 444.560000  30.825000 ;
      RECT 423.230000  23.295000 447.625000  23.420000 ;
      RECT 423.230000  23.295000 447.625000  30.825000 ;
      RECT 445.240000   0.000000 447.765000  22.245000 ;
      RECT 445.240000  22.245000 447.765000  22.315000 ;
      RECT 445.310000  22.315000 447.765000  23.155000 ;
      RECT 445.380000   0.000000 447.625000  22.190000 ;
      RECT 445.415000  22.190000 447.625000  22.225000 ;
      RECT 445.450000  22.225000 447.625000  22.260000 ;
      RECT 445.450000  22.260000 447.625000  23.295000 ;
      RECT 447.485000  86.005000 450.015000 235.840000 ;
      RECT 447.485000 235.840000 447.605000 238.250000 ;
      RECT 447.485000 238.250000 447.605000 244.110000 ;
      RECT 447.485000 244.110000 447.605000 244.215000 ;
      RECT 447.625000  86.060000 449.875000 235.785000 ;
      RECT 447.625000 235.785000 449.805000 235.855000 ;
      RECT 447.625000 235.855000 449.735000 235.925000 ;
      RECT 447.625000 235.925000 449.665000 235.995000 ;
      RECT 447.625000 235.995000 449.595000 236.065000 ;
      RECT 447.625000 236.065000 449.525000 236.135000 ;
      RECT 447.625000 236.135000 449.455000 236.205000 ;
      RECT 447.625000 236.205000 449.385000 236.275000 ;
      RECT 447.625000 236.275000 449.315000 236.345000 ;
      RECT 447.625000 236.345000 449.245000 236.415000 ;
      RECT 447.625000 236.415000 449.175000 236.485000 ;
      RECT 447.625000 236.485000 449.105000 236.555000 ;
      RECT 447.625000 236.555000 449.035000 236.625000 ;
      RECT 447.625000 236.625000 448.965000 236.695000 ;
      RECT 447.625000 236.695000 448.895000 236.765000 ;
      RECT 447.625000 236.765000 448.825000 236.835000 ;
      RECT 447.625000 236.835000 448.755000 236.905000 ;
      RECT 447.625000 236.905000 448.685000 236.975000 ;
      RECT 447.625000 236.975000 448.615000 237.045000 ;
      RECT 447.625000 237.045000 448.545000 237.115000 ;
      RECT 447.625000 237.115000 448.475000 237.185000 ;
      RECT 447.625000 237.185000 448.405000 237.255000 ;
      RECT 447.625000 237.255000 448.335000 237.325000 ;
      RECT 447.625000 237.325000 448.265000 237.395000 ;
      RECT 447.625000 237.395000 448.195000 237.465000 ;
      RECT 447.625000 237.465000 448.125000 237.535000 ;
      RECT 447.625000 237.535000 448.055000 237.605000 ;
      RECT 447.625000 237.605000 447.985000 237.675000 ;
      RECT 447.625000 237.675000 447.915000 237.745000 ;
      RECT 447.625000 237.745000 447.845000 237.815000 ;
      RECT 447.625000 237.815000 447.775000 237.885000 ;
      RECT 447.625000 237.885000 447.705000 237.955000 ;
      RECT 447.625000 237.955000 447.635000 238.025000 ;
      RECT 447.635000  86.050000 449.875000  86.060000 ;
      RECT 447.705000  85.980000 449.875000  86.050000 ;
      RECT 447.775000  85.910000 449.875000  85.980000 ;
      RECT 447.845000  85.840000 449.875000  85.910000 ;
      RECT 447.915000  85.770000 449.875000  85.840000 ;
      RECT 447.985000  85.700000 449.875000  85.770000 ;
      RECT 448.055000  85.630000 449.875000  85.700000 ;
      RECT 448.125000  85.560000 449.875000  85.630000 ;
      RECT 448.145000 238.480000 448.355000 238.570000 ;
      RECT 448.145000 238.570000 448.355000 245.155000 ;
      RECT 448.195000  85.490000 449.875000  85.560000 ;
      RECT 448.265000  85.420000 449.875000  85.490000 ;
      RECT 448.305000   0.000000 448.515000  83.500000 ;
      RECT 448.335000  85.350000 449.875000  85.420000 ;
      RECT 448.405000  85.280000 449.875000  85.350000 ;
      RECT 448.475000  85.210000 449.875000  85.280000 ;
      RECT 448.545000  85.140000 449.875000  85.210000 ;
      RECT 448.615000  85.070000 449.875000  85.140000 ;
      RECT 448.685000  85.000000 449.875000  85.070000 ;
      RECT 448.755000  84.930000 449.875000  85.000000 ;
      RECT 448.825000  84.860000 449.875000  84.930000 ;
      RECT 448.895000  84.790000 449.875000  84.860000 ;
      RECT 448.895000 238.800000 449.105000 238.890000 ;
      RECT 448.895000 238.890000 449.105000 245.555000 ;
      RECT 448.965000  84.720000 449.875000  84.790000 ;
      RECT 449.035000  84.650000 449.875000  84.720000 ;
      RECT 449.055000   0.000000 449.265000  83.455000 ;
      RECT 449.055000  83.455000 449.220000  83.500000 ;
      RECT 449.105000  84.580000 449.875000  84.650000 ;
      RECT 449.175000  84.510000 449.875000  84.580000 ;
      RECT 449.245000  84.440000 449.875000  84.510000 ;
      RECT 449.315000  84.370000 449.875000  84.440000 ;
      RECT 449.385000  84.300000 449.875000  84.370000 ;
      RECT 449.455000  84.230000 449.875000  84.300000 ;
      RECT 449.525000  84.160000 449.875000  84.230000 ;
      RECT 449.595000  84.090000 449.875000  84.160000 ;
      RECT 449.645000 239.120000 449.855000 239.210000 ;
      RECT 449.645000 239.210000 449.855000 240.855000 ;
      RECT 449.645000 240.855000 450.605000 241.925000 ;
      RECT 449.645000 241.925000 450.975000 242.365000 ;
      RECT 449.645000 242.365000 480.000000 245.955000 ;
      RECT 449.665000  84.020000 449.875000  84.090000 ;
      RECT 449.735000  83.950000 449.875000  84.020000 ;
      RECT 449.785000 240.995000 450.465000 242.065000 ;
      RECT 449.785000 242.065000 450.835000 242.505000 ;
      RECT 449.785000 242.505000 480.000000 246.095000 ;
      RECT 449.785000 242.505000 480.000000 253.715000 ;
      RECT 449.785000 242.505000 480.000000 253.715000 ;
      RECT 449.785000 242.505000 480.000000 253.715000 ;
      RECT 449.805000   0.000000 450.015000  83.685000 ;
      RECT 449.805000  83.685000 450.015000  86.005000 ;
      RECT 449.805000  83.880000 449.875000  83.950000 ;
      RECT 450.395000 239.440000 450.605000 239.530000 ;
      RECT 450.395000 239.530000 450.605000 240.855000 ;
      RECT 450.555000   0.000000 450.765000 236.070000 ;
      RECT 450.555000 236.070000 450.765000 236.160000 ;
      RECT 451.145000 239.760000 451.355000 239.850000 ;
      RECT 451.145000 239.850000 451.355000 241.700000 ;
      RECT 451.145000 241.700000 451.230000 241.825000 ;
      RECT 451.305000   0.000000 451.515000 236.390000 ;
      RECT 451.305000 236.390000 451.515000 236.480000 ;
      RECT 451.895000 240.080000 480.000000 242.365000 ;
      RECT 452.035000 240.135000 480.000000 242.505000 ;
      RECT 452.055000   0.000000 452.265000 236.710000 ;
      RECT 452.055000 236.710000 452.265000 236.800000 ;
      RECT 452.065000 240.105000 480.000000 240.135000 ;
      RECT 452.065000 240.105000 480.000000 240.135000 ;
      RECT 452.135000 240.035000 480.000000 240.105000 ;
      RECT 452.135000 240.035000 480.000000 240.105000 ;
      RECT 452.205000 239.965000 480.000000 240.035000 ;
      RECT 452.205000 239.965000 480.000000 240.035000 ;
      RECT 452.275000 239.895000 480.000000 239.965000 ;
      RECT 452.275000 239.895000 480.000000 239.965000 ;
      RECT 452.345000 239.825000 480.000000 239.895000 ;
      RECT 452.345000 239.825000 480.000000 239.895000 ;
      RECT 452.415000 239.755000 480.000000 239.825000 ;
      RECT 452.415000 239.755000 480.000000 239.825000 ;
      RECT 452.485000 239.685000 480.000000 239.755000 ;
      RECT 452.485000 239.685000 480.000000 239.755000 ;
      RECT 452.555000 239.615000 480.000000 239.685000 ;
      RECT 452.555000 239.615000 480.000000 239.685000 ;
      RECT 452.625000 239.545000 480.000000 239.615000 ;
      RECT 452.625000 239.545000 480.000000 239.615000 ;
      RECT 452.695000 239.475000 480.000000 239.545000 ;
      RECT 452.695000 239.475000 480.000000 239.545000 ;
      RECT 452.765000 239.405000 480.000000 239.475000 ;
      RECT 452.765000 239.405000 480.000000 239.475000 ;
      RECT 452.805000   0.000000 453.015000 237.030000 ;
      RECT 452.805000 237.030000 453.015000 237.120000 ;
      RECT 452.835000 239.335000 480.000000 239.405000 ;
      RECT 452.835000 239.335000 480.000000 239.405000 ;
      RECT 452.905000 239.265000 480.000000 239.335000 ;
      RECT 452.905000 239.265000 480.000000 239.335000 ;
      RECT 452.975000 239.195000 480.000000 239.265000 ;
      RECT 452.975000 239.195000 480.000000 239.265000 ;
      RECT 453.045000 239.125000 480.000000 239.195000 ;
      RECT 453.045000 239.125000 480.000000 239.195000 ;
      RECT 453.115000 239.055000 480.000000 239.125000 ;
      RECT 453.115000 239.055000 480.000000 239.125000 ;
      RECT 453.185000 238.985000 480.000000 239.055000 ;
      RECT 453.185000 238.985000 480.000000 239.055000 ;
      RECT 453.255000 238.915000 480.000000 238.985000 ;
      RECT 453.255000 238.915000 480.000000 238.985000 ;
      RECT 453.325000 238.845000 480.000000 238.915000 ;
      RECT 453.325000 238.845000 480.000000 238.915000 ;
      RECT 453.395000 238.775000 480.000000 238.845000 ;
      RECT 453.395000 238.775000 480.000000 238.845000 ;
      RECT 453.465000 238.705000 480.000000 238.775000 ;
      RECT 453.465000 238.705000 480.000000 238.775000 ;
      RECT 453.535000 238.635000 480.000000 238.705000 ;
      RECT 453.535000 238.635000 480.000000 238.705000 ;
      RECT 453.555000   0.000000 453.765000 237.350000 ;
      RECT 453.555000 237.350000 453.765000 237.440000 ;
      RECT 453.605000 238.565000 480.000000 238.635000 ;
      RECT 453.605000 238.565000 480.000000 238.635000 ;
      RECT 453.675000 238.495000 480.000000 238.565000 ;
      RECT 453.675000 238.495000 480.000000 238.565000 ;
      RECT 453.745000 238.425000 480.000000 238.495000 ;
      RECT 453.745000 238.425000 480.000000 238.495000 ;
      RECT 453.815000 238.355000 480.000000 238.425000 ;
      RECT 453.815000 238.355000 480.000000 238.425000 ;
      RECT 453.885000 238.285000 480.000000 238.355000 ;
      RECT 453.885000 238.285000 480.000000 238.355000 ;
      RECT 453.955000 238.215000 480.000000 238.285000 ;
      RECT 453.955000 238.215000 480.000000 238.285000 ;
      RECT 454.025000 238.145000 480.000000 238.215000 ;
      RECT 454.025000 238.145000 480.000000 238.215000 ;
      RECT 454.095000 238.075000 480.000000 238.145000 ;
      RECT 454.095000 238.075000 480.000000 238.145000 ;
      RECT 454.165000 238.005000 480.000000 238.075000 ;
      RECT 454.165000 238.005000 480.000000 238.075000 ;
      RECT 454.235000 237.935000 480.000000 238.005000 ;
      RECT 454.235000 237.935000 480.000000 238.005000 ;
      RECT 454.305000   0.000000 464.390000  60.435000 ;
      RECT 454.305000  60.435000 480.000000 237.670000 ;
      RECT 454.305000 237.670000 480.000000 240.080000 ;
      RECT 454.305000 237.865000 480.000000 237.935000 ;
      RECT 454.305000 237.865000 480.000000 237.935000 ;
      RECT 454.375000 237.795000 480.000000 237.865000 ;
      RECT 454.375000 237.795000 480.000000 237.865000 ;
      RECT 454.445000   0.000000 464.250000  60.575000 ;
      RECT 454.445000  60.575000 480.000000 237.725000 ;
      RECT 454.445000  60.575000 480.000000 242.505000 ;
      RECT 454.445000 237.725000 480.000000 237.795000 ;
      RECT 454.445000 237.725000 480.000000 237.795000 ;
      RECT 465.310000   0.000000 465.890000  60.435000 ;
      RECT 465.450000   0.000000 465.750000  60.575000 ;
      RECT 466.810000   0.000000 480.000000  60.435000 ;
      RECT 466.950000   0.000000 480.000000  60.575000 ;
    LAYER met3 ;
      RECT 0.000000 0.000000 480.000000 253.715000 ;
    LAYER met4 ;
      RECT   0.000000   0.000000 480.000000  55.350000 ;
      RECT   0.000000   0.000000 480.000000  55.350000 ;
      RECT   0.000000  61.600000 480.000000  62.200000 ;
      RECT   0.000000  61.600000 480.000000  62.200000 ;
      RECT   0.000000  67.650000 480.000000  68.250000 ;
      RECT   0.000000  67.650000 480.000000  68.250000 ;
      RECT   0.000000  72.500000 480.000000  73.015000 ;
      RECT   0.000000  72.500000 480.000000  73.115000 ;
      RECT   0.000000  73.015000   9.460000  73.055000 ;
      RECT   0.000000  73.055000   9.420000  73.095000 ;
      RECT   0.000000  73.095000   9.415000  73.100000 ;
      RECT   0.000000  73.115000   9.455000  73.200000 ;
      RECT   0.000000  78.450000 480.000000  79.150000 ;
      RECT   0.000000  78.550000 480.000000  79.150000 ;
      RECT   0.000000  84.600000 480.000000  85.200000 ;
      RECT   0.000000  84.600000 480.000000  85.200000 ;
      RECT   0.000000  89.450000 480.000000  90.050000 ;
      RECT   0.000000  89.450000 480.000000  90.050000 ;
      RECT   0.000000  94.300000 480.000000  94.900000 ;
      RECT   0.000000  94.300000 480.000000  94.900000 ;
      RECT   0.000000 100.350000 480.000000 101.050000 ;
      RECT   0.000000 100.350000 480.000000 101.150000 ;
      RECT   0.000000 110.750000 480.000000 111.550000 ;
      RECT   0.000000 110.850000 480.000000 111.550000 ;
      RECT   0.000000 116.800000 480.000000 117.400000 ;
      RECT   0.000000 116.800000 480.000000 117.400000 ;
      RECT   0.000000 122.650000 480.000000 123.350000 ;
      RECT   0.000000 122.650000 480.000000 123.450000 ;
      RECT   0.000000 149.015000  28.960000 159.510000 ;
      RECT   0.000000 149.115000  18.425000 149.265000 ;
      RECT   0.000000 149.115000  18.425000 149.265000 ;
      RECT   0.000000 149.265000  18.575000 149.415000 ;
      RECT   0.000000 149.265000  18.575000 149.415000 ;
      RECT   0.000000 149.415000  18.725000 149.565000 ;
      RECT   0.000000 149.415000  18.725000 149.565000 ;
      RECT   0.000000 149.565000  18.875000 149.715000 ;
      RECT   0.000000 149.565000  18.875000 149.715000 ;
      RECT   0.000000 149.715000  19.025000 149.865000 ;
      RECT   0.000000 149.715000  19.025000 149.865000 ;
      RECT   0.000000 149.865000  19.175000 150.015000 ;
      RECT   0.000000 149.865000  19.175000 150.015000 ;
      RECT   0.000000 150.015000  19.325000 150.165000 ;
      RECT   0.000000 150.015000  19.325000 150.165000 ;
      RECT   0.000000 150.165000  19.475000 150.315000 ;
      RECT   0.000000 150.165000  19.475000 150.315000 ;
      RECT   0.000000 150.315000  19.625000 150.465000 ;
      RECT   0.000000 150.315000  19.625000 150.465000 ;
      RECT   0.000000 150.465000  19.775000 150.615000 ;
      RECT   0.000000 150.465000  19.775000 150.615000 ;
      RECT   0.000000 150.615000  19.925000 150.765000 ;
      RECT   0.000000 150.615000  19.925000 150.765000 ;
      RECT   0.000000 150.765000  20.075000 150.915000 ;
      RECT   0.000000 150.765000  20.075000 150.915000 ;
      RECT   0.000000 150.915000  20.225000 151.065000 ;
      RECT   0.000000 150.915000  20.225000 151.065000 ;
      RECT   0.000000 151.065000  20.375000 151.215000 ;
      RECT   0.000000 151.065000  20.375000 151.215000 ;
      RECT   0.000000 151.215000  20.525000 151.365000 ;
      RECT   0.000000 151.215000  20.525000 151.365000 ;
      RECT   0.000000 151.365000  20.675000 151.515000 ;
      RECT   0.000000 151.365000  20.675000 151.515000 ;
      RECT   0.000000 151.515000  20.825000 151.665000 ;
      RECT   0.000000 151.515000  20.825000 151.665000 ;
      RECT   0.000000 151.665000  20.975000 151.815000 ;
      RECT   0.000000 151.665000  20.975000 151.815000 ;
      RECT   0.000000 151.815000  21.125000 151.965000 ;
      RECT   0.000000 151.815000  21.125000 151.965000 ;
      RECT   0.000000 151.965000  21.275000 152.115000 ;
      RECT   0.000000 151.965000  21.275000 152.115000 ;
      RECT   0.000000 152.115000  21.425000 152.265000 ;
      RECT   0.000000 152.115000  21.425000 152.265000 ;
      RECT   0.000000 152.265000  21.575000 152.415000 ;
      RECT   0.000000 152.265000  21.575000 152.415000 ;
      RECT   0.000000 152.415000  21.725000 152.565000 ;
      RECT   0.000000 152.415000  21.725000 152.565000 ;
      RECT   0.000000 152.565000  21.875000 152.715000 ;
      RECT   0.000000 152.565000  21.875000 152.715000 ;
      RECT   0.000000 152.715000  22.025000 152.865000 ;
      RECT   0.000000 152.715000  22.025000 152.865000 ;
      RECT   0.000000 152.865000  22.175000 153.015000 ;
      RECT   0.000000 152.865000  22.175000 153.015000 ;
      RECT   0.000000 153.015000  22.325000 153.165000 ;
      RECT   0.000000 153.015000  22.325000 153.165000 ;
      RECT   0.000000 153.165000  22.475000 153.315000 ;
      RECT   0.000000 153.165000  22.475000 153.315000 ;
      RECT   0.000000 153.315000  22.625000 153.465000 ;
      RECT   0.000000 153.315000  22.625000 153.465000 ;
      RECT   0.000000 153.465000  22.775000 153.615000 ;
      RECT   0.000000 153.465000  22.775000 153.615000 ;
      RECT   0.000000 153.615000  22.925000 153.765000 ;
      RECT   0.000000 153.615000  22.925000 153.765000 ;
      RECT   0.000000 153.765000  23.075000 153.915000 ;
      RECT   0.000000 153.765000  23.075000 153.915000 ;
      RECT   0.000000 153.915000  23.225000 154.065000 ;
      RECT   0.000000 153.915000  23.225000 154.065000 ;
      RECT   0.000000 154.065000  23.375000 154.215000 ;
      RECT   0.000000 154.065000  23.375000 154.215000 ;
      RECT   0.000000 154.215000  23.525000 154.365000 ;
      RECT   0.000000 154.215000  23.525000 154.365000 ;
      RECT   0.000000 154.365000  23.675000 154.515000 ;
      RECT   0.000000 154.365000  23.675000 154.515000 ;
      RECT   0.000000 154.515000  23.825000 154.665000 ;
      RECT   0.000000 154.515000  23.825000 154.665000 ;
      RECT   0.000000 154.665000  23.975000 154.815000 ;
      RECT   0.000000 154.665000  23.975000 154.815000 ;
      RECT   0.000000 154.815000  24.125000 154.965000 ;
      RECT   0.000000 154.815000  24.125000 154.965000 ;
      RECT   0.000000 154.965000  24.275000 155.115000 ;
      RECT   0.000000 154.965000  24.275000 155.115000 ;
      RECT   0.000000 155.115000  24.425000 155.265000 ;
      RECT   0.000000 155.115000  24.425000 155.265000 ;
      RECT   0.000000 155.265000  24.575000 155.415000 ;
      RECT   0.000000 155.265000  24.575000 155.415000 ;
      RECT   0.000000 155.415000  24.725000 155.565000 ;
      RECT   0.000000 155.415000  24.725000 155.565000 ;
      RECT   0.000000 155.565000  24.875000 155.715000 ;
      RECT   0.000000 155.565000  24.875000 155.715000 ;
      RECT   0.000000 155.715000  25.025000 155.865000 ;
      RECT   0.000000 155.715000  25.025000 155.865000 ;
      RECT   0.000000 155.865000  25.175000 156.015000 ;
      RECT   0.000000 155.865000  25.175000 156.015000 ;
      RECT   0.000000 156.015000  25.325000 156.165000 ;
      RECT   0.000000 156.015000  25.325000 156.165000 ;
      RECT   0.000000 156.165000  25.475000 156.315000 ;
      RECT   0.000000 156.165000  25.475000 156.315000 ;
      RECT   0.000000 156.315000  25.625000 156.465000 ;
      RECT   0.000000 156.315000  25.625000 156.465000 ;
      RECT   0.000000 156.465000  25.775000 156.615000 ;
      RECT   0.000000 156.465000  25.775000 156.615000 ;
      RECT   0.000000 156.615000  25.925000 156.765000 ;
      RECT   0.000000 156.615000  25.925000 156.765000 ;
      RECT   0.000000 156.765000  26.075000 156.915000 ;
      RECT   0.000000 156.765000  26.075000 156.915000 ;
      RECT   0.000000 156.915000  26.225000 157.065000 ;
      RECT   0.000000 156.915000  26.225000 157.065000 ;
      RECT   0.000000 157.065000  26.375000 157.215000 ;
      RECT   0.000000 157.065000  26.375000 157.215000 ;
      RECT   0.000000 157.215000  26.525000 157.365000 ;
      RECT   0.000000 157.215000  26.525000 157.365000 ;
      RECT   0.000000 157.365000  26.675000 157.515000 ;
      RECT   0.000000 157.365000  26.675000 157.515000 ;
      RECT   0.000000 157.515000  26.825000 157.665000 ;
      RECT   0.000000 157.515000  26.825000 157.665000 ;
      RECT   0.000000 157.665000  26.975000 157.815000 ;
      RECT   0.000000 157.665000  26.975000 157.815000 ;
      RECT   0.000000 157.815000  27.125000 157.965000 ;
      RECT   0.000000 157.815000  27.125000 157.965000 ;
      RECT   0.000000 157.965000  27.275000 158.115000 ;
      RECT   0.000000 157.965000  27.275000 158.115000 ;
      RECT   0.000000 158.115000  27.425000 158.265000 ;
      RECT   0.000000 158.115000  27.425000 158.265000 ;
      RECT   0.000000 158.265000  27.575000 158.415000 ;
      RECT   0.000000 158.265000  27.575000 158.415000 ;
      RECT   0.000000 158.415000  27.725000 158.565000 ;
      RECT   0.000000 158.415000  27.725000 158.565000 ;
      RECT   0.000000 158.565000  27.875000 158.715000 ;
      RECT   0.000000 158.565000  27.875000 158.715000 ;
      RECT   0.000000 158.715000  28.025000 158.865000 ;
      RECT   0.000000 158.715000  28.025000 158.865000 ;
      RECT   0.000000 158.865000  28.175000 159.015000 ;
      RECT   0.000000 158.865000  28.175000 159.015000 ;
      RECT   0.000000 159.015000  28.325000 159.165000 ;
      RECT   0.000000 159.015000  28.325000 159.165000 ;
      RECT   0.000000 159.165000  28.475000 159.315000 ;
      RECT   0.000000 159.165000  28.475000 159.315000 ;
      RECT   0.000000 159.315000  28.625000 159.465000 ;
      RECT   0.000000 159.315000  28.625000 159.465000 ;
      RECT   0.000000 159.465000  28.775000 159.550000 ;
      RECT   0.000000 159.465000  28.775000 159.550000 ;
      RECT   0.000000 159.510000  28.960000 207.450000 ;
      RECT   0.000000 159.550000  28.860000 207.490000 ;
      RECT   0.000000 207.450000  49.710000 228.200000 ;
      RECT   0.000000 207.490000  28.860000 207.640000 ;
      RECT   0.000000 207.490000  28.860000 207.640000 ;
      RECT   0.000000 207.640000  29.010000 207.790000 ;
      RECT   0.000000 207.640000  29.010000 207.790000 ;
      RECT   0.000000 207.790000  29.160000 207.940000 ;
      RECT   0.000000 207.790000  29.160000 207.940000 ;
      RECT   0.000000 207.940000  29.310000 208.090000 ;
      RECT   0.000000 207.940000  29.310000 208.090000 ;
      RECT   0.000000 208.090000  29.460000 208.240000 ;
      RECT   0.000000 208.090000  29.460000 208.240000 ;
      RECT   0.000000 208.240000  29.610000 208.390000 ;
      RECT   0.000000 208.240000  29.610000 208.390000 ;
      RECT   0.000000 208.390000  29.760000 208.540000 ;
      RECT   0.000000 208.390000  29.760000 208.540000 ;
      RECT   0.000000 208.540000  29.910000 208.690000 ;
      RECT   0.000000 208.540000  29.910000 208.690000 ;
      RECT   0.000000 208.690000  30.060000 208.840000 ;
      RECT   0.000000 208.690000  30.060000 208.840000 ;
      RECT   0.000000 208.840000  30.210000 208.990000 ;
      RECT   0.000000 208.840000  30.210000 208.990000 ;
      RECT   0.000000 208.990000  30.360000 209.140000 ;
      RECT   0.000000 208.990000  30.360000 209.140000 ;
      RECT   0.000000 209.140000  30.510000 209.290000 ;
      RECT   0.000000 209.140000  30.510000 209.290000 ;
      RECT   0.000000 209.290000  30.660000 209.440000 ;
      RECT   0.000000 209.290000  30.660000 209.440000 ;
      RECT   0.000000 209.440000  30.810000 209.590000 ;
      RECT   0.000000 209.440000  30.810000 209.590000 ;
      RECT   0.000000 209.590000  30.960000 209.740000 ;
      RECT   0.000000 209.590000  30.960000 209.740000 ;
      RECT   0.000000 209.740000  31.110000 209.890000 ;
      RECT   0.000000 209.740000  31.110000 209.890000 ;
      RECT   0.000000 209.890000  31.260000 210.040000 ;
      RECT   0.000000 209.890000  31.260000 210.040000 ;
      RECT   0.000000 210.040000  31.410000 210.190000 ;
      RECT   0.000000 210.040000  31.410000 210.190000 ;
      RECT   0.000000 210.190000  31.560000 210.340000 ;
      RECT   0.000000 210.190000  31.560000 210.340000 ;
      RECT   0.000000 210.340000  31.710000 210.490000 ;
      RECT   0.000000 210.340000  31.710000 210.490000 ;
      RECT   0.000000 210.490000  31.860000 210.640000 ;
      RECT   0.000000 210.490000  31.860000 210.640000 ;
      RECT   0.000000 210.640000  32.010000 210.790000 ;
      RECT   0.000000 210.640000  32.010000 210.790000 ;
      RECT   0.000000 210.790000  32.160000 210.940000 ;
      RECT   0.000000 210.790000  32.160000 210.940000 ;
      RECT   0.000000 210.940000  32.310000 211.090000 ;
      RECT   0.000000 210.940000  32.310000 211.090000 ;
      RECT   0.000000 211.090000  32.460000 211.240000 ;
      RECT   0.000000 211.090000  32.460000 211.240000 ;
      RECT   0.000000 211.240000  32.610000 211.390000 ;
      RECT   0.000000 211.240000  32.610000 211.390000 ;
      RECT   0.000000 211.390000  32.760000 211.540000 ;
      RECT   0.000000 211.390000  32.760000 211.540000 ;
      RECT   0.000000 211.540000  32.910000 211.690000 ;
      RECT   0.000000 211.540000  32.910000 211.690000 ;
      RECT   0.000000 211.690000  33.060000 211.840000 ;
      RECT   0.000000 211.690000  33.060000 211.840000 ;
      RECT   0.000000 211.840000  33.210000 211.990000 ;
      RECT   0.000000 211.840000  33.210000 211.990000 ;
      RECT   0.000000 211.990000  33.360000 212.140000 ;
      RECT   0.000000 211.990000  33.360000 212.140000 ;
      RECT   0.000000 212.140000  33.510000 212.290000 ;
      RECT   0.000000 212.140000  33.510000 212.290000 ;
      RECT   0.000000 212.290000  33.660000 212.440000 ;
      RECT   0.000000 212.290000  33.660000 212.440000 ;
      RECT   0.000000 212.440000  33.810000 212.590000 ;
      RECT   0.000000 212.440000  33.810000 212.590000 ;
      RECT   0.000000 212.590000  33.960000 212.740000 ;
      RECT   0.000000 212.590000  33.960000 212.740000 ;
      RECT   0.000000 212.740000  34.110000 212.890000 ;
      RECT   0.000000 212.740000  34.110000 212.890000 ;
      RECT   0.000000 212.890000  34.260000 213.040000 ;
      RECT   0.000000 212.890000  34.260000 213.040000 ;
      RECT   0.000000 213.040000  34.410000 213.190000 ;
      RECT   0.000000 213.040000  34.410000 213.190000 ;
      RECT   0.000000 213.190000  34.560000 213.340000 ;
      RECT   0.000000 213.190000  34.560000 213.340000 ;
      RECT   0.000000 213.340000  34.710000 213.490000 ;
      RECT   0.000000 213.340000  34.710000 213.490000 ;
      RECT   0.000000 213.490000  34.860000 213.640000 ;
      RECT   0.000000 213.490000  34.860000 213.640000 ;
      RECT   0.000000 213.640000  35.010000 213.790000 ;
      RECT   0.000000 213.640000  35.010000 213.790000 ;
      RECT   0.000000 213.790000  35.160000 213.940000 ;
      RECT   0.000000 213.790000  35.160000 213.940000 ;
      RECT   0.000000 213.940000  35.310000 214.090000 ;
      RECT   0.000000 213.940000  35.310000 214.090000 ;
      RECT   0.000000 214.090000  35.460000 214.240000 ;
      RECT   0.000000 214.090000  35.460000 214.240000 ;
      RECT   0.000000 214.240000  35.610000 214.390000 ;
      RECT   0.000000 214.240000  35.610000 214.390000 ;
      RECT   0.000000 214.390000  35.760000 214.540000 ;
      RECT   0.000000 214.390000  35.760000 214.540000 ;
      RECT   0.000000 214.540000  35.910000 214.690000 ;
      RECT   0.000000 214.540000  35.910000 214.690000 ;
      RECT   0.000000 214.690000  36.060000 214.840000 ;
      RECT   0.000000 214.690000  36.060000 214.840000 ;
      RECT   0.000000 214.840000  36.210000 214.990000 ;
      RECT   0.000000 214.840000  36.210000 214.990000 ;
      RECT   0.000000 214.990000  36.360000 215.140000 ;
      RECT   0.000000 214.990000  36.360000 215.140000 ;
      RECT   0.000000 215.140000  36.510000 215.290000 ;
      RECT   0.000000 215.140000  36.510000 215.290000 ;
      RECT   0.000000 215.290000  36.660000 215.440000 ;
      RECT   0.000000 215.290000  36.660000 215.440000 ;
      RECT   0.000000 215.440000  36.810000 215.590000 ;
      RECT   0.000000 215.440000  36.810000 215.590000 ;
      RECT   0.000000 215.590000  36.960000 215.740000 ;
      RECT   0.000000 215.590000  36.960000 215.740000 ;
      RECT   0.000000 215.740000  37.110000 215.890000 ;
      RECT   0.000000 215.740000  37.110000 215.890000 ;
      RECT   0.000000 215.890000  37.260000 216.040000 ;
      RECT   0.000000 215.890000  37.260000 216.040000 ;
      RECT   0.000000 216.040000  37.410000 216.190000 ;
      RECT   0.000000 216.040000  37.410000 216.190000 ;
      RECT   0.000000 216.190000  37.560000 216.340000 ;
      RECT   0.000000 216.190000  37.560000 216.340000 ;
      RECT   0.000000 216.340000  37.710000 216.490000 ;
      RECT   0.000000 216.340000  37.710000 216.490000 ;
      RECT   0.000000 216.490000  37.860000 216.640000 ;
      RECT   0.000000 216.490000  37.860000 216.640000 ;
      RECT   0.000000 216.640000  38.010000 216.790000 ;
      RECT   0.000000 216.640000  38.010000 216.790000 ;
      RECT   0.000000 216.790000  38.160000 216.940000 ;
      RECT   0.000000 216.790000  38.160000 216.940000 ;
      RECT   0.000000 216.940000  38.310000 217.090000 ;
      RECT   0.000000 216.940000  38.310000 217.090000 ;
      RECT   0.000000 217.090000  38.460000 217.240000 ;
      RECT   0.000000 217.090000  38.460000 217.240000 ;
      RECT   0.000000 217.240000  38.610000 217.390000 ;
      RECT   0.000000 217.240000  38.610000 217.390000 ;
      RECT   0.000000 217.390000  38.760000 217.540000 ;
      RECT   0.000000 217.390000  38.760000 217.540000 ;
      RECT   0.000000 217.540000  38.910000 217.690000 ;
      RECT   0.000000 217.540000  38.910000 217.690000 ;
      RECT   0.000000 217.690000  39.060000 217.840000 ;
      RECT   0.000000 217.690000  39.060000 217.840000 ;
      RECT   0.000000 217.840000  39.210000 217.990000 ;
      RECT   0.000000 217.840000  39.210000 217.990000 ;
      RECT   0.000000 217.990000  39.360000 218.140000 ;
      RECT   0.000000 217.990000  39.360000 218.140000 ;
      RECT   0.000000 218.140000  39.510000 218.290000 ;
      RECT   0.000000 218.140000  39.510000 218.290000 ;
      RECT   0.000000 218.290000  39.660000 218.440000 ;
      RECT   0.000000 218.290000  39.660000 218.440000 ;
      RECT   0.000000 218.440000  39.810000 218.590000 ;
      RECT   0.000000 218.440000  39.810000 218.590000 ;
      RECT   0.000000 218.590000  39.960000 218.740000 ;
      RECT   0.000000 218.590000  39.960000 218.740000 ;
      RECT   0.000000 218.740000  40.110000 218.890000 ;
      RECT   0.000000 218.740000  40.110000 218.890000 ;
      RECT   0.000000 218.890000  40.260000 219.040000 ;
      RECT   0.000000 218.890000  40.260000 219.040000 ;
      RECT   0.000000 219.040000  40.410000 219.190000 ;
      RECT   0.000000 219.040000  40.410000 219.190000 ;
      RECT   0.000000 219.190000  40.560000 219.340000 ;
      RECT   0.000000 219.190000  40.560000 219.340000 ;
      RECT   0.000000 219.340000  40.710000 219.490000 ;
      RECT   0.000000 219.340000  40.710000 219.490000 ;
      RECT   0.000000 219.490000  40.860000 219.640000 ;
      RECT   0.000000 219.490000  40.860000 219.640000 ;
      RECT   0.000000 219.640000  41.010000 219.790000 ;
      RECT   0.000000 219.640000  41.010000 219.790000 ;
      RECT   0.000000 219.790000  41.160000 219.940000 ;
      RECT   0.000000 219.790000  41.160000 219.940000 ;
      RECT   0.000000 219.940000  41.310000 220.090000 ;
      RECT   0.000000 219.940000  41.310000 220.090000 ;
      RECT   0.000000 220.090000  41.460000 220.240000 ;
      RECT   0.000000 220.090000  41.460000 220.240000 ;
      RECT   0.000000 220.240000  41.610000 220.390000 ;
      RECT   0.000000 220.240000  41.610000 220.390000 ;
      RECT   0.000000 220.390000  41.760000 220.540000 ;
      RECT   0.000000 220.390000  41.760000 220.540000 ;
      RECT   0.000000 220.540000  41.910000 220.690000 ;
      RECT   0.000000 220.540000  41.910000 220.690000 ;
      RECT   0.000000 220.690000  42.060000 220.840000 ;
      RECT   0.000000 220.690000  42.060000 220.840000 ;
      RECT   0.000000 220.840000  42.210000 220.990000 ;
      RECT   0.000000 220.840000  42.210000 220.990000 ;
      RECT   0.000000 220.990000  42.360000 221.140000 ;
      RECT   0.000000 220.990000  42.360000 221.140000 ;
      RECT   0.000000 221.140000  42.510000 221.290000 ;
      RECT   0.000000 221.140000  42.510000 221.290000 ;
      RECT   0.000000 221.290000  42.660000 221.440000 ;
      RECT   0.000000 221.290000  42.660000 221.440000 ;
      RECT   0.000000 221.440000  42.810000 221.590000 ;
      RECT   0.000000 221.440000  42.810000 221.590000 ;
      RECT   0.000000 221.590000  42.960000 221.740000 ;
      RECT   0.000000 221.590000  42.960000 221.740000 ;
      RECT   0.000000 221.740000  43.110000 221.890000 ;
      RECT   0.000000 221.740000  43.110000 221.890000 ;
      RECT   0.000000 221.890000  43.260000 222.040000 ;
      RECT   0.000000 221.890000  43.260000 222.040000 ;
      RECT   0.000000 222.040000  43.410000 222.190000 ;
      RECT   0.000000 222.040000  43.410000 222.190000 ;
      RECT   0.000000 222.190000  43.560000 222.340000 ;
      RECT   0.000000 222.190000  43.560000 222.340000 ;
      RECT   0.000000 222.340000  43.710000 222.490000 ;
      RECT   0.000000 222.340000  43.710000 222.490000 ;
      RECT   0.000000 222.490000  43.860000 222.640000 ;
      RECT   0.000000 222.490000  43.860000 222.640000 ;
      RECT   0.000000 222.640000  44.010000 222.790000 ;
      RECT   0.000000 222.640000  44.010000 222.790000 ;
      RECT   0.000000 222.790000  44.160000 222.940000 ;
      RECT   0.000000 222.790000  44.160000 222.940000 ;
      RECT   0.000000 222.940000  44.310000 223.090000 ;
      RECT   0.000000 222.940000  44.310000 223.090000 ;
      RECT   0.000000 223.090000  44.460000 223.240000 ;
      RECT   0.000000 223.090000  44.460000 223.240000 ;
      RECT   0.000000 223.240000  44.610000 223.390000 ;
      RECT   0.000000 223.240000  44.610000 223.390000 ;
      RECT   0.000000 223.390000  44.760000 223.540000 ;
      RECT   0.000000 223.390000  44.760000 223.540000 ;
      RECT   0.000000 223.540000  44.910000 223.690000 ;
      RECT   0.000000 223.540000  44.910000 223.690000 ;
      RECT   0.000000 223.690000  45.060000 223.840000 ;
      RECT   0.000000 223.690000  45.060000 223.840000 ;
      RECT   0.000000 223.840000  45.210000 223.990000 ;
      RECT   0.000000 223.840000  45.210000 223.990000 ;
      RECT   0.000000 223.990000  45.360000 224.140000 ;
      RECT   0.000000 223.990000  45.360000 224.140000 ;
      RECT   0.000000 224.140000  45.510000 224.290000 ;
      RECT   0.000000 224.140000  45.510000 224.290000 ;
      RECT   0.000000 224.290000  45.660000 224.440000 ;
      RECT   0.000000 224.290000  45.660000 224.440000 ;
      RECT   0.000000 224.440000  45.810000 224.590000 ;
      RECT   0.000000 224.440000  45.810000 224.590000 ;
      RECT   0.000000 224.590000  45.960000 224.740000 ;
      RECT   0.000000 224.590000  45.960000 224.740000 ;
      RECT   0.000000 224.740000  46.110000 224.890000 ;
      RECT   0.000000 224.740000  46.110000 224.890000 ;
      RECT   0.000000 224.890000  46.260000 225.040000 ;
      RECT   0.000000 224.890000  46.260000 225.040000 ;
      RECT   0.000000 225.040000  46.410000 225.190000 ;
      RECT   0.000000 225.040000  46.410000 225.190000 ;
      RECT   0.000000 225.190000  46.560000 225.340000 ;
      RECT   0.000000 225.190000  46.560000 225.340000 ;
      RECT   0.000000 225.340000  46.710000 225.490000 ;
      RECT   0.000000 225.340000  46.710000 225.490000 ;
      RECT   0.000000 225.490000  46.860000 225.640000 ;
      RECT   0.000000 225.490000  46.860000 225.640000 ;
      RECT   0.000000 225.640000  47.010000 225.790000 ;
      RECT   0.000000 225.640000  47.010000 225.790000 ;
      RECT   0.000000 225.790000  47.160000 225.940000 ;
      RECT   0.000000 225.790000  47.160000 225.940000 ;
      RECT   0.000000 225.940000  47.310000 226.090000 ;
      RECT   0.000000 225.940000  47.310000 226.090000 ;
      RECT   0.000000 226.090000  47.460000 226.240000 ;
      RECT   0.000000 226.090000  47.460000 226.240000 ;
      RECT   0.000000 226.240000  47.610000 226.390000 ;
      RECT   0.000000 226.240000  47.610000 226.390000 ;
      RECT   0.000000 226.390000  47.760000 226.540000 ;
      RECT   0.000000 226.390000  47.760000 226.540000 ;
      RECT   0.000000 226.540000  47.910000 226.690000 ;
      RECT   0.000000 226.540000  47.910000 226.690000 ;
      RECT   0.000000 226.690000  48.060000 226.840000 ;
      RECT   0.000000 226.690000  48.060000 226.840000 ;
      RECT   0.000000 226.840000  48.210000 226.990000 ;
      RECT   0.000000 226.840000  48.210000 226.990000 ;
      RECT   0.000000 226.990000  48.360000 227.140000 ;
      RECT   0.000000 226.990000  48.360000 227.140000 ;
      RECT   0.000000 227.140000  48.510000 227.290000 ;
      RECT   0.000000 227.140000  48.510000 227.290000 ;
      RECT   0.000000 227.290000  48.660000 227.440000 ;
      RECT   0.000000 227.290000  48.660000 227.440000 ;
      RECT   0.000000 227.440000  48.810000 227.590000 ;
      RECT   0.000000 227.440000  48.810000 227.590000 ;
      RECT   0.000000 227.590000  48.960000 227.740000 ;
      RECT   0.000000 227.590000  48.960000 227.740000 ;
      RECT   0.000000 227.740000  49.110000 227.890000 ;
      RECT   0.000000 227.740000  49.110000 227.890000 ;
      RECT   0.000000 227.890000  49.260000 228.040000 ;
      RECT   0.000000 227.890000  49.260000 228.040000 ;
      RECT   0.000000 228.040000  49.410000 228.190000 ;
      RECT   0.000000 228.040000  49.410000 228.190000 ;
      RECT   0.000000 228.190000  49.560000 228.340000 ;
      RECT   0.000000 228.190000  49.560000 228.340000 ;
      RECT   0.000000 228.200000 480.000000 229.100000 ;
      RECT   0.000000 228.340000  49.710000 228.490000 ;
      RECT   0.000000 228.340000  49.710000 228.490000 ;
      RECT   0.000000 228.490000  49.860000 228.640000 ;
      RECT   0.000000 228.490000  49.860000 228.640000 ;
      RECT   0.000000 228.640000  50.010000 228.790000 ;
      RECT   0.000000 228.640000  50.010000 228.790000 ;
      RECT   0.000000 228.790000  50.160000 228.940000 ;
      RECT   0.000000 228.790000  50.160000 228.940000 ;
      RECT   0.000000 228.940000  50.310000 229.090000 ;
      RECT   0.000000 228.940000  50.310000 229.090000 ;
      RECT   0.000000 229.090000  50.460000 229.100000 ;
      RECT   0.000000 229.090000  50.460000 229.100000 ;
      RECT  28.940000 123.450000 468.500000 123.550000 ;
      RECT  29.030000 123.350000 468.510000 123.400000 ;
      RECT  29.080000 123.400000 468.460000 123.450000 ;
      RECT  29.230000 123.550000 468.310000 123.740000 ;
      RECT  29.230000 123.740000 443.095000 148.955000 ;
      RECT  29.330000 123.450000 468.335000 123.575000 ;
      RECT  29.330000 123.575000 468.210000 123.700000 ;
      RECT  29.480000 123.700000 468.060000 123.850000 ;
      RECT  29.630000 123.850000 467.910000 124.000000 ;
      RECT  29.780000 124.000000 467.760000 124.150000 ;
      RECT  29.930000 124.150000 467.610000 124.300000 ;
      RECT  30.080000 124.300000 467.460000 124.450000 ;
      RECT  30.230000 124.450000 467.310000 124.600000 ;
      RECT  30.380000 124.600000 467.160000 124.750000 ;
      RECT  30.530000 124.750000 467.010000 124.900000 ;
      RECT  30.680000 124.900000 466.860000 125.050000 ;
      RECT  30.830000 125.050000 466.710000 125.200000 ;
      RECT  30.980000 125.200000 466.560000 125.350000 ;
      RECT  31.130000 125.350000 466.410000 125.500000 ;
      RECT  31.280000 125.500000 466.260000 125.650000 ;
      RECT  31.430000 125.650000 466.110000 125.800000 ;
      RECT  31.580000 125.800000 465.960000 125.950000 ;
      RECT  31.730000 125.950000 465.810000 126.100000 ;
      RECT  31.880000 126.100000 465.660000 126.250000 ;
      RECT  32.030000 126.250000 465.510000 126.400000 ;
      RECT  32.180000 126.400000 465.360000 126.550000 ;
      RECT  32.330000 126.550000 465.210000 126.700000 ;
      RECT  32.480000 126.700000 465.060000 126.850000 ;
      RECT  32.630000 126.850000 464.910000 127.000000 ;
      RECT  32.780000 127.000000 464.760000 127.150000 ;
      RECT  32.930000 127.150000 464.610000 127.300000 ;
      RECT  33.080000 127.300000 464.460000 127.450000 ;
      RECT  33.230000 127.450000 464.310000 127.600000 ;
      RECT  33.380000 127.600000 464.160000 127.750000 ;
      RECT  33.530000 127.750000 464.010000 127.900000 ;
      RECT  33.680000 127.900000 463.860000 128.050000 ;
      RECT  33.830000 128.050000 463.710000 128.200000 ;
      RECT  33.980000 128.200000 463.560000 128.350000 ;
      RECT  34.130000 128.350000 463.410000 128.500000 ;
      RECT  34.280000 128.500000 463.260000 128.650000 ;
      RECT  34.430000 128.650000 463.110000 128.800000 ;
      RECT  34.580000 128.800000 462.960000 128.950000 ;
      RECT  34.730000 128.950000 462.810000 129.100000 ;
      RECT  34.880000 129.100000 462.660000 129.250000 ;
      RECT  35.030000 129.250000 462.510000 129.400000 ;
      RECT  35.180000 129.400000 462.360000 129.550000 ;
      RECT  35.330000 129.550000 462.210000 129.700000 ;
      RECT  35.480000 129.700000 462.060000 129.850000 ;
      RECT  35.630000 129.850000 461.910000 130.000000 ;
      RECT  35.780000 130.000000 461.760000 130.150000 ;
      RECT  35.930000 130.150000 461.610000 130.300000 ;
      RECT  36.080000 130.300000 461.460000 130.450000 ;
      RECT  36.230000 130.450000 461.310000 130.600000 ;
      RECT  36.380000 130.600000 461.160000 130.750000 ;
      RECT  36.530000 130.750000 461.010000 130.900000 ;
      RECT  36.680000 130.900000 460.860000 131.050000 ;
      RECT  36.830000 131.050000 460.710000 131.200000 ;
      RECT  36.980000 131.200000 460.560000 131.350000 ;
      RECT  37.130000 131.350000 460.410000 131.500000 ;
      RECT  37.280000 131.500000 460.260000 131.650000 ;
      RECT  37.430000 131.650000 460.110000 131.800000 ;
      RECT  37.580000 131.800000 459.960000 131.950000 ;
      RECT  37.730000 131.950000 459.810000 132.100000 ;
      RECT  37.880000 132.100000 459.660000 132.250000 ;
      RECT  38.030000 132.250000 459.510000 132.400000 ;
      RECT  38.180000 132.400000 459.360000 132.550000 ;
      RECT  38.330000 132.550000 459.210000 132.700000 ;
      RECT  38.480000 132.700000 459.060000 132.850000 ;
      RECT  38.630000 132.850000 458.910000 133.000000 ;
      RECT  38.780000 133.000000 458.760000 133.150000 ;
      RECT  38.930000 133.150000 458.610000 133.300000 ;
      RECT  39.080000 133.300000 458.460000 133.450000 ;
      RECT  39.230000 133.450000 458.310000 133.600000 ;
      RECT  39.380000 133.600000 458.160000 133.750000 ;
      RECT  39.530000 133.750000 458.010000 133.900000 ;
      RECT  39.680000 133.900000 457.860000 134.050000 ;
      RECT  39.830000 134.050000 457.710000 134.200000 ;
      RECT  39.980000 134.200000 457.560000 134.350000 ;
      RECT  40.130000 134.350000 457.410000 134.500000 ;
      RECT  40.280000 134.500000 457.260000 134.650000 ;
      RECT  40.430000 134.650000 457.110000 134.800000 ;
      RECT  40.580000 134.800000 456.960000 134.950000 ;
      RECT  40.730000 134.950000 456.810000 135.100000 ;
      RECT  40.880000 135.100000 456.660000 135.250000 ;
      RECT  41.030000 135.250000 456.510000 135.400000 ;
      RECT  41.180000 135.400000 456.360000 135.550000 ;
      RECT  41.330000 135.550000 456.210000 135.700000 ;
      RECT  41.480000 135.700000 456.060000 135.850000 ;
      RECT  41.630000 135.850000 455.910000 136.000000 ;
      RECT  41.780000 136.000000 455.760000 136.150000 ;
      RECT  41.930000 136.150000 455.610000 136.300000 ;
      RECT  42.080000 136.300000 455.460000 136.450000 ;
      RECT  42.230000 136.450000 455.310000 136.600000 ;
      RECT  42.380000 136.600000 455.160000 136.750000 ;
      RECT  42.530000 136.750000 455.010000 136.900000 ;
      RECT  42.680000 136.900000 454.860000 137.050000 ;
      RECT  42.830000 137.050000 454.710000 137.200000 ;
      RECT  42.980000 137.200000 454.560000 137.350000 ;
      RECT  43.130000 137.350000 454.410000 137.500000 ;
      RECT  43.280000 137.500000 454.260000 137.650000 ;
      RECT  43.430000 137.650000 454.110000 137.800000 ;
      RECT  43.580000 137.800000 453.960000 137.950000 ;
      RECT  43.730000 137.950000 453.810000 138.100000 ;
      RECT  43.880000 138.100000 453.660000 138.250000 ;
      RECT  44.030000 138.250000 453.510000 138.400000 ;
      RECT  44.180000 138.400000 453.360000 138.550000 ;
      RECT  44.330000 138.550000 453.210000 138.700000 ;
      RECT  44.480000 138.700000 453.060000 138.850000 ;
      RECT  44.630000 138.850000 452.910000 139.000000 ;
      RECT  44.780000 139.000000 452.760000 139.150000 ;
      RECT  44.930000 139.150000 452.610000 139.300000 ;
      RECT  45.080000 139.300000 452.460000 139.450000 ;
      RECT  45.230000 139.450000 452.310000 139.600000 ;
      RECT  45.380000 139.600000 452.160000 139.750000 ;
      RECT  45.530000 139.750000 452.010000 139.900000 ;
      RECT  45.680000 139.900000 451.860000 140.050000 ;
      RECT  45.830000 140.050000 451.710000 140.200000 ;
      RECT  45.980000 140.200000 451.560000 140.350000 ;
      RECT  46.130000 140.350000 451.410000 140.500000 ;
      RECT  46.280000 140.500000 451.260000 140.650000 ;
      RECT  46.430000 140.650000 451.110000 140.800000 ;
      RECT  46.580000 140.800000 450.960000 140.950000 ;
      RECT  46.730000 140.950000 450.810000 141.100000 ;
      RECT  46.880000 141.100000 450.660000 141.250000 ;
      RECT  47.030000 141.250000 450.510000 141.400000 ;
      RECT  47.180000 141.400000 450.360000 141.550000 ;
      RECT  47.330000 141.550000 450.210000 141.700000 ;
      RECT  47.480000 141.700000 450.060000 141.850000 ;
      RECT  47.630000 141.850000 449.910000 142.000000 ;
      RECT  47.780000 142.000000 449.760000 142.150000 ;
      RECT  47.930000 142.150000 449.610000 142.300000 ;
      RECT  48.080000 142.300000 449.460000 142.450000 ;
      RECT  48.230000 142.450000 449.310000 142.600000 ;
      RECT  48.380000 142.600000 449.160000 142.750000 ;
      RECT  48.530000 142.750000 449.010000 142.900000 ;
      RECT  48.680000 142.900000 448.860000 143.050000 ;
      RECT  48.830000 143.050000 448.710000 143.200000 ;
      RECT  48.980000 143.200000 448.560000 143.350000 ;
      RECT  49.130000 143.350000 448.410000 143.500000 ;
      RECT  49.280000 143.500000 448.260000 143.650000 ;
      RECT  49.430000 143.650000 448.110000 143.800000 ;
      RECT  49.580000 143.800000 447.960000 143.950000 ;
      RECT  49.730000 143.950000 447.810000 144.100000 ;
      RECT  49.820000 228.300000 399.300000 228.450000 ;
      RECT  49.880000 144.100000 447.660000 144.250000 ;
      RECT  49.970000 228.450000 399.150000 228.600000 ;
      RECT  50.030000 144.250000 447.510000 144.400000 ;
      RECT  50.120000 228.600000 399.000000 228.750000 ;
      RECT  50.180000 144.400000 447.360000 144.550000 ;
      RECT  50.270000 228.750000 398.850000 228.900000 ;
      RECT  50.330000 144.550000 447.210000 144.700000 ;
      RECT  50.420000 228.900000 398.700000 229.050000 ;
      RECT  50.470000 229.050000 398.650000 229.100000 ;
      RECT  50.480000 144.700000 447.060000 144.850000 ;
      RECT  50.630000 144.850000 446.910000 145.000000 ;
      RECT  50.780000 145.000000 446.760000 145.150000 ;
      RECT  50.930000 145.150000 446.610000 145.300000 ;
      RECT  51.080000 145.300000 446.460000 145.450000 ;
      RECT  51.230000 145.450000 446.310000 145.600000 ;
      RECT  51.380000 145.600000 446.160000 145.750000 ;
      RECT  51.530000 145.750000 446.010000 145.900000 ;
      RECT  51.680000 145.900000 445.860000 146.050000 ;
      RECT  51.830000 146.050000 445.710000 146.200000 ;
      RECT  51.980000 146.200000 445.560000 146.350000 ;
      RECT  52.130000 146.350000 445.410000 146.500000 ;
      RECT  52.280000 146.500000 445.260000 146.650000 ;
      RECT  52.430000 146.650000 445.110000 146.800000 ;
      RECT  52.580000 146.800000 444.960000 146.950000 ;
      RECT  52.730000 146.950000 444.810000 147.100000 ;
      RECT  52.880000 147.100000 444.660000 147.250000 ;
      RECT  53.030000 147.250000 444.510000 147.400000 ;
      RECT  53.180000 147.400000 444.360000 147.550000 ;
      RECT  53.330000 147.550000 444.210000 147.700000 ;
      RECT  53.480000 147.700000 444.060000 147.850000 ;
      RECT  53.630000 147.850000 443.910000 148.000000 ;
      RECT  53.780000 148.000000 443.760000 148.150000 ;
      RECT  53.930000 148.150000 443.610000 148.300000 ;
      RECT  54.080000 148.300000 443.460000 148.450000 ;
      RECT  54.230000 148.450000 443.310000 148.600000 ;
      RECT  54.380000 148.600000 443.160000 148.750000 ;
      RECT  54.445000 148.955000 394.575000 197.475000 ;
      RECT  54.445000 197.475000 387.845000 204.205000 ;
      RECT  54.530000 148.750000 443.010000 148.900000 ;
      RECT  54.545000 148.900000 442.995000 148.915000 ;
      RECT  54.545000 148.915000 442.845000 149.065000 ;
      RECT  54.545000 149.065000 442.695000 149.215000 ;
      RECT  54.545000 149.215000 442.545000 149.365000 ;
      RECT  54.545000 149.365000 442.395000 149.515000 ;
      RECT  54.545000 149.515000 442.245000 149.665000 ;
      RECT  54.545000 149.665000 442.095000 149.815000 ;
      RECT  54.545000 149.815000 441.945000 149.965000 ;
      RECT  54.545000 149.965000 441.795000 150.115000 ;
      RECT  54.545000 150.115000 441.645000 150.265000 ;
      RECT  54.545000 150.265000 441.495000 150.415000 ;
      RECT  54.545000 150.415000 441.345000 150.565000 ;
      RECT  54.545000 150.565000 441.195000 150.715000 ;
      RECT  54.545000 150.715000 441.045000 150.865000 ;
      RECT  54.545000 150.865000 440.895000 151.015000 ;
      RECT  54.545000 151.015000 440.745000 151.165000 ;
      RECT  54.545000 151.165000 440.595000 151.315000 ;
      RECT  54.545000 151.315000 440.445000 151.465000 ;
      RECT  54.545000 151.465000 440.295000 151.615000 ;
      RECT  54.545000 151.615000 440.145000 151.765000 ;
      RECT  54.545000 151.765000 439.995000 151.915000 ;
      RECT  54.545000 151.915000 439.845000 152.065000 ;
      RECT  54.545000 152.065000 439.695000 152.215000 ;
      RECT  54.545000 152.215000 439.545000 152.365000 ;
      RECT  54.545000 152.365000 439.395000 152.515000 ;
      RECT  54.545000 152.515000 439.245000 152.665000 ;
      RECT  54.545000 152.665000 439.095000 152.815000 ;
      RECT  54.545000 152.815000 438.945000 152.965000 ;
      RECT  54.545000 152.965000 438.795000 153.115000 ;
      RECT  54.545000 153.115000 438.645000 153.265000 ;
      RECT  54.545000 153.265000 438.495000 153.415000 ;
      RECT  54.545000 153.415000 438.345000 153.565000 ;
      RECT  54.545000 153.565000 438.195000 153.715000 ;
      RECT  54.545000 153.715000 438.045000 153.865000 ;
      RECT  54.545000 153.865000 437.895000 154.015000 ;
      RECT  54.545000 154.015000 437.745000 154.165000 ;
      RECT  54.545000 154.165000 437.595000 154.315000 ;
      RECT  54.545000 154.315000 437.445000 154.465000 ;
      RECT  54.545000 154.465000 437.295000 154.615000 ;
      RECT  54.545000 154.615000 437.145000 154.765000 ;
      RECT  54.545000 154.765000 436.995000 154.915000 ;
      RECT  54.545000 154.915000 436.845000 155.065000 ;
      RECT  54.545000 155.065000 436.695000 155.215000 ;
      RECT  54.545000 155.215000 436.545000 155.365000 ;
      RECT  54.545000 155.365000 436.395000 155.515000 ;
      RECT  54.545000 155.515000 436.245000 155.665000 ;
      RECT  54.545000 155.665000 436.095000 155.815000 ;
      RECT  54.545000 155.815000 435.945000 155.965000 ;
      RECT  54.545000 155.965000 435.795000 156.115000 ;
      RECT  54.545000 156.115000 435.645000 156.265000 ;
      RECT  54.545000 156.265000 435.495000 156.415000 ;
      RECT  54.545000 156.415000 435.345000 156.565000 ;
      RECT  54.545000 156.565000 435.195000 156.715000 ;
      RECT  54.545000 156.715000 435.045000 156.865000 ;
      RECT  54.545000 156.865000 434.895000 157.015000 ;
      RECT  54.545000 157.015000 434.745000 157.165000 ;
      RECT  54.545000 157.165000 434.595000 157.315000 ;
      RECT  54.545000 157.315000 434.445000 157.465000 ;
      RECT  54.545000 157.465000 434.295000 157.615000 ;
      RECT  54.545000 157.615000 434.145000 157.765000 ;
      RECT  54.545000 157.765000 433.995000 157.915000 ;
      RECT  54.545000 157.915000 433.845000 158.065000 ;
      RECT  54.545000 158.065000 433.695000 158.215000 ;
      RECT  54.545000 158.215000 433.545000 158.365000 ;
      RECT  54.545000 158.365000 433.395000 158.515000 ;
      RECT  54.545000 158.515000 433.245000 158.665000 ;
      RECT  54.545000 158.665000 433.095000 158.815000 ;
      RECT  54.545000 158.815000 432.945000 158.965000 ;
      RECT  54.545000 158.965000 432.795000 159.115000 ;
      RECT  54.545000 159.115000 432.645000 159.265000 ;
      RECT  54.545000 159.265000 432.495000 159.415000 ;
      RECT  54.545000 159.415000 432.345000 159.565000 ;
      RECT  54.545000 159.565000 432.195000 159.715000 ;
      RECT  54.545000 159.715000 432.045000 159.865000 ;
      RECT  54.545000 159.865000 431.895000 160.015000 ;
      RECT  54.545000 160.015000 431.745000 160.165000 ;
      RECT  54.545000 160.165000 431.595000 160.315000 ;
      RECT  54.545000 160.315000 431.445000 160.465000 ;
      RECT  54.545000 160.465000 431.295000 160.615000 ;
      RECT  54.545000 160.615000 431.145000 160.765000 ;
      RECT  54.545000 160.765000 430.995000 160.915000 ;
      RECT  54.545000 160.915000 430.845000 161.065000 ;
      RECT  54.545000 161.065000 430.695000 161.215000 ;
      RECT  54.545000 161.215000 430.545000 161.365000 ;
      RECT  54.545000 161.365000 430.395000 161.515000 ;
      RECT  54.545000 161.515000 430.245000 161.665000 ;
      RECT  54.545000 161.665000 430.095000 161.815000 ;
      RECT  54.545000 161.815000 429.945000 161.965000 ;
      RECT  54.545000 161.965000 429.795000 162.115000 ;
      RECT  54.545000 162.115000 429.645000 162.265000 ;
      RECT  54.545000 162.265000 429.495000 162.415000 ;
      RECT  54.545000 162.415000 429.345000 162.565000 ;
      RECT  54.545000 162.565000 429.195000 162.715000 ;
      RECT  54.545000 162.715000 429.045000 162.865000 ;
      RECT  54.545000 162.865000 428.895000 163.015000 ;
      RECT  54.545000 163.015000 428.745000 163.165000 ;
      RECT  54.545000 163.165000 428.595000 163.315000 ;
      RECT  54.545000 163.315000 428.445000 163.465000 ;
      RECT  54.545000 163.465000 428.295000 163.615000 ;
      RECT  54.545000 163.615000 428.145000 163.765000 ;
      RECT  54.545000 163.765000 427.995000 163.915000 ;
      RECT  54.545000 163.915000 427.845000 164.065000 ;
      RECT  54.545000 164.065000 427.695000 164.215000 ;
      RECT  54.545000 164.215000 427.545000 164.365000 ;
      RECT  54.545000 164.365000 427.395000 164.515000 ;
      RECT  54.545000 164.515000 427.245000 164.665000 ;
      RECT  54.545000 164.665000 427.095000 164.815000 ;
      RECT  54.545000 164.815000 426.945000 164.965000 ;
      RECT  54.545000 164.965000 426.795000 165.115000 ;
      RECT  54.545000 165.115000 426.645000 165.265000 ;
      RECT  54.545000 165.265000 426.495000 165.415000 ;
      RECT  54.545000 165.415000 426.345000 165.565000 ;
      RECT  54.545000 165.565000 426.195000 165.715000 ;
      RECT  54.545000 165.715000 426.045000 165.865000 ;
      RECT  54.545000 165.865000 425.895000 166.015000 ;
      RECT  54.545000 166.015000 425.745000 166.165000 ;
      RECT  54.545000 166.165000 425.595000 166.315000 ;
      RECT  54.545000 166.315000 425.445000 166.465000 ;
      RECT  54.545000 166.465000 425.295000 166.615000 ;
      RECT  54.545000 166.615000 425.145000 166.765000 ;
      RECT  54.545000 166.765000 424.995000 166.915000 ;
      RECT  54.545000 166.915000 424.845000 167.065000 ;
      RECT  54.545000 167.065000 424.695000 167.215000 ;
      RECT  54.545000 167.215000 424.545000 167.365000 ;
      RECT  54.545000 167.365000 424.395000 167.515000 ;
      RECT  54.545000 167.515000 424.245000 167.665000 ;
      RECT  54.545000 167.665000 424.095000 167.815000 ;
      RECT  54.545000 167.815000 423.945000 167.965000 ;
      RECT  54.545000 167.965000 423.795000 168.115000 ;
      RECT  54.545000 168.115000 423.645000 168.265000 ;
      RECT  54.545000 168.265000 423.495000 168.415000 ;
      RECT  54.545000 168.415000 423.345000 168.565000 ;
      RECT  54.545000 168.565000 423.195000 168.715000 ;
      RECT  54.545000 168.715000 423.045000 168.865000 ;
      RECT  54.545000 168.865000 422.895000 169.015000 ;
      RECT  54.545000 169.015000 422.745000 169.165000 ;
      RECT  54.545000 169.165000 422.595000 169.315000 ;
      RECT  54.545000 169.315000 422.445000 169.465000 ;
      RECT  54.545000 169.465000 422.295000 169.615000 ;
      RECT  54.545000 169.615000 422.145000 169.765000 ;
      RECT  54.545000 169.765000 421.995000 169.915000 ;
      RECT  54.545000 169.915000 421.845000 170.065000 ;
      RECT  54.545000 170.065000 421.695000 170.215000 ;
      RECT  54.545000 170.215000 421.545000 170.365000 ;
      RECT  54.545000 170.365000 421.395000 170.515000 ;
      RECT  54.545000 170.515000 421.245000 170.665000 ;
      RECT  54.545000 170.665000 421.095000 170.815000 ;
      RECT  54.545000 170.815000 420.945000 170.965000 ;
      RECT  54.545000 170.965000 420.795000 171.115000 ;
      RECT  54.545000 171.115000 420.645000 171.265000 ;
      RECT  54.545000 171.265000 420.495000 171.415000 ;
      RECT  54.545000 171.415000 420.345000 171.565000 ;
      RECT  54.545000 171.565000 420.195000 171.715000 ;
      RECT  54.545000 171.715000 420.045000 171.865000 ;
      RECT  54.545000 171.865000 419.895000 172.015000 ;
      RECT  54.545000 172.015000 419.745000 172.165000 ;
      RECT  54.545000 172.165000 419.595000 172.315000 ;
      RECT  54.545000 172.315000 419.445000 172.465000 ;
      RECT  54.545000 172.465000 419.295000 172.615000 ;
      RECT  54.545000 172.615000 419.145000 172.765000 ;
      RECT  54.545000 172.765000 418.995000 172.915000 ;
      RECT  54.545000 172.915000 418.845000 173.065000 ;
      RECT  54.545000 173.065000 418.695000 173.215000 ;
      RECT  54.545000 173.215000 418.545000 173.365000 ;
      RECT  54.545000 173.365000 418.395000 173.515000 ;
      RECT  54.545000 173.515000 418.245000 173.665000 ;
      RECT  54.545000 173.665000 418.095000 173.815000 ;
      RECT  54.545000 173.815000 417.945000 173.965000 ;
      RECT  54.545000 173.965000 417.795000 174.115000 ;
      RECT  54.545000 174.115000 417.645000 174.265000 ;
      RECT  54.545000 174.265000 417.495000 174.415000 ;
      RECT  54.545000 174.415000 417.345000 174.565000 ;
      RECT  54.545000 174.565000 417.195000 174.715000 ;
      RECT  54.545000 174.715000 417.045000 174.865000 ;
      RECT  54.545000 174.865000 416.895000 175.015000 ;
      RECT  54.545000 175.015000 416.745000 175.165000 ;
      RECT  54.545000 175.165000 416.595000 175.315000 ;
      RECT  54.545000 175.315000 416.445000 175.465000 ;
      RECT  54.545000 175.465000 416.295000 175.615000 ;
      RECT  54.545000 175.615000 416.145000 175.765000 ;
      RECT  54.545000 175.765000 415.995000 175.915000 ;
      RECT  54.545000 175.915000 415.845000 176.065000 ;
      RECT  54.545000 176.065000 415.695000 176.215000 ;
      RECT  54.545000 176.215000 415.545000 176.365000 ;
      RECT  54.545000 176.365000 415.395000 176.515000 ;
      RECT  54.545000 176.515000 415.245000 176.665000 ;
      RECT  54.545000 176.665000 415.095000 176.815000 ;
      RECT  54.545000 176.815000 414.945000 176.965000 ;
      RECT  54.545000 176.965000 414.795000 177.115000 ;
      RECT  54.545000 177.115000 414.645000 177.265000 ;
      RECT  54.545000 177.265000 414.495000 177.415000 ;
      RECT  54.545000 177.415000 414.345000 177.565000 ;
      RECT  54.545000 177.565000 414.195000 177.715000 ;
      RECT  54.545000 177.715000 414.045000 177.865000 ;
      RECT  54.545000 177.865000 413.895000 178.015000 ;
      RECT  54.545000 178.015000 413.745000 178.165000 ;
      RECT  54.545000 178.165000 413.595000 178.315000 ;
      RECT  54.545000 178.315000 413.445000 178.465000 ;
      RECT  54.545000 178.465000 413.295000 178.615000 ;
      RECT  54.545000 178.615000 413.145000 178.765000 ;
      RECT  54.545000 178.765000 412.995000 178.915000 ;
      RECT  54.545000 178.915000 412.845000 179.065000 ;
      RECT  54.545000 179.065000 412.695000 179.215000 ;
      RECT  54.545000 179.215000 412.545000 179.365000 ;
      RECT  54.545000 179.365000 412.395000 179.515000 ;
      RECT  54.545000 179.515000 412.245000 179.665000 ;
      RECT  54.545000 179.665000 412.095000 179.815000 ;
      RECT  54.545000 179.815000 411.945000 179.965000 ;
      RECT  54.545000 179.965000 411.795000 180.115000 ;
      RECT  54.545000 180.115000 411.645000 180.265000 ;
      RECT  54.545000 180.265000 411.495000 180.415000 ;
      RECT  54.545000 180.415000 411.345000 180.565000 ;
      RECT  54.545000 180.565000 411.195000 180.715000 ;
      RECT  54.545000 180.715000 411.045000 180.865000 ;
      RECT  54.545000 180.865000 410.895000 181.015000 ;
      RECT  54.545000 181.015000 410.745000 181.165000 ;
      RECT  54.545000 181.165000 410.595000 181.315000 ;
      RECT  54.545000 181.315000 410.445000 181.465000 ;
      RECT  54.545000 181.465000 410.295000 181.615000 ;
      RECT  54.545000 181.615000 410.145000 181.765000 ;
      RECT  54.545000 181.765000 409.995000 181.915000 ;
      RECT  54.545000 181.915000 409.845000 182.065000 ;
      RECT  54.545000 182.065000 409.695000 182.215000 ;
      RECT  54.545000 182.215000 409.545000 182.365000 ;
      RECT  54.545000 182.365000 409.395000 182.515000 ;
      RECT  54.545000 182.515000 409.245000 182.665000 ;
      RECT  54.545000 182.665000 409.095000 182.815000 ;
      RECT  54.545000 182.815000 408.945000 182.965000 ;
      RECT  54.545000 182.965000 408.795000 183.115000 ;
      RECT  54.545000 183.115000 408.645000 183.265000 ;
      RECT  54.545000 183.265000 408.495000 183.415000 ;
      RECT  54.545000 183.415000 408.345000 183.565000 ;
      RECT  54.545000 183.565000 408.195000 183.715000 ;
      RECT  54.545000 183.715000 408.045000 183.865000 ;
      RECT  54.545000 183.865000 407.895000 184.015000 ;
      RECT  54.545000 184.015000 407.745000 184.165000 ;
      RECT  54.545000 184.165000 407.595000 184.315000 ;
      RECT  54.545000 184.315000 407.445000 184.465000 ;
      RECT  54.545000 184.465000 407.295000 184.615000 ;
      RECT  54.545000 184.615000 407.145000 184.765000 ;
      RECT  54.545000 184.765000 406.995000 184.915000 ;
      RECT  54.545000 184.915000 406.845000 185.065000 ;
      RECT  54.545000 185.065000 406.695000 185.215000 ;
      RECT  54.545000 185.215000 406.545000 185.365000 ;
      RECT  54.545000 185.365000 406.395000 185.515000 ;
      RECT  54.545000 185.515000 406.245000 185.665000 ;
      RECT  54.545000 185.665000 406.095000 185.815000 ;
      RECT  54.545000 185.815000 405.945000 185.965000 ;
      RECT  54.545000 185.965000 405.795000 186.115000 ;
      RECT  54.545000 186.115000 405.645000 186.265000 ;
      RECT  54.545000 186.265000 405.495000 186.415000 ;
      RECT  54.545000 186.415000 405.345000 186.565000 ;
      RECT  54.545000 186.565000 405.195000 186.715000 ;
      RECT  54.545000 186.715000 405.045000 186.865000 ;
      RECT  54.545000 186.865000 404.895000 187.015000 ;
      RECT  54.545000 187.015000 404.745000 187.165000 ;
      RECT  54.545000 187.165000 404.595000 187.315000 ;
      RECT  54.545000 187.315000 404.445000 187.465000 ;
      RECT  54.545000 187.465000 404.295000 187.615000 ;
      RECT  54.545000 187.615000 404.145000 187.765000 ;
      RECT  54.545000 187.765000 403.995000 187.915000 ;
      RECT  54.545000 187.915000 403.845000 188.065000 ;
      RECT  54.545000 188.065000 403.695000 188.215000 ;
      RECT  54.545000 188.215000 403.545000 188.365000 ;
      RECT  54.545000 188.365000 403.395000 188.515000 ;
      RECT  54.545000 188.515000 403.245000 188.665000 ;
      RECT  54.545000 188.665000 403.095000 188.815000 ;
      RECT  54.545000 188.815000 402.945000 188.965000 ;
      RECT  54.545000 188.965000 402.795000 189.115000 ;
      RECT  54.545000 189.115000 402.645000 189.265000 ;
      RECT  54.545000 189.265000 402.495000 189.415000 ;
      RECT  54.545000 189.415000 402.345000 189.565000 ;
      RECT  54.545000 189.565000 402.195000 189.715000 ;
      RECT  54.545000 189.715000 402.045000 189.865000 ;
      RECT  54.545000 189.865000 401.895000 190.015000 ;
      RECT  54.545000 190.015000 401.745000 190.165000 ;
      RECT  54.545000 190.165000 401.595000 190.315000 ;
      RECT  54.545000 190.315000 401.445000 190.465000 ;
      RECT  54.545000 190.465000 401.295000 190.615000 ;
      RECT  54.545000 190.615000 401.145000 190.765000 ;
      RECT  54.545000 190.765000 400.995000 190.915000 ;
      RECT  54.545000 190.915000 400.845000 191.065000 ;
      RECT  54.545000 191.065000 400.695000 191.215000 ;
      RECT  54.545000 191.215000 400.545000 191.365000 ;
      RECT  54.545000 191.365000 400.395000 191.515000 ;
      RECT  54.545000 191.515000 400.245000 191.665000 ;
      RECT  54.545000 191.665000 400.095000 191.815000 ;
      RECT  54.545000 191.815000 399.945000 191.965000 ;
      RECT  54.545000 191.965000 399.795000 192.115000 ;
      RECT  54.545000 192.115000 399.645000 192.265000 ;
      RECT  54.545000 192.265000 399.495000 192.415000 ;
      RECT  54.545000 192.415000 399.345000 192.565000 ;
      RECT  54.545000 192.565000 399.195000 192.715000 ;
      RECT  54.545000 192.715000 399.045000 192.865000 ;
      RECT  54.545000 192.865000 398.895000 193.015000 ;
      RECT  54.545000 193.015000 398.745000 193.165000 ;
      RECT  54.545000 193.165000 398.595000 193.315000 ;
      RECT  54.545000 193.315000 398.445000 193.465000 ;
      RECT  54.545000 193.465000 398.295000 193.615000 ;
      RECT  54.545000 193.615000 398.145000 193.765000 ;
      RECT  54.545000 193.765000 397.995000 193.915000 ;
      RECT  54.545000 193.915000 397.845000 194.065000 ;
      RECT  54.545000 194.065000 397.695000 194.215000 ;
      RECT  54.545000 194.215000 397.545000 194.365000 ;
      RECT  54.545000 194.365000 397.395000 194.515000 ;
      RECT  54.545000 194.515000 397.245000 194.665000 ;
      RECT  54.545000 194.665000 397.095000 194.815000 ;
      RECT  54.545000 194.815000 396.945000 194.965000 ;
      RECT  54.545000 194.965000 396.795000 195.115000 ;
      RECT  54.545000 195.115000 396.645000 195.265000 ;
      RECT  54.545000 195.265000 396.495000 195.415000 ;
      RECT  54.545000 195.415000 396.345000 195.565000 ;
      RECT  54.545000 195.565000 396.195000 195.715000 ;
      RECT  54.545000 195.715000 396.045000 195.865000 ;
      RECT  54.545000 195.865000 395.895000 196.015000 ;
      RECT  54.545000 196.015000 395.745000 196.165000 ;
      RECT  54.545000 196.165000 395.595000 196.315000 ;
      RECT  54.545000 196.315000 395.445000 196.465000 ;
      RECT  54.545000 196.465000 395.295000 196.615000 ;
      RECT  54.545000 196.615000 395.145000 196.765000 ;
      RECT  54.545000 196.765000 394.995000 196.915000 ;
      RECT  54.545000 196.915000 394.845000 197.065000 ;
      RECT  54.545000 197.065000 394.695000 197.215000 ;
      RECT  54.545000 197.215000 394.545000 197.365000 ;
      RECT  54.545000 197.365000 394.475000 197.435000 ;
      RECT  54.695000 197.435000 394.325000 197.585000 ;
      RECT  54.845000 197.585000 394.175000 197.735000 ;
      RECT  54.995000 197.735000 394.025000 197.885000 ;
      RECT  55.145000 197.885000 393.875000 198.035000 ;
      RECT  55.295000 198.035000 393.725000 198.185000 ;
      RECT  55.445000 198.185000 393.575000 198.335000 ;
      RECT  55.595000 198.335000 393.425000 198.485000 ;
      RECT  55.745000 198.485000 393.275000 198.635000 ;
      RECT  55.895000 198.635000 393.125000 198.785000 ;
      RECT  56.045000 198.785000 392.975000 198.935000 ;
      RECT  56.195000 198.935000 392.825000 199.085000 ;
      RECT  56.345000 199.085000 392.675000 199.235000 ;
      RECT  56.495000 199.235000 392.525000 199.385000 ;
      RECT  56.645000 199.385000 392.375000 199.535000 ;
      RECT  56.795000 199.535000 392.225000 199.685000 ;
      RECT  56.945000 199.685000 392.075000 199.835000 ;
      RECT  57.095000 199.835000 391.925000 199.985000 ;
      RECT  57.245000 199.985000 391.775000 200.135000 ;
      RECT  57.395000 200.135000 391.625000 200.285000 ;
      RECT  57.545000 200.285000 391.475000 200.435000 ;
      RECT  57.695000 200.435000 391.325000 200.585000 ;
      RECT  57.845000 200.585000 391.175000 200.735000 ;
      RECT  57.995000 200.735000 391.025000 200.885000 ;
      RECT  58.145000 200.885000 390.875000 201.035000 ;
      RECT  58.295000 201.035000 390.725000 201.185000 ;
      RECT  58.445000 201.185000 390.575000 201.335000 ;
      RECT  58.595000 201.335000 390.425000 201.485000 ;
      RECT  58.745000 201.485000 390.275000 201.635000 ;
      RECT  58.895000 201.635000 390.125000 201.785000 ;
      RECT  59.045000 201.785000 389.975000 201.935000 ;
      RECT  59.195000 201.935000 389.825000 202.085000 ;
      RECT  59.345000 202.085000 389.675000 202.235000 ;
      RECT  59.495000 202.235000 389.525000 202.385000 ;
      RECT  59.645000 202.385000 389.375000 202.535000 ;
      RECT  59.795000 202.535000 389.225000 202.685000 ;
      RECT  59.945000 202.685000 389.075000 202.835000 ;
      RECT  60.095000 202.835000 388.925000 202.985000 ;
      RECT  60.245000 202.985000 388.775000 203.135000 ;
      RECT  60.395000 203.135000 388.625000 203.285000 ;
      RECT  60.545000 203.285000 388.475000 203.435000 ;
      RECT  60.695000 203.435000 388.325000 203.585000 ;
      RECT  60.845000 203.585000 388.175000 203.735000 ;
      RECT  60.995000 203.735000 388.025000 203.885000 ;
      RECT  61.145000 203.885000 387.875000 204.035000 ;
      RECT  61.215000 204.035000 387.805000 204.105000 ;
      RECT 398.700000 229.050000 480.000000 229.100000 ;
      RECT 398.700000 229.050000 480.000000 229.100000 ;
      RECT 398.850000 228.900000 480.000000 229.050000 ;
      RECT 398.850000 228.900000 480.000000 229.050000 ;
      RECT 399.000000 228.750000 480.000000 228.900000 ;
      RECT 399.000000 228.750000 480.000000 228.900000 ;
      RECT 399.150000 228.600000 480.000000 228.750000 ;
      RECT 399.150000 228.600000 480.000000 228.750000 ;
      RECT 399.300000 228.450000 480.000000 228.600000 ;
      RECT 399.300000 228.450000 480.000000 228.600000 ;
      RECT 399.450000 228.300000 480.000000 228.450000 ;
      RECT 399.450000 228.300000 480.000000 228.450000 ;
      RECT 399.585000 228.165000 480.000000 228.300000 ;
      RECT 399.600000 228.150000 480.000000 228.300000 ;
      RECT 399.600000 228.150000 480.000000 228.300000 ;
      RECT 399.735000 228.015000 480.000000 228.165000 ;
      RECT 399.750000 228.000000 480.000000 228.150000 ;
      RECT 399.750000 228.000000 480.000000 228.150000 ;
      RECT 399.885000 227.865000 480.000000 228.015000 ;
      RECT 399.900000 227.850000 480.000000 228.000000 ;
      RECT 399.900000 227.850000 480.000000 228.000000 ;
      RECT 400.035000 227.715000 480.000000 227.865000 ;
      RECT 400.050000 227.700000 480.000000 227.850000 ;
      RECT 400.050000 227.700000 480.000000 227.850000 ;
      RECT 400.185000 227.565000 480.000000 227.715000 ;
      RECT 400.200000 227.550000 480.000000 227.700000 ;
      RECT 400.200000 227.550000 480.000000 227.700000 ;
      RECT 400.335000 227.415000 480.000000 227.565000 ;
      RECT 400.350000 227.400000 480.000000 227.550000 ;
      RECT 400.350000 227.400000 480.000000 227.550000 ;
      RECT 400.485000 227.265000 480.000000 227.415000 ;
      RECT 400.500000 227.250000 480.000000 227.400000 ;
      RECT 400.500000 227.250000 480.000000 227.400000 ;
      RECT 400.635000 227.115000 480.000000 227.265000 ;
      RECT 400.650000 227.100000 480.000000 227.250000 ;
      RECT 400.650000 227.100000 480.000000 227.250000 ;
      RECT 400.785000 226.965000 480.000000 227.115000 ;
      RECT 400.800000 226.950000 480.000000 227.100000 ;
      RECT 400.800000 226.950000 480.000000 227.100000 ;
      RECT 400.935000 226.815000 480.000000 226.965000 ;
      RECT 400.950000 226.800000 480.000000 226.950000 ;
      RECT 400.950000 226.800000 480.000000 226.950000 ;
      RECT 401.085000 226.665000 480.000000 226.815000 ;
      RECT 401.100000 226.650000 480.000000 226.800000 ;
      RECT 401.100000 226.650000 480.000000 226.800000 ;
      RECT 401.235000 226.515000 480.000000 226.665000 ;
      RECT 401.250000 226.500000 480.000000 226.650000 ;
      RECT 401.250000 226.500000 480.000000 226.650000 ;
      RECT 401.385000 226.365000 480.000000 226.515000 ;
      RECT 401.400000 226.350000 480.000000 226.500000 ;
      RECT 401.400000 226.350000 480.000000 226.500000 ;
      RECT 401.535000 226.215000 480.000000 226.365000 ;
      RECT 401.550000 226.200000 480.000000 226.350000 ;
      RECT 401.550000 226.200000 480.000000 226.350000 ;
      RECT 401.685000 226.065000 480.000000 226.215000 ;
      RECT 401.700000 226.050000 480.000000 226.200000 ;
      RECT 401.700000 226.050000 480.000000 226.200000 ;
      RECT 401.835000 225.915000 480.000000 226.065000 ;
      RECT 401.850000 225.900000 480.000000 226.050000 ;
      RECT 401.850000 225.900000 480.000000 226.050000 ;
      RECT 401.985000 225.765000 480.000000 225.915000 ;
      RECT 402.000000 225.750000 480.000000 225.900000 ;
      RECT 402.000000 225.750000 480.000000 225.900000 ;
      RECT 402.135000 225.615000 480.000000 225.765000 ;
      RECT 402.150000 225.600000 480.000000 225.750000 ;
      RECT 402.150000 225.600000 480.000000 225.750000 ;
      RECT 402.285000 225.465000 480.000000 225.615000 ;
      RECT 402.300000 225.450000 480.000000 225.600000 ;
      RECT 402.300000 225.450000 480.000000 225.600000 ;
      RECT 402.435000 225.315000 480.000000 225.465000 ;
      RECT 402.450000 225.300000 480.000000 225.450000 ;
      RECT 402.450000 225.300000 480.000000 225.450000 ;
      RECT 402.585000 225.165000 480.000000 225.315000 ;
      RECT 402.600000 225.150000 480.000000 225.300000 ;
      RECT 402.600000 225.150000 480.000000 225.300000 ;
      RECT 402.735000 225.015000 480.000000 225.165000 ;
      RECT 402.750000 225.000000 480.000000 225.150000 ;
      RECT 402.750000 225.000000 480.000000 225.150000 ;
      RECT 402.885000 224.865000 480.000000 225.015000 ;
      RECT 402.900000 224.850000 480.000000 225.000000 ;
      RECT 402.900000 224.850000 480.000000 225.000000 ;
      RECT 403.035000 224.715000 480.000000 224.865000 ;
      RECT 403.050000 224.700000 480.000000 224.850000 ;
      RECT 403.050000 224.700000 480.000000 224.850000 ;
      RECT 403.185000 224.565000 480.000000 224.715000 ;
      RECT 403.200000 224.550000 480.000000 224.700000 ;
      RECT 403.200000 224.550000 480.000000 224.700000 ;
      RECT 403.335000 224.415000 480.000000 224.565000 ;
      RECT 403.350000 224.400000 480.000000 224.550000 ;
      RECT 403.350000 224.400000 480.000000 224.550000 ;
      RECT 403.485000 224.265000 480.000000 224.415000 ;
      RECT 403.500000 224.250000 480.000000 224.400000 ;
      RECT 403.500000 224.250000 480.000000 224.400000 ;
      RECT 403.635000 224.115000 480.000000 224.265000 ;
      RECT 403.650000 224.100000 480.000000 224.250000 ;
      RECT 403.650000 224.100000 480.000000 224.250000 ;
      RECT 403.785000 223.965000 480.000000 224.115000 ;
      RECT 403.800000 223.950000 480.000000 224.100000 ;
      RECT 403.800000 223.950000 480.000000 224.100000 ;
      RECT 403.935000 223.815000 480.000000 223.965000 ;
      RECT 403.950000 223.800000 480.000000 223.950000 ;
      RECT 403.950000 223.800000 480.000000 223.950000 ;
      RECT 404.085000 223.665000 480.000000 223.815000 ;
      RECT 404.100000 223.650000 480.000000 223.800000 ;
      RECT 404.100000 223.650000 480.000000 223.800000 ;
      RECT 404.235000 223.515000 480.000000 223.665000 ;
      RECT 404.250000 223.500000 480.000000 223.650000 ;
      RECT 404.250000 223.500000 480.000000 223.650000 ;
      RECT 404.385000 223.365000 480.000000 223.515000 ;
      RECT 404.400000 223.350000 480.000000 223.500000 ;
      RECT 404.400000 223.350000 480.000000 223.500000 ;
      RECT 404.535000 223.215000 480.000000 223.365000 ;
      RECT 404.550000 223.200000 480.000000 223.350000 ;
      RECT 404.550000 223.200000 480.000000 223.350000 ;
      RECT 404.685000 223.065000 480.000000 223.215000 ;
      RECT 404.700000 223.050000 480.000000 223.200000 ;
      RECT 404.700000 223.050000 480.000000 223.200000 ;
      RECT 404.835000 222.915000 480.000000 223.065000 ;
      RECT 404.850000 222.900000 480.000000 223.050000 ;
      RECT 404.850000 222.900000 480.000000 223.050000 ;
      RECT 404.985000 222.765000 480.000000 222.915000 ;
      RECT 405.000000 222.750000 480.000000 222.900000 ;
      RECT 405.000000 222.750000 480.000000 222.900000 ;
      RECT 405.135000 222.615000 480.000000 222.765000 ;
      RECT 405.150000 222.600000 480.000000 222.750000 ;
      RECT 405.150000 222.600000 480.000000 222.750000 ;
      RECT 405.285000 222.465000 480.000000 222.615000 ;
      RECT 405.300000 222.450000 480.000000 222.600000 ;
      RECT 405.300000 222.450000 480.000000 222.600000 ;
      RECT 405.435000 222.315000 480.000000 222.465000 ;
      RECT 405.450000 222.300000 480.000000 222.450000 ;
      RECT 405.450000 222.300000 480.000000 222.450000 ;
      RECT 405.585000 222.165000 480.000000 222.315000 ;
      RECT 405.600000 222.150000 480.000000 222.300000 ;
      RECT 405.600000 222.150000 480.000000 222.300000 ;
      RECT 405.735000 222.015000 480.000000 222.165000 ;
      RECT 405.750000 222.000000 480.000000 222.150000 ;
      RECT 405.750000 222.000000 480.000000 222.150000 ;
      RECT 405.885000 221.865000 480.000000 222.015000 ;
      RECT 405.900000 221.850000 480.000000 222.000000 ;
      RECT 405.900000 221.850000 480.000000 222.000000 ;
      RECT 406.035000 221.715000 480.000000 221.865000 ;
      RECT 406.050000 221.700000 480.000000 221.850000 ;
      RECT 406.050000 221.700000 480.000000 221.850000 ;
      RECT 406.185000 221.565000 480.000000 221.715000 ;
      RECT 406.200000 221.550000 480.000000 221.700000 ;
      RECT 406.200000 221.550000 480.000000 221.700000 ;
      RECT 406.335000 221.415000 480.000000 221.565000 ;
      RECT 406.350000 221.400000 480.000000 221.550000 ;
      RECT 406.350000 221.400000 480.000000 221.550000 ;
      RECT 406.485000 221.265000 480.000000 221.415000 ;
      RECT 406.500000 221.250000 480.000000 221.400000 ;
      RECT 406.500000 221.250000 480.000000 221.400000 ;
      RECT 406.635000 221.115000 480.000000 221.265000 ;
      RECT 406.650000 221.100000 480.000000 221.250000 ;
      RECT 406.650000 221.100000 480.000000 221.250000 ;
      RECT 406.785000 220.965000 480.000000 221.115000 ;
      RECT 406.800000 220.950000 480.000000 221.100000 ;
      RECT 406.800000 220.950000 480.000000 221.100000 ;
      RECT 406.935000 220.815000 480.000000 220.965000 ;
      RECT 406.950000 220.800000 480.000000 220.950000 ;
      RECT 406.950000 220.800000 480.000000 220.950000 ;
      RECT 407.085000 220.665000 480.000000 220.815000 ;
      RECT 407.100000 220.650000 480.000000 220.800000 ;
      RECT 407.100000 220.650000 480.000000 220.800000 ;
      RECT 407.235000 220.515000 480.000000 220.665000 ;
      RECT 407.250000 220.500000 480.000000 220.650000 ;
      RECT 407.250000 220.500000 480.000000 220.650000 ;
      RECT 407.385000 220.365000 480.000000 220.515000 ;
      RECT 407.400000 220.350000 480.000000 220.500000 ;
      RECT 407.400000 220.350000 480.000000 220.500000 ;
      RECT 407.535000 220.215000 480.000000 220.365000 ;
      RECT 407.550000 220.200000 480.000000 220.350000 ;
      RECT 407.550000 220.200000 480.000000 220.350000 ;
      RECT 407.685000 220.065000 480.000000 220.215000 ;
      RECT 407.700000 220.050000 480.000000 220.200000 ;
      RECT 407.700000 220.050000 480.000000 220.200000 ;
      RECT 407.835000 219.915000 480.000000 220.065000 ;
      RECT 407.850000 219.900000 480.000000 220.050000 ;
      RECT 407.850000 219.900000 480.000000 220.050000 ;
      RECT 407.985000 219.765000 480.000000 219.915000 ;
      RECT 408.000000 219.750000 480.000000 219.900000 ;
      RECT 408.000000 219.750000 480.000000 219.900000 ;
      RECT 408.135000 219.615000 480.000000 219.765000 ;
      RECT 408.150000 219.600000 480.000000 219.750000 ;
      RECT 408.150000 219.600000 480.000000 219.750000 ;
      RECT 408.285000 219.465000 480.000000 219.615000 ;
      RECT 408.300000 219.450000 480.000000 219.600000 ;
      RECT 408.300000 219.450000 480.000000 219.600000 ;
      RECT 408.435000 219.315000 480.000000 219.465000 ;
      RECT 408.450000 219.300000 480.000000 219.450000 ;
      RECT 408.450000 219.300000 480.000000 219.450000 ;
      RECT 408.585000 219.165000 480.000000 219.315000 ;
      RECT 408.600000 219.150000 480.000000 219.300000 ;
      RECT 408.600000 219.150000 480.000000 219.300000 ;
      RECT 408.735000 219.015000 480.000000 219.165000 ;
      RECT 408.750000 219.000000 480.000000 219.150000 ;
      RECT 408.750000 219.000000 480.000000 219.150000 ;
      RECT 408.885000 218.865000 480.000000 219.015000 ;
      RECT 408.900000 218.850000 480.000000 219.000000 ;
      RECT 408.900000 218.850000 480.000000 219.000000 ;
      RECT 409.035000 218.715000 480.000000 218.865000 ;
      RECT 409.050000 218.700000 480.000000 218.850000 ;
      RECT 409.050000 218.700000 480.000000 218.850000 ;
      RECT 409.185000 218.565000 480.000000 218.715000 ;
      RECT 409.200000 218.550000 480.000000 218.700000 ;
      RECT 409.200000 218.550000 480.000000 218.700000 ;
      RECT 409.335000 218.415000 480.000000 218.565000 ;
      RECT 409.350000 218.400000 480.000000 218.550000 ;
      RECT 409.350000 218.400000 480.000000 218.550000 ;
      RECT 409.485000 218.265000 480.000000 218.415000 ;
      RECT 409.500000 218.250000 480.000000 218.400000 ;
      RECT 409.500000 218.250000 480.000000 218.400000 ;
      RECT 409.635000 218.115000 480.000000 218.265000 ;
      RECT 409.650000 218.100000 480.000000 218.250000 ;
      RECT 409.650000 218.100000 480.000000 218.250000 ;
      RECT 409.785000 217.965000 480.000000 218.115000 ;
      RECT 409.800000 217.950000 480.000000 218.100000 ;
      RECT 409.800000 217.950000 480.000000 218.100000 ;
      RECT 409.935000 217.815000 480.000000 217.965000 ;
      RECT 409.950000 217.800000 480.000000 217.950000 ;
      RECT 409.950000 217.800000 480.000000 217.950000 ;
      RECT 410.085000 217.665000 480.000000 217.815000 ;
      RECT 410.100000 217.650000 480.000000 217.800000 ;
      RECT 410.100000 217.650000 480.000000 217.800000 ;
      RECT 410.235000 217.515000 480.000000 217.665000 ;
      RECT 410.250000 217.500000 480.000000 217.650000 ;
      RECT 410.250000 217.500000 480.000000 217.650000 ;
      RECT 410.385000 217.365000 480.000000 217.515000 ;
      RECT 410.400000 217.350000 480.000000 217.500000 ;
      RECT 410.400000 217.350000 480.000000 217.500000 ;
      RECT 410.535000 217.215000 480.000000 217.365000 ;
      RECT 410.550000 217.200000 480.000000 217.350000 ;
      RECT 410.550000 217.200000 480.000000 217.350000 ;
      RECT 410.685000 217.065000 480.000000 217.215000 ;
      RECT 410.700000 217.050000 480.000000 217.200000 ;
      RECT 410.700000 217.050000 480.000000 217.200000 ;
      RECT 410.835000 216.915000 480.000000 217.065000 ;
      RECT 410.850000 216.900000 480.000000 217.050000 ;
      RECT 410.850000 216.900000 480.000000 217.050000 ;
      RECT 410.985000 216.765000 480.000000 216.915000 ;
      RECT 411.000000 216.750000 480.000000 216.900000 ;
      RECT 411.000000 216.750000 480.000000 216.900000 ;
      RECT 411.135000 216.615000 480.000000 216.765000 ;
      RECT 411.150000 216.600000 480.000000 216.750000 ;
      RECT 411.150000 216.600000 480.000000 216.750000 ;
      RECT 411.285000 216.465000 480.000000 216.615000 ;
      RECT 411.300000 216.450000 480.000000 216.600000 ;
      RECT 411.300000 216.450000 480.000000 216.600000 ;
      RECT 411.435000 216.315000 480.000000 216.465000 ;
      RECT 411.450000 216.300000 480.000000 216.450000 ;
      RECT 411.450000 216.300000 480.000000 216.450000 ;
      RECT 411.585000 216.165000 480.000000 216.315000 ;
      RECT 411.600000 216.150000 480.000000 216.300000 ;
      RECT 411.600000 216.150000 480.000000 216.300000 ;
      RECT 411.735000 216.015000 480.000000 216.165000 ;
      RECT 411.750000 216.000000 480.000000 216.150000 ;
      RECT 411.750000 216.000000 480.000000 216.150000 ;
      RECT 411.885000 215.865000 480.000000 216.015000 ;
      RECT 411.900000 215.850000 480.000000 216.000000 ;
      RECT 411.900000 215.850000 480.000000 216.000000 ;
      RECT 412.035000 215.715000 480.000000 215.865000 ;
      RECT 412.050000 215.700000 480.000000 215.850000 ;
      RECT 412.050000 215.700000 480.000000 215.850000 ;
      RECT 412.185000 215.565000 480.000000 215.715000 ;
      RECT 412.200000 215.550000 480.000000 215.700000 ;
      RECT 412.200000 215.550000 480.000000 215.700000 ;
      RECT 412.335000 215.415000 480.000000 215.565000 ;
      RECT 412.350000 215.400000 480.000000 215.550000 ;
      RECT 412.350000 215.400000 480.000000 215.550000 ;
      RECT 412.485000 215.265000 480.000000 215.415000 ;
      RECT 412.500000 215.250000 480.000000 215.400000 ;
      RECT 412.500000 215.250000 480.000000 215.400000 ;
      RECT 412.635000 215.115000 480.000000 215.265000 ;
      RECT 412.650000 215.100000 480.000000 215.250000 ;
      RECT 412.650000 215.100000 480.000000 215.250000 ;
      RECT 412.785000 214.965000 480.000000 215.115000 ;
      RECT 412.800000 214.950000 480.000000 215.100000 ;
      RECT 412.800000 214.950000 480.000000 215.100000 ;
      RECT 412.935000 214.815000 480.000000 214.965000 ;
      RECT 412.950000 214.800000 480.000000 214.950000 ;
      RECT 412.950000 214.800000 480.000000 214.950000 ;
      RECT 413.085000 214.665000 480.000000 214.815000 ;
      RECT 413.100000 214.650000 480.000000 214.800000 ;
      RECT 413.100000 214.650000 480.000000 214.800000 ;
      RECT 413.235000 214.515000 480.000000 214.665000 ;
      RECT 413.250000 214.500000 480.000000 214.650000 ;
      RECT 413.250000 214.500000 480.000000 214.650000 ;
      RECT 413.385000 214.365000 480.000000 214.515000 ;
      RECT 413.400000 214.350000 480.000000 214.500000 ;
      RECT 413.400000 214.350000 480.000000 214.500000 ;
      RECT 413.535000 214.215000 480.000000 214.365000 ;
      RECT 413.550000 214.200000 480.000000 214.350000 ;
      RECT 413.550000 214.200000 480.000000 214.350000 ;
      RECT 413.685000 214.065000 480.000000 214.215000 ;
      RECT 413.700000 214.050000 480.000000 214.200000 ;
      RECT 413.700000 214.050000 480.000000 214.200000 ;
      RECT 413.835000 213.915000 480.000000 214.065000 ;
      RECT 413.850000 213.900000 480.000000 214.050000 ;
      RECT 413.850000 213.900000 480.000000 214.050000 ;
      RECT 413.985000 213.765000 480.000000 213.915000 ;
      RECT 414.000000 213.750000 480.000000 213.900000 ;
      RECT 414.000000 213.750000 480.000000 213.900000 ;
      RECT 414.135000 213.615000 480.000000 213.765000 ;
      RECT 414.150000 213.600000 480.000000 213.750000 ;
      RECT 414.150000 213.600000 480.000000 213.750000 ;
      RECT 414.285000 213.465000 480.000000 213.615000 ;
      RECT 414.300000 213.450000 480.000000 213.600000 ;
      RECT 414.300000 213.450000 480.000000 213.600000 ;
      RECT 414.435000 213.315000 480.000000 213.465000 ;
      RECT 414.450000 213.300000 480.000000 213.450000 ;
      RECT 414.450000 213.300000 480.000000 213.450000 ;
      RECT 414.585000 213.165000 480.000000 213.315000 ;
      RECT 414.600000 213.150000 480.000000 213.300000 ;
      RECT 414.600000 213.150000 480.000000 213.300000 ;
      RECT 414.735000 213.015000 480.000000 213.165000 ;
      RECT 414.750000 213.000000 480.000000 213.150000 ;
      RECT 414.750000 213.000000 480.000000 213.150000 ;
      RECT 414.885000 212.865000 480.000000 213.015000 ;
      RECT 414.900000 212.850000 480.000000 213.000000 ;
      RECT 414.900000 212.850000 480.000000 213.000000 ;
      RECT 415.035000 212.715000 480.000000 212.865000 ;
      RECT 415.050000 212.700000 480.000000 212.850000 ;
      RECT 415.050000 212.700000 480.000000 212.850000 ;
      RECT 415.185000 212.565000 480.000000 212.715000 ;
      RECT 415.200000 212.550000 480.000000 212.700000 ;
      RECT 415.200000 212.550000 480.000000 212.700000 ;
      RECT 415.335000 212.415000 480.000000 212.565000 ;
      RECT 415.350000 212.400000 480.000000 212.550000 ;
      RECT 415.350000 212.400000 480.000000 212.550000 ;
      RECT 415.485000 212.265000 480.000000 212.415000 ;
      RECT 415.500000 212.250000 480.000000 212.400000 ;
      RECT 415.500000 212.250000 480.000000 212.400000 ;
      RECT 415.635000 212.115000 480.000000 212.265000 ;
      RECT 415.650000 212.100000 480.000000 212.250000 ;
      RECT 415.650000 212.100000 480.000000 212.250000 ;
      RECT 415.785000 211.965000 480.000000 212.115000 ;
      RECT 415.800000 211.950000 480.000000 212.100000 ;
      RECT 415.800000 211.950000 480.000000 212.100000 ;
      RECT 415.935000 211.815000 480.000000 211.965000 ;
      RECT 415.950000 211.800000 480.000000 211.950000 ;
      RECT 415.950000 211.800000 480.000000 211.950000 ;
      RECT 416.085000 211.665000 480.000000 211.815000 ;
      RECT 416.100000 211.650000 480.000000 211.800000 ;
      RECT 416.100000 211.650000 480.000000 211.800000 ;
      RECT 416.235000 211.515000 480.000000 211.665000 ;
      RECT 416.250000 211.500000 480.000000 211.650000 ;
      RECT 416.250000 211.500000 480.000000 211.650000 ;
      RECT 416.385000 211.365000 480.000000 211.515000 ;
      RECT 416.400000 211.350000 480.000000 211.500000 ;
      RECT 416.400000 211.350000 480.000000 211.500000 ;
      RECT 416.535000 211.215000 480.000000 211.365000 ;
      RECT 416.550000 211.200000 480.000000 211.350000 ;
      RECT 416.550000 211.200000 480.000000 211.350000 ;
      RECT 416.685000 211.065000 480.000000 211.215000 ;
      RECT 416.700000 211.050000 480.000000 211.200000 ;
      RECT 416.700000 211.050000 480.000000 211.200000 ;
      RECT 416.835000 210.915000 480.000000 211.065000 ;
      RECT 416.850000 210.900000 480.000000 211.050000 ;
      RECT 416.850000 210.900000 480.000000 211.050000 ;
      RECT 416.985000 210.765000 480.000000 210.915000 ;
      RECT 417.000000 210.750000 480.000000 210.900000 ;
      RECT 417.000000 210.750000 480.000000 210.900000 ;
      RECT 417.135000 210.615000 480.000000 210.765000 ;
      RECT 417.150000 210.600000 480.000000 210.750000 ;
      RECT 417.150000 210.600000 480.000000 210.750000 ;
      RECT 417.285000 210.465000 480.000000 210.615000 ;
      RECT 417.300000 210.450000 480.000000 210.600000 ;
      RECT 417.300000 210.450000 480.000000 210.600000 ;
      RECT 417.435000 210.315000 480.000000 210.465000 ;
      RECT 417.450000 210.300000 480.000000 210.450000 ;
      RECT 417.450000 210.300000 480.000000 210.450000 ;
      RECT 417.585000 210.165000 480.000000 210.315000 ;
      RECT 417.600000 210.150000 480.000000 210.300000 ;
      RECT 417.600000 210.150000 480.000000 210.300000 ;
      RECT 417.735000 210.015000 480.000000 210.165000 ;
      RECT 417.750000 210.000000 480.000000 210.150000 ;
      RECT 417.750000 210.000000 480.000000 210.150000 ;
      RECT 417.885000 209.865000 480.000000 210.015000 ;
      RECT 417.900000 209.850000 480.000000 210.000000 ;
      RECT 417.900000 209.850000 480.000000 210.000000 ;
      RECT 418.035000 209.715000 480.000000 209.865000 ;
      RECT 418.050000 209.700000 480.000000 209.850000 ;
      RECT 418.050000 209.700000 480.000000 209.850000 ;
      RECT 418.185000 209.565000 480.000000 209.715000 ;
      RECT 418.200000 209.550000 480.000000 209.700000 ;
      RECT 418.200000 209.550000 480.000000 209.700000 ;
      RECT 418.335000 209.415000 480.000000 209.565000 ;
      RECT 418.350000 209.400000 480.000000 209.550000 ;
      RECT 418.350000 209.400000 480.000000 209.550000 ;
      RECT 418.485000 209.265000 480.000000 209.415000 ;
      RECT 418.500000 209.250000 480.000000 209.400000 ;
      RECT 418.500000 209.250000 480.000000 209.400000 ;
      RECT 418.635000 209.115000 480.000000 209.265000 ;
      RECT 418.650000 209.100000 480.000000 209.250000 ;
      RECT 418.650000 209.100000 480.000000 209.250000 ;
      RECT 418.785000 208.965000 480.000000 209.115000 ;
      RECT 418.800000 208.950000 480.000000 209.100000 ;
      RECT 418.800000 208.950000 480.000000 209.100000 ;
      RECT 418.935000 208.815000 480.000000 208.965000 ;
      RECT 418.950000 208.800000 480.000000 208.950000 ;
      RECT 418.950000 208.800000 480.000000 208.950000 ;
      RECT 419.085000 208.665000 480.000000 208.815000 ;
      RECT 419.100000 208.650000 480.000000 208.800000 ;
      RECT 419.100000 208.650000 480.000000 208.800000 ;
      RECT 419.235000 208.515000 480.000000 208.665000 ;
      RECT 419.250000 208.500000 480.000000 208.650000 ;
      RECT 419.250000 208.500000 480.000000 208.650000 ;
      RECT 419.385000 208.365000 480.000000 208.515000 ;
      RECT 419.400000 208.350000 480.000000 208.500000 ;
      RECT 419.400000 208.350000 480.000000 208.500000 ;
      RECT 419.535000 208.215000 480.000000 208.365000 ;
      RECT 419.550000 208.200000 480.000000 208.350000 ;
      RECT 419.550000 208.200000 480.000000 208.350000 ;
      RECT 419.685000 208.065000 480.000000 208.215000 ;
      RECT 419.700000 208.050000 480.000000 208.200000 ;
      RECT 419.700000 208.050000 480.000000 208.200000 ;
      RECT 419.835000 207.915000 480.000000 208.065000 ;
      RECT 419.850000 207.900000 480.000000 208.050000 ;
      RECT 419.850000 207.900000 480.000000 208.050000 ;
      RECT 419.985000 207.765000 480.000000 207.915000 ;
      RECT 420.000000 207.750000 480.000000 207.900000 ;
      RECT 420.000000 207.750000 480.000000 207.900000 ;
      RECT 420.135000 207.615000 480.000000 207.765000 ;
      RECT 420.150000 207.600000 480.000000 207.750000 ;
      RECT 420.150000 207.600000 480.000000 207.750000 ;
      RECT 420.285000 207.465000 480.000000 207.615000 ;
      RECT 420.300000 207.450000 480.000000 207.600000 ;
      RECT 420.300000 207.450000 480.000000 207.600000 ;
      RECT 420.435000 207.315000 480.000000 207.465000 ;
      RECT 420.450000 207.300000 480.000000 207.450000 ;
      RECT 420.450000 207.300000 480.000000 207.450000 ;
      RECT 420.585000 207.165000 480.000000 207.315000 ;
      RECT 420.600000 207.150000 480.000000 207.300000 ;
      RECT 420.600000 207.150000 480.000000 207.300000 ;
      RECT 420.735000 207.015000 480.000000 207.165000 ;
      RECT 420.750000 207.000000 480.000000 207.150000 ;
      RECT 420.750000 207.000000 480.000000 207.150000 ;
      RECT 420.885000 206.865000 480.000000 207.015000 ;
      RECT 420.900000 206.850000 480.000000 207.000000 ;
      RECT 420.900000 206.850000 480.000000 207.000000 ;
      RECT 421.035000 206.715000 480.000000 206.865000 ;
      RECT 421.050000 206.700000 480.000000 206.850000 ;
      RECT 421.050000 206.700000 480.000000 206.850000 ;
      RECT 421.185000 206.565000 480.000000 206.715000 ;
      RECT 421.200000 206.550000 480.000000 206.700000 ;
      RECT 421.200000 206.550000 480.000000 206.700000 ;
      RECT 421.335000 206.415000 480.000000 206.565000 ;
      RECT 421.350000 206.400000 480.000000 206.550000 ;
      RECT 421.350000 206.400000 480.000000 206.550000 ;
      RECT 421.485000 206.265000 480.000000 206.415000 ;
      RECT 421.500000 206.250000 480.000000 206.400000 ;
      RECT 421.500000 206.250000 480.000000 206.400000 ;
      RECT 421.635000 206.115000 480.000000 206.265000 ;
      RECT 421.650000 206.100000 480.000000 206.250000 ;
      RECT 421.650000 206.100000 480.000000 206.250000 ;
      RECT 421.785000 205.965000 480.000000 206.115000 ;
      RECT 421.800000 205.950000 480.000000 206.100000 ;
      RECT 421.800000 205.950000 480.000000 206.100000 ;
      RECT 421.935000 205.815000 480.000000 205.965000 ;
      RECT 421.950000 205.800000 480.000000 205.950000 ;
      RECT 421.950000 205.800000 480.000000 205.950000 ;
      RECT 422.085000 205.665000 480.000000 205.815000 ;
      RECT 422.100000 205.650000 480.000000 205.800000 ;
      RECT 422.100000 205.650000 480.000000 205.800000 ;
      RECT 422.235000 205.515000 480.000000 205.665000 ;
      RECT 422.250000 205.500000 480.000000 205.650000 ;
      RECT 422.250000 205.500000 480.000000 205.650000 ;
      RECT 422.385000 205.365000 480.000000 205.515000 ;
      RECT 422.400000 205.350000 480.000000 205.500000 ;
      RECT 422.400000 205.350000 480.000000 205.500000 ;
      RECT 422.535000 205.215000 480.000000 205.365000 ;
      RECT 422.550000 205.200000 480.000000 205.350000 ;
      RECT 422.550000 205.200000 480.000000 205.350000 ;
      RECT 422.685000 205.065000 480.000000 205.215000 ;
      RECT 422.700000 205.050000 480.000000 205.200000 ;
      RECT 422.700000 205.050000 480.000000 205.200000 ;
      RECT 422.835000 204.915000 480.000000 205.065000 ;
      RECT 422.850000 204.900000 480.000000 205.050000 ;
      RECT 422.850000 204.900000 480.000000 205.050000 ;
      RECT 422.985000 204.765000 480.000000 204.915000 ;
      RECT 423.000000 204.750000 480.000000 204.900000 ;
      RECT 423.000000 204.750000 480.000000 204.900000 ;
      RECT 423.135000 204.615000 480.000000 204.765000 ;
      RECT 423.150000 204.600000 480.000000 204.750000 ;
      RECT 423.150000 204.600000 480.000000 204.750000 ;
      RECT 423.285000 204.465000 480.000000 204.615000 ;
      RECT 423.300000 204.450000 480.000000 204.600000 ;
      RECT 423.300000 204.450000 480.000000 204.600000 ;
      RECT 423.435000 204.315000 480.000000 204.465000 ;
      RECT 423.450000 204.300000 480.000000 204.450000 ;
      RECT 423.450000 204.300000 480.000000 204.450000 ;
      RECT 423.585000 204.165000 480.000000 204.315000 ;
      RECT 423.600000 204.150000 480.000000 204.300000 ;
      RECT 423.600000 204.150000 480.000000 204.300000 ;
      RECT 423.735000 204.015000 480.000000 204.165000 ;
      RECT 423.750000 204.000000 480.000000 204.150000 ;
      RECT 423.750000 204.000000 480.000000 204.150000 ;
      RECT 423.885000 203.865000 480.000000 204.015000 ;
      RECT 423.900000 203.850000 480.000000 204.000000 ;
      RECT 423.900000 203.850000 480.000000 204.000000 ;
      RECT 424.035000 203.715000 480.000000 203.865000 ;
      RECT 424.050000 203.700000 480.000000 203.850000 ;
      RECT 424.050000 203.700000 480.000000 203.850000 ;
      RECT 424.185000 203.565000 480.000000 203.715000 ;
      RECT 424.200000 203.550000 480.000000 203.700000 ;
      RECT 424.200000 203.550000 480.000000 203.700000 ;
      RECT 424.335000 203.415000 480.000000 203.565000 ;
      RECT 424.350000 203.400000 480.000000 203.550000 ;
      RECT 424.350000 203.400000 480.000000 203.550000 ;
      RECT 424.485000 203.265000 480.000000 203.415000 ;
      RECT 424.500000 203.250000 480.000000 203.400000 ;
      RECT 424.500000 203.250000 480.000000 203.400000 ;
      RECT 424.635000 203.115000 480.000000 203.265000 ;
      RECT 424.650000 203.100000 480.000000 203.250000 ;
      RECT 424.650000 203.100000 480.000000 203.250000 ;
      RECT 424.785000 202.965000 480.000000 203.115000 ;
      RECT 424.800000 202.950000 480.000000 203.100000 ;
      RECT 424.800000 202.950000 480.000000 203.100000 ;
      RECT 424.935000 202.815000 480.000000 202.965000 ;
      RECT 424.950000 202.800000 480.000000 202.950000 ;
      RECT 424.950000 202.800000 480.000000 202.950000 ;
      RECT 425.085000 202.665000 480.000000 202.815000 ;
      RECT 425.100000 202.650000 480.000000 202.800000 ;
      RECT 425.100000 202.650000 480.000000 202.800000 ;
      RECT 425.235000 202.515000 480.000000 202.665000 ;
      RECT 425.250000 202.500000 480.000000 202.650000 ;
      RECT 425.250000 202.500000 480.000000 202.650000 ;
      RECT 425.385000 202.365000 480.000000 202.515000 ;
      RECT 425.400000 202.350000 480.000000 202.500000 ;
      RECT 425.400000 202.350000 480.000000 202.500000 ;
      RECT 425.535000 202.215000 480.000000 202.365000 ;
      RECT 425.550000 202.200000 480.000000 202.350000 ;
      RECT 425.550000 202.200000 480.000000 202.350000 ;
      RECT 425.685000 202.065000 480.000000 202.215000 ;
      RECT 425.700000 202.050000 480.000000 202.200000 ;
      RECT 425.700000 202.050000 480.000000 202.200000 ;
      RECT 425.835000 201.915000 480.000000 202.065000 ;
      RECT 425.850000 201.900000 480.000000 202.050000 ;
      RECT 425.850000 201.900000 480.000000 202.050000 ;
      RECT 425.985000 201.765000 480.000000 201.915000 ;
      RECT 426.000000 201.750000 480.000000 201.900000 ;
      RECT 426.000000 201.750000 480.000000 201.900000 ;
      RECT 426.135000 201.615000 480.000000 201.765000 ;
      RECT 426.150000 201.600000 480.000000 201.750000 ;
      RECT 426.150000 201.600000 480.000000 201.750000 ;
      RECT 426.285000 201.465000 480.000000 201.615000 ;
      RECT 426.300000 201.450000 480.000000 201.600000 ;
      RECT 426.300000 201.450000 480.000000 201.600000 ;
      RECT 426.435000 201.315000 480.000000 201.465000 ;
      RECT 426.450000 201.300000 480.000000 201.450000 ;
      RECT 426.450000 201.300000 480.000000 201.450000 ;
      RECT 426.585000 201.165000 480.000000 201.315000 ;
      RECT 426.600000 201.150000 480.000000 201.300000 ;
      RECT 426.600000 201.150000 480.000000 201.300000 ;
      RECT 426.735000 201.015000 480.000000 201.165000 ;
      RECT 426.750000 201.000000 480.000000 201.150000 ;
      RECT 426.750000 201.000000 480.000000 201.150000 ;
      RECT 426.885000 200.865000 480.000000 201.015000 ;
      RECT 426.900000 200.850000 480.000000 201.000000 ;
      RECT 426.900000 200.850000 480.000000 201.000000 ;
      RECT 427.035000 200.715000 480.000000 200.865000 ;
      RECT 427.050000 200.700000 480.000000 200.850000 ;
      RECT 427.050000 200.700000 480.000000 200.850000 ;
      RECT 427.185000 200.565000 480.000000 200.715000 ;
      RECT 427.200000 200.550000 480.000000 200.700000 ;
      RECT 427.200000 200.550000 480.000000 200.700000 ;
      RECT 427.335000 200.415000 480.000000 200.565000 ;
      RECT 427.350000 200.400000 480.000000 200.550000 ;
      RECT 427.350000 200.400000 480.000000 200.550000 ;
      RECT 427.485000 200.265000 480.000000 200.415000 ;
      RECT 427.500000 200.250000 480.000000 200.400000 ;
      RECT 427.500000 200.250000 480.000000 200.400000 ;
      RECT 427.635000 200.115000 480.000000 200.265000 ;
      RECT 427.650000 200.100000 480.000000 200.250000 ;
      RECT 427.650000 200.100000 480.000000 200.250000 ;
      RECT 427.785000 199.965000 480.000000 200.115000 ;
      RECT 427.800000 199.950000 480.000000 200.100000 ;
      RECT 427.800000 199.950000 480.000000 200.100000 ;
      RECT 427.935000 199.815000 480.000000 199.965000 ;
      RECT 427.950000 199.800000 480.000000 199.950000 ;
      RECT 427.950000 199.800000 480.000000 199.950000 ;
      RECT 428.085000 199.665000 480.000000 199.815000 ;
      RECT 428.100000 199.650000 480.000000 199.800000 ;
      RECT 428.100000 199.650000 480.000000 199.800000 ;
      RECT 428.235000 199.515000 480.000000 199.665000 ;
      RECT 428.250000 199.500000 480.000000 199.650000 ;
      RECT 428.250000 199.500000 480.000000 199.650000 ;
      RECT 428.385000 199.365000 480.000000 199.515000 ;
      RECT 428.400000 199.350000 480.000000 199.500000 ;
      RECT 428.400000 199.350000 480.000000 199.500000 ;
      RECT 428.535000 199.215000 480.000000 199.365000 ;
      RECT 428.550000 199.200000 480.000000 199.350000 ;
      RECT 428.550000 199.200000 480.000000 199.350000 ;
      RECT 428.685000 199.065000 480.000000 199.215000 ;
      RECT 428.700000 199.050000 480.000000 199.200000 ;
      RECT 428.700000 199.050000 480.000000 199.200000 ;
      RECT 428.835000 198.915000 480.000000 199.065000 ;
      RECT 428.850000 198.900000 480.000000 199.050000 ;
      RECT 428.850000 198.900000 480.000000 199.050000 ;
      RECT 428.985000 198.765000 480.000000 198.915000 ;
      RECT 429.000000 198.750000 480.000000 198.900000 ;
      RECT 429.000000 198.750000 480.000000 198.900000 ;
      RECT 429.135000 198.615000 480.000000 198.765000 ;
      RECT 429.150000 198.600000 480.000000 198.750000 ;
      RECT 429.150000 198.600000 480.000000 198.750000 ;
      RECT 429.285000 198.465000 480.000000 198.615000 ;
      RECT 429.300000 198.450000 480.000000 198.600000 ;
      RECT 429.300000 198.450000 480.000000 198.600000 ;
      RECT 429.435000 198.315000 480.000000 198.465000 ;
      RECT 429.450000 198.300000 480.000000 198.450000 ;
      RECT 429.450000 198.300000 480.000000 198.450000 ;
      RECT 429.585000 198.165000 480.000000 198.315000 ;
      RECT 429.600000 198.150000 480.000000 198.300000 ;
      RECT 429.600000 198.150000 480.000000 198.300000 ;
      RECT 429.735000 198.015000 480.000000 198.165000 ;
      RECT 429.750000 198.000000 480.000000 198.150000 ;
      RECT 429.750000 198.000000 480.000000 198.150000 ;
      RECT 429.885000 197.865000 480.000000 198.015000 ;
      RECT 429.900000 197.850000 480.000000 198.000000 ;
      RECT 429.900000 197.850000 480.000000 198.000000 ;
      RECT 430.035000 197.715000 480.000000 197.865000 ;
      RECT 430.050000 197.700000 480.000000 197.850000 ;
      RECT 430.050000 197.700000 480.000000 197.850000 ;
      RECT 430.185000 197.565000 480.000000 197.715000 ;
      RECT 430.200000 197.550000 480.000000 197.700000 ;
      RECT 430.200000 197.550000 480.000000 197.700000 ;
      RECT 430.335000 197.415000 480.000000 197.565000 ;
      RECT 430.350000 197.400000 480.000000 197.550000 ;
      RECT 430.350000 197.400000 480.000000 197.550000 ;
      RECT 430.485000 197.265000 480.000000 197.415000 ;
      RECT 430.500000 197.250000 480.000000 197.400000 ;
      RECT 430.500000 197.250000 480.000000 197.400000 ;
      RECT 430.635000 197.115000 480.000000 197.265000 ;
      RECT 430.650000 197.100000 480.000000 197.250000 ;
      RECT 430.650000 197.100000 480.000000 197.250000 ;
      RECT 430.785000 196.965000 480.000000 197.115000 ;
      RECT 430.800000 196.950000 480.000000 197.100000 ;
      RECT 430.800000 196.950000 480.000000 197.100000 ;
      RECT 430.935000 196.815000 480.000000 196.965000 ;
      RECT 430.950000 196.800000 480.000000 196.950000 ;
      RECT 430.950000 196.800000 480.000000 196.950000 ;
      RECT 431.085000 196.665000 480.000000 196.815000 ;
      RECT 431.100000 196.650000 480.000000 196.800000 ;
      RECT 431.100000 196.650000 480.000000 196.800000 ;
      RECT 431.235000 196.515000 480.000000 196.665000 ;
      RECT 431.250000 196.500000 480.000000 196.650000 ;
      RECT 431.250000 196.500000 480.000000 196.650000 ;
      RECT 431.385000 196.365000 480.000000 196.515000 ;
      RECT 431.400000 196.350000 480.000000 196.500000 ;
      RECT 431.400000 196.350000 480.000000 196.500000 ;
      RECT 431.535000 196.215000 480.000000 196.365000 ;
      RECT 431.550000 196.200000 480.000000 196.350000 ;
      RECT 431.550000 196.200000 480.000000 196.350000 ;
      RECT 431.685000 196.065000 480.000000 196.215000 ;
      RECT 431.700000 196.050000 480.000000 196.200000 ;
      RECT 431.700000 196.050000 480.000000 196.200000 ;
      RECT 431.835000 195.915000 480.000000 196.065000 ;
      RECT 431.850000 195.900000 480.000000 196.050000 ;
      RECT 431.850000 195.900000 480.000000 196.050000 ;
      RECT 431.985000 195.765000 480.000000 195.915000 ;
      RECT 432.000000 195.750000 480.000000 195.900000 ;
      RECT 432.000000 195.750000 480.000000 195.900000 ;
      RECT 432.135000 195.615000 480.000000 195.765000 ;
      RECT 432.150000 195.600000 480.000000 195.750000 ;
      RECT 432.150000 195.600000 480.000000 195.750000 ;
      RECT 432.285000 195.465000 480.000000 195.615000 ;
      RECT 432.300000 195.450000 480.000000 195.600000 ;
      RECT 432.300000 195.450000 480.000000 195.600000 ;
      RECT 432.435000 195.315000 480.000000 195.465000 ;
      RECT 432.450000 195.300000 480.000000 195.450000 ;
      RECT 432.450000 195.300000 480.000000 195.450000 ;
      RECT 432.585000 195.165000 480.000000 195.315000 ;
      RECT 432.600000 195.150000 480.000000 195.300000 ;
      RECT 432.600000 195.150000 480.000000 195.300000 ;
      RECT 432.735000 195.015000 480.000000 195.165000 ;
      RECT 432.750000 195.000000 480.000000 195.150000 ;
      RECT 432.750000 195.000000 480.000000 195.150000 ;
      RECT 432.885000 194.865000 480.000000 195.015000 ;
      RECT 432.900000 194.850000 480.000000 195.000000 ;
      RECT 432.900000 194.850000 480.000000 195.000000 ;
      RECT 433.035000 194.715000 480.000000 194.865000 ;
      RECT 433.050000 194.700000 480.000000 194.850000 ;
      RECT 433.050000 194.700000 480.000000 194.850000 ;
      RECT 433.185000 194.565000 480.000000 194.715000 ;
      RECT 433.200000 194.550000 480.000000 194.700000 ;
      RECT 433.200000 194.550000 480.000000 194.700000 ;
      RECT 433.335000 194.415000 480.000000 194.565000 ;
      RECT 433.350000 194.400000 480.000000 194.550000 ;
      RECT 433.350000 194.400000 480.000000 194.550000 ;
      RECT 433.485000 194.265000 480.000000 194.415000 ;
      RECT 433.500000 194.250000 480.000000 194.400000 ;
      RECT 433.500000 194.250000 480.000000 194.400000 ;
      RECT 433.635000 194.115000 480.000000 194.265000 ;
      RECT 433.650000 194.100000 480.000000 194.250000 ;
      RECT 433.650000 194.100000 480.000000 194.250000 ;
      RECT 433.785000 193.965000 480.000000 194.115000 ;
      RECT 433.800000 193.950000 480.000000 194.100000 ;
      RECT 433.800000 193.950000 480.000000 194.100000 ;
      RECT 433.935000 193.815000 480.000000 193.965000 ;
      RECT 433.950000 193.800000 480.000000 193.950000 ;
      RECT 433.950000 193.800000 480.000000 193.950000 ;
      RECT 434.085000 193.665000 480.000000 193.815000 ;
      RECT 434.100000 193.650000 480.000000 193.800000 ;
      RECT 434.100000 193.650000 480.000000 193.800000 ;
      RECT 434.235000 193.515000 480.000000 193.665000 ;
      RECT 434.250000 193.500000 480.000000 193.650000 ;
      RECT 434.250000 193.500000 480.000000 193.650000 ;
      RECT 434.385000 193.365000 480.000000 193.515000 ;
      RECT 434.400000 193.350000 480.000000 193.500000 ;
      RECT 434.400000 193.350000 480.000000 193.500000 ;
      RECT 434.535000 193.215000 480.000000 193.365000 ;
      RECT 434.550000 193.200000 480.000000 193.350000 ;
      RECT 434.550000 193.200000 480.000000 193.350000 ;
      RECT 434.685000 193.065000 480.000000 193.215000 ;
      RECT 434.700000 193.050000 480.000000 193.200000 ;
      RECT 434.700000 193.050000 480.000000 193.200000 ;
      RECT 434.835000 192.915000 480.000000 193.065000 ;
      RECT 434.850000 192.900000 480.000000 193.050000 ;
      RECT 434.850000 192.900000 480.000000 193.050000 ;
      RECT 434.985000 192.765000 480.000000 192.915000 ;
      RECT 435.000000 192.750000 480.000000 192.900000 ;
      RECT 435.000000 192.750000 480.000000 192.900000 ;
      RECT 435.135000 192.615000 480.000000 192.765000 ;
      RECT 435.150000 192.600000 480.000000 192.750000 ;
      RECT 435.150000 192.600000 480.000000 192.750000 ;
      RECT 435.285000 192.465000 480.000000 192.615000 ;
      RECT 435.300000 192.450000 480.000000 192.600000 ;
      RECT 435.300000 192.450000 480.000000 192.600000 ;
      RECT 435.435000 192.315000 480.000000 192.465000 ;
      RECT 435.450000 192.300000 480.000000 192.450000 ;
      RECT 435.450000 192.300000 480.000000 192.450000 ;
      RECT 435.585000 192.165000 480.000000 192.315000 ;
      RECT 435.600000 192.150000 480.000000 192.300000 ;
      RECT 435.600000 192.150000 480.000000 192.300000 ;
      RECT 435.735000 192.015000 480.000000 192.165000 ;
      RECT 435.750000 192.000000 480.000000 192.150000 ;
      RECT 435.750000 192.000000 480.000000 192.150000 ;
      RECT 435.885000 191.865000 480.000000 192.015000 ;
      RECT 435.900000 191.850000 480.000000 192.000000 ;
      RECT 435.900000 191.850000 480.000000 192.000000 ;
      RECT 436.035000 191.715000 480.000000 191.865000 ;
      RECT 436.050000 191.700000 480.000000 191.850000 ;
      RECT 436.050000 191.700000 480.000000 191.850000 ;
      RECT 436.185000 191.565000 480.000000 191.715000 ;
      RECT 436.200000 191.550000 480.000000 191.700000 ;
      RECT 436.200000 191.550000 480.000000 191.700000 ;
      RECT 436.335000 191.415000 480.000000 191.565000 ;
      RECT 436.350000 191.400000 480.000000 191.550000 ;
      RECT 436.350000 191.400000 480.000000 191.550000 ;
      RECT 436.485000 191.265000 480.000000 191.415000 ;
      RECT 436.500000 191.250000 480.000000 191.400000 ;
      RECT 436.500000 191.250000 480.000000 191.400000 ;
      RECT 436.635000 191.115000 480.000000 191.265000 ;
      RECT 436.650000 191.100000 480.000000 191.250000 ;
      RECT 436.650000 191.100000 480.000000 191.250000 ;
      RECT 436.785000 190.965000 480.000000 191.115000 ;
      RECT 436.800000 190.950000 480.000000 191.100000 ;
      RECT 436.800000 190.950000 480.000000 191.100000 ;
      RECT 436.935000 190.815000 480.000000 190.965000 ;
      RECT 436.950000 190.800000 480.000000 190.950000 ;
      RECT 436.950000 190.800000 480.000000 190.950000 ;
      RECT 437.085000 190.665000 480.000000 190.815000 ;
      RECT 437.100000 190.650000 480.000000 190.800000 ;
      RECT 437.100000 190.650000 480.000000 190.800000 ;
      RECT 437.235000 190.515000 480.000000 190.665000 ;
      RECT 437.250000 190.500000 480.000000 190.650000 ;
      RECT 437.250000 190.500000 480.000000 190.650000 ;
      RECT 437.385000 190.365000 480.000000 190.515000 ;
      RECT 437.400000 190.350000 480.000000 190.500000 ;
      RECT 437.400000 190.350000 480.000000 190.500000 ;
      RECT 437.535000 190.215000 480.000000 190.365000 ;
      RECT 437.550000 190.200000 480.000000 190.350000 ;
      RECT 437.550000 190.200000 480.000000 190.350000 ;
      RECT 437.685000 190.065000 480.000000 190.215000 ;
      RECT 437.700000 190.050000 480.000000 190.200000 ;
      RECT 437.700000 190.050000 480.000000 190.200000 ;
      RECT 437.835000 189.915000 480.000000 190.065000 ;
      RECT 437.850000 189.900000 480.000000 190.050000 ;
      RECT 437.850000 189.900000 480.000000 190.050000 ;
      RECT 437.985000 189.765000 480.000000 189.915000 ;
      RECT 438.000000 189.750000 480.000000 189.900000 ;
      RECT 438.000000 189.750000 480.000000 189.900000 ;
      RECT 438.135000 189.615000 480.000000 189.765000 ;
      RECT 438.150000 189.600000 480.000000 189.750000 ;
      RECT 438.150000 189.600000 480.000000 189.750000 ;
      RECT 438.285000 189.465000 480.000000 189.615000 ;
      RECT 438.300000 189.450000 480.000000 189.600000 ;
      RECT 438.300000 189.450000 480.000000 189.600000 ;
      RECT 438.435000 189.315000 480.000000 189.465000 ;
      RECT 438.450000 189.300000 480.000000 189.450000 ;
      RECT 438.450000 189.300000 480.000000 189.450000 ;
      RECT 438.585000 189.165000 480.000000 189.315000 ;
      RECT 438.600000 189.150000 480.000000 189.300000 ;
      RECT 438.600000 189.150000 480.000000 189.300000 ;
      RECT 438.735000 189.015000 480.000000 189.165000 ;
      RECT 438.750000 189.000000 480.000000 189.150000 ;
      RECT 438.750000 189.000000 480.000000 189.150000 ;
      RECT 438.885000 188.865000 480.000000 189.015000 ;
      RECT 438.900000 188.850000 480.000000 189.000000 ;
      RECT 438.900000 188.850000 480.000000 189.000000 ;
      RECT 439.035000 188.715000 480.000000 188.865000 ;
      RECT 439.050000 188.700000 480.000000 188.850000 ;
      RECT 439.050000 188.700000 480.000000 188.850000 ;
      RECT 439.185000 188.565000 480.000000 188.715000 ;
      RECT 439.200000 188.550000 480.000000 188.700000 ;
      RECT 439.200000 188.550000 480.000000 188.700000 ;
      RECT 439.335000 188.415000 480.000000 188.565000 ;
      RECT 439.350000 188.400000 480.000000 188.550000 ;
      RECT 439.350000 188.400000 480.000000 188.550000 ;
      RECT 439.485000 188.265000 480.000000 188.415000 ;
      RECT 439.500000 188.250000 480.000000 188.400000 ;
      RECT 439.500000 188.250000 480.000000 188.400000 ;
      RECT 439.635000 188.115000 480.000000 188.265000 ;
      RECT 439.650000 188.100000 480.000000 188.250000 ;
      RECT 439.650000 188.100000 480.000000 188.250000 ;
      RECT 439.785000 187.965000 480.000000 188.115000 ;
      RECT 439.800000 187.950000 480.000000 188.100000 ;
      RECT 439.800000 187.950000 480.000000 188.100000 ;
      RECT 439.935000 187.815000 480.000000 187.965000 ;
      RECT 439.950000 187.800000 480.000000 187.950000 ;
      RECT 439.950000 187.800000 480.000000 187.950000 ;
      RECT 440.085000 187.665000 480.000000 187.815000 ;
      RECT 440.100000 187.650000 480.000000 187.800000 ;
      RECT 440.100000 187.650000 480.000000 187.800000 ;
      RECT 440.235000 187.515000 480.000000 187.665000 ;
      RECT 440.250000 187.500000 480.000000 187.650000 ;
      RECT 440.250000 187.500000 480.000000 187.650000 ;
      RECT 440.385000 187.365000 480.000000 187.515000 ;
      RECT 440.400000 187.350000 480.000000 187.500000 ;
      RECT 440.400000 187.350000 480.000000 187.500000 ;
      RECT 440.535000 187.215000 480.000000 187.365000 ;
      RECT 440.550000 187.200000 480.000000 187.350000 ;
      RECT 440.550000 187.200000 480.000000 187.350000 ;
      RECT 440.685000 187.065000 480.000000 187.215000 ;
      RECT 440.700000 187.050000 480.000000 187.200000 ;
      RECT 440.700000 187.050000 480.000000 187.200000 ;
      RECT 440.835000 186.915000 480.000000 187.065000 ;
      RECT 440.850000 186.900000 480.000000 187.050000 ;
      RECT 440.850000 186.900000 480.000000 187.050000 ;
      RECT 440.985000 186.765000 480.000000 186.915000 ;
      RECT 441.000000 186.750000 480.000000 186.900000 ;
      RECT 441.000000 186.750000 480.000000 186.900000 ;
      RECT 441.135000 186.615000 480.000000 186.765000 ;
      RECT 441.150000 186.600000 480.000000 186.750000 ;
      RECT 441.150000 186.600000 480.000000 186.750000 ;
      RECT 441.285000 186.465000 480.000000 186.615000 ;
      RECT 441.300000 186.450000 480.000000 186.600000 ;
      RECT 441.300000 186.450000 480.000000 186.600000 ;
      RECT 441.435000 186.315000 480.000000 186.465000 ;
      RECT 441.450000 186.300000 480.000000 186.450000 ;
      RECT 441.450000 186.300000 480.000000 186.450000 ;
      RECT 441.585000 186.165000 480.000000 186.315000 ;
      RECT 441.600000 186.150000 480.000000 186.300000 ;
      RECT 441.600000 186.150000 480.000000 186.300000 ;
      RECT 441.735000 186.015000 480.000000 186.165000 ;
      RECT 441.750000 186.000000 480.000000 186.150000 ;
      RECT 441.750000 186.000000 480.000000 186.150000 ;
      RECT 441.885000 185.865000 480.000000 186.015000 ;
      RECT 441.900000 185.850000 480.000000 186.000000 ;
      RECT 441.900000 185.850000 480.000000 186.000000 ;
      RECT 442.035000 185.715000 480.000000 185.865000 ;
      RECT 442.050000 185.700000 480.000000 185.850000 ;
      RECT 442.050000 185.700000 480.000000 185.850000 ;
      RECT 442.185000 185.565000 480.000000 185.715000 ;
      RECT 442.200000 185.550000 480.000000 185.700000 ;
      RECT 442.200000 185.550000 480.000000 185.700000 ;
      RECT 442.335000 185.415000 480.000000 185.565000 ;
      RECT 442.350000 185.400000 480.000000 185.550000 ;
      RECT 442.350000 185.400000 480.000000 185.550000 ;
      RECT 442.485000 185.265000 480.000000 185.415000 ;
      RECT 442.500000 185.250000 480.000000 185.400000 ;
      RECT 442.500000 185.250000 480.000000 185.400000 ;
      RECT 442.635000 185.115000 480.000000 185.265000 ;
      RECT 442.650000 185.100000 480.000000 185.250000 ;
      RECT 442.650000 185.100000 480.000000 185.250000 ;
      RECT 442.785000 184.965000 480.000000 185.115000 ;
      RECT 442.800000 184.950000 480.000000 185.100000 ;
      RECT 442.800000 184.950000 480.000000 185.100000 ;
      RECT 442.935000 184.815000 480.000000 184.965000 ;
      RECT 442.950000 184.800000 480.000000 184.950000 ;
      RECT 442.950000 184.800000 480.000000 184.950000 ;
      RECT 443.085000 184.665000 480.000000 184.815000 ;
      RECT 443.100000 184.650000 480.000000 184.800000 ;
      RECT 443.100000 184.650000 480.000000 184.800000 ;
      RECT 443.235000 184.515000 480.000000 184.665000 ;
      RECT 443.250000 184.500000 480.000000 184.650000 ;
      RECT 443.250000 184.500000 480.000000 184.650000 ;
      RECT 443.385000 184.365000 480.000000 184.515000 ;
      RECT 443.400000 184.350000 480.000000 184.500000 ;
      RECT 443.400000 184.350000 480.000000 184.500000 ;
      RECT 443.535000 184.215000 480.000000 184.365000 ;
      RECT 443.550000 184.200000 480.000000 184.350000 ;
      RECT 443.550000 184.200000 480.000000 184.350000 ;
      RECT 443.685000 184.065000 480.000000 184.215000 ;
      RECT 443.700000 184.050000 480.000000 184.200000 ;
      RECT 443.700000 184.050000 480.000000 184.200000 ;
      RECT 443.835000 183.915000 480.000000 184.065000 ;
      RECT 443.850000 183.900000 480.000000 184.050000 ;
      RECT 443.850000 183.900000 480.000000 184.050000 ;
      RECT 443.985000 183.765000 480.000000 183.915000 ;
      RECT 444.000000 183.750000 480.000000 183.900000 ;
      RECT 444.000000 183.750000 480.000000 183.900000 ;
      RECT 444.135000 183.615000 480.000000 183.765000 ;
      RECT 444.150000 183.600000 480.000000 183.750000 ;
      RECT 444.150000 183.600000 480.000000 183.750000 ;
      RECT 444.285000 183.465000 480.000000 183.615000 ;
      RECT 444.300000 183.450000 480.000000 183.600000 ;
      RECT 444.300000 183.450000 480.000000 183.600000 ;
      RECT 444.435000 183.315000 480.000000 183.465000 ;
      RECT 444.450000 183.300000 480.000000 183.450000 ;
      RECT 444.450000 183.300000 480.000000 183.450000 ;
      RECT 444.585000 183.165000 480.000000 183.315000 ;
      RECT 444.600000 183.150000 480.000000 183.300000 ;
      RECT 444.600000 183.150000 480.000000 183.300000 ;
      RECT 444.735000 183.015000 480.000000 183.165000 ;
      RECT 444.750000 183.000000 480.000000 183.150000 ;
      RECT 444.750000 183.000000 480.000000 183.150000 ;
      RECT 444.885000 182.865000 480.000000 183.015000 ;
      RECT 444.900000 182.850000 480.000000 183.000000 ;
      RECT 444.900000 182.850000 480.000000 183.000000 ;
      RECT 445.035000 182.715000 480.000000 182.865000 ;
      RECT 445.050000 182.700000 480.000000 182.850000 ;
      RECT 445.050000 182.700000 480.000000 182.850000 ;
      RECT 445.185000 182.565000 480.000000 182.715000 ;
      RECT 445.200000 182.550000 480.000000 182.700000 ;
      RECT 445.200000 182.550000 480.000000 182.700000 ;
      RECT 445.335000 182.415000 480.000000 182.565000 ;
      RECT 445.350000 182.400000 480.000000 182.550000 ;
      RECT 445.350000 182.400000 480.000000 182.550000 ;
      RECT 445.485000 182.265000 480.000000 182.415000 ;
      RECT 445.500000 182.250000 480.000000 182.400000 ;
      RECT 445.500000 182.250000 480.000000 182.400000 ;
      RECT 445.635000 182.115000 480.000000 182.265000 ;
      RECT 445.650000 182.100000 480.000000 182.250000 ;
      RECT 445.650000 182.100000 480.000000 182.250000 ;
      RECT 445.785000 181.965000 480.000000 182.115000 ;
      RECT 445.800000 181.950000 480.000000 182.100000 ;
      RECT 445.800000 181.950000 480.000000 182.100000 ;
      RECT 445.935000 181.815000 480.000000 181.965000 ;
      RECT 445.950000 181.800000 480.000000 181.950000 ;
      RECT 445.950000 181.800000 480.000000 181.950000 ;
      RECT 446.085000 181.665000 480.000000 181.815000 ;
      RECT 446.100000 181.650000 480.000000 181.800000 ;
      RECT 446.100000 181.650000 480.000000 181.800000 ;
      RECT 446.235000 181.515000 480.000000 181.665000 ;
      RECT 446.250000 181.500000 480.000000 181.650000 ;
      RECT 446.250000 181.500000 480.000000 181.650000 ;
      RECT 446.385000 181.365000 480.000000 181.515000 ;
      RECT 446.400000 181.350000 480.000000 181.500000 ;
      RECT 446.400000 181.350000 480.000000 181.500000 ;
      RECT 446.535000 181.215000 480.000000 181.365000 ;
      RECT 446.550000 181.200000 480.000000 181.350000 ;
      RECT 446.550000 181.200000 480.000000 181.350000 ;
      RECT 446.685000 181.065000 480.000000 181.215000 ;
      RECT 446.700000 181.050000 480.000000 181.200000 ;
      RECT 446.700000 181.050000 480.000000 181.200000 ;
      RECT 446.835000 180.915000 480.000000 181.065000 ;
      RECT 446.850000 180.900000 480.000000 181.050000 ;
      RECT 446.850000 180.900000 480.000000 181.050000 ;
      RECT 446.985000 180.765000 480.000000 180.915000 ;
      RECT 447.000000 180.750000 480.000000 180.900000 ;
      RECT 447.000000 180.750000 480.000000 180.900000 ;
      RECT 447.135000 180.615000 480.000000 180.765000 ;
      RECT 447.150000 180.600000 480.000000 180.750000 ;
      RECT 447.150000 180.600000 480.000000 180.750000 ;
      RECT 447.285000 180.465000 480.000000 180.615000 ;
      RECT 447.300000 180.450000 480.000000 180.600000 ;
      RECT 447.300000 180.450000 480.000000 180.600000 ;
      RECT 447.435000 180.315000 480.000000 180.465000 ;
      RECT 447.450000 180.300000 480.000000 180.450000 ;
      RECT 447.450000 180.300000 480.000000 180.450000 ;
      RECT 447.585000 180.165000 480.000000 180.315000 ;
      RECT 447.600000 180.150000 480.000000 180.300000 ;
      RECT 447.600000 180.150000 480.000000 180.300000 ;
      RECT 447.735000 180.015000 480.000000 180.165000 ;
      RECT 447.750000 180.000000 480.000000 180.150000 ;
      RECT 447.750000 180.000000 480.000000 180.150000 ;
      RECT 447.885000 179.865000 480.000000 180.015000 ;
      RECT 447.900000 179.850000 480.000000 180.000000 ;
      RECT 447.900000 179.850000 480.000000 180.000000 ;
      RECT 448.035000 179.715000 480.000000 179.865000 ;
      RECT 448.050000 179.700000 480.000000 179.850000 ;
      RECT 448.050000 179.700000 480.000000 179.850000 ;
      RECT 448.185000 179.565000 480.000000 179.715000 ;
      RECT 448.200000 179.550000 480.000000 179.700000 ;
      RECT 448.200000 179.550000 480.000000 179.700000 ;
      RECT 448.335000 179.415000 480.000000 179.565000 ;
      RECT 448.350000 179.400000 480.000000 179.550000 ;
      RECT 448.350000 179.400000 480.000000 179.550000 ;
      RECT 448.485000 179.265000 480.000000 179.415000 ;
      RECT 448.500000 179.250000 480.000000 179.400000 ;
      RECT 448.500000 179.250000 480.000000 179.400000 ;
      RECT 448.635000 179.115000 480.000000 179.265000 ;
      RECT 448.650000 179.100000 480.000000 179.250000 ;
      RECT 448.650000 179.100000 480.000000 179.250000 ;
      RECT 448.785000 178.965000 480.000000 179.115000 ;
      RECT 448.800000 178.950000 480.000000 179.100000 ;
      RECT 448.800000 178.950000 480.000000 179.100000 ;
      RECT 448.935000 178.815000 480.000000 178.965000 ;
      RECT 448.950000 178.800000 480.000000 178.950000 ;
      RECT 448.950000 178.800000 480.000000 178.950000 ;
      RECT 449.085000 178.665000 480.000000 178.815000 ;
      RECT 449.100000 178.650000 480.000000 178.800000 ;
      RECT 449.100000 178.650000 480.000000 178.800000 ;
      RECT 449.235000 178.515000 480.000000 178.665000 ;
      RECT 449.250000 178.500000 480.000000 178.650000 ;
      RECT 449.250000 178.500000 480.000000 178.650000 ;
      RECT 449.385000 178.365000 480.000000 178.515000 ;
      RECT 449.400000 178.350000 480.000000 178.500000 ;
      RECT 449.400000 178.350000 480.000000 178.500000 ;
      RECT 449.535000 178.215000 480.000000 178.365000 ;
      RECT 449.550000 178.200000 480.000000 178.350000 ;
      RECT 449.550000 178.200000 480.000000 178.350000 ;
      RECT 449.685000 178.065000 480.000000 178.215000 ;
      RECT 449.700000 178.050000 480.000000 178.200000 ;
      RECT 449.700000 178.050000 480.000000 178.200000 ;
      RECT 449.835000 177.915000 480.000000 178.065000 ;
      RECT 449.850000 177.900000 480.000000 178.050000 ;
      RECT 449.850000 177.900000 480.000000 178.050000 ;
      RECT 449.985000 177.765000 480.000000 177.915000 ;
      RECT 450.000000 177.750000 480.000000 177.900000 ;
      RECT 450.000000 177.750000 480.000000 177.900000 ;
      RECT 450.135000 177.615000 480.000000 177.765000 ;
      RECT 450.150000 177.600000 480.000000 177.750000 ;
      RECT 450.150000 177.600000 480.000000 177.750000 ;
      RECT 450.285000 177.465000 480.000000 177.615000 ;
      RECT 450.300000 177.450000 480.000000 177.600000 ;
      RECT 450.300000 177.450000 480.000000 177.600000 ;
      RECT 450.435000 177.315000 480.000000 177.465000 ;
      RECT 450.450000 177.300000 480.000000 177.450000 ;
      RECT 450.450000 177.300000 480.000000 177.450000 ;
      RECT 450.585000 177.165000 480.000000 177.315000 ;
      RECT 450.600000 177.150000 480.000000 177.300000 ;
      RECT 450.600000 177.150000 480.000000 177.300000 ;
      RECT 450.735000 177.015000 480.000000 177.165000 ;
      RECT 450.750000 177.000000 480.000000 177.150000 ;
      RECT 450.750000 177.000000 480.000000 177.150000 ;
      RECT 450.885000 176.865000 480.000000 177.015000 ;
      RECT 450.900000 176.850000 480.000000 177.000000 ;
      RECT 450.900000 176.850000 480.000000 177.000000 ;
      RECT 451.035000 176.715000 480.000000 176.865000 ;
      RECT 451.050000 176.700000 480.000000 176.850000 ;
      RECT 451.050000 176.700000 480.000000 176.850000 ;
      RECT 451.185000 176.565000 480.000000 176.715000 ;
      RECT 451.200000 176.550000 480.000000 176.700000 ;
      RECT 451.200000 176.550000 480.000000 176.700000 ;
      RECT 451.335000 176.415000 480.000000 176.565000 ;
      RECT 451.350000 176.400000 480.000000 176.550000 ;
      RECT 451.350000 176.400000 480.000000 176.550000 ;
      RECT 451.485000 176.265000 480.000000 176.415000 ;
      RECT 451.500000 176.250000 480.000000 176.400000 ;
      RECT 451.500000 176.250000 480.000000 176.400000 ;
      RECT 451.635000 176.115000 480.000000 176.265000 ;
      RECT 451.650000 176.100000 480.000000 176.250000 ;
      RECT 451.650000 176.100000 480.000000 176.250000 ;
      RECT 451.785000 175.965000 480.000000 176.115000 ;
      RECT 451.800000 175.950000 480.000000 176.100000 ;
      RECT 451.800000 175.950000 480.000000 176.100000 ;
      RECT 451.935000 175.815000 480.000000 175.965000 ;
      RECT 451.950000 175.800000 480.000000 175.950000 ;
      RECT 451.950000 175.800000 480.000000 175.950000 ;
      RECT 452.085000 175.665000 480.000000 175.815000 ;
      RECT 452.100000 175.650000 480.000000 175.800000 ;
      RECT 452.100000 175.650000 480.000000 175.800000 ;
      RECT 452.235000 175.515000 480.000000 175.665000 ;
      RECT 452.250000 175.500000 480.000000 175.650000 ;
      RECT 452.250000 175.500000 480.000000 175.650000 ;
      RECT 452.385000 175.365000 480.000000 175.515000 ;
      RECT 452.400000 175.350000 480.000000 175.500000 ;
      RECT 452.400000 175.350000 480.000000 175.500000 ;
      RECT 452.535000 175.215000 480.000000 175.365000 ;
      RECT 452.550000 175.200000 480.000000 175.350000 ;
      RECT 452.550000 175.200000 480.000000 175.350000 ;
      RECT 452.685000 175.065000 480.000000 175.215000 ;
      RECT 452.700000 175.050000 480.000000 175.200000 ;
      RECT 452.700000 175.050000 480.000000 175.200000 ;
      RECT 452.835000 174.915000 480.000000 175.065000 ;
      RECT 452.850000 174.900000 480.000000 175.050000 ;
      RECT 452.850000 174.900000 480.000000 175.050000 ;
      RECT 452.985000 174.765000 480.000000 174.915000 ;
      RECT 453.000000 174.750000 480.000000 174.900000 ;
      RECT 453.000000 174.750000 480.000000 174.900000 ;
      RECT 453.135000 174.615000 480.000000 174.765000 ;
      RECT 453.150000 174.600000 480.000000 174.750000 ;
      RECT 453.150000 174.600000 480.000000 174.750000 ;
      RECT 453.285000 174.465000 480.000000 174.615000 ;
      RECT 453.300000 174.450000 480.000000 174.600000 ;
      RECT 453.300000 174.450000 480.000000 174.600000 ;
      RECT 453.435000 174.315000 480.000000 174.465000 ;
      RECT 453.450000 174.300000 480.000000 174.450000 ;
      RECT 453.450000 174.300000 480.000000 174.450000 ;
      RECT 453.585000 174.165000 480.000000 174.315000 ;
      RECT 453.600000 174.150000 480.000000 174.300000 ;
      RECT 453.600000 174.150000 480.000000 174.300000 ;
      RECT 453.735000 174.015000 480.000000 174.165000 ;
      RECT 453.750000 174.000000 480.000000 174.150000 ;
      RECT 453.750000 174.000000 480.000000 174.150000 ;
      RECT 453.885000 173.865000 480.000000 174.015000 ;
      RECT 453.900000 173.850000 480.000000 174.000000 ;
      RECT 453.900000 173.850000 480.000000 174.000000 ;
      RECT 454.035000 173.715000 480.000000 173.865000 ;
      RECT 454.050000 173.700000 480.000000 173.850000 ;
      RECT 454.050000 173.700000 480.000000 173.850000 ;
      RECT 454.185000 173.565000 480.000000 173.715000 ;
      RECT 454.200000 173.550000 480.000000 173.700000 ;
      RECT 454.200000 173.550000 480.000000 173.700000 ;
      RECT 454.335000 173.415000 480.000000 173.565000 ;
      RECT 454.350000 173.400000 480.000000 173.550000 ;
      RECT 454.350000 173.400000 480.000000 173.550000 ;
      RECT 454.485000 173.265000 480.000000 173.415000 ;
      RECT 454.500000 173.250000 480.000000 173.400000 ;
      RECT 454.500000 173.250000 480.000000 173.400000 ;
      RECT 454.635000 173.115000 480.000000 173.265000 ;
      RECT 454.650000 173.100000 480.000000 173.250000 ;
      RECT 454.650000 173.100000 480.000000 173.250000 ;
      RECT 454.785000 172.965000 480.000000 173.115000 ;
      RECT 454.800000 172.950000 480.000000 173.100000 ;
      RECT 454.800000 172.950000 480.000000 173.100000 ;
      RECT 454.935000 172.815000 480.000000 172.965000 ;
      RECT 454.950000 172.800000 480.000000 172.950000 ;
      RECT 454.950000 172.800000 480.000000 172.950000 ;
      RECT 455.085000 172.665000 480.000000 172.815000 ;
      RECT 455.100000 172.650000 480.000000 172.800000 ;
      RECT 455.100000 172.650000 480.000000 172.800000 ;
      RECT 455.235000 172.515000 480.000000 172.665000 ;
      RECT 455.250000 172.500000 480.000000 172.650000 ;
      RECT 455.250000 172.500000 480.000000 172.650000 ;
      RECT 455.385000 172.365000 480.000000 172.515000 ;
      RECT 455.400000 172.350000 480.000000 172.500000 ;
      RECT 455.400000 172.350000 480.000000 172.500000 ;
      RECT 455.535000 172.215000 480.000000 172.365000 ;
      RECT 455.550000 172.200000 480.000000 172.350000 ;
      RECT 455.550000 172.200000 480.000000 172.350000 ;
      RECT 455.685000 172.065000 480.000000 172.215000 ;
      RECT 455.700000 172.050000 480.000000 172.200000 ;
      RECT 455.700000 172.050000 480.000000 172.200000 ;
      RECT 455.835000 171.915000 480.000000 172.065000 ;
      RECT 455.850000 171.900000 480.000000 172.050000 ;
      RECT 455.850000 171.900000 480.000000 172.050000 ;
      RECT 455.985000 171.765000 480.000000 171.915000 ;
      RECT 456.000000 171.750000 480.000000 171.900000 ;
      RECT 456.000000 171.750000 480.000000 171.900000 ;
      RECT 456.135000 171.615000 480.000000 171.765000 ;
      RECT 456.150000 171.600000 480.000000 171.750000 ;
      RECT 456.150000 171.600000 480.000000 171.750000 ;
      RECT 456.285000 171.465000 480.000000 171.615000 ;
      RECT 456.300000 171.450000 480.000000 171.600000 ;
      RECT 456.300000 171.450000 480.000000 171.600000 ;
      RECT 456.435000 171.315000 480.000000 171.465000 ;
      RECT 456.450000 171.300000 480.000000 171.450000 ;
      RECT 456.450000 171.300000 480.000000 171.450000 ;
      RECT 456.585000 171.165000 480.000000 171.315000 ;
      RECT 456.600000 171.150000 480.000000 171.300000 ;
      RECT 456.600000 171.150000 480.000000 171.300000 ;
      RECT 456.735000 171.015000 480.000000 171.165000 ;
      RECT 456.750000 171.000000 480.000000 171.150000 ;
      RECT 456.750000 171.000000 480.000000 171.150000 ;
      RECT 456.885000 170.865000 480.000000 171.015000 ;
      RECT 456.900000 170.850000 480.000000 171.000000 ;
      RECT 456.900000 170.850000 480.000000 171.000000 ;
      RECT 457.035000 170.715000 480.000000 170.865000 ;
      RECT 457.050000 170.700000 480.000000 170.850000 ;
      RECT 457.050000 170.700000 480.000000 170.850000 ;
      RECT 457.185000 170.565000 480.000000 170.715000 ;
      RECT 457.200000 170.550000 480.000000 170.700000 ;
      RECT 457.200000 170.550000 480.000000 170.700000 ;
      RECT 457.335000 170.415000 480.000000 170.565000 ;
      RECT 457.350000 170.400000 480.000000 170.550000 ;
      RECT 457.350000 170.400000 480.000000 170.550000 ;
      RECT 457.485000 170.265000 480.000000 170.415000 ;
      RECT 457.500000 170.250000 480.000000 170.400000 ;
      RECT 457.500000 170.250000 480.000000 170.400000 ;
      RECT 457.635000 170.115000 480.000000 170.265000 ;
      RECT 457.650000 170.100000 480.000000 170.250000 ;
      RECT 457.650000 170.100000 480.000000 170.250000 ;
      RECT 457.785000 169.965000 480.000000 170.115000 ;
      RECT 457.800000 169.950000 480.000000 170.100000 ;
      RECT 457.800000 169.950000 480.000000 170.100000 ;
      RECT 457.935000 169.815000 480.000000 169.965000 ;
      RECT 457.950000 169.800000 480.000000 169.950000 ;
      RECT 457.950000 169.800000 480.000000 169.950000 ;
      RECT 458.050000  73.115000 480.000000  73.200000 ;
      RECT 458.085000 169.665000 480.000000 169.815000 ;
      RECT 458.100000 169.650000 480.000000 169.800000 ;
      RECT 458.100000 169.650000 480.000000 169.800000 ;
      RECT 458.130000  73.015000 480.000000  73.055000 ;
      RECT 458.170000  73.055000 480.000000  73.095000 ;
      RECT 458.175000  73.095000 480.000000  73.100000 ;
      RECT 458.235000 169.515000 480.000000 169.665000 ;
      RECT 458.250000 169.500000 480.000000 169.650000 ;
      RECT 458.250000 169.500000 480.000000 169.650000 ;
      RECT 458.385000 169.365000 480.000000 169.515000 ;
      RECT 458.400000 169.350000 480.000000 169.500000 ;
      RECT 458.400000 169.350000 480.000000 169.500000 ;
      RECT 458.535000 169.215000 480.000000 169.365000 ;
      RECT 458.550000 169.200000 480.000000 169.350000 ;
      RECT 458.550000 169.200000 480.000000 169.350000 ;
      RECT 458.685000 169.065000 480.000000 169.215000 ;
      RECT 458.700000 169.050000 480.000000 169.200000 ;
      RECT 458.700000 169.050000 480.000000 169.200000 ;
      RECT 458.835000 168.915000 480.000000 169.065000 ;
      RECT 458.850000 168.900000 480.000000 169.050000 ;
      RECT 458.850000 168.900000 480.000000 169.050000 ;
      RECT 458.985000 168.765000 480.000000 168.915000 ;
      RECT 459.000000 168.750000 480.000000 168.900000 ;
      RECT 459.000000 168.750000 480.000000 168.900000 ;
      RECT 459.135000 168.615000 480.000000 168.765000 ;
      RECT 459.150000 168.600000 480.000000 168.750000 ;
      RECT 459.150000 168.600000 480.000000 168.750000 ;
      RECT 459.285000 168.465000 480.000000 168.615000 ;
      RECT 459.300000 168.450000 480.000000 168.600000 ;
      RECT 459.300000 168.450000 480.000000 168.600000 ;
      RECT 459.435000 168.315000 480.000000 168.465000 ;
      RECT 459.450000 168.300000 480.000000 168.450000 ;
      RECT 459.450000 168.300000 480.000000 168.450000 ;
      RECT 459.585000 168.165000 480.000000 168.315000 ;
      RECT 459.600000 168.150000 480.000000 168.300000 ;
      RECT 459.600000 168.150000 480.000000 168.300000 ;
      RECT 459.735000 168.015000 480.000000 168.165000 ;
      RECT 459.750000 168.000000 480.000000 168.150000 ;
      RECT 459.750000 168.000000 480.000000 168.150000 ;
      RECT 459.885000 167.865000 480.000000 168.015000 ;
      RECT 459.900000 167.850000 480.000000 168.000000 ;
      RECT 459.900000 167.850000 480.000000 168.000000 ;
      RECT 460.035000 167.715000 480.000000 167.865000 ;
      RECT 460.050000 167.700000 480.000000 167.850000 ;
      RECT 460.050000 167.700000 480.000000 167.850000 ;
      RECT 460.185000 167.565000 480.000000 167.715000 ;
      RECT 460.200000 167.550000 480.000000 167.700000 ;
      RECT 460.200000 167.550000 480.000000 167.700000 ;
      RECT 460.335000 167.415000 480.000000 167.565000 ;
      RECT 460.350000 167.400000 480.000000 167.550000 ;
      RECT 460.350000 167.400000 480.000000 167.550000 ;
      RECT 460.485000 167.265000 480.000000 167.415000 ;
      RECT 460.500000 167.250000 480.000000 167.400000 ;
      RECT 460.500000 167.250000 480.000000 167.400000 ;
      RECT 460.635000 167.115000 480.000000 167.265000 ;
      RECT 460.650000 167.100000 480.000000 167.250000 ;
      RECT 460.650000 167.100000 480.000000 167.250000 ;
      RECT 460.785000 166.965000 480.000000 167.115000 ;
      RECT 460.800000 166.950000 480.000000 167.100000 ;
      RECT 460.800000 166.950000 480.000000 167.100000 ;
      RECT 460.935000 166.815000 480.000000 166.965000 ;
      RECT 460.950000 166.800000 480.000000 166.950000 ;
      RECT 460.950000 166.800000 480.000000 166.950000 ;
      RECT 461.085000 166.665000 480.000000 166.815000 ;
      RECT 461.100000 166.650000 480.000000 166.800000 ;
      RECT 461.100000 166.650000 480.000000 166.800000 ;
      RECT 461.235000 166.515000 480.000000 166.665000 ;
      RECT 461.250000 166.500000 480.000000 166.650000 ;
      RECT 461.250000 166.500000 480.000000 166.650000 ;
      RECT 461.385000 166.365000 480.000000 166.515000 ;
      RECT 461.400000 166.350000 480.000000 166.500000 ;
      RECT 461.400000 166.350000 480.000000 166.500000 ;
      RECT 461.535000 166.215000 480.000000 166.365000 ;
      RECT 461.550000 166.200000 480.000000 166.350000 ;
      RECT 461.550000 166.200000 480.000000 166.350000 ;
      RECT 461.685000 166.065000 480.000000 166.215000 ;
      RECT 461.700000 166.050000 480.000000 166.200000 ;
      RECT 461.700000 166.050000 480.000000 166.200000 ;
      RECT 461.835000 165.915000 480.000000 166.065000 ;
      RECT 461.850000 165.900000 480.000000 166.050000 ;
      RECT 461.850000 165.900000 480.000000 166.050000 ;
      RECT 461.985000 165.765000 480.000000 165.915000 ;
      RECT 462.000000 165.750000 480.000000 165.900000 ;
      RECT 462.000000 165.750000 480.000000 165.900000 ;
      RECT 462.135000 165.615000 480.000000 165.765000 ;
      RECT 462.150000 165.600000 480.000000 165.750000 ;
      RECT 462.150000 165.600000 480.000000 165.750000 ;
      RECT 462.285000 165.465000 480.000000 165.615000 ;
      RECT 462.300000 165.450000 480.000000 165.600000 ;
      RECT 462.300000 165.450000 480.000000 165.600000 ;
      RECT 462.435000 165.315000 480.000000 165.465000 ;
      RECT 462.450000 165.300000 480.000000 165.450000 ;
      RECT 462.450000 165.300000 480.000000 165.450000 ;
      RECT 462.585000 165.165000 480.000000 165.315000 ;
      RECT 462.600000 165.150000 480.000000 165.300000 ;
      RECT 462.600000 165.150000 480.000000 165.300000 ;
      RECT 462.735000 165.015000 480.000000 165.165000 ;
      RECT 462.750000 165.000000 480.000000 165.150000 ;
      RECT 462.750000 165.000000 480.000000 165.150000 ;
      RECT 462.885000 164.865000 480.000000 165.015000 ;
      RECT 462.900000 164.850000 480.000000 165.000000 ;
      RECT 462.900000 164.850000 480.000000 165.000000 ;
      RECT 463.035000 164.715000 480.000000 164.865000 ;
      RECT 463.050000 164.700000 480.000000 164.850000 ;
      RECT 463.050000 164.700000 480.000000 164.850000 ;
      RECT 463.185000 164.565000 480.000000 164.715000 ;
      RECT 463.200000 164.550000 480.000000 164.700000 ;
      RECT 463.200000 164.550000 480.000000 164.700000 ;
      RECT 463.335000 164.415000 480.000000 164.565000 ;
      RECT 463.350000 164.400000 480.000000 164.550000 ;
      RECT 463.350000 164.400000 480.000000 164.550000 ;
      RECT 463.485000 164.265000 480.000000 164.415000 ;
      RECT 463.500000 164.250000 480.000000 164.400000 ;
      RECT 463.500000 164.250000 480.000000 164.400000 ;
      RECT 463.635000 164.115000 480.000000 164.265000 ;
      RECT 463.650000 164.100000 480.000000 164.250000 ;
      RECT 463.650000 164.100000 480.000000 164.250000 ;
      RECT 463.785000 163.965000 480.000000 164.115000 ;
      RECT 463.800000 163.950000 480.000000 164.100000 ;
      RECT 463.800000 163.950000 480.000000 164.100000 ;
      RECT 463.935000 163.815000 480.000000 163.965000 ;
      RECT 463.950000 163.800000 480.000000 163.950000 ;
      RECT 463.950000 163.800000 480.000000 163.950000 ;
      RECT 464.085000 163.665000 480.000000 163.815000 ;
      RECT 464.100000 163.650000 480.000000 163.800000 ;
      RECT 464.100000 163.650000 480.000000 163.800000 ;
      RECT 464.235000 163.515000 480.000000 163.665000 ;
      RECT 464.250000 163.500000 480.000000 163.650000 ;
      RECT 464.250000 163.500000 480.000000 163.650000 ;
      RECT 464.385000 163.365000 480.000000 163.515000 ;
      RECT 464.400000 163.350000 480.000000 163.500000 ;
      RECT 464.400000 163.350000 480.000000 163.500000 ;
      RECT 464.535000 163.215000 480.000000 163.365000 ;
      RECT 464.550000 163.200000 480.000000 163.350000 ;
      RECT 464.550000 163.200000 480.000000 163.350000 ;
      RECT 464.685000 163.065000 480.000000 163.215000 ;
      RECT 464.700000 163.050000 480.000000 163.200000 ;
      RECT 464.700000 163.050000 480.000000 163.200000 ;
      RECT 464.835000 162.915000 480.000000 163.065000 ;
      RECT 464.850000 162.900000 480.000000 163.050000 ;
      RECT 464.850000 162.900000 480.000000 163.050000 ;
      RECT 464.985000 162.765000 480.000000 162.915000 ;
      RECT 465.000000 162.750000 480.000000 162.900000 ;
      RECT 465.000000 162.750000 480.000000 162.900000 ;
      RECT 465.135000 162.615000 480.000000 162.765000 ;
      RECT 465.150000 162.600000 480.000000 162.750000 ;
      RECT 465.150000 162.600000 480.000000 162.750000 ;
      RECT 465.285000 162.465000 480.000000 162.615000 ;
      RECT 465.300000 162.450000 480.000000 162.600000 ;
      RECT 465.300000 162.450000 480.000000 162.600000 ;
      RECT 465.435000 162.315000 480.000000 162.465000 ;
      RECT 465.450000 162.300000 480.000000 162.450000 ;
      RECT 465.450000 162.300000 480.000000 162.450000 ;
      RECT 465.585000 162.165000 480.000000 162.315000 ;
      RECT 465.600000 162.150000 480.000000 162.300000 ;
      RECT 465.600000 162.150000 480.000000 162.300000 ;
      RECT 465.735000 162.015000 480.000000 162.165000 ;
      RECT 465.750000 162.000000 480.000000 162.150000 ;
      RECT 465.750000 162.000000 480.000000 162.150000 ;
      RECT 465.885000 161.865000 480.000000 162.015000 ;
      RECT 465.900000 161.850000 480.000000 162.000000 ;
      RECT 465.900000 161.850000 480.000000 162.000000 ;
      RECT 466.035000 161.715000 480.000000 161.865000 ;
      RECT 466.050000 161.700000 480.000000 161.850000 ;
      RECT 466.050000 161.700000 480.000000 161.850000 ;
      RECT 466.185000 161.565000 480.000000 161.715000 ;
      RECT 466.200000 161.550000 480.000000 161.700000 ;
      RECT 466.200000 161.550000 480.000000 161.700000 ;
      RECT 466.335000 161.415000 480.000000 161.565000 ;
      RECT 466.350000 161.400000 480.000000 161.550000 ;
      RECT 466.350000 161.400000 480.000000 161.550000 ;
      RECT 466.485000 161.265000 480.000000 161.415000 ;
      RECT 466.500000 161.250000 480.000000 161.400000 ;
      RECT 466.500000 161.250000 480.000000 161.400000 ;
      RECT 466.635000 161.115000 480.000000 161.265000 ;
      RECT 466.650000 161.100000 480.000000 161.250000 ;
      RECT 466.650000 161.100000 480.000000 161.250000 ;
      RECT 466.785000 160.965000 480.000000 161.115000 ;
      RECT 466.800000 160.950000 480.000000 161.100000 ;
      RECT 466.800000 160.950000 480.000000 161.100000 ;
      RECT 466.935000 160.815000 480.000000 160.965000 ;
      RECT 466.950000 160.800000 480.000000 160.950000 ;
      RECT 466.950000 160.800000 480.000000 160.950000 ;
      RECT 467.085000 160.665000 480.000000 160.815000 ;
      RECT 467.100000 160.650000 480.000000 160.800000 ;
      RECT 467.100000 160.650000 480.000000 160.800000 ;
      RECT 467.235000 160.515000 480.000000 160.665000 ;
      RECT 467.250000 160.500000 480.000000 160.650000 ;
      RECT 467.250000 160.500000 480.000000 160.650000 ;
      RECT 467.385000 160.365000 480.000000 160.515000 ;
      RECT 467.400000 160.350000 480.000000 160.500000 ;
      RECT 467.400000 160.350000 480.000000 160.500000 ;
      RECT 467.535000 160.215000 480.000000 160.365000 ;
      RECT 467.550000 160.200000 480.000000 160.350000 ;
      RECT 467.550000 160.200000 480.000000 160.350000 ;
      RECT 467.685000 160.065000 480.000000 160.215000 ;
      RECT 467.700000 160.050000 480.000000 160.200000 ;
      RECT 467.700000 160.050000 480.000000 160.200000 ;
      RECT 467.835000 159.915000 480.000000 160.065000 ;
      RECT 467.850000 159.900000 480.000000 160.050000 ;
      RECT 467.850000 159.900000 480.000000 160.050000 ;
      RECT 467.985000 159.765000 480.000000 159.915000 ;
      RECT 468.000000 159.750000 480.000000 159.900000 ;
      RECT 468.000000 159.750000 480.000000 159.900000 ;
      RECT 468.135000 159.615000 480.000000 159.765000 ;
      RECT 468.150000 159.600000 480.000000 159.750000 ;
      RECT 468.150000 159.600000 480.000000 159.750000 ;
      RECT 468.285000 159.465000 480.000000 159.615000 ;
      RECT 468.300000 159.450000 480.000000 159.600000 ;
      RECT 468.300000 159.450000 480.000000 159.600000 ;
      RECT 468.435000 159.315000 480.000000 159.465000 ;
      RECT 468.450000 159.300000 480.000000 159.450000 ;
      RECT 468.450000 159.300000 480.000000 159.450000 ;
      RECT 468.585000 159.165000 480.000000 159.315000 ;
      RECT 468.600000 159.150000 480.000000 159.300000 ;
      RECT 468.600000 159.150000 480.000000 159.300000 ;
      RECT 468.735000 159.015000 480.000000 159.165000 ;
      RECT 468.750000 159.000000 480.000000 159.150000 ;
      RECT 468.750000 159.000000 480.000000 159.150000 ;
      RECT 468.885000 158.865000 480.000000 159.015000 ;
      RECT 468.900000 158.850000 480.000000 159.000000 ;
      RECT 468.900000 158.850000 480.000000 159.000000 ;
      RECT 469.035000 158.715000 480.000000 158.865000 ;
      RECT 469.050000 158.700000 480.000000 158.850000 ;
      RECT 469.050000 158.700000 480.000000 158.850000 ;
      RECT 469.185000 158.565000 480.000000 158.715000 ;
      RECT 469.200000 158.550000 480.000000 158.700000 ;
      RECT 469.200000 158.550000 480.000000 158.700000 ;
      RECT 469.335000 158.415000 480.000000 158.565000 ;
      RECT 469.350000 158.400000 480.000000 158.550000 ;
      RECT 469.350000 158.400000 480.000000 158.550000 ;
      RECT 469.485000 158.265000 480.000000 158.415000 ;
      RECT 469.500000 158.250000 480.000000 158.400000 ;
      RECT 469.500000 158.250000 480.000000 158.400000 ;
      RECT 469.635000 158.115000 480.000000 158.265000 ;
      RECT 469.650000 158.100000 480.000000 158.250000 ;
      RECT 469.650000 158.100000 480.000000 158.250000 ;
      RECT 469.785000 157.965000 480.000000 158.115000 ;
      RECT 469.800000 157.950000 480.000000 158.100000 ;
      RECT 469.800000 157.950000 480.000000 158.100000 ;
      RECT 469.935000 157.815000 480.000000 157.965000 ;
      RECT 469.950000 157.800000 480.000000 157.950000 ;
      RECT 469.950000 157.800000 480.000000 157.950000 ;
      RECT 470.085000 157.665000 480.000000 157.815000 ;
      RECT 470.100000 157.650000 480.000000 157.800000 ;
      RECT 470.100000 157.650000 480.000000 157.800000 ;
      RECT 470.235000 157.515000 480.000000 157.665000 ;
      RECT 470.250000 157.500000 480.000000 157.650000 ;
      RECT 470.250000 157.500000 480.000000 157.650000 ;
      RECT 470.385000 157.365000 480.000000 157.515000 ;
      RECT 470.400000 157.350000 480.000000 157.500000 ;
      RECT 470.400000 157.350000 480.000000 157.500000 ;
      RECT 470.535000 157.215000 480.000000 157.365000 ;
      RECT 470.550000 157.200000 480.000000 157.350000 ;
      RECT 470.550000 157.200000 480.000000 157.350000 ;
      RECT 470.685000 157.065000 480.000000 157.215000 ;
      RECT 470.700000 157.050000 480.000000 157.200000 ;
      RECT 470.700000 157.050000 480.000000 157.200000 ;
      RECT 470.835000 156.915000 480.000000 157.065000 ;
      RECT 470.850000 156.900000 480.000000 157.050000 ;
      RECT 470.850000 156.900000 480.000000 157.050000 ;
      RECT 470.985000 156.765000 480.000000 156.915000 ;
      RECT 471.000000 156.750000 480.000000 156.900000 ;
      RECT 471.000000 156.750000 480.000000 156.900000 ;
      RECT 471.135000 156.615000 480.000000 156.765000 ;
      RECT 471.150000 156.600000 480.000000 156.750000 ;
      RECT 471.150000 156.600000 480.000000 156.750000 ;
      RECT 471.285000 156.465000 480.000000 156.615000 ;
      RECT 471.300000 156.450000 480.000000 156.600000 ;
      RECT 471.300000 156.450000 480.000000 156.600000 ;
      RECT 471.435000 156.315000 480.000000 156.465000 ;
      RECT 471.450000 156.300000 480.000000 156.450000 ;
      RECT 471.450000 156.300000 480.000000 156.450000 ;
      RECT 471.585000 156.165000 480.000000 156.315000 ;
      RECT 471.600000 156.150000 480.000000 156.300000 ;
      RECT 471.600000 156.150000 480.000000 156.300000 ;
      RECT 471.735000 156.015000 480.000000 156.165000 ;
      RECT 471.750000 156.000000 480.000000 156.150000 ;
      RECT 471.750000 156.000000 480.000000 156.150000 ;
      RECT 471.885000 155.865000 480.000000 156.015000 ;
      RECT 471.900000 155.850000 480.000000 156.000000 ;
      RECT 471.900000 155.850000 480.000000 156.000000 ;
      RECT 472.035000 155.715000 480.000000 155.865000 ;
      RECT 472.050000 155.700000 480.000000 155.850000 ;
      RECT 472.050000 155.700000 480.000000 155.850000 ;
      RECT 472.185000 155.565000 480.000000 155.715000 ;
      RECT 472.200000 155.550000 480.000000 155.700000 ;
      RECT 472.200000 155.550000 480.000000 155.700000 ;
      RECT 472.335000 155.415000 480.000000 155.565000 ;
      RECT 472.350000 155.400000 480.000000 155.550000 ;
      RECT 472.350000 155.400000 480.000000 155.550000 ;
      RECT 472.485000 155.265000 480.000000 155.415000 ;
      RECT 472.500000 155.250000 480.000000 155.400000 ;
      RECT 472.500000 155.250000 480.000000 155.400000 ;
      RECT 472.635000 155.115000 480.000000 155.265000 ;
      RECT 472.650000 155.100000 480.000000 155.250000 ;
      RECT 472.650000 155.100000 480.000000 155.250000 ;
      RECT 472.785000 154.965000 480.000000 155.115000 ;
      RECT 472.800000 154.950000 480.000000 155.100000 ;
      RECT 472.800000 154.950000 480.000000 155.100000 ;
      RECT 472.935000 154.815000 480.000000 154.965000 ;
      RECT 472.950000 154.800000 480.000000 154.950000 ;
      RECT 472.950000 154.800000 480.000000 154.950000 ;
      RECT 473.085000 154.665000 480.000000 154.815000 ;
      RECT 473.100000 154.650000 480.000000 154.800000 ;
      RECT 473.100000 154.650000 480.000000 154.800000 ;
      RECT 473.235000 154.515000 480.000000 154.665000 ;
      RECT 473.250000 154.500000 480.000000 154.650000 ;
      RECT 473.250000 154.500000 480.000000 154.650000 ;
      RECT 473.385000 154.365000 480.000000 154.515000 ;
      RECT 473.400000 154.350000 480.000000 154.500000 ;
      RECT 473.400000 154.350000 480.000000 154.500000 ;
      RECT 473.535000 154.215000 480.000000 154.365000 ;
      RECT 473.550000 154.200000 480.000000 154.350000 ;
      RECT 473.550000 154.200000 480.000000 154.350000 ;
      RECT 473.685000 154.065000 480.000000 154.215000 ;
      RECT 473.700000 154.050000 480.000000 154.200000 ;
      RECT 473.700000 154.050000 480.000000 154.200000 ;
      RECT 473.835000 153.915000 480.000000 154.065000 ;
      RECT 473.850000 153.900000 480.000000 154.050000 ;
      RECT 473.850000 153.900000 480.000000 154.050000 ;
      RECT 473.985000 153.765000 480.000000 153.915000 ;
      RECT 474.000000 153.750000 480.000000 153.900000 ;
      RECT 474.000000 153.750000 480.000000 153.900000 ;
      RECT 474.135000 153.615000 480.000000 153.765000 ;
      RECT 474.150000 153.600000 480.000000 153.750000 ;
      RECT 474.150000 153.600000 480.000000 153.750000 ;
      RECT 474.285000 153.465000 480.000000 153.615000 ;
      RECT 474.300000 153.450000 480.000000 153.600000 ;
      RECT 474.300000 153.450000 480.000000 153.600000 ;
      RECT 474.435000 153.315000 480.000000 153.465000 ;
      RECT 474.450000 153.300000 480.000000 153.450000 ;
      RECT 474.450000 153.300000 480.000000 153.450000 ;
      RECT 474.585000 153.165000 480.000000 153.315000 ;
      RECT 474.600000 153.150000 480.000000 153.300000 ;
      RECT 474.600000 153.150000 480.000000 153.300000 ;
      RECT 474.735000 153.015000 480.000000 153.165000 ;
      RECT 474.750000 153.000000 480.000000 153.150000 ;
      RECT 474.750000 153.000000 480.000000 153.150000 ;
      RECT 474.885000 152.865000 480.000000 153.015000 ;
      RECT 474.900000 152.850000 480.000000 153.000000 ;
      RECT 474.900000 152.850000 480.000000 153.000000 ;
      RECT 475.035000 152.715000 480.000000 152.865000 ;
      RECT 475.050000 152.700000 480.000000 152.850000 ;
      RECT 475.050000 152.700000 480.000000 152.850000 ;
      RECT 475.185000 152.565000 480.000000 152.715000 ;
      RECT 475.200000 152.550000 480.000000 152.700000 ;
      RECT 475.200000 152.550000 480.000000 152.700000 ;
      RECT 475.335000 152.415000 480.000000 152.565000 ;
      RECT 475.350000 152.400000 480.000000 152.550000 ;
      RECT 475.350000 152.400000 480.000000 152.550000 ;
      RECT 475.485000 152.265000 480.000000 152.415000 ;
      RECT 475.500000 152.250000 480.000000 152.400000 ;
      RECT 475.500000 152.250000 480.000000 152.400000 ;
      RECT 475.635000 152.115000 480.000000 152.265000 ;
      RECT 475.650000 152.100000 480.000000 152.250000 ;
      RECT 475.650000 152.100000 480.000000 152.250000 ;
      RECT 475.785000 151.965000 480.000000 152.115000 ;
      RECT 475.800000 151.950000 480.000000 152.100000 ;
      RECT 475.800000 151.950000 480.000000 152.100000 ;
      RECT 475.935000 151.815000 480.000000 151.965000 ;
      RECT 475.950000 151.800000 480.000000 151.950000 ;
      RECT 475.950000 151.800000 480.000000 151.950000 ;
      RECT 476.085000 151.665000 480.000000 151.815000 ;
      RECT 476.100000 151.650000 480.000000 151.800000 ;
      RECT 476.100000 151.650000 480.000000 151.800000 ;
      RECT 476.235000 151.515000 480.000000 151.665000 ;
      RECT 476.250000 151.500000 480.000000 151.650000 ;
      RECT 476.250000 151.500000 480.000000 151.650000 ;
      RECT 476.385000 151.365000 480.000000 151.515000 ;
      RECT 476.400000 151.350000 480.000000 151.500000 ;
      RECT 476.400000 151.350000 480.000000 151.500000 ;
      RECT 476.535000 151.215000 480.000000 151.365000 ;
      RECT 476.550000 151.200000 480.000000 151.350000 ;
      RECT 476.550000 151.200000 480.000000 151.350000 ;
      RECT 476.685000 151.065000 480.000000 151.215000 ;
      RECT 476.700000 151.050000 480.000000 151.200000 ;
      RECT 476.700000 151.050000 480.000000 151.200000 ;
      RECT 476.835000 150.915000 480.000000 151.065000 ;
      RECT 476.850000 150.900000 480.000000 151.050000 ;
      RECT 476.850000 150.900000 480.000000 151.050000 ;
      RECT 476.985000 150.765000 480.000000 150.915000 ;
      RECT 477.000000 150.750000 480.000000 150.900000 ;
      RECT 477.000000 150.750000 480.000000 150.900000 ;
      RECT 477.135000 150.615000 480.000000 150.765000 ;
      RECT 477.150000 150.600000 480.000000 150.750000 ;
      RECT 477.150000 150.600000 480.000000 150.750000 ;
      RECT 477.285000 150.465000 480.000000 150.615000 ;
      RECT 477.300000 150.450000 480.000000 150.600000 ;
      RECT 477.300000 150.450000 480.000000 150.600000 ;
      RECT 477.435000 150.315000 480.000000 150.465000 ;
      RECT 477.450000 150.300000 480.000000 150.450000 ;
      RECT 477.450000 150.300000 480.000000 150.450000 ;
      RECT 477.585000 150.165000 480.000000 150.315000 ;
      RECT 477.600000 150.150000 480.000000 150.300000 ;
      RECT 477.600000 150.150000 480.000000 150.300000 ;
      RECT 477.735000 150.015000 480.000000 150.165000 ;
      RECT 477.750000 150.000000 480.000000 150.150000 ;
      RECT 477.750000 150.000000 480.000000 150.150000 ;
      RECT 477.885000 149.865000 480.000000 150.015000 ;
      RECT 477.900000 149.850000 480.000000 150.000000 ;
      RECT 477.900000 149.850000 480.000000 150.000000 ;
      RECT 478.035000 149.715000 480.000000 149.865000 ;
      RECT 478.050000 149.700000 480.000000 149.850000 ;
      RECT 478.050000 149.700000 480.000000 149.850000 ;
      RECT 478.185000 149.565000 480.000000 149.715000 ;
      RECT 478.200000 149.550000 480.000000 149.700000 ;
      RECT 478.200000 149.550000 480.000000 149.700000 ;
      RECT 478.335000 149.415000 480.000000 149.565000 ;
      RECT 478.350000 149.400000 480.000000 149.550000 ;
      RECT 478.350000 149.400000 480.000000 149.550000 ;
      RECT 478.485000 149.265000 480.000000 149.415000 ;
      RECT 478.500000 149.250000 480.000000 149.400000 ;
      RECT 478.500000 149.250000 480.000000 149.400000 ;
      RECT 478.595000 149.015000 480.000000 228.200000 ;
      RECT 478.635000 149.115000 480.000000 149.265000 ;
      RECT 478.650000 149.100000 480.000000 149.250000 ;
      RECT 478.650000 149.100000 480.000000 149.250000 ;
      RECT 478.800000 148.950000 480.000000 149.100000 ;
      RECT 478.800000 148.950000 480.000000 149.100000 ;
      RECT 478.950000 148.800000 480.000000 148.950000 ;
      RECT 478.950000 148.800000 480.000000 148.950000 ;
      RECT 479.100000 148.650000 480.000000 148.800000 ;
      RECT 479.100000 148.650000 480.000000 148.800000 ;
      RECT 479.250000 148.500000 480.000000 148.650000 ;
      RECT 479.250000 148.500000 480.000000 148.650000 ;
      RECT 479.400000 148.350000 480.000000 148.500000 ;
      RECT 479.400000 148.350000 480.000000 148.500000 ;
      RECT 479.550000 148.200000 480.000000 148.350000 ;
      RECT 479.550000 148.200000 480.000000 148.350000 ;
      RECT 479.700000 148.050000 480.000000 148.200000 ;
      RECT 479.700000 148.050000 480.000000 148.200000 ;
      RECT 479.850000 147.900000 480.000000 148.050000 ;
      RECT 479.850000 147.900000 480.000000 148.050000 ;
    LAYER met5 ;
      RECT   0.000000   0.000000 480.000000  55.050000 ;
      RECT   0.000000   0.000000 480.000000  55.050000 ;
      RECT   0.000000 149.515000  18.260000 149.915000 ;
      RECT   0.000000 149.515000  28.460000 159.715000 ;
      RECT   0.000000 149.915000  18.660000 150.315000 ;
      RECT   0.000000 150.315000  19.060000 150.715000 ;
      RECT   0.000000 150.715000  19.460000 151.115000 ;
      RECT   0.000000 151.115000  19.860000 151.515000 ;
      RECT   0.000000 151.515000  20.260000 151.915000 ;
      RECT   0.000000 151.915000  20.660000 152.315000 ;
      RECT   0.000000 152.315000  21.060000 152.715000 ;
      RECT   0.000000 152.715000  21.460000 153.115000 ;
      RECT   0.000000 153.115000  21.860000 153.515000 ;
      RECT   0.000000 153.515000  22.260000 153.915000 ;
      RECT   0.000000 153.915000  22.660000 154.315000 ;
      RECT   0.000000 154.315000  23.060000 154.715000 ;
      RECT   0.000000 154.715000  23.460000 155.115000 ;
      RECT   0.000000 155.115000  23.860000 155.515000 ;
      RECT   0.000000 155.515000  24.260000 155.915000 ;
      RECT   0.000000 155.915000  24.660000 156.315000 ;
      RECT   0.000000 156.315000  25.060000 156.715000 ;
      RECT   0.000000 156.715000  25.460000 157.115000 ;
      RECT   0.000000 157.115000  25.860000 157.515000 ;
      RECT   0.000000 157.515000  26.260000 157.915000 ;
      RECT   0.000000 157.915000  26.660000 158.315000 ;
      RECT   0.000000 158.315000  27.060000 158.715000 ;
      RECT   0.000000 158.715000  27.460000 159.115000 ;
      RECT   0.000000 159.115000  27.860000 159.515000 ;
      RECT   0.000000 159.515000  28.260000 159.715000 ;
      RECT   0.000000 159.715000  28.460000 207.655000 ;
      RECT   0.000000 159.715000  28.460000 207.655000 ;
      RECT   0.000000 207.655000  28.460000 208.055000 ;
      RECT   0.000000 207.655000  49.505000 228.700000 ;
      RECT   0.000000 208.055000  28.860000 208.455000 ;
      RECT   0.000000 208.455000  29.260000 208.855000 ;
      RECT   0.000000 208.855000  29.660000 209.255000 ;
      RECT   0.000000 209.255000  30.060000 209.655000 ;
      RECT   0.000000 209.655000  30.460000 210.055000 ;
      RECT   0.000000 210.055000  30.860000 210.455000 ;
      RECT   0.000000 210.455000  31.260000 210.855000 ;
      RECT   0.000000 210.855000  31.660000 211.255000 ;
      RECT   0.000000 211.255000  32.060000 211.655000 ;
      RECT   0.000000 211.655000  32.460000 212.055000 ;
      RECT   0.000000 212.055000  32.860000 212.455000 ;
      RECT   0.000000 212.455000  33.260000 212.855000 ;
      RECT   0.000000 212.855000  33.660000 213.255000 ;
      RECT   0.000000 213.255000  34.060000 213.655000 ;
      RECT   0.000000 213.655000  34.460000 214.055000 ;
      RECT   0.000000 214.055000  34.860000 214.455000 ;
      RECT   0.000000 214.455000  35.260000 214.855000 ;
      RECT   0.000000 214.855000  35.660000 215.255000 ;
      RECT   0.000000 215.255000  36.060000 215.655000 ;
      RECT   0.000000 215.655000  36.460000 216.055000 ;
      RECT   0.000000 216.055000  36.860000 216.455000 ;
      RECT   0.000000 216.455000  37.260000 216.855000 ;
      RECT   0.000000 216.855000  37.660000 217.255000 ;
      RECT   0.000000 217.255000  38.060000 217.655000 ;
      RECT   0.000000 217.655000  38.460000 218.055000 ;
      RECT   0.000000 218.055000  38.860000 218.455000 ;
      RECT   0.000000 218.455000  39.260000 218.855000 ;
      RECT   0.000000 218.855000  39.660000 219.255000 ;
      RECT   0.000000 219.255000  40.060000 219.655000 ;
      RECT   0.000000 219.655000  40.460000 220.055000 ;
      RECT   0.000000 220.055000  40.860000 220.455000 ;
      RECT   0.000000 220.455000  41.260000 220.855000 ;
      RECT   0.000000 220.855000  41.660000 221.255000 ;
      RECT   0.000000 221.255000  42.060000 221.655000 ;
      RECT   0.000000 221.655000  42.460000 222.055000 ;
      RECT   0.000000 222.055000  42.860000 222.455000 ;
      RECT   0.000000 222.455000  43.260000 222.855000 ;
      RECT   0.000000 222.855000  43.660000 223.255000 ;
      RECT   0.000000 223.255000  44.060000 223.655000 ;
      RECT   0.000000 223.655000  44.460000 224.055000 ;
      RECT   0.000000 224.055000  44.860000 224.455000 ;
      RECT   0.000000 224.455000  45.260000 224.855000 ;
      RECT   0.000000 224.855000  45.660000 225.255000 ;
      RECT   0.000000 225.255000  46.060000 225.655000 ;
      RECT   0.000000 225.655000  46.460000 226.055000 ;
      RECT   0.000000 226.055000  46.860000 226.455000 ;
      RECT   0.000000 226.455000  47.260000 226.855000 ;
      RECT   0.000000 226.855000  47.660000 227.255000 ;
      RECT   0.000000 227.255000  48.060000 227.655000 ;
      RECT   0.000000 227.655000  48.460000 228.055000 ;
      RECT   0.000000 228.055000  48.860000 228.455000 ;
      RECT   0.000000 228.455000  49.260000 228.700000 ;
      RECT  29.145000 122.950000 466.455000 124.875000 ;
      RECT  29.545000 122.950000 467.980000 123.350000 ;
      RECT  29.945000 123.350000 467.580000 123.750000 ;
      RECT  30.345000 123.750000 467.180000 124.150000 ;
      RECT  30.745000 124.150000 466.780000 124.550000 ;
      RECT  31.070000 124.550000 466.455000 124.875000 ;
      RECT  31.070000 124.875000 104.990000 131.875000 ;
      RECT  31.470000 124.875000 111.590000 125.275000 ;
      RECT  31.870000 125.275000 111.190000 125.675000 ;
      RECT  32.270000 125.675000 110.790000 126.075000 ;
      RECT  32.670000 126.075000 110.390000 126.475000 ;
      RECT  33.070000 126.475000 109.990000 126.875000 ;
      RECT  33.470000 126.875000 109.590000 127.275000 ;
      RECT  33.870000 127.275000 109.190000 127.675000 ;
      RECT  34.270000 127.675000 108.790000 128.075000 ;
      RECT  34.670000 128.075000 108.390000 128.475000 ;
      RECT  35.070000 128.475000 107.990000 128.875000 ;
      RECT  35.470000 128.875000 107.590000 129.275000 ;
      RECT  35.870000 129.275000 107.190000 129.675000 ;
      RECT  36.270000 129.675000 106.790000 130.075000 ;
      RECT  36.670000 130.075000 106.390000 130.475000 ;
      RECT  37.070000 130.475000 105.990000 130.875000 ;
      RECT  37.470000 130.875000 105.590000 131.275000 ;
      RECT  37.870000 131.275000 105.190000 131.675000 ;
      RECT  38.070000 131.675000 104.990000 131.875000 ;
      RECT  38.070000 131.875000 104.990000 132.550000 ;
      RECT  38.405000 131.875000 104.990000 132.210000 ;
      RECT  38.745000 132.210000 104.990000 132.550000 ;
      RECT  39.280000 132.550000 104.990000 133.085000 ;
      RECT  39.280000 132.550000 104.990000 133.085000 ;
      RECT  39.280000 133.085000 104.990000 145.105000 ;
      RECT  39.680000 133.085000 104.990000 133.485000 ;
      RECT  40.080000 133.485000 104.990000 133.885000 ;
      RECT  40.480000 133.885000 104.990000 134.285000 ;
      RECT  40.880000 134.285000 104.990000 134.685000 ;
      RECT  41.280000 134.685000 104.990000 135.085000 ;
      RECT  41.680000 135.085000 104.990000 135.485000 ;
      RECT  42.080000 135.485000 104.990000 135.885000 ;
      RECT  42.480000 135.885000 104.990000 136.285000 ;
      RECT  42.880000 136.285000 104.990000 136.685000 ;
      RECT  43.280000 136.685000 104.990000 137.085000 ;
      RECT  43.680000 137.085000 104.990000 137.485000 ;
      RECT  44.080000 137.485000 104.990000 137.885000 ;
      RECT  44.480000 137.885000 104.990000 138.285000 ;
      RECT  44.880000 138.285000 104.990000 138.685000 ;
      RECT  45.280000 138.685000 104.990000 139.085000 ;
      RECT  45.680000 139.085000 104.990000 139.485000 ;
      RECT  46.080000 139.485000 104.990000 139.885000 ;
      RECT  46.480000 139.885000 104.990000 140.285000 ;
      RECT  46.880000 140.285000 104.990000 140.685000 ;
      RECT  47.280000 140.685000 104.990000 141.085000 ;
      RECT  47.680000 141.085000 104.990000 141.485000 ;
      RECT  48.080000 141.485000 104.990000 141.885000 ;
      RECT  48.480000 141.885000 104.990000 142.285000 ;
      RECT  48.880000 142.285000 104.990000 142.685000 ;
      RECT  49.280000 142.685000 104.990000 143.085000 ;
      RECT  49.680000 143.085000 104.990000 143.485000 ;
      RECT  50.080000 143.485000 104.990000 143.885000 ;
      RECT  50.480000 143.885000 104.990000 144.285000 ;
      RECT  50.880000 144.285000 104.990000 144.685000 ;
      RECT  51.280000 144.685000 104.990000 145.085000 ;
      RECT  51.300000 145.085000 104.990000 145.105000 ;
      RECT  51.790000 145.105000 104.990000 145.595000 ;
      RECT  51.790000 145.105000 104.990000 145.595000 ;
      RECT  51.790000 145.595000 104.990000 148.750000 ;
      RECT  52.190000 145.595000 104.990000 145.995000 ;
      RECT  52.590000 145.995000 104.990000 146.395000 ;
      RECT  52.990000 146.395000 104.990000 146.795000 ;
      RECT  53.390000 146.795000 104.990000 147.195000 ;
      RECT  53.790000 147.195000 104.990000 147.595000 ;
      RECT  54.190000 147.595000 104.990000 147.995000 ;
      RECT  54.590000 147.995000 104.990000 148.395000 ;
      RECT  54.945000 148.395000 104.990000 148.750000 ;
      RECT  54.945000 148.750000 104.990000 194.875000 ;
      RECT  54.945000 148.750000 104.990000 194.875000 ;
      RECT  54.945000 194.875000 104.990000 195.275000 ;
      RECT  54.945000 194.875000 107.380000 197.270000 ;
      RECT  54.945000 195.275000 105.390000 195.675000 ;
      RECT  54.945000 195.675000 105.790000 196.075000 ;
      RECT  54.945000 196.075000 106.190000 196.475000 ;
      RECT  54.945000 196.475000 106.590000 196.875000 ;
      RECT  54.945000 196.875000 106.990000 197.270000 ;
      RECT  54.945000 197.270000 111.990000 201.875000 ;
      RECT  55.345000 197.270000 107.380000 197.670000 ;
      RECT  55.745000 197.670000 107.785000 198.070000 ;
      RECT  56.145000 198.070000 108.185000 198.470000 ;
      RECT  56.545000 198.470000 108.585000 198.870000 ;
      RECT  56.945000 198.870000 108.985000 199.270000 ;
      RECT  57.345000 199.270000 109.385000 199.670000 ;
      RECT  57.745000 199.670000 109.785000 200.070000 ;
      RECT  58.145000 200.070000 110.185000 200.470000 ;
      RECT  58.545000 200.470000 110.585000 200.870000 ;
      RECT  58.945000 200.870000 110.985000 201.270000 ;
      RECT  59.345000 201.270000 111.385000 201.670000 ;
      RECT  59.550000 201.670000 111.785000 201.875000 ;
      RECT  59.550000 201.875000 387.640000 203.690000 ;
      RECT  59.950000 201.875000 389.055000 202.275000 ;
      RECT  60.350000 202.275000 388.655000 202.675000 ;
      RECT  60.750000 202.675000 388.255000 203.075000 ;
      RECT  61.150000 203.075000 387.855000 203.475000 ;
      RECT  61.365000 203.475000 387.640000 203.690000 ;
      RECT 164.990000 124.875000 218.015000 131.875000 ;
      RECT 165.190000 201.675000 224.815000 201.875000 ;
      RECT 165.390000 124.875000 224.615000 125.275000 ;
      RECT 165.590000 201.275000 224.415000 201.675000 ;
      RECT 165.790000 125.275000 224.215000 125.675000 ;
      RECT 165.990000 200.875000 224.015000 201.275000 ;
      RECT 166.190000 125.675000 223.815000 126.075000 ;
      RECT 166.390000 200.475000 223.615000 200.875000 ;
      RECT 166.590000 126.075000 223.415000 126.475000 ;
      RECT 166.790000 200.075000 223.215000 200.475000 ;
      RECT 166.990000 126.475000 223.015000 126.875000 ;
      RECT 167.190000 199.675000 222.815000 200.075000 ;
      RECT 167.390000 126.875000 222.615000 127.275000 ;
      RECT 167.590000 199.275000 222.415000 199.675000 ;
      RECT 167.790000 127.275000 222.215000 127.675000 ;
      RECT 167.990000 198.875000 222.015000 199.275000 ;
      RECT 168.190000 127.675000 221.815000 128.075000 ;
      RECT 168.390000 198.475000 221.615000 198.875000 ;
      RECT 168.590000 128.075000 221.415000 128.475000 ;
      RECT 168.790000 198.075000 221.215000 198.475000 ;
      RECT 168.990000 128.475000 221.015000 128.875000 ;
      RECT 169.190000 197.675000 220.815000 198.075000 ;
      RECT 169.390000 128.875000 220.615000 129.275000 ;
      RECT 169.590000 197.275000 220.415000 197.675000 ;
      RECT 169.790000 129.275000 220.215000 129.675000 ;
      RECT 169.990000 196.875000 220.015000 197.275000 ;
      RECT 170.190000 129.675000 219.815000 130.075000 ;
      RECT 170.390000 196.475000 219.615000 196.875000 ;
      RECT 170.590000 130.075000 219.415000 130.475000 ;
      RECT 170.790000 196.075000 219.215000 196.475000 ;
      RECT 170.990000 130.475000 219.015000 130.875000 ;
      RECT 171.190000 195.675000 218.815000 196.075000 ;
      RECT 171.390000 130.875000 218.615000 131.275000 ;
      RECT 171.590000 195.275000 218.415000 195.675000 ;
      RECT 171.790000 131.275000 218.215000 131.675000 ;
      RECT 171.990000 131.675000 218.015000 131.875000 ;
      RECT 171.990000 131.875000 218.015000 194.875000 ;
      RECT 171.990000 131.875000 218.015000 194.875000 ;
      RECT 171.990000 194.875000 218.015000 195.275000 ;
      RECT 171.990000 194.875000 225.015000 201.875000 ;
      RECT 278.015000 124.875000 459.455000 131.875000 ;
      RECT 278.215000 201.675000 389.455000 201.875000 ;
      RECT 278.415000 124.875000 466.055000 125.275000 ;
      RECT 278.615000 201.275000 389.655000 201.675000 ;
      RECT 278.815000 125.275000 465.655000 125.675000 ;
      RECT 279.015000 200.875000 390.055000 201.275000 ;
      RECT 279.215000 125.675000 465.255000 126.075000 ;
      RECT 279.415000 200.475000 390.455000 200.875000 ;
      RECT 279.615000 126.075000 464.855000 126.475000 ;
      RECT 279.815000 200.075000 390.855000 200.475000 ;
      RECT 280.015000 126.475000 464.455000 126.875000 ;
      RECT 280.215000 199.675000 391.255000 200.075000 ;
      RECT 280.415000 126.875000 464.055000 127.275000 ;
      RECT 280.615000 199.275000 391.655000 199.675000 ;
      RECT 280.815000 127.275000 463.655000 127.675000 ;
      RECT 281.015000 198.875000 392.055000 199.275000 ;
      RECT 281.215000 127.675000 463.255000 128.075000 ;
      RECT 281.415000 198.475000 392.455000 198.875000 ;
      RECT 281.615000 128.075000 462.855000 128.475000 ;
      RECT 281.815000 198.075000 392.855000 198.475000 ;
      RECT 282.015000 128.475000 462.455000 128.875000 ;
      RECT 282.215000 197.675000 393.255000 198.075000 ;
      RECT 282.415000 128.875000 462.055000 129.275000 ;
      RECT 282.615000 197.275000 393.655000 197.675000 ;
      RECT 282.815000 129.275000 461.655000 129.675000 ;
      RECT 283.015000 196.875000 394.055000 197.275000 ;
      RECT 283.215000 129.675000 461.255000 130.075000 ;
      RECT 283.415000 196.475000 394.455000 196.875000 ;
      RECT 283.615000 130.075000 460.855000 130.475000 ;
      RECT 283.815000 196.075000 394.855000 196.475000 ;
      RECT 284.015000 130.475000 460.455000 130.875000 ;
      RECT 284.215000 195.675000 395.255000 196.075000 ;
      RECT 284.415000 130.875000 460.055000 131.275000 ;
      RECT 284.615000 195.275000 395.655000 195.675000 ;
      RECT 284.815000 131.275000 459.655000 131.675000 ;
      RECT 285.015000 131.675000 459.455000 131.875000 ;
      RECT 285.015000 131.875000 446.620000 144.710000 ;
      RECT 285.015000 131.875000 459.055000 132.275000 ;
      RECT 285.015000 132.275000 458.655000 132.675000 ;
      RECT 285.015000 132.675000 458.255000 133.075000 ;
      RECT 285.015000 133.075000 457.855000 133.475000 ;
      RECT 285.015000 133.475000 457.455000 133.875000 ;
      RECT 285.015000 133.875000 457.055000 134.275000 ;
      RECT 285.015000 134.275000 456.655000 134.675000 ;
      RECT 285.015000 134.675000 456.255000 135.075000 ;
      RECT 285.015000 135.075000 455.855000 135.475000 ;
      RECT 285.015000 135.475000 455.455000 135.875000 ;
      RECT 285.015000 135.875000 455.055000 136.275000 ;
      RECT 285.015000 136.275000 454.655000 136.675000 ;
      RECT 285.015000 136.675000 454.255000 137.075000 ;
      RECT 285.015000 137.075000 453.855000 137.475000 ;
      RECT 285.015000 137.475000 453.455000 137.875000 ;
      RECT 285.015000 137.875000 453.055000 138.275000 ;
      RECT 285.015000 138.275000 452.655000 138.675000 ;
      RECT 285.015000 138.675000 452.255000 139.075000 ;
      RECT 285.015000 139.075000 451.855000 139.475000 ;
      RECT 285.015000 139.475000 451.455000 139.875000 ;
      RECT 285.015000 139.875000 451.055000 140.275000 ;
      RECT 285.015000 140.275000 450.655000 140.675000 ;
      RECT 285.015000 140.675000 450.255000 141.075000 ;
      RECT 285.015000 141.075000 449.855000 141.475000 ;
      RECT 285.015000 141.475000 449.455000 141.875000 ;
      RECT 285.015000 141.875000 449.055000 142.275000 ;
      RECT 285.015000 142.275000 448.655000 142.675000 ;
      RECT 285.015000 142.675000 448.255000 143.075000 ;
      RECT 285.015000 143.075000 447.855000 143.475000 ;
      RECT 285.015000 143.475000 447.455000 143.875000 ;
      RECT 285.015000 143.875000 447.055000 144.275000 ;
      RECT 285.015000 144.275000 446.655000 144.675000 ;
      RECT 285.015000 144.675000 446.620000 144.710000 ;
      RECT 285.015000 144.710000 446.090000 145.240000 ;
      RECT 285.015000 144.710000 446.090000 145.240000 ;
      RECT 285.015000 145.240000 440.380000 150.950000 ;
      RECT 285.015000 145.240000 445.690000 145.640000 ;
      RECT 285.015000 145.640000 445.290000 146.040000 ;
      RECT 285.015000 146.040000 444.890000 146.440000 ;
      RECT 285.015000 146.440000 444.490000 146.840000 ;
      RECT 285.015000 146.840000 444.090000 147.240000 ;
      RECT 285.015000 147.240000 443.690000 147.640000 ;
      RECT 285.015000 147.640000 443.290000 148.040000 ;
      RECT 285.015000 148.040000 442.890000 148.440000 ;
      RECT 285.015000 148.440000 442.490000 148.840000 ;
      RECT 285.015000 148.840000 442.090000 149.240000 ;
      RECT 285.015000 149.240000 441.690000 149.640000 ;
      RECT 285.015000 149.640000 441.290000 150.040000 ;
      RECT 285.015000 150.040000 440.890000 150.440000 ;
      RECT 285.015000 150.440000 440.490000 150.840000 ;
      RECT 285.015000 150.840000 440.380000 150.950000 ;
      RECT 285.015000 150.950000 439.890000 151.440000 ;
      RECT 285.015000 150.950000 439.890000 151.440000 ;
      RECT 285.015000 151.440000 396.455000 194.875000 ;
      RECT 285.015000 151.440000 439.490000 151.840000 ;
      RECT 285.015000 151.840000 439.090000 152.240000 ;
      RECT 285.015000 152.240000 438.690000 152.640000 ;
      RECT 285.015000 152.640000 438.290000 153.040000 ;
      RECT 285.015000 153.040000 437.890000 153.440000 ;
      RECT 285.015000 153.440000 437.490000 153.840000 ;
      RECT 285.015000 153.840000 437.090000 154.240000 ;
      RECT 285.015000 154.240000 436.690000 154.640000 ;
      RECT 285.015000 154.640000 436.290000 155.040000 ;
      RECT 285.015000 155.040000 435.890000 155.440000 ;
      RECT 285.015000 155.440000 435.490000 155.840000 ;
      RECT 285.015000 155.840000 435.090000 156.240000 ;
      RECT 285.015000 156.240000 434.690000 156.640000 ;
      RECT 285.015000 156.640000 434.290000 157.040000 ;
      RECT 285.015000 157.040000 433.890000 157.440000 ;
      RECT 285.015000 157.440000 433.490000 157.840000 ;
      RECT 285.015000 157.840000 433.090000 158.240000 ;
      RECT 285.015000 158.240000 432.690000 158.640000 ;
      RECT 285.015000 158.640000 432.290000 159.040000 ;
      RECT 285.015000 159.040000 431.890000 159.440000 ;
      RECT 285.015000 159.440000 431.490000 159.840000 ;
      RECT 285.015000 159.840000 431.090000 160.240000 ;
      RECT 285.015000 160.240000 430.690000 160.640000 ;
      RECT 285.015000 160.640000 430.290000 161.040000 ;
      RECT 285.015000 161.040000 429.890000 161.440000 ;
      RECT 285.015000 161.440000 429.490000 161.840000 ;
      RECT 285.015000 161.840000 429.090000 162.240000 ;
      RECT 285.015000 162.240000 428.690000 162.640000 ;
      RECT 285.015000 162.640000 428.290000 163.040000 ;
      RECT 285.015000 163.040000 427.890000 163.440000 ;
      RECT 285.015000 163.440000 427.490000 163.840000 ;
      RECT 285.015000 163.840000 427.090000 164.240000 ;
      RECT 285.015000 164.240000 426.690000 164.640000 ;
      RECT 285.015000 164.640000 426.290000 165.040000 ;
      RECT 285.015000 165.040000 425.890000 165.440000 ;
      RECT 285.015000 165.440000 425.490000 165.840000 ;
      RECT 285.015000 165.840000 425.090000 166.240000 ;
      RECT 285.015000 166.240000 424.690000 166.640000 ;
      RECT 285.015000 166.640000 424.290000 167.040000 ;
      RECT 285.015000 167.040000 423.890000 167.440000 ;
      RECT 285.015000 167.440000 423.490000 167.840000 ;
      RECT 285.015000 167.840000 423.090000 168.240000 ;
      RECT 285.015000 168.240000 422.690000 168.640000 ;
      RECT 285.015000 168.640000 422.290000 169.040000 ;
      RECT 285.015000 169.040000 421.890000 169.440000 ;
      RECT 285.015000 169.440000 421.490000 169.840000 ;
      RECT 285.015000 169.840000 421.090000 170.240000 ;
      RECT 285.015000 170.240000 420.690000 170.640000 ;
      RECT 285.015000 170.640000 420.290000 171.040000 ;
      RECT 285.015000 171.040000 419.890000 171.440000 ;
      RECT 285.015000 171.440000 419.490000 171.840000 ;
      RECT 285.015000 171.840000 419.090000 172.240000 ;
      RECT 285.015000 172.240000 418.690000 172.640000 ;
      RECT 285.015000 172.640000 418.290000 173.040000 ;
      RECT 285.015000 173.040000 417.890000 173.440000 ;
      RECT 285.015000 173.440000 417.490000 173.840000 ;
      RECT 285.015000 173.840000 417.090000 174.240000 ;
      RECT 285.015000 174.240000 416.690000 174.640000 ;
      RECT 285.015000 174.640000 416.290000 175.040000 ;
      RECT 285.015000 175.040000 415.890000 175.440000 ;
      RECT 285.015000 175.440000 415.490000 175.840000 ;
      RECT 285.015000 175.840000 415.090000 176.240000 ;
      RECT 285.015000 176.240000 414.690000 176.640000 ;
      RECT 285.015000 176.640000 414.290000 177.040000 ;
      RECT 285.015000 177.040000 413.890000 177.440000 ;
      RECT 285.015000 177.440000 413.490000 177.840000 ;
      RECT 285.015000 177.840000 413.090000 178.240000 ;
      RECT 285.015000 178.240000 412.690000 178.640000 ;
      RECT 285.015000 178.640000 412.290000 179.040000 ;
      RECT 285.015000 179.040000 411.890000 179.440000 ;
      RECT 285.015000 179.440000 411.490000 179.840000 ;
      RECT 285.015000 179.840000 411.090000 180.240000 ;
      RECT 285.015000 180.240000 410.690000 180.640000 ;
      RECT 285.015000 180.640000 410.290000 181.040000 ;
      RECT 285.015000 181.040000 409.890000 181.440000 ;
      RECT 285.015000 181.440000 409.490000 181.840000 ;
      RECT 285.015000 181.840000 409.090000 182.240000 ;
      RECT 285.015000 182.240000 408.690000 182.640000 ;
      RECT 285.015000 182.640000 408.290000 183.040000 ;
      RECT 285.015000 183.040000 407.890000 183.440000 ;
      RECT 285.015000 183.440000 407.490000 183.840000 ;
      RECT 285.015000 183.840000 407.090000 184.240000 ;
      RECT 285.015000 184.240000 406.690000 184.640000 ;
      RECT 285.015000 184.640000 406.290000 185.040000 ;
      RECT 285.015000 185.040000 405.890000 185.440000 ;
      RECT 285.015000 185.440000 405.490000 185.840000 ;
      RECT 285.015000 185.840000 405.090000 186.240000 ;
      RECT 285.015000 186.240000 404.690000 186.640000 ;
      RECT 285.015000 186.640000 404.290000 187.040000 ;
      RECT 285.015000 187.040000 403.890000 187.440000 ;
      RECT 285.015000 187.440000 403.490000 187.840000 ;
      RECT 285.015000 187.840000 403.090000 188.240000 ;
      RECT 285.015000 188.240000 402.690000 188.640000 ;
      RECT 285.015000 188.640000 402.290000 189.040000 ;
      RECT 285.015000 189.040000 401.890000 189.440000 ;
      RECT 285.015000 189.440000 401.490000 189.840000 ;
      RECT 285.015000 189.840000 401.090000 190.240000 ;
      RECT 285.015000 190.240000 400.690000 190.640000 ;
      RECT 285.015000 190.640000 400.290000 191.040000 ;
      RECT 285.015000 191.040000 399.890000 191.440000 ;
      RECT 285.015000 191.440000 399.490000 191.840000 ;
      RECT 285.015000 191.840000 399.090000 192.240000 ;
      RECT 285.015000 192.240000 398.690000 192.640000 ;
      RECT 285.015000 192.640000 398.290000 193.040000 ;
      RECT 285.015000 193.040000 397.890000 193.440000 ;
      RECT 285.015000 193.440000 397.490000 193.840000 ;
      RECT 285.015000 193.840000 397.090000 194.240000 ;
      RECT 285.015000 194.240000 396.690000 194.640000 ;
      RECT 285.015000 194.640000 396.455000 194.875000 ;
      RECT 285.015000 194.875000 389.455000 201.875000 ;
      RECT 285.015000 194.875000 396.055000 195.275000 ;
      RECT 400.015000 228.300000 480.000000 228.700000 ;
      RECT 400.415000 227.900000 480.000000 228.300000 ;
      RECT 400.815000 227.500000 480.000000 227.900000 ;
      RECT 401.215000 227.100000 480.000000 227.500000 ;
      RECT 401.615000 226.700000 480.000000 227.100000 ;
      RECT 402.015000 226.300000 480.000000 226.700000 ;
      RECT 402.415000 225.900000 480.000000 226.300000 ;
      RECT 402.815000 225.500000 480.000000 225.900000 ;
      RECT 403.215000 225.100000 480.000000 225.500000 ;
      RECT 403.615000 224.700000 480.000000 225.100000 ;
      RECT 404.015000 224.300000 480.000000 224.700000 ;
      RECT 404.415000 223.900000 480.000000 224.300000 ;
      RECT 404.815000 223.500000 480.000000 223.900000 ;
      RECT 405.215000 223.100000 480.000000 223.500000 ;
      RECT 405.615000 222.700000 480.000000 223.100000 ;
      RECT 406.015000 222.300000 480.000000 222.700000 ;
      RECT 406.415000 221.900000 480.000000 222.300000 ;
      RECT 406.815000 221.500000 480.000000 221.900000 ;
      RECT 407.215000 221.100000 480.000000 221.500000 ;
      RECT 407.615000 220.700000 480.000000 221.100000 ;
      RECT 408.015000 220.300000 480.000000 220.700000 ;
      RECT 408.415000 219.900000 480.000000 220.300000 ;
      RECT 408.815000 219.500000 480.000000 219.900000 ;
      RECT 409.215000 219.100000 480.000000 219.500000 ;
      RECT 409.615000 218.700000 480.000000 219.100000 ;
      RECT 410.015000 218.300000 480.000000 218.700000 ;
      RECT 410.415000 217.900000 480.000000 218.300000 ;
      RECT 410.815000 217.500000 480.000000 217.900000 ;
      RECT 411.215000 217.100000 480.000000 217.500000 ;
      RECT 411.615000 216.700000 480.000000 217.100000 ;
      RECT 412.015000 216.300000 480.000000 216.700000 ;
      RECT 412.415000 215.900000 480.000000 216.300000 ;
      RECT 412.815000 215.500000 480.000000 215.900000 ;
      RECT 413.215000 215.100000 480.000000 215.500000 ;
      RECT 413.615000 214.700000 480.000000 215.100000 ;
      RECT 414.015000 214.300000 480.000000 214.700000 ;
      RECT 414.415000 213.900000 480.000000 214.300000 ;
      RECT 414.815000 213.500000 480.000000 213.900000 ;
      RECT 415.215000 213.100000 480.000000 213.500000 ;
      RECT 415.615000 212.700000 480.000000 213.100000 ;
      RECT 416.015000 212.300000 480.000000 212.700000 ;
      RECT 416.415000 211.900000 480.000000 212.300000 ;
      RECT 416.815000 211.500000 480.000000 211.900000 ;
      RECT 417.215000 211.100000 480.000000 211.500000 ;
      RECT 417.615000 210.700000 480.000000 211.100000 ;
      RECT 418.015000 210.300000 480.000000 210.700000 ;
      RECT 418.415000 209.900000 480.000000 210.300000 ;
      RECT 418.815000 209.500000 480.000000 209.900000 ;
      RECT 419.215000 209.100000 480.000000 209.500000 ;
      RECT 419.615000 208.700000 480.000000 209.100000 ;
      RECT 420.015000 208.300000 480.000000 208.700000 ;
      RECT 420.415000 207.900000 480.000000 208.300000 ;
      RECT 420.815000 207.500000 480.000000 207.900000 ;
      RECT 421.215000 207.100000 480.000000 207.500000 ;
      RECT 421.615000 206.700000 480.000000 207.100000 ;
      RECT 422.015000 206.300000 480.000000 206.700000 ;
      RECT 422.415000 205.900000 480.000000 206.300000 ;
      RECT 422.815000 205.500000 480.000000 205.900000 ;
      RECT 423.215000 205.100000 480.000000 205.500000 ;
      RECT 423.615000 204.700000 480.000000 205.100000 ;
      RECT 424.015000 204.300000 480.000000 204.700000 ;
      RECT 424.415000 203.900000 480.000000 204.300000 ;
      RECT 424.815000 203.500000 480.000000 203.900000 ;
      RECT 425.215000 203.100000 480.000000 203.500000 ;
      RECT 425.615000 202.700000 480.000000 203.100000 ;
      RECT 426.015000 202.300000 480.000000 202.700000 ;
      RECT 426.415000 201.900000 480.000000 202.300000 ;
      RECT 426.815000 201.500000 480.000000 201.900000 ;
      RECT 427.215000 201.100000 480.000000 201.500000 ;
      RECT 427.615000 200.700000 480.000000 201.100000 ;
      RECT 428.015000 200.300000 480.000000 200.700000 ;
      RECT 428.415000 199.900000 480.000000 200.300000 ;
      RECT 428.815000 199.500000 480.000000 199.900000 ;
      RECT 429.215000 199.100000 480.000000 199.500000 ;
      RECT 429.615000 198.700000 480.000000 199.100000 ;
      RECT 430.015000 198.300000 480.000000 198.700000 ;
      RECT 430.415000 197.900000 480.000000 198.300000 ;
      RECT 430.815000 197.500000 480.000000 197.900000 ;
      RECT 431.215000 197.100000 480.000000 197.500000 ;
      RECT 431.615000 196.700000 480.000000 197.100000 ;
      RECT 432.015000 196.300000 480.000000 196.700000 ;
      RECT 432.415000 195.900000 480.000000 196.300000 ;
      RECT 432.815000 195.500000 480.000000 195.900000 ;
      RECT 433.215000 195.100000 480.000000 195.500000 ;
      RECT 433.615000 194.700000 480.000000 195.100000 ;
      RECT 434.015000 194.300000 480.000000 194.700000 ;
      RECT 434.415000 193.900000 480.000000 194.300000 ;
      RECT 434.815000 193.500000 480.000000 193.900000 ;
      RECT 435.215000 193.100000 480.000000 193.500000 ;
      RECT 435.615000 192.700000 480.000000 193.100000 ;
      RECT 436.015000 192.300000 480.000000 192.700000 ;
      RECT 436.415000 191.900000 480.000000 192.300000 ;
      RECT 436.815000 191.500000 480.000000 191.900000 ;
      RECT 437.215000 191.100000 480.000000 191.500000 ;
      RECT 437.615000 190.700000 480.000000 191.100000 ;
      RECT 438.015000 190.300000 480.000000 190.700000 ;
      RECT 438.415000 189.900000 480.000000 190.300000 ;
      RECT 438.815000 189.500000 480.000000 189.900000 ;
      RECT 439.215000 189.100000 480.000000 189.500000 ;
      RECT 439.615000 188.700000 480.000000 189.100000 ;
      RECT 440.015000 188.300000 480.000000 188.700000 ;
      RECT 440.415000 187.900000 480.000000 188.300000 ;
      RECT 440.815000 187.500000 480.000000 187.900000 ;
      RECT 441.215000 187.100000 480.000000 187.500000 ;
      RECT 441.615000 186.700000 480.000000 187.100000 ;
      RECT 442.015000 186.300000 480.000000 186.700000 ;
      RECT 442.415000 185.900000 480.000000 186.300000 ;
      RECT 442.815000 185.500000 480.000000 185.900000 ;
      RECT 443.215000 185.100000 480.000000 185.500000 ;
      RECT 443.615000 184.700000 480.000000 185.100000 ;
      RECT 444.015000 184.300000 480.000000 184.700000 ;
      RECT 444.415000 183.900000 480.000000 184.300000 ;
      RECT 444.815000 183.500000 480.000000 183.900000 ;
      RECT 445.215000 183.100000 480.000000 183.500000 ;
      RECT 445.615000 182.700000 480.000000 183.100000 ;
      RECT 446.015000 182.300000 480.000000 182.700000 ;
      RECT 446.415000 181.900000 480.000000 182.300000 ;
      RECT 446.815000 181.500000 480.000000 181.900000 ;
      RECT 447.215000 181.100000 480.000000 181.500000 ;
      RECT 447.615000 180.700000 480.000000 181.100000 ;
      RECT 448.015000 180.300000 480.000000 180.700000 ;
      RECT 448.415000 179.900000 480.000000 180.300000 ;
      RECT 448.815000 179.500000 480.000000 179.900000 ;
      RECT 449.215000 179.100000 480.000000 179.500000 ;
      RECT 449.615000 178.700000 480.000000 179.100000 ;
      RECT 450.015000 178.300000 480.000000 178.700000 ;
      RECT 450.415000 177.900000 480.000000 178.300000 ;
      RECT 450.815000 177.500000 480.000000 177.900000 ;
      RECT 451.215000 177.100000 480.000000 177.500000 ;
      RECT 451.615000 176.700000 480.000000 177.100000 ;
      RECT 452.015000 176.300000 480.000000 176.700000 ;
      RECT 452.415000 175.900000 480.000000 176.300000 ;
      RECT 452.815000 175.500000 480.000000 175.900000 ;
      RECT 453.215000 175.100000 480.000000 175.500000 ;
      RECT 453.615000 174.700000 480.000000 175.100000 ;
      RECT 454.015000 174.300000 480.000000 174.700000 ;
      RECT 454.415000 173.900000 480.000000 174.300000 ;
      RECT 454.815000 173.500000 480.000000 173.900000 ;
      RECT 455.215000 173.100000 480.000000 173.500000 ;
      RECT 455.615000 172.700000 480.000000 173.100000 ;
      RECT 456.015000 172.300000 480.000000 172.700000 ;
      RECT 456.415000 171.900000 480.000000 172.300000 ;
      RECT 456.815000 171.500000 480.000000 171.900000 ;
      RECT 457.215000 171.100000 480.000000 171.500000 ;
      RECT 457.615000 170.700000 480.000000 171.100000 ;
      RECT 458.015000 170.300000 480.000000 170.700000 ;
      RECT 458.415000 169.900000 480.000000 170.300000 ;
      RECT 458.815000 169.500000 480.000000 169.900000 ;
      RECT 459.215000 169.100000 480.000000 169.500000 ;
      RECT 459.615000 168.700000 480.000000 169.100000 ;
      RECT 460.015000 168.300000 480.000000 168.700000 ;
      RECT 460.415000 167.900000 480.000000 168.300000 ;
      RECT 460.815000 167.500000 480.000000 167.900000 ;
      RECT 461.215000 167.100000 480.000000 167.500000 ;
      RECT 461.615000 166.700000 480.000000 167.100000 ;
      RECT 462.015000 166.300000 480.000000 166.700000 ;
      RECT 462.415000 165.900000 480.000000 166.300000 ;
      RECT 462.815000 165.500000 480.000000 165.900000 ;
      RECT 463.215000 165.100000 480.000000 165.500000 ;
      RECT 463.615000 164.700000 480.000000 165.100000 ;
      RECT 464.015000 164.300000 480.000000 164.700000 ;
      RECT 464.415000 163.900000 480.000000 164.300000 ;
      RECT 464.815000 163.500000 480.000000 163.900000 ;
      RECT 465.215000 163.100000 480.000000 163.500000 ;
      RECT 465.615000 162.700000 480.000000 163.100000 ;
      RECT 466.015000 162.300000 480.000000 162.700000 ;
      RECT 466.415000 161.900000 480.000000 162.300000 ;
      RECT 466.815000 161.500000 480.000000 161.900000 ;
      RECT 467.215000 161.100000 480.000000 161.500000 ;
      RECT 467.615000 160.700000 480.000000 161.100000 ;
      RECT 468.015000 160.300000 480.000000 160.700000 ;
      RECT 468.415000 159.900000 480.000000 160.300000 ;
      RECT 468.815000 159.500000 480.000000 159.900000 ;
      RECT 469.215000 159.100000 480.000000 159.500000 ;
      RECT 469.615000 158.700000 480.000000 159.100000 ;
      RECT 470.015000 158.300000 480.000000 158.700000 ;
      RECT 470.415000 157.900000 480.000000 158.300000 ;
      RECT 470.815000 157.500000 480.000000 157.900000 ;
      RECT 471.215000 157.100000 480.000000 157.500000 ;
      RECT 471.615000 156.700000 480.000000 157.100000 ;
      RECT 472.015000 156.300000 480.000000 156.700000 ;
      RECT 472.415000 155.900000 480.000000 156.300000 ;
      RECT 472.815000 155.500000 480.000000 155.900000 ;
      RECT 473.215000 155.100000 480.000000 155.500000 ;
      RECT 473.615000 154.700000 480.000000 155.100000 ;
      RECT 474.015000 154.300000 480.000000 154.700000 ;
      RECT 474.415000 153.900000 480.000000 154.300000 ;
      RECT 474.815000 153.500000 480.000000 153.900000 ;
      RECT 475.215000 153.100000 480.000000 153.500000 ;
      RECT 475.615000 152.700000 480.000000 153.100000 ;
      RECT 476.015000 152.300000 480.000000 152.700000 ;
      RECT 476.415000 151.900000 480.000000 152.300000 ;
      RECT 476.815000 151.500000 480.000000 151.900000 ;
      RECT 477.215000 151.100000 480.000000 151.500000 ;
      RECT 477.615000 150.700000 480.000000 151.100000 ;
      RECT 478.015000 150.300000 480.000000 150.700000 ;
      RECT 478.415000 149.900000 480.000000 150.300000 ;
      RECT 478.815000 149.500000 480.000000 149.900000 ;
      RECT 478.815000 149.500000 480.000000 228.700000 ;
  END
END sky130_fd_io__top_sio_macro
END LIBRARY
