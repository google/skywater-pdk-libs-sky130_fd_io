# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sky130_fd_io__top_sio_macro
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 480 BY 253.715 ;
  SYMMETRY R90 ;

  PIN vreg_en_refgen
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.84 22.305 445.1 22.34 ;
        RECT 444.84 22.34 445.135 22.375 ;
        RECT 444.84 22.375 445.17 23.015 ;
        RECT 444.84 0 445.1 22.305 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.0156 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END vreg_en_refgen

  PIN hld_h_n_refgen
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.955 14.81 405.595 15.07 ;
        RECT 404.995 14.685 405.255 14.725 ;
        RECT 404.995 14.725 405.295 14.765 ;
        RECT 404.995 14.765 405.335 14.77 ;
        RECT 404.995 14.77 405.34 14.79 ;
        RECT 404.975 14.79 405.36 14.81 ;
        RECT 404.995 0 405.255 14.685 ;
    END
    ANTENNAGATEAREA 2.4 LAYER met1 ;
    ANTENNAGATEAREA 2.4 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.6307 LAYER met2 ;
    ANTENNAGATEAREA 2.4 LAYER met3 ;
    ANTENNAGATEAREA 2.4 LAYER met4 ;
    ANTENNAGATEAREA 2.4 LAYER met5 ;
  END hld_h_n_refgen

  PIN voh_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.405 0 449.665 83.515 ;
        RECT 449.405 83.515 449.665 83.57 ;
        RECT 449.35 83.57 449.665 83.625 ;
        RECT 449.295 83.625 449.595 83.695 ;
        RECT 449.225 83.695 449.525 83.765 ;
        RECT 449.155 83.765 449.455 83.835 ;
        RECT 449.085 83.835 449.385 83.905 ;
        RECT 449.015 83.905 449.315 83.975 ;
        RECT 448.945 83.975 449.245 84.045 ;
        RECT 448.875 84.045 449.175 84.115 ;
        RECT 448.805 84.115 449.105 84.185 ;
        RECT 448.735 84.185 449.035 84.255 ;
        RECT 448.665 84.255 448.965 84.325 ;
        RECT 448.595 84.325 448.895 84.395 ;
        RECT 448.525 84.395 448.825 84.465 ;
        RECT 448.455 84.465 448.755 84.535 ;
        RECT 448.385 84.535 448.685 84.605 ;
        RECT 448.315 84.605 448.615 84.675 ;
        RECT 448.245 84.675 448.545 84.745 ;
        RECT 448.175 84.745 448.475 84.815 ;
        RECT 448.105 84.815 448.405 84.885 ;
        RECT 448.035 84.885 448.335 84.955 ;
        RECT 447.965 84.955 448.265 85.025 ;
        RECT 447.895 85.025 448.195 85.095 ;
        RECT 447.825 85.095 448.125 85.165 ;
        RECT 447.755 85.165 448.055 85.235 ;
        RECT 447.685 85.235 447.985 85.305 ;
        RECT 447.615 85.305 447.915 85.375 ;
        RECT 447.545 85.375 447.845 85.445 ;
        RECT 447.475 85.445 447.775 85.515 ;
        RECT 447.405 85.515 447.705 85.585 ;
        RECT 447.335 85.585 447.635 85.655 ;
        RECT 447.265 85.655 447.565 85.725 ;
        RECT 447.195 85.725 447.495 85.795 ;
        RECT 447.125 85.795 447.455 85.835 ;
        RECT 447.085 85.835 447.4 85.89 ;
        RECT 447.085 85.89 447.345 85.945 ;
        RECT 446.92 244.355 447.56 244.615 ;
        RECT 447.085 244.19 447.365 244.26 ;
        RECT 447.015 244.26 447.435 244.33 ;
        RECT 446.945 244.33 447.505 244.355 ;
        RECT 447.085 244.17 447.345 244.18 ;
        RECT 447.085 244.18 447.355 244.19 ;
        RECT 447.085 85.945 447.345 244.17 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 171.999 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END voh_sel[0]

  PIN voh_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.155 0 450.415 235.9 ;
        RECT 450.155 235.9 450.415 235.955 ;
        RECT 450.1 235.955 450.415 236.01 ;
        RECT 450.045 236.01 450.345 236.08 ;
        RECT 449.975 236.08 450.275 236.15 ;
        RECT 449.905 236.15 450.205 236.22 ;
        RECT 449.835 236.22 450.135 236.29 ;
        RECT 449.765 236.29 450.065 236.36 ;
        RECT 449.695 236.36 449.995 236.43 ;
        RECT 449.625 236.43 449.925 236.5 ;
        RECT 449.555 236.5 449.855 236.57 ;
        RECT 449.485 236.57 449.785 236.64 ;
        RECT 449.415 236.64 449.715 236.71 ;
        RECT 449.345 236.71 449.645 236.78 ;
        RECT 449.275 236.78 449.575 236.85 ;
        RECT 449.205 236.85 449.505 236.92 ;
        RECT 449.135 236.92 449.435 236.99 ;
        RECT 449.065 236.99 449.365 237.06 ;
        RECT 448.995 237.06 449.295 237.13 ;
        RECT 448.925 237.13 449.225 237.2 ;
        RECT 448.855 237.2 449.155 237.27 ;
        RECT 448.785 237.27 449.085 237.34 ;
        RECT 448.715 237.34 449.015 237.41 ;
        RECT 448.645 237.41 448.945 237.48 ;
        RECT 448.575 237.48 448.875 237.55 ;
        RECT 448.505 237.55 448.805 237.62 ;
        RECT 448.435 237.62 448.735 237.69 ;
        RECT 448.365 237.69 448.665 237.76 ;
        RECT 448.295 237.76 448.595 237.83 ;
        RECT 448.225 237.83 448.525 237.9 ;
        RECT 448.155 237.9 448.455 237.97 ;
        RECT 448.085 237.97 448.385 238.04 ;
        RECT 448.015 238.04 448.315 238.11 ;
        RECT 447.945 238.11 448.245 238.18 ;
        RECT 447.875 238.18 448.175 238.25 ;
        RECT 447.805 238.25 448.115 238.31 ;
        RECT 447.745 238.31 448.06 238.365 ;
        RECT 447.745 238.365 448.005 238.42 ;
        RECT 447.745 238.42 448.005 245.015 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 172.136 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END voh_sel[1]

  PIN voutref_dft
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.53 0 465.17 60.295 ;
    END
    ANTENNADIFFAREA 2.65 LAYER met1 ;
    ANTENNADIFFAREA 2.65 LAYER met2 ;
    ANTENNADIFFAREA 2.65 LAYER met3 ;
    ANTENNADIFFAREA 2.65 LAYER met4 ;
    ANTENNADIFFAREA 2.65 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 42.1365 LAYER met2 ;
  END voutref_dft

  PIN ibuf_sel_refgen
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.69 0 422.95 23.14 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.044 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END ibuf_sel_refgen

  PIN vref_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.155 0 453.415 237.18 ;
        RECT 453.155 237.18 453.415 237.235 ;
        RECT 453.1 237.235 453.415 237.29 ;
        RECT 453.045 237.29 453.345 237.36 ;
        RECT 452.975 237.36 453.275 237.43 ;
        RECT 452.905 237.43 453.205 237.5 ;
        RECT 452.835 237.5 453.135 237.57 ;
        RECT 452.765 237.57 453.065 237.64 ;
        RECT 452.695 237.64 452.995 237.71 ;
        RECT 452.625 237.71 452.925 237.78 ;
        RECT 452.555 237.78 452.855 237.85 ;
        RECT 452.485 237.85 452.785 237.92 ;
        RECT 452.415 237.92 452.715 237.99 ;
        RECT 452.345 237.99 452.645 238.06 ;
        RECT 452.275 238.06 452.575 238.13 ;
        RECT 452.205 238.13 452.505 238.2 ;
        RECT 452.135 238.2 452.435 238.27 ;
        RECT 452.065 238.27 452.365 238.34 ;
        RECT 451.995 238.34 452.295 238.41 ;
        RECT 451.925 238.41 452.225 238.48 ;
        RECT 451.855 238.48 452.155 238.55 ;
        RECT 451.785 238.55 452.085 238.62 ;
        RECT 451.715 238.62 452.015 238.69 ;
        RECT 451.645 238.69 451.945 238.76 ;
        RECT 451.575 238.76 451.875 238.83 ;
        RECT 451.505 238.83 451.805 238.9 ;
        RECT 451.435 238.9 451.735 238.97 ;
        RECT 451.365 238.97 451.665 239.04 ;
        RECT 451.295 239.04 451.595 239.11 ;
        RECT 451.225 239.11 451.525 239.18 ;
        RECT 451.155 239.18 451.455 239.25 ;
        RECT 451.085 239.25 451.385 239.32 ;
        RECT 451.015 239.32 451.315 239.39 ;
        RECT 450.945 239.39 451.245 239.46 ;
        RECT 450.875 239.46 451.175 239.53 ;
        RECT 450.805 239.53 451.115 239.59 ;
        RECT 450.745 239.59 451.06 239.645 ;
        RECT 450.745 239.645 451.005 239.7 ;
        RECT 450.745 239.7 451.005 241.785 ;
    END
    ANTENNAGATEAREA 0.999 LAYER met1 ;
    ANTENNAGATEAREA 0.999 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 172.049 LAYER met2 ;
    ANTENNAGATEAREA 0.999 LAYER met3 ;
    ANTENNAGATEAREA 0.999 LAYER met4 ;
    ANTENNAGATEAREA 0.999 LAYER met5 ;
  END vref_sel[0]

  PIN voh_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.905 0 451.165 236.22 ;
        RECT 450.905 236.22 451.165 236.275 ;
        RECT 450.85 236.275 451.165 236.33 ;
        RECT 450.795 236.33 451.095 236.4 ;
        RECT 450.725 236.4 451.025 236.47 ;
        RECT 450.655 236.47 450.955 236.54 ;
        RECT 450.585 236.54 450.885 236.61 ;
        RECT 450.515 236.61 450.815 236.68 ;
        RECT 450.445 236.68 450.745 236.75 ;
        RECT 450.375 236.75 450.675 236.82 ;
        RECT 450.305 236.82 450.605 236.89 ;
        RECT 450.235 236.89 450.535 236.96 ;
        RECT 450.165 236.96 450.465 237.03 ;
        RECT 450.095 237.03 450.395 237.1 ;
        RECT 450.025 237.1 450.325 237.17 ;
        RECT 449.955 237.17 450.255 237.24 ;
        RECT 449.885 237.24 450.185 237.31 ;
        RECT 449.815 237.31 450.115 237.38 ;
        RECT 449.745 237.38 450.045 237.45 ;
        RECT 449.675 237.45 449.975 237.52 ;
        RECT 449.605 237.52 449.905 237.59 ;
        RECT 449.535 237.59 449.835 237.66 ;
        RECT 449.465 237.66 449.765 237.73 ;
        RECT 449.395 237.73 449.695 237.8 ;
        RECT 449.325 237.8 449.625 237.87 ;
        RECT 449.255 237.87 449.555 237.94 ;
        RECT 449.185 237.94 449.485 238.01 ;
        RECT 449.115 238.01 449.415 238.08 ;
        RECT 449.045 238.08 449.345 238.15 ;
        RECT 448.975 238.15 449.275 238.22 ;
        RECT 448.905 238.22 449.205 238.29 ;
        RECT 448.835 238.29 449.135 238.36 ;
        RECT 448.765 238.36 449.065 238.43 ;
        RECT 448.695 238.43 448.995 238.5 ;
        RECT 448.625 238.5 448.925 238.57 ;
        RECT 448.555 238.57 448.865 238.63 ;
        RECT 448.495 238.63 448.81 238.685 ;
        RECT 448.495 238.685 448.755 238.74 ;
        RECT 448.495 238.74 448.755 245.415 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 172.395 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END voh_sel[2]

  PIN vohref
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.445 0 419.705 5.035 ;
    END
    ANTENNADIFFAREA 2.65 LAYER met1 ;
    ANTENNADIFFAREA 2.65 LAYER met2 ;
    ANTENNADIFFAREA 2.65 LAYER met3 ;
    ANTENNADIFFAREA 2.65 LAYER met4 ;
    ANTENNADIFFAREA 2.65 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 58.065 LAYER met2 ;
  END vohref

  PIN pad_a_esd_1_h[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.99 0 178.99 24.23 ;
    END
    ANTENNAPARTIALMETALSIDEAREA 16.7475 LAYER met2 ;
  END pad_a_esd_1_h[0]

  PIN ibuf_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.57 0 254.83 28.84 ;
        RECT 254.57 28.84 254.83 28.895 ;
        RECT 254.57 28.895 254.885 28.95 ;
        RECT 254.64 28.95 254.94 29.02 ;
        RECT 254.71 29.02 255.01 29.09 ;
        RECT 254.78 29.09 255.08 29.16 ;
        RECT 254.85 29.16 255.15 29.23 ;
        RECT 254.92 29.23 255.22 29.3 ;
        RECT 254.99 29.3 255.29 29.37 ;
        RECT 255.045 29.37 255.36 29.425 ;
        RECT 255.1 29.425 255.36 29.48 ;
        RECT 255.1 29.48 255.36 29.86 ;
        RECT 255.1 29.86 255.36 29.915 ;
        RECT 255.1 29.915 255.415 29.97 ;
        RECT 255.105 29.97 255.47 29.975 ;
        RECT 255.11 29.975 255.475 29.98 ;
        RECT 255.115 29.98 255.48 29.985 ;
        RECT 255.185 29.985 256.25 30.055 ;
        RECT 255.255 30.055 256.25 30.125 ;
        RECT 255.325 30.125 256.25 30.195 ;
        RECT 255.375 30.195 256.25 30.245 ;
        RECT 255.545 30.245 255.935 30.305 ;
        RECT 255.605 30.305 255.875 30.365 ;
        RECT 255.61 30.365 255.87 30.37 ;
        RECT 255.61 30.37 255.87 42.74 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.3479 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END ibuf_sel[1]

  PIN enable_vdda_h
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.405 0 452.665 236.86 ;
        RECT 452.405 236.86 452.665 236.915 ;
        RECT 452.35 236.915 452.665 236.97 ;
        RECT 452.295 236.97 452.595 237.04 ;
        RECT 452.225 237.04 452.525 237.11 ;
        RECT 452.155 237.11 452.455 237.18 ;
        RECT 452.085 237.18 452.385 237.25 ;
        RECT 452.015 237.25 452.315 237.32 ;
        RECT 451.945 237.32 452.245 237.39 ;
        RECT 451.875 237.39 452.175 237.46 ;
        RECT 451.805 237.46 452.105 237.53 ;
        RECT 451.735 237.53 452.035 237.6 ;
        RECT 451.665 237.6 451.965 237.67 ;
        RECT 451.595 237.67 451.895 237.74 ;
        RECT 451.525 237.74 451.825 237.81 ;
        RECT 451.455 237.81 451.755 237.88 ;
        RECT 451.385 237.88 451.685 237.95 ;
        RECT 451.315 237.95 451.615 238.02 ;
        RECT 451.245 238.02 451.545 238.09 ;
        RECT 451.175 238.09 451.475 238.16 ;
        RECT 451.105 238.16 451.405 238.23 ;
        RECT 451.035 238.23 451.335 238.3 ;
        RECT 450.965 238.3 451.265 238.37 ;
        RECT 450.895 238.37 451.195 238.44 ;
        RECT 450.825 238.44 451.125 238.51 ;
        RECT 450.755 238.51 451.055 238.58 ;
        RECT 450.685 238.58 450.985 238.65 ;
        RECT 450.615 238.65 450.915 238.72 ;
        RECT 450.545 238.72 450.845 238.79 ;
        RECT 450.475 238.79 450.775 238.86 ;
        RECT 450.405 238.86 450.705 238.93 ;
        RECT 450.335 238.93 450.635 239 ;
        RECT 450.265 239 450.565 239.07 ;
        RECT 450.195 239.07 450.495 239.14 ;
        RECT 450.125 239.14 450.425 239.21 ;
        RECT 450.055 239.21 450.365 239.27 ;
        RECT 449.995 239.27 450.31 239.325 ;
        RECT 449.995 239.325 450.255 239.38 ;
        RECT 449.995 239.38 450.255 240.715 ;
    END
    ANTENNAGATEAREA 19.2 LAYER met1 ;
    ANTENNAGATEAREA 19.2 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 171.065 LAYER met2 ;
    ANTENNAGATEAREA 19.2 LAYER met3 ;
    ANTENNAGATEAREA 19.2 LAYER met4 ;
    ANTENNAGATEAREA 19.2 LAYER met5 ;
  END enable_vdda_h

  PIN vinref_dft
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.03 0 466.67 60.295 ;
    END
    ANTENNADIFFAREA 2.65 LAYER met1 ;
    ANTENNADIFFAREA 2.65 LAYER met2 ;
    ANTENNADIFFAREA 2.65 LAYER met3 ;
    ANTENNADIFFAREA 2.65 LAYER met4 ;
    ANTENNADIFFAREA 2.65 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 42.1365 LAYER met2 ;
  END vinref_dft

  PIN vtrip_sel_refgen
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.84 0 403.1 23.14 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.0545 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END vtrip_sel_refgen

  PIN dft_refgen
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.655 0 451.915 236.54 ;
        RECT 451.655 236.54 451.915 236.595 ;
        RECT 451.6 236.595 451.915 236.65 ;
        RECT 451.545 236.65 451.845 236.72 ;
        RECT 451.475 236.72 451.775 236.79 ;
        RECT 451.405 236.79 451.705 236.86 ;
        RECT 451.335 236.86 451.635 236.93 ;
        RECT 451.265 236.93 451.565 237 ;
        RECT 451.195 237 451.495 237.07 ;
        RECT 451.125 237.07 451.425 237.14 ;
        RECT 451.055 237.14 451.355 237.21 ;
        RECT 450.985 237.21 451.285 237.28 ;
        RECT 450.915 237.28 451.215 237.35 ;
        RECT 450.845 237.35 451.145 237.42 ;
        RECT 450.775 237.42 451.075 237.49 ;
        RECT 450.705 237.49 451.005 237.56 ;
        RECT 450.635 237.56 450.935 237.63 ;
        RECT 450.565 237.63 450.865 237.7 ;
        RECT 450.495 237.7 450.795 237.77 ;
        RECT 450.425 237.77 450.725 237.84 ;
        RECT 450.355 237.84 450.655 237.91 ;
        RECT 450.285 237.91 450.585 237.98 ;
        RECT 450.215 237.98 450.515 238.05 ;
        RECT 450.145 238.05 450.445 238.12 ;
        RECT 450.075 238.12 450.375 238.19 ;
        RECT 450.005 238.19 450.305 238.26 ;
        RECT 449.935 238.26 450.235 238.33 ;
        RECT 449.865 238.33 450.165 238.4 ;
        RECT 449.795 238.4 450.095 238.47 ;
        RECT 449.725 238.47 450.025 238.54 ;
        RECT 449.655 238.54 449.955 238.61 ;
        RECT 449.585 238.61 449.885 238.68 ;
        RECT 449.515 238.68 449.815 238.75 ;
        RECT 449.445 238.75 449.745 238.82 ;
        RECT 449.375 238.82 449.675 238.89 ;
        RECT 449.305 238.89 449.615 238.95 ;
        RECT 449.245 238.95 449.56 239.005 ;
        RECT 449.245 239.005 449.505 239.06 ;
        RECT 449.245 239.06 449.505 245.815 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 172.587 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END dft_refgen

  PIN pad_a_esd_1_h[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.015 0 213.015 24.23 ;
    END
    ANTENNAPARTIALMETALSIDEAREA 16.7475 LAYER met2 ;
  END pad_a_esd_1_h[1]

  PIN pad_a_esd_0_h[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.9 0 304.745 30.545 ;
    END
    ANTENNAPARTIALMETALSIDEAREA 21.168 LAYER met2 ;
  END pad_a_esd_0_h[1]

  PIN vref_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.905 0 454.165 237.5 ;
        RECT 453.905 237.5 454.165 237.555 ;
        RECT 453.85 237.555 454.165 237.61 ;
        RECT 453.795 237.61 454.095 237.68 ;
        RECT 453.725 237.68 454.025 237.75 ;
        RECT 453.655 237.75 453.955 237.82 ;
        RECT 453.585 237.82 453.885 237.89 ;
        RECT 453.515 237.89 453.815 237.96 ;
        RECT 453.445 237.96 453.745 238.03 ;
        RECT 453.375 238.03 453.675 238.1 ;
        RECT 453.305 238.1 453.605 238.17 ;
        RECT 453.235 238.17 453.535 238.24 ;
        RECT 453.165 238.24 453.465 238.31 ;
        RECT 453.095 238.31 453.395 238.38 ;
        RECT 453.025 238.38 453.325 238.45 ;
        RECT 452.955 238.45 453.255 238.52 ;
        RECT 452.885 238.52 453.185 238.59 ;
        RECT 452.815 238.59 453.115 238.66 ;
        RECT 452.745 238.66 453.045 238.73 ;
        RECT 452.675 238.73 452.975 238.8 ;
        RECT 452.605 238.8 452.905 238.87 ;
        RECT 452.535 238.87 452.835 238.94 ;
        RECT 452.465 238.94 452.765 239.01 ;
        RECT 452.395 239.01 452.695 239.08 ;
        RECT 452.325 239.08 452.625 239.15 ;
        RECT 452.255 239.15 452.555 239.22 ;
        RECT 452.185 239.22 452.485 239.29 ;
        RECT 452.115 239.29 452.415 239.36 ;
        RECT 452.045 239.36 452.345 239.43 ;
        RECT 451.975 239.43 452.275 239.5 ;
        RECT 451.905 239.5 452.205 239.57 ;
        RECT 451.835 239.57 452.135 239.64 ;
        RECT 451.765 239.64 452.065 239.71 ;
        RECT 451.695 239.71 451.995 239.78 ;
        RECT 451.625 239.78 451.925 239.85 ;
        RECT 451.555 239.85 451.865 239.91 ;
        RECT 451.495 239.91 451.81 239.965 ;
        RECT 451.495 239.965 451.755 240.02 ;
        RECT 451.115 241.965 451.755 242.225 ;
        RECT 451.495 241.76 451.755 241.83 ;
        RECT 451.425 241.83 451.755 241.9 ;
        RECT 451.355 241.9 451.755 241.965 ;
        RECT 451.495 240.02 451.755 241.76 ;
    END
    ANTENNAGATEAREA 0.999 LAYER met1 ;
    ANTENNAGATEAREA 0.999 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 179.002 LAYER met2 ;
    ANTENNAGATEAREA 0.999 LAYER met3 ;
    ANTENNAGATEAREA 0.999 LAYER met4 ;
    ANTENNAGATEAREA 0.999 LAYER met5 ;
  END vref_sel[1]

  PIN pad_a_esd_0_h[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.26 0 86.105 30.545 ;
    END
    ANTENNAPARTIALMETALSIDEAREA 21.168 LAYER met2 ;
  END pad_a_esd_0_h[0]

  PIN pad_a_noesd_h[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.245 0 87.095 33.235 ;
    END
    ANTENNAPARTIALMETALSIDEAREA 23.051 LAYER met2 ;
  END pad_a_noesd_h[0]

  PIN pad_a_noesd_h[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.91 0 303.76 33.235 ;
    END
    ANTENNAPARTIALMETALSIDEAREA 23.0545 LAYER met2 ;
  END pad_a_noesd_h[1]

  PIN inp_dis[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.035 0 283.295 1.24 ;
        RECT 283.035 1.24 283.295 1.295 ;
        RECT 282.98 1.295 283.295 1.35 ;
        RECT 282.925 1.35 283.225 1.42 ;
        RECT 282.855 1.42 283.155 1.49 ;
        RECT 282.785 1.49 283.085 1.56 ;
        RECT 282.715 1.56 283.015 1.63 ;
        RECT 282.645 1.63 282.945 1.7 ;
        RECT 282.575 1.7 282.875 1.77 ;
        RECT 282.505 1.77 282.805 1.84 ;
        RECT 282.435 1.84 282.735 1.91 ;
        RECT 282.365 1.91 282.69 1.955 ;
        RECT 282.32 1.955 282.635 2.01 ;
        RECT 282.32 2.01 282.58 2.065 ;
        RECT 282.32 2.065 282.58 18.155 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.7529 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END inp_dis[1]

  PIN inp_dis[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.71 0 106.97 1.24 ;
        RECT 106.71 1.24 106.97 1.295 ;
        RECT 106.71 1.295 107.025 1.35 ;
        RECT 106.78 1.35 107.08 1.42 ;
        RECT 106.85 1.42 107.15 1.49 ;
        RECT 106.92 1.49 107.22 1.56 ;
        RECT 106.99 1.56 107.29 1.63 ;
        RECT 107.06 1.63 107.36 1.7 ;
        RECT 107.13 1.7 107.43 1.77 ;
        RECT 107.2 1.77 107.5 1.84 ;
        RECT 107.27 1.84 107.57 1.91 ;
        RECT 107.315 1.91 107.64 1.955 ;
        RECT 107.37 1.955 107.685 2.01 ;
        RECT 107.425 2.01 107.685 2.065 ;
        RECT 107.425 2.065 107.685 18.155 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.7529 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END inp_dis[0]

  PIN tie_lo_esd[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.09 0 110.35 17.355 ;
        RECT 110.09 17.355 110.35 17.41 ;
        RECT 110.035 17.41 110.35 17.465 ;
        RECT 109.98 17.465 110.28 17.535 ;
        RECT 109.91 17.535 110.21 17.605 ;
        RECT 109.84 17.605 110.185 17.63 ;
        RECT 109.815 17.63 110.13 17.685 ;
        RECT 109.815 17.685 110.075 17.74 ;
        RECT 109.815 17.74 110.075 36.3 ;
        RECT 109.815 36.3 110.075 36.31 ;
        RECT 109.815 36.31 110.085 36.32 ;
        RECT 109.815 36.32 110.095 36.41 ;
        RECT 109.825 36.41 110.095 36.42 ;
        RECT 109.835 36.42 110.095 36.43 ;
        RECT 109.835 36.43 110.095 45.48 ;
        RECT 109.835 45.48 110.095 45.535 ;
        RECT 109.78 45.535 110.095 45.59 ;
        RECT 109.725 45.59 110.025 45.66 ;
        RECT 109.655 45.66 109.955 45.73 ;
        RECT 109.585 45.73 109.885 45.8 ;
        RECT 109.515 45.8 109.835 45.85 ;
        RECT 109.465 45.85 109.78 45.905 ;
        RECT 109.465 45.905 109.725 45.96 ;
        RECT 109.465 45.96 109.725 46.565 ;
        RECT 109.465 46.565 109.725 46.62 ;
        RECT 109.41 46.62 109.725 46.675 ;
        RECT 109.355 46.675 109.655 46.745 ;
        RECT 109.285 46.745 109.585 46.815 ;
        RECT 109.215 46.815 109.515 46.885 ;
        RECT 109.145 46.885 109.445 46.955 ;
        RECT 109.075 46.955 109.375 47.025 ;
        RECT 109.005 47.025 109.305 47.095 ;
        RECT 108.935 47.095 109.235 47.165 ;
        RECT 108.865 47.165 109.165 47.235 ;
        RECT 108.795 47.235 109.095 47.305 ;
        RECT 108.725 47.305 109.025 47.375 ;
        RECT 108.655 47.375 108.955 47.445 ;
        RECT 108.585 47.445 108.94 47.46 ;
        RECT 108.57 47.46 108.885 47.515 ;
        RECT 108.57 47.515 108.83 47.57 ;
        RECT 108.57 56.455 108.83 56.51 ;
        RECT 108.57 56.51 108.885 56.565 ;
        RECT 108.64 56.565 108.94 56.635 ;
        RECT 108.71 56.635 109.01 56.705 ;
        RECT 108.78 56.705 109.08 56.775 ;
        RECT 108.85 56.775 109.15 56.845 ;
        RECT 108.92 56.845 109.22 56.915 ;
        RECT 108.99 56.915 109.29 56.985 ;
        RECT 109.06 56.985 109.36 57.055 ;
        RECT 109.13 57.055 109.43 57.125 ;
        RECT 109.2 57.125 109.5 57.195 ;
        RECT 109.27 57.195 109.57 57.265 ;
        RECT 109.325 57.265 109.64 57.32 ;
        RECT 109.38 57.32 109.64 57.375 ;
        RECT 109.38 57.375 109.64 74.88 ;
        RECT 109.38 74.88 109.64 74.935 ;
        RECT 109.325 74.935 109.64 74.99 ;
        RECT 109.27 74.99 109.57 75.06 ;
        RECT 109.2 75.06 109.5 75.13 ;
        RECT 109.13 75.13 109.43 75.2 ;
        RECT 109.06 75.2 109.36 75.27 ;
        RECT 108.99 75.27 109.29 75.34 ;
        RECT 108.92 75.34 109.22 75.41 ;
        RECT 108.85 75.41 109.15 75.48 ;
        RECT 108.78 75.48 109.08 75.55 ;
        RECT 108.71 75.55 109.01 75.62 ;
        RECT 108.64 75.62 108.94 75.69 ;
        RECT 108.57 75.69 108.87 75.76 ;
        RECT 108.5 75.76 108.8 75.83 ;
        RECT 108.43 75.83 108.73 75.9 ;
        RECT 108.36 75.9 108.66 75.97 ;
        RECT 108.29 75.97 108.59 76.04 ;
        RECT 108.22 76.04 108.52 76.11 ;
        RECT 108.15 76.11 108.45 76.18 ;
        RECT 108.08 76.18 108.38 76.25 ;
        RECT 108.01 76.25 108.31 76.32 ;
        RECT 107.94 76.32 108.24 76.39 ;
        RECT 107.87 76.39 108.17 76.46 ;
        RECT 107.8 76.46 108.12 76.51 ;
        RECT 107.75 76.51 108.065 76.565 ;
        RECT 107.75 76.565 108.01 76.62 ;
        RECT 107.75 76.62 108.01 87.54 ;
        RECT 107.75 87.54 108.01 87.595 ;
        RECT 107.695 87.595 108.01 87.65 ;
        RECT 107.64 87.65 107.94 87.72 ;
        RECT 107.57 87.72 107.87 87.79 ;
        RECT 107.5 87.79 107.8 87.86 ;
        RECT 107.43 87.86 107.73 87.93 ;
        RECT 107.36 87.93 107.66 88 ;
        RECT 107.29 88 107.59 88.07 ;
        RECT 107.22 88.07 107.52 88.14 ;
        RECT 107.15 88.14 107.45 88.21 ;
        RECT 107.08 88.21 107.38 88.28 ;
        RECT 107.01 88.28 107.31 88.35 ;
        RECT 106.94 88.35 107.24 88.42 ;
        RECT 106.87 88.42 107.17 88.49 ;
        RECT 106.8 88.49 107.1 88.56 ;
        RECT 106.73 88.56 107.03 88.63 ;
        RECT 106.66 88.63 106.96 88.7 ;
        RECT 106.59 88.7 106.89 88.77 ;
        RECT 106.52 88.77 106.82 88.84 ;
        RECT 106.45 88.84 106.75 88.91 ;
        RECT 106.38 88.91 106.68 88.98 ;
        RECT 106.31 88.98 106.61 89.05 ;
        RECT 106.24 89.05 106.54 89.12 ;
        RECT 106.17 89.12 106.47 89.19 ;
        RECT 106.1 89.19 106.4 89.26 ;
        RECT 106.03 89.26 106.33 89.33 ;
        RECT 105.96 89.33 106.26 89.4 ;
        RECT 105.89 89.4 106.19 89.47 ;
        RECT 105.82 89.47 106.18 89.48 ;
        RECT 105.81 89.48 106.14 89.52 ;
        RECT 105.81 89.52 106.1 89.56 ;
        RECT 105.81 89.56 106.095 89.565 ;
        RECT 105.81 89.565 106.095 94.165 ;
        RECT 105.81 94.165 106.095 94.205 ;
        RECT 105.77 94.205 106.095 94.245 ;
        RECT 105.73 94.245 106.095 94.25 ;
        RECT 105.725 94.25 106.025 94.32 ;
        RECT 105.655 94.32 105.955 94.39 ;
        RECT 105.585 94.39 105.885 94.46 ;
        RECT 105.515 94.46 105.815 94.53 ;
        RECT 105.445 94.53 105.745 94.6 ;
        RECT 105.375 94.6 105.675 94.67 ;
        RECT 105.305 94.67 105.645 94.7 ;
        RECT 100.59 94.7 105.575 94.77 ;
        RECT 100.52 94.77 105.505 94.84 ;
        RECT 100.45 94.84 105.435 94.91 ;
        RECT 100.38 94.91 105.385 94.96 ;
        RECT 92.35 102.94 92.675 102.985 ;
        RECT 92.42 102.87 92.72 102.94 ;
        RECT 92.49 102.8 92.79 102.87 ;
        RECT 92.56 102.73 92.86 102.8 ;
        RECT 92.63 102.66 92.93 102.73 ;
        RECT 92.7 102.59 93 102.66 ;
        RECT 92.77 102.52 93.07 102.59 ;
        RECT 92.84 102.45 93.14 102.52 ;
        RECT 92.91 102.38 93.21 102.45 ;
        RECT 92.98 102.31 93.28 102.38 ;
        RECT 93.05 102.24 93.35 102.31 ;
        RECT 93.12 102.17 93.42 102.24 ;
        RECT 93.19 102.1 93.49 102.17 ;
        RECT 93.26 102.03 93.56 102.1 ;
        RECT 93.33 101.96 93.63 102.03 ;
        RECT 93.4 101.89 93.7 101.96 ;
        RECT 93.47 101.82 93.77 101.89 ;
        RECT 93.54 101.75 93.84 101.82 ;
        RECT 93.61 101.68 93.91 101.75 ;
        RECT 93.68 101.61 93.98 101.68 ;
        RECT 93.75 101.54 94.05 101.61 ;
        RECT 93.82 101.47 94.12 101.54 ;
        RECT 93.89 101.4 94.19 101.47 ;
        RECT 93.96 101.33 94.26 101.4 ;
        RECT 94.03 101.26 94.33 101.33 ;
        RECT 94.1 101.19 94.4 101.26 ;
        RECT 94.17 101.12 94.47 101.19 ;
        RECT 94.24 101.05 94.54 101.12 ;
        RECT 94.31 100.98 94.61 101.05 ;
        RECT 94.38 100.91 94.68 100.98 ;
        RECT 94.45 100.84 94.75 100.91 ;
        RECT 94.52 100.77 94.82 100.84 ;
        RECT 94.59 100.7 94.89 100.77 ;
        RECT 94.66 100.63 94.96 100.7 ;
        RECT 94.73 100.56 95.03 100.63 ;
        RECT 94.8 100.49 95.1 100.56 ;
        RECT 94.87 100.42 95.17 100.49 ;
        RECT 94.94 100.35 95.24 100.42 ;
        RECT 95.01 100.28 95.31 100.35 ;
        RECT 95.08 100.21 95.38 100.28 ;
        RECT 95.15 100.14 95.45 100.21 ;
        RECT 95.22 100.07 95.52 100.14 ;
        RECT 95.29 100 95.59 100.07 ;
        RECT 95.36 99.93 95.66 100 ;
        RECT 95.43 99.86 95.73 99.93 ;
        RECT 95.5 99.79 95.8 99.86 ;
        RECT 95.57 99.72 95.87 99.79 ;
        RECT 95.64 99.65 95.94 99.72 ;
        RECT 95.71 99.58 96.01 99.65 ;
        RECT 95.78 99.51 96.08 99.58 ;
        RECT 95.85 99.44 96.15 99.51 ;
        RECT 95.92 99.37 96.22 99.44 ;
        RECT 95.99 99.3 96.29 99.37 ;
        RECT 96.06 99.23 96.36 99.3 ;
        RECT 96.13 99.16 96.43 99.23 ;
        RECT 96.2 99.09 96.5 99.16 ;
        RECT 96.27 99.02 96.57 99.09 ;
        RECT 96.34 98.95 96.64 99.02 ;
        RECT 96.41 98.88 96.71 98.95 ;
        RECT 96.48 98.81 96.78 98.88 ;
        RECT 96.55 98.74 96.85 98.81 ;
        RECT 96.62 98.67 96.92 98.74 ;
        RECT 96.69 98.6 96.99 98.67 ;
        RECT 96.76 98.53 97.06 98.6 ;
        RECT 96.83 98.46 97.13 98.53 ;
        RECT 96.9 98.39 97.2 98.46 ;
        RECT 96.97 98.32 97.27 98.39 ;
        RECT 97.04 98.25 97.34 98.32 ;
        RECT 97.11 98.18 97.41 98.25 ;
        RECT 97.18 98.11 97.48 98.18 ;
        RECT 97.25 98.04 97.55 98.11 ;
        RECT 97.32 97.97 97.62 98.04 ;
        RECT 97.39 97.9 97.69 97.97 ;
        RECT 97.46 97.83 97.76 97.9 ;
        RECT 97.53 97.76 97.83 97.83 ;
        RECT 97.6 97.69 97.9 97.76 ;
        RECT 97.67 97.62 97.97 97.69 ;
        RECT 97.74 97.55 98.04 97.62 ;
        RECT 97.81 97.48 98.11 97.55 ;
        RECT 97.88 97.41 98.18 97.48 ;
        RECT 97.95 97.34 98.25 97.41 ;
        RECT 98.02 97.27 98.32 97.34 ;
        RECT 98.09 97.2 98.39 97.27 ;
        RECT 98.16 97.13 98.46 97.2 ;
        RECT 98.23 97.06 98.53 97.13 ;
        RECT 98.3 96.99 98.6 97.06 ;
        RECT 98.37 96.92 98.67 96.99 ;
        RECT 98.44 96.85 98.74 96.92 ;
        RECT 98.51 96.78 98.81 96.85 ;
        RECT 98.58 96.71 98.88 96.78 ;
        RECT 98.65 96.64 98.95 96.71 ;
        RECT 98.72 96.57 99.02 96.64 ;
        RECT 98.79 96.5 99.09 96.57 ;
        RECT 98.86 96.43 99.16 96.5 ;
        RECT 98.93 96.36 99.23 96.43 ;
        RECT 99 96.29 99.3 96.36 ;
        RECT 99.07 96.22 99.37 96.29 ;
        RECT 99.14 96.15 99.44 96.22 ;
        RECT 99.21 96.08 99.51 96.15 ;
        RECT 99.28 96.01 99.58 96.08 ;
        RECT 99.35 95.94 99.65 96.01 ;
        RECT 99.42 95.87 99.72 95.94 ;
        RECT 99.49 95.8 99.79 95.87 ;
        RECT 99.56 95.73 99.86 95.8 ;
        RECT 99.63 95.66 99.93 95.73 ;
        RECT 99.7 95.59 100 95.66 ;
        RECT 99.77 95.52 100.07 95.59 ;
        RECT 99.84 95.45 100.14 95.52 ;
        RECT 99.91 95.38 100.21 95.45 ;
        RECT 99.98 95.31 100.28 95.38 ;
        RECT 100.05 95.24 100.35 95.31 ;
        RECT 100.12 95.17 100.42 95.24 ;
        RECT 100.19 95.1 100.49 95.17 ;
        RECT 100.26 95.03 100.56 95.1 ;
        RECT 100.33 94.96 100.63 95.03 ;
        RECT 92.305 102.985 92.635 103.025 ;
        RECT 92.305 103.025 92.595 103.065 ;
        RECT 92.305 111.375 92.595 111.435 ;
        RECT 92.305 111.435 92.655 111.495 ;
        RECT 92.305 111.495 92.715 111.5 ;
        RECT 108.57 47.57 108.83 56.455 ;
        RECT 92.305 111.5 93.345 111.6 ;
        RECT 92.375 111.6 93.345 111.67 ;
        RECT 92.445 111.67 93.345 111.74 ;
        RECT 92.465 111.74 93.345 111.76 ;
        RECT 93.085 111.9 93.345 112.14 ;
        RECT 93.015 111.76 93.345 111.83 ;
        RECT 93.085 111.83 93.345 111.9 ;
        RECT 92.305 103.065 92.595 111.375 ;
    END
    ANTENNAGATEAREA 2.4 LAYER met1 ;
    ANTENNAGATEAREA 2.4 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 186.303 LAYER met2 ;
    ANTENNAGATEAREA 2.4 LAYER met3 ;
    ANTENNAGATEAREA 2.4 LAYER met4 ;
    ANTENNAGATEAREA 2.4 LAYER met5 ;
  END tie_lo_esd[0]

  PIN tie_lo_esd[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.655 0 279.915 17.355 ;
        RECT 279.655 17.355 279.915 17.41 ;
        RECT 279.655 17.41 279.97 17.465 ;
        RECT 279.725 17.465 280.025 17.535 ;
        RECT 279.795 17.535 280.095 17.605 ;
        RECT 279.82 17.605 280.165 17.63 ;
        RECT 279.875 17.63 280.19 17.685 ;
        RECT 279.93 17.685 280.19 17.74 ;
        RECT 279.93 17.74 280.19 36.3 ;
        RECT 279.93 36.3 280.19 36.31 ;
        RECT 279.92 36.31 280.19 36.32 ;
        RECT 279.91 36.32 280.19 36.41 ;
        RECT 279.91 36.41 280.18 36.42 ;
        RECT 279.91 36.42 280.17 36.43 ;
        RECT 279.91 36.43 280.17 45.48 ;
        RECT 279.91 45.48 280.17 45.535 ;
        RECT 279.91 45.535 280.225 45.59 ;
        RECT 279.98 45.59 280.28 45.66 ;
        RECT 280.05 45.66 280.35 45.73 ;
        RECT 280.12 45.73 280.42 45.8 ;
        RECT 280.17 45.8 280.49 45.85 ;
        RECT 280.225 45.85 280.54 45.905 ;
        RECT 280.28 45.905 280.54 45.96 ;
        RECT 280.28 45.96 280.54 46.565 ;
        RECT 280.28 46.565 280.54 46.62 ;
        RECT 280.28 46.62 280.595 46.675 ;
        RECT 280.35 46.675 280.65 46.745 ;
        RECT 280.42 46.745 280.72 46.815 ;
        RECT 280.49 46.815 280.79 46.885 ;
        RECT 280.56 46.885 280.86 46.955 ;
        RECT 280.63 46.955 280.93 47.025 ;
        RECT 280.7 47.025 281 47.095 ;
        RECT 280.77 47.095 281.07 47.165 ;
        RECT 280.84 47.165 281.14 47.235 ;
        RECT 280.91 47.235 281.21 47.305 ;
        RECT 280.98 47.305 281.28 47.375 ;
        RECT 281.05 47.375 281.35 47.445 ;
        RECT 281.065 47.445 281.42 47.46 ;
        RECT 281.12 47.46 281.435 47.515 ;
        RECT 281.175 47.515 281.435 47.57 ;
        RECT 281.175 56.455 281.435 56.51 ;
        RECT 281.12 56.51 281.435 56.565 ;
        RECT 281.065 56.565 281.365 56.635 ;
        RECT 280.995 56.635 281.295 56.705 ;
        RECT 280.925 56.705 281.225 56.775 ;
        RECT 280.855 56.775 281.155 56.845 ;
        RECT 280.785 56.845 281.085 56.915 ;
        RECT 280.715 56.915 281.015 56.985 ;
        RECT 280.645 56.985 280.945 57.055 ;
        RECT 280.575 57.055 280.875 57.125 ;
        RECT 280.505 57.125 280.805 57.195 ;
        RECT 280.435 57.195 280.735 57.265 ;
        RECT 280.365 57.265 280.68 57.32 ;
        RECT 280.365 57.32 280.625 57.375 ;
        RECT 280.365 57.375 280.625 74.88 ;
        RECT 280.365 74.88 280.625 74.935 ;
        RECT 280.365 74.935 280.68 74.99 ;
        RECT 280.435 74.99 280.735 75.06 ;
        RECT 280.505 75.06 280.805 75.13 ;
        RECT 280.575 75.13 280.875 75.2 ;
        RECT 280.645 75.2 280.945 75.27 ;
        RECT 280.715 75.27 281.015 75.34 ;
        RECT 280.785 75.34 281.085 75.41 ;
        RECT 280.855 75.41 281.155 75.48 ;
        RECT 280.925 75.48 281.225 75.55 ;
        RECT 280.995 75.55 281.295 75.62 ;
        RECT 281.065 75.62 281.365 75.69 ;
        RECT 281.135 75.69 281.435 75.76 ;
        RECT 281.205 75.76 281.505 75.83 ;
        RECT 281.275 75.83 281.575 75.9 ;
        RECT 281.345 75.9 281.645 75.97 ;
        RECT 281.415 75.97 281.715 76.04 ;
        RECT 281.485 76.04 281.785 76.11 ;
        RECT 281.555 76.11 281.855 76.18 ;
        RECT 281.625 76.18 281.925 76.25 ;
        RECT 281.695 76.25 281.995 76.32 ;
        RECT 281.765 76.32 282.065 76.39 ;
        RECT 281.835 76.39 282.135 76.46 ;
        RECT 281.885 76.46 282.205 76.51 ;
        RECT 281.94 76.51 282.255 76.565 ;
        RECT 281.995 76.565 282.255 76.62 ;
        RECT 281.995 76.62 282.255 87.54 ;
        RECT 281.995 87.54 282.255 87.595 ;
        RECT 281.995 87.595 282.31 87.65 ;
        RECT 282.065 87.65 282.365 87.72 ;
        RECT 282.135 87.72 282.435 87.79 ;
        RECT 282.205 87.79 282.505 87.86 ;
        RECT 282.275 87.86 282.575 87.93 ;
        RECT 282.345 87.93 282.645 88 ;
        RECT 282.415 88 282.715 88.07 ;
        RECT 282.485 88.07 282.785 88.14 ;
        RECT 282.555 88.14 282.855 88.21 ;
        RECT 282.625 88.21 282.925 88.28 ;
        RECT 282.695 88.28 282.995 88.35 ;
        RECT 282.765 88.35 283.065 88.42 ;
        RECT 282.835 88.42 283.135 88.49 ;
        RECT 282.905 88.49 283.205 88.56 ;
        RECT 282.975 88.56 283.275 88.63 ;
        RECT 283.045 88.63 283.345 88.7 ;
        RECT 283.115 88.7 283.415 88.77 ;
        RECT 283.185 88.77 283.485 88.84 ;
        RECT 283.255 88.84 283.555 88.91 ;
        RECT 283.325 88.91 283.625 88.98 ;
        RECT 283.395 88.98 283.695 89.05 ;
        RECT 283.465 89.05 283.765 89.12 ;
        RECT 283.535 89.12 283.835 89.19 ;
        RECT 283.605 89.19 283.905 89.26 ;
        RECT 283.675 89.26 283.975 89.33 ;
        RECT 283.745 89.33 284.045 89.4 ;
        RECT 283.815 89.4 284.115 89.47 ;
        RECT 283.825 89.47 284.185 89.48 ;
        RECT 283.865 89.48 284.195 89.52 ;
        RECT 283.905 89.52 284.195 89.56 ;
        RECT 283.91 89.56 284.195 89.565 ;
        RECT 283.91 89.565 284.195 94.165 ;
        RECT 283.91 94.165 284.195 94.205 ;
        RECT 283.91 94.205 284.235 94.245 ;
        RECT 283.91 94.245 284.275 94.25 ;
        RECT 283.98 94.25 284.28 94.32 ;
        RECT 284.05 94.32 284.35 94.39 ;
        RECT 284.12 94.39 284.42 94.46 ;
        RECT 284.19 94.46 284.49 94.53 ;
        RECT 284.26 94.53 284.56 94.6 ;
        RECT 284.33 94.6 284.63 94.67 ;
        RECT 284.36 94.67 284.7 94.7 ;
        RECT 284.43 94.7 289.415 94.77 ;
        RECT 284.5 94.77 289.485 94.84 ;
        RECT 284.57 94.84 289.555 94.91 ;
        RECT 284.62 94.91 289.625 94.96 ;
        RECT 297.33 102.94 297.655 102.985 ;
        RECT 297.285 102.87 297.585 102.94 ;
        RECT 297.215 102.8 297.515 102.87 ;
        RECT 297.145 102.73 297.445 102.8 ;
        RECT 297.075 102.66 297.375 102.73 ;
        RECT 297.005 102.59 297.305 102.66 ;
        RECT 296.935 102.52 297.235 102.59 ;
        RECT 296.865 102.45 297.165 102.52 ;
        RECT 296.795 102.38 297.095 102.45 ;
        RECT 296.725 102.31 297.025 102.38 ;
        RECT 296.655 102.24 296.955 102.31 ;
        RECT 296.585 102.17 296.885 102.24 ;
        RECT 296.515 102.1 296.815 102.17 ;
        RECT 296.445 102.03 296.745 102.1 ;
        RECT 296.375 101.96 296.675 102.03 ;
        RECT 296.305 101.89 296.605 101.96 ;
        RECT 296.235 101.82 296.535 101.89 ;
        RECT 296.165 101.75 296.465 101.82 ;
        RECT 296.095 101.68 296.395 101.75 ;
        RECT 296.025 101.61 296.325 101.68 ;
        RECT 295.955 101.54 296.255 101.61 ;
        RECT 295.885 101.47 296.185 101.54 ;
        RECT 295.815 101.4 296.115 101.47 ;
        RECT 295.745 101.33 296.045 101.4 ;
        RECT 295.675 101.26 295.975 101.33 ;
        RECT 295.605 101.19 295.905 101.26 ;
        RECT 295.535 101.12 295.835 101.19 ;
        RECT 295.465 101.05 295.765 101.12 ;
        RECT 295.395 100.98 295.695 101.05 ;
        RECT 295.325 100.91 295.625 100.98 ;
        RECT 295.255 100.84 295.555 100.91 ;
        RECT 295.185 100.77 295.485 100.84 ;
        RECT 295.115 100.7 295.415 100.77 ;
        RECT 295.045 100.63 295.345 100.7 ;
        RECT 294.975 100.56 295.275 100.63 ;
        RECT 294.905 100.49 295.205 100.56 ;
        RECT 294.835 100.42 295.135 100.49 ;
        RECT 294.765 100.35 295.065 100.42 ;
        RECT 294.695 100.28 294.995 100.35 ;
        RECT 294.625 100.21 294.925 100.28 ;
        RECT 294.555 100.14 294.855 100.21 ;
        RECT 294.485 100.07 294.785 100.14 ;
        RECT 294.415 100 294.715 100.07 ;
        RECT 294.345 99.93 294.645 100 ;
        RECT 294.275 99.86 294.575 99.93 ;
        RECT 294.205 99.79 294.505 99.86 ;
        RECT 294.135 99.72 294.435 99.79 ;
        RECT 294.065 99.65 294.365 99.72 ;
        RECT 293.995 99.58 294.295 99.65 ;
        RECT 293.925 99.51 294.225 99.58 ;
        RECT 293.855 99.44 294.155 99.51 ;
        RECT 293.785 99.37 294.085 99.44 ;
        RECT 293.715 99.3 294.015 99.37 ;
        RECT 293.645 99.23 293.945 99.3 ;
        RECT 293.575 99.16 293.875 99.23 ;
        RECT 293.505 99.09 293.805 99.16 ;
        RECT 293.435 99.02 293.735 99.09 ;
        RECT 293.365 98.95 293.665 99.02 ;
        RECT 293.295 98.88 293.595 98.95 ;
        RECT 293.225 98.81 293.525 98.88 ;
        RECT 293.155 98.74 293.455 98.81 ;
        RECT 293.085 98.67 293.385 98.74 ;
        RECT 293.015 98.6 293.315 98.67 ;
        RECT 292.945 98.53 293.245 98.6 ;
        RECT 292.875 98.46 293.175 98.53 ;
        RECT 292.805 98.39 293.105 98.46 ;
        RECT 292.735 98.32 293.035 98.39 ;
        RECT 292.665 98.25 292.965 98.32 ;
        RECT 292.595 98.18 292.895 98.25 ;
        RECT 292.525 98.11 292.825 98.18 ;
        RECT 292.455 98.04 292.755 98.11 ;
        RECT 292.385 97.97 292.685 98.04 ;
        RECT 292.315 97.9 292.615 97.97 ;
        RECT 292.245 97.83 292.545 97.9 ;
        RECT 292.175 97.76 292.475 97.83 ;
        RECT 292.105 97.69 292.405 97.76 ;
        RECT 292.035 97.62 292.335 97.69 ;
        RECT 291.965 97.55 292.265 97.62 ;
        RECT 291.895 97.48 292.195 97.55 ;
        RECT 291.825 97.41 292.125 97.48 ;
        RECT 291.755 97.34 292.055 97.41 ;
        RECT 291.685 97.27 291.985 97.34 ;
        RECT 291.615 97.2 291.915 97.27 ;
        RECT 291.545 97.13 291.845 97.2 ;
        RECT 291.475 97.06 291.775 97.13 ;
        RECT 291.405 96.99 291.705 97.06 ;
        RECT 291.335 96.92 291.635 96.99 ;
        RECT 291.265 96.85 291.565 96.92 ;
        RECT 291.195 96.78 291.495 96.85 ;
        RECT 291.125 96.71 291.425 96.78 ;
        RECT 291.055 96.64 291.355 96.71 ;
        RECT 290.985 96.57 291.285 96.64 ;
        RECT 290.915 96.5 291.215 96.57 ;
        RECT 290.845 96.43 291.145 96.5 ;
        RECT 290.775 96.36 291.075 96.43 ;
        RECT 290.705 96.29 291.005 96.36 ;
        RECT 290.635 96.22 290.935 96.29 ;
        RECT 290.565 96.15 290.865 96.22 ;
        RECT 290.495 96.08 290.795 96.15 ;
        RECT 290.425 96.01 290.725 96.08 ;
        RECT 290.355 95.94 290.655 96.01 ;
        RECT 290.285 95.87 290.585 95.94 ;
        RECT 290.215 95.8 290.515 95.87 ;
        RECT 290.145 95.73 290.445 95.8 ;
        RECT 290.075 95.66 290.375 95.73 ;
        RECT 290.005 95.59 290.305 95.66 ;
        RECT 289.935 95.52 290.235 95.59 ;
        RECT 289.865 95.45 290.165 95.52 ;
        RECT 289.795 95.38 290.095 95.45 ;
        RECT 289.725 95.31 290.025 95.38 ;
        RECT 289.655 95.24 289.955 95.31 ;
        RECT 289.585 95.17 289.885 95.24 ;
        RECT 289.515 95.1 289.815 95.17 ;
        RECT 289.445 95.03 289.745 95.1 ;
        RECT 289.375 94.96 289.675 95.03 ;
        RECT 297.37 102.985 297.7 103.025 ;
        RECT 297.41 103.025 297.7 103.065 ;
        RECT 297.41 111.375 297.7 111.435 ;
        RECT 297.35 111.435 297.7 111.495 ;
        RECT 297.29 111.495 297.7 111.5 ;
        RECT 281.175 47.57 281.435 56.455 ;
        RECT 296.66 111.5 297.7 111.6 ;
        RECT 296.66 111.6 297.63 111.67 ;
        RECT 296.66 111.67 297.56 111.74 ;
        RECT 296.66 111.74 297.54 111.76 ;
        RECT 296.66 111.9 296.92 112.14 ;
        RECT 296.66 111.76 296.99 111.83 ;
        RECT 296.66 111.83 296.92 111.9 ;
        RECT 297.41 103.065 297.7 111.375 ;
    END
    ANTENNAGATEAREA 2.4 LAYER met1 ;
    ANTENNAGATEAREA 2.4 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 186.303 LAYER met2 ;
    ANTENNAGATEAREA 2.4 LAYER met3 ;
    ANTENNAGATEAREA 2.4 LAYER met4 ;
    ANTENNAGATEAREA 2.4 LAYER met5 ;
  END tie_lo_esd[1]

  PIN out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.17 46.28 265.47 46.35 ;
        RECT 265.1 46.35 265.4 46.42 ;
        RECT 265.03 46.42 265.33 46.49 ;
        RECT 264.96 46.49 265.26 46.56 ;
        RECT 264.89 46.56 265.19 46.63 ;
        RECT 264.82 46.63 265.12 46.7 ;
        RECT 264.75 46.7 265.05 46.77 ;
        RECT 264.68 46.77 264.98 46.84 ;
        RECT 264.61 46.84 264.91 46.91 ;
        RECT 264.54 46.91 264.84 46.98 ;
        RECT 264.47 46.98 264.77 47.05 ;
        RECT 264.4 47.05 264.7 47.12 ;
        RECT 264.33 47.12 264.63 47.19 ;
        RECT 264.26 47.19 264.56 47.26 ;
        RECT 264.19 47.26 264.49 47.33 ;
        RECT 264.12 47.33 264.46 47.36 ;
        RECT 264.09 47.36 264.405 47.415 ;
        RECT 264.09 47.415 264.35 47.47 ;
        RECT 265.43 46.02 268.55 46.09 ;
        RECT 265.36 46.09 268.55 46.16 ;
        RECT 265.29 46.16 268.55 46.23 ;
        RECT 265.22 46.23 268.55 46.28 ;
        RECT 268.29 0 268.55 45.84 ;
        RECT 268.29 45.84 268.55 45.91 ;
        RECT 268.22 45.91 268.55 45.98 ;
        RECT 268.15 45.98 268.55 46.02 ;
        RECT 264.09 47.47 264.35 48.665 ;
        RECT 264.09 48.665 264.35 48.735 ;
        RECT 264.09 48.735 264.42 48.805 ;
        RECT 264.09 48.805 264.49 48.83 ;
        RECT 264.09 48.83 264.515 48.9 ;
        RECT 264.02 48.9 264.585 48.97 ;
        RECT 263.95 48.97 264.655 51.845 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 38.6826 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END out[1]

  PIN out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.535 46.28 124.835 46.35 ;
        RECT 124.605 46.35 124.905 46.42 ;
        RECT 124.675 46.42 124.975 46.49 ;
        RECT 124.745 46.49 125.045 46.56 ;
        RECT 124.815 46.56 125.115 46.63 ;
        RECT 124.885 46.63 125.185 46.7 ;
        RECT 124.955 46.7 125.255 46.77 ;
        RECT 125.025 46.77 125.325 46.84 ;
        RECT 125.095 46.84 125.395 46.91 ;
        RECT 125.165 46.91 125.465 46.98 ;
        RECT 125.235 46.98 125.535 47.05 ;
        RECT 125.305 47.05 125.605 47.12 ;
        RECT 125.375 47.12 125.675 47.19 ;
        RECT 125.445 47.19 125.745 47.26 ;
        RECT 125.515 47.26 125.815 47.33 ;
        RECT 125.545 47.33 125.885 47.36 ;
        RECT 125.6 47.36 125.915 47.415 ;
        RECT 125.655 47.415 125.915 47.47 ;
        RECT 121.455 46.02 124.575 46.09 ;
        RECT 121.455 46.09 124.645 46.16 ;
        RECT 121.455 46.16 124.715 46.23 ;
        RECT 121.455 46.23 124.785 46.28 ;
        RECT 121.455 0 121.715 45.84 ;
        RECT 121.455 45.84 121.715 45.91 ;
        RECT 121.455 45.91 121.785 45.98 ;
        RECT 121.455 45.98 121.855 46.02 ;
        RECT 125.655 47.47 125.915 48.665 ;
        RECT 125.655 48.665 125.915 48.735 ;
        RECT 125.585 48.735 125.915 48.805 ;
        RECT 125.515 48.805 125.915 48.83 ;
        RECT 125.49 48.83 125.915 48.9 ;
        RECT 125.42 48.9 125.985 48.97 ;
        RECT 125.35 48.97 126.055 51.845 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 38.6826 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END out[0]

  PIN vtrip_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.125 0 128.385 10.065 ;
        RECT 128.125 10.065 128.385 10.12 ;
        RECT 128.07 10.12 128.385 10.175 ;
        RECT 128.015 10.175 128.315 10.245 ;
        RECT 127.945 10.245 128.245 10.315 ;
        RECT 127.875 10.315 128.175 10.385 ;
        RECT 127.805 10.385 128.105 10.455 ;
        RECT 127.735 10.455 128.035 10.525 ;
        RECT 127.665 10.525 127.965 10.595 ;
        RECT 127.595 10.595 127.895 10.665 ;
        RECT 127.525 10.665 127.825 10.735 ;
        RECT 127.455 10.735 127.755 10.805 ;
        RECT 127.385 10.805 127.685 10.875 ;
        RECT 127.315 10.875 127.63 10.93 ;
        RECT 127.26 10.93 127.575 10.985 ;
        RECT 127.26 10.985 127.52 11.04 ;
        RECT 127.26 11.04 127.52 23.665 ;
        RECT 127.26 23.665 127.52 23.72 ;
        RECT 127.26 23.72 127.575 23.775 ;
        RECT 127.33 23.775 127.63 23.845 ;
        RECT 127.4 23.845 127.7 23.915 ;
        RECT 127.47 23.915 127.77 23.985 ;
        RECT 127.54 23.985 127.84 24.055 ;
        RECT 127.61 24.055 127.91 24.125 ;
        RECT 127.68 24.125 127.98 24.195 ;
        RECT 127.75 24.195 128.05 24.265 ;
        RECT 127.805 24.265 128.12 24.32 ;
        RECT 127.86 24.32 128.12 24.375 ;
        RECT 127.86 42.525 128.12 42.585 ;
        RECT 127.86 42.585 128.18 42.645 ;
        RECT 127.86 42.645 128.24 42.65 ;
        RECT 127.86 42.65 128.88 42.91 ;
        RECT 127.86 24.375 128.12 42.525 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.7546 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END vtrip_sel[0]

  PIN vtrip_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.62 0 261.88 10.065 ;
        RECT 261.62 10.065 261.88 10.12 ;
        RECT 261.62 10.12 261.935 10.175 ;
        RECT 261.69 10.175 261.99 10.245 ;
        RECT 261.76 10.245 262.06 10.315 ;
        RECT 261.83 10.315 262.13 10.385 ;
        RECT 261.9 10.385 262.2 10.455 ;
        RECT 261.97 10.455 262.27 10.525 ;
        RECT 262.04 10.525 262.34 10.595 ;
        RECT 262.11 10.595 262.41 10.665 ;
        RECT 262.18 10.665 262.48 10.735 ;
        RECT 262.25 10.735 262.55 10.805 ;
        RECT 262.32 10.805 262.62 10.875 ;
        RECT 262.375 10.875 262.69 10.93 ;
        RECT 262.43 10.93 262.745 10.985 ;
        RECT 262.485 10.985 262.745 11.04 ;
        RECT 262.485 11.04 262.745 23.665 ;
        RECT 262.485 23.665 262.745 23.72 ;
        RECT 262.43 23.72 262.745 23.775 ;
        RECT 262.375 23.775 262.675 23.845 ;
        RECT 262.305 23.845 262.605 23.915 ;
        RECT 262.235 23.915 262.535 23.985 ;
        RECT 262.165 23.985 262.465 24.055 ;
        RECT 262.095 24.055 262.395 24.125 ;
        RECT 262.025 24.125 262.325 24.195 ;
        RECT 261.955 24.195 262.255 24.265 ;
        RECT 261.885 24.265 262.2 24.32 ;
        RECT 261.885 24.32 262.145 24.375 ;
        RECT 261.885 42.525 262.145 42.585 ;
        RECT 261.825 42.585 262.145 42.645 ;
        RECT 261.765 42.645 262.145 42.65 ;
        RECT 261.125 42.65 262.145 42.91 ;
        RECT 261.885 24.375 262.145 42.525 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.7546 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END vtrip_sel[1]

  PIN dm1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.765 0 234.025 33.835 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.6449 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END dm1[1]

  PIN dm1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.935 41.985 236.195 41.99 ;
        RECT 235.93 41.99 236.195 41.995 ;
        RECT 235.925 41.995 236.195 42.095 ;
        RECT 235.925 42.095 236.19 42.1 ;
        RECT 235.925 42.1 236.185 42.105 ;
        RECT 235.935 0 236.195 41.985 ;
        RECT 235.925 42.105 236.185 42.91 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.7774 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END dm1[2]

  PIN dm1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.365 0 233.625 33.095 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.6139 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END dm1[0]

  PIN enable_h
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.335 2.19 236.595 2.21 ;
        RECT 236.335 2.21 236.615 2.23 ;
        RECT 236.335 2.23 236.635 2.235 ;
        RECT 236.335 0 236.595 2.19 ;
        RECT 236.335 2.235 236.64 3.005 ;
        RECT 236.335 3.005 236.62 3.025 ;
        RECT 236.335 3.025 236.6 3.045 ;
        RECT 236.335 3.045 236.595 3.05 ;
        RECT 236.335 3.05 236.595 34.945 ;
    END
    PORT
      LAYER met2 ;
        RECT 153.39 2.235 153.67 3.005 ;
        RECT 153.41 2.215 153.67 2.225 ;
        RECT 153.4 2.225 153.67 2.235 ;
        RECT 153.41 0 153.67 2.215 ;
        RECT 153.4 3.005 153.67 3.015 ;
        RECT 153.41 3.015 153.67 3.025 ;
        RECT 153.41 3.025 153.67 34.945 ;
    END
    ANTENNAGATEAREA 10.8 LAYER met1 ;
    ANTENNAGATEAREA 10.8 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.2048 LAYER met2 ;
    ANTENNAGATEAREA 29.4 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 484.29 LAYER met3 ;
    ANTENNAGATEAREA 10.8 LAYER met4 ;
    ANTENNAGATEAREA 10.8 LAYER met5 ;
    ANTENNAPARTIALCUTAREA 0.24 LAYER via2 ;
  END enable_h

  PIN vreg_en[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.805 0 150.065 27.875 ;
        RECT 149.805 27.875 150.065 27.945 ;
        RECT 149.805 27.945 150.135 28.015 ;
        RECT 149.805 28.015 150.205 28.085 ;
        RECT 149.805 28.085 150.275 28.155 ;
        RECT 149.805 28.155 150.345 28.225 ;
        RECT 149.805 28.225 150.415 28.25 ;
        RECT 149.875 28.25 150.44 28.32 ;
        RECT 149.945 28.32 150.51 28.39 ;
        RECT 149.97 28.39 150.58 28.415 ;
        RECT 150.04 28.415 150.605 28.485 ;
        RECT 150.11 28.485 150.605 28.555 ;
        RECT 150.18 28.555 150.605 28.625 ;
        RECT 150.25 28.625 150.605 28.695 ;
        RECT 150.32 28.695 150.605 28.765 ;
        RECT 150.345 28.765 150.605 28.79 ;
        RECT 150.345 28.79 150.605 30.725 ;
        RECT 150.345 30.725 150.605 30.795 ;
        RECT 150.275 30.795 150.605 30.865 ;
        RECT 150.205 30.865 150.605 30.935 ;
        RECT 150.135 30.935 150.605 31.005 ;
        RECT 150.065 31.005 150.605 31.075 ;
        RECT 149.995 31.075 150.605 31.1 ;
        RECT 149.97 31.1 150.535 31.17 ;
        RECT 149.9 31.17 150.465 31.24 ;
        RECT 149.83 31.24 150.44 31.265 ;
        RECT 149.805 31.265 150.37 31.335 ;
        RECT 149.805 31.335 150.3 31.405 ;
        RECT 149.805 31.405 150.23 31.475 ;
        RECT 149.805 31.475 150.16 31.545 ;
        RECT 149.805 31.545 150.09 31.615 ;
        RECT 149.805 31.615 150.065 31.64 ;
        RECT 149.805 31.64 150.065 58.14 ;
        RECT 149.805 58.14 150.065 58.2 ;
        RECT 149.805 58.2 150.125 58.26 ;
        RECT 149.805 58.26 150.185 58.265 ;
        RECT 149.805 58.265 150.445 58.525 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 43.929 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END vreg_en[0]

  PIN vreg_en[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.94 0 240.2 27.875 ;
        RECT 239.94 27.875 240.2 27.945 ;
        RECT 239.87 27.945 240.2 28.015 ;
        RECT 239.8 28.015 240.2 28.085 ;
        RECT 239.73 28.085 240.2 28.155 ;
        RECT 239.66 28.155 240.2 28.225 ;
        RECT 239.59 28.225 240.2 28.25 ;
        RECT 239.565 28.25 240.13 28.32 ;
        RECT 239.495 28.32 240.06 28.39 ;
        RECT 239.425 28.39 240.035 28.415 ;
        RECT 239.4 28.415 239.965 28.485 ;
        RECT 239.4 28.485 239.895 28.555 ;
        RECT 239.4 28.555 239.825 28.625 ;
        RECT 239.4 28.625 239.755 28.695 ;
        RECT 239.4 28.695 239.685 28.765 ;
        RECT 239.4 28.765 239.66 28.79 ;
        RECT 239.4 28.79 239.66 30.725 ;
        RECT 239.4 30.725 239.66 30.795 ;
        RECT 239.4 30.795 239.73 30.865 ;
        RECT 239.4 30.865 239.8 30.935 ;
        RECT 239.4 30.935 239.87 31.005 ;
        RECT 239.4 31.005 239.94 31.075 ;
        RECT 239.4 31.075 240.01 31.1 ;
        RECT 239.47 31.1 240.035 31.17 ;
        RECT 239.54 31.17 240.105 31.24 ;
        RECT 239.565 31.24 240.175 31.265 ;
        RECT 239.635 31.265 240.2 31.335 ;
        RECT 239.705 31.335 240.2 31.405 ;
        RECT 239.775 31.405 240.2 31.475 ;
        RECT 239.845 31.475 240.2 31.545 ;
        RECT 239.915 31.545 240.2 31.615 ;
        RECT 239.94 31.615 240.2 31.64 ;
        RECT 239.94 31.64 240.2 58.14 ;
        RECT 239.94 58.14 240.2 58.2 ;
        RECT 239.88 58.2 240.2 58.26 ;
        RECT 239.82 58.26 240.2 58.265 ;
        RECT 239.56 58.265 240.2 58.525 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 43.929 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END vreg_en[1]

  PIN slow[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.13 0 242.39 46.135 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 40.264 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END slow[1]

  PIN slow[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.615 0 147.875 46.135 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 40.264 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END slow[0]

  PIN oe_n[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.215 0 147.475 26.81 ;
        RECT 147.215 26.81 147.475 26.865 ;
        RECT 147.16 26.865 147.475 26.92 ;
        RECT 147.105 26.92 147.405 26.99 ;
        RECT 147.035 26.99 147.335 27.06 ;
        RECT 146.965 27.06 147.265 27.13 ;
        RECT 146.895 27.13 147.195 27.2 ;
        RECT 146.825 27.2 147.125 27.27 ;
        RECT 146.755 27.27 147.055 27.34 ;
        RECT 146.685 27.34 146.985 27.41 ;
        RECT 146.615 27.41 146.915 27.48 ;
        RECT 146.545 27.48 146.845 27.55 ;
        RECT 146.475 27.55 146.775 27.62 ;
        RECT 146.405 27.62 146.705 27.69 ;
        RECT 146.335 27.69 146.635 27.76 ;
        RECT 146.265 27.76 146.565 27.83 ;
        RECT 146.195 27.83 146.495 27.9 ;
        RECT 146.125 27.9 146.425 27.97 ;
        RECT 146.055 27.97 146.355 28.04 ;
        RECT 145.985 28.04 146.285 28.11 ;
        RECT 145.915 28.11 146.215 28.18 ;
        RECT 145.845 28.18 146.145 28.25 ;
        RECT 145.775 28.25 146.075 28.32 ;
        RECT 145.705 28.32 146.005 28.39 ;
        RECT 145.635 28.39 145.95 28.445 ;
        RECT 145.635 28.445 145.895 28.5 ;
        RECT 145.635 28.5 145.895 49.23 ;
        RECT 145.635 49.23 145.895 49.29 ;
        RECT 145.575 49.29 145.895 49.35 ;
        RECT 145.515 49.35 145.895 49.355 ;
        RECT 145.255 49.355 145.895 49.615 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 37.6305 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END oe_n[0]

  PIN oe_n[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.53 0 242.79 26.81 ;
        RECT 242.53 26.81 242.79 26.865 ;
        RECT 242.53 26.865 242.845 26.92 ;
        RECT 242.6 26.92 242.9 26.99 ;
        RECT 242.67 26.99 242.97 27.06 ;
        RECT 242.74 27.06 243.04 27.13 ;
        RECT 242.81 27.13 243.11 27.2 ;
        RECT 242.88 27.2 243.18 27.27 ;
        RECT 242.95 27.27 243.25 27.34 ;
        RECT 243.02 27.34 243.32 27.41 ;
        RECT 243.09 27.41 243.39 27.48 ;
        RECT 243.16 27.48 243.46 27.55 ;
        RECT 243.23 27.55 243.53 27.62 ;
        RECT 243.3 27.62 243.6 27.69 ;
        RECT 243.37 27.69 243.67 27.76 ;
        RECT 243.44 27.76 243.74 27.83 ;
        RECT 243.51 27.83 243.81 27.9 ;
        RECT 243.58 27.9 243.88 27.97 ;
        RECT 243.65 27.97 243.95 28.04 ;
        RECT 243.72 28.04 244.02 28.11 ;
        RECT 243.79 28.11 244.09 28.18 ;
        RECT 243.86 28.18 244.16 28.25 ;
        RECT 243.93 28.25 244.23 28.32 ;
        RECT 244 28.32 244.3 28.39 ;
        RECT 244.055 28.39 244.37 28.445 ;
        RECT 244.11 28.445 244.37 28.5 ;
        RECT 244.11 28.5 244.37 49.23 ;
        RECT 244.11 49.23 244.37 49.29 ;
        RECT 244.11 49.29 244.43 49.35 ;
        RECT 244.11 49.35 244.49 49.355 ;
        RECT 244.11 49.355 244.75 49.615 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 37.6305 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END oe_n[1]

  PIN dm0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.38 0 156.64 33.095 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.6139 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END dm0[0]

  PIN dm0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.98 0 156.24 33.835 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.6449 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END dm0[1]

  PIN dm0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.81 41.985 154.07 41.99 ;
        RECT 153.81 41.99 154.075 41.995 ;
        RECT 153.81 41.995 154.08 42.095 ;
        RECT 153.815 42.095 154.08 42.1 ;
        RECT 153.82 42.1 154.08 42.105 ;
        RECT 153.81 0 154.07 41.985 ;
        RECT 153.82 42.105 154.08 42.91 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.7774 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END dm0[2]

  PIN in_h[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.34 0 247.6 10.59 ;
    END
    ANTENNADIFFAREA 4.435 LAYER met1 ;
    ANTENNADIFFAREA 4.435 LAYER met2 ;
    ANTENNADIFFAREA 4.435 LAYER met3 ;
    ANTENNADIFFAREA 4.435 LAYER met4 ;
    ANTENNADIFFAREA 4.435 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1995 LAYER met2 ;
  END in_h[1]

  PIN in_h[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.405 0 142.665 10.59 ;
    END
    ANTENNADIFFAREA 4.435 LAYER met1 ;
    ANTENNADIFFAREA 4.435 LAYER met2 ;
    ANTENNADIFFAREA 4.435 LAYER met3 ;
    ANTENNADIFFAREA 4.435 LAYER met4 ;
    ANTENNADIFFAREA 4.435 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.1995 LAYER met2 ;
  END in_h[0]

  PIN in[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.005 0 142.265 7.58 ;
    END
    ANTENNADIFFAREA 2.225 LAYER met1 ;
    ANTENNADIFFAREA 2.225 LAYER met2 ;
    ANTENNADIFFAREA 2.225 LAYER met3 ;
    ANTENNADIFFAREA 2.225 LAYER met4 ;
    ANTENNADIFFAREA 2.225 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 11.3144 LAYER met2 ;
  END in[0]

  PIN in[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.74 0 248 7.58 ;
    END
    ANTENNADIFFAREA 2.225 LAYER met1 ;
    ANTENNADIFFAREA 2.225 LAYER met2 ;
    ANTENNADIFFAREA 2.225 LAYER met3 ;
    ANTENNADIFFAREA 2.225 LAYER met4 ;
    ANTENNADIFFAREA 2.225 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 11.3144 LAYER met2 ;
  END in[1]

  PIN hld_ovr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.46 0 248.805 1.88 ;
        RECT 248.46 1.88 248.805 1.935 ;
        RECT 248.46 1.935 248.86 1.99 ;
        RECT 248.46 1.99 248.915 1.995 ;
        RECT 248.46 1.995 248.92 2.04 ;
        RECT 248.415 2.04 248.965 2.085 ;
        RECT 248.37 2.085 249.01 2.345 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.7736 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END hld_ovr[1]

  PIN hld_ovr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.2 0 141.545 1.88 ;
        RECT 141.2 1.88 141.545 1.935 ;
        RECT 141.145 1.935 141.545 1.99 ;
        RECT 141.09 1.99 141.545 1.995 ;
        RECT 141.085 1.995 141.545 2.04 ;
        RECT 141.04 2.04 141.59 2.085 ;
        RECT 140.995 2.085 141.635 2.345 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.7736 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END hld_ovr[0]

  PIN hld_h_n[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.17 36.69 254.81 36.95 ;
        RECT 254.17 36.565 254.43 36.625 ;
        RECT 254.17 36.625 254.49 36.685 ;
        RECT 254.17 36.685 254.55 36.69 ;
        RECT 254.17 0 254.43 36.565 ;
    END
    ANTENNAGATEAREA 2.4 LAYER met1 ;
    ANTENNAGATEAREA 2.4 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.8919 LAYER met2 ;
    ANTENNAGATEAREA 2.4 LAYER met3 ;
    ANTENNAGATEAREA 2.4 LAYER met4 ;
    ANTENNAGATEAREA 2.4 LAYER met5 ;
  END hld_h_n[1]

  PIN hld_h_n[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.195 36.69 135.835 36.95 ;
        RECT 135.575 36.565 135.835 36.625 ;
        RECT 135.515 36.625 135.835 36.685 ;
        RECT 135.455 36.685 135.835 36.69 ;
        RECT 135.575 0 135.835 36.565 ;
    END
    ANTENNAGATEAREA 2.4 LAYER met1 ;
    ANTENNAGATEAREA 2.4 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 25.8919 LAYER met2 ;
    ANTENNAGATEAREA 2.4 LAYER met3 ;
    ANTENNAGATEAREA 2.4 LAYER met4 ;
    ANTENNAGATEAREA 2.4 LAYER met5 ;
  END hld_h_n[0]

  PIN ibuf_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.175 0 135.435 28.84 ;
        RECT 135.175 28.84 135.435 28.895 ;
        RECT 135.12 28.895 135.435 28.95 ;
        RECT 135.065 28.95 135.365 29.02 ;
        RECT 134.995 29.02 135.295 29.09 ;
        RECT 134.925 29.09 135.225 29.16 ;
        RECT 134.855 29.16 135.155 29.23 ;
        RECT 134.785 29.23 135.085 29.3 ;
        RECT 134.715 29.3 135.015 29.37 ;
        RECT 134.645 29.37 134.96 29.425 ;
        RECT 134.645 29.425 134.905 29.48 ;
        RECT 134.645 29.48 134.905 29.86 ;
        RECT 134.645 29.86 134.905 29.915 ;
        RECT 134.59 29.915 134.905 29.97 ;
        RECT 134.535 29.97 134.9 29.975 ;
        RECT 134.53 29.975 134.895 29.98 ;
        RECT 134.525 29.98 134.89 29.985 ;
        RECT 133.755 29.985 134.82 30.055 ;
        RECT 133.755 30.055 134.75 30.125 ;
        RECT 133.755 30.125 134.68 30.195 ;
        RECT 133.755 30.195 134.63 30.245 ;
        RECT 134.07 30.245 134.46 30.305 ;
        RECT 134.13 30.305 134.4 30.365 ;
        RECT 134.135 30.365 134.395 30.37 ;
        RECT 134.135 30.37 134.395 42.74 ;
    END
    ANTENNAGATEAREA 0.72 LAYER met1 ;
    ANTENNAGATEAREA 0.72 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.3479 LAYER met2 ;
    ANTENNAGATEAREA 0.72 LAYER met3 ;
    ANTENNAGATEAREA 0.72 LAYER met4 ;
    ANTENNAGATEAREA 0.72 LAYER met5 ;
  END ibuf_sel[0]

  PIN amuxbus_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0 102.08 480 105.06 ;
    END
    PORT
      LAYER met2 ;
        RECT 448.655 0 448.915 83.36 ;
    END
    ANTENNADIFFAREA 2.65 LAYER met1 ;
    ANTENNADIFFAREA 2.65 LAYER met2 ;
    ANTENNADIFFAREA 2.65 LAYER met3 ;
    ANTENNADIFFAREA 2.65 LAYER met4 ;
    ANTENNADIFFAREA 2.65 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 72.1229 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.775 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 772.768 LAYER met4 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3 ;
  END amuxbus_b

  PIN amuxbus_a
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0 106.84 480 109.82 ;
    END
    PORT
      LAYER met2 ;
        RECT 447.905 0 448.165 83.36 ;
    END
    ANTENNADIFFAREA 2.65 LAYER met1 ;
    ANTENNADIFFAREA 2.65 LAYER met2 ;
    ANTENNADIFFAREA 2.65 LAYER met3 ;
    ANTENNADIFFAREA 2.65 LAYER met4 ;
    ANTENNADIFFAREA 2.65 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 75.4549 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.256 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 772.768 LAYER met4 ;
    ANTENNAPARTIALCUTAREA 0.28 LAYER via2 ;
    ANTENNAPARTIALCUTAREA 0.28 LAYER via3 ;
  END amuxbus_a

  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 62.7 480 67.15 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 62.6 480 67.25 ;
    END
  END vccd

  PIN vcchib
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 55.85 480 61.1 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 55.75 480 61.2 ;
    END
  END vcchib

  PIN vdda
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 68.75 480 72 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 68.65 480 72.1 ;
    END
  END vdda

  PIN vddio
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 73.6 480 78.05 ;
    END
    PORT
      LAYER met5 ;
        RECT 18.77 148.715 53.78 148.895 ;
        RECT 18.95 148.895 53.96 149.075 ;
        RECT 18.955 149.075 54.14 149.08 ;
        RECT 19.355 149.08 54.145 149.48 ;
        RECT 19.755 149.48 54.145 149.88 ;
        RECT 20.155 149.88 54.145 150.28 ;
        RECT 20.555 150.28 54.145 150.68 ;
        RECT 20.955 150.68 54.145 151.08 ;
        RECT 21.355 151.08 54.145 151.48 ;
        RECT 21.755 151.48 54.145 151.88 ;
        RECT 22.155 151.88 54.145 152.28 ;
        RECT 22.555 152.28 54.145 152.68 ;
        RECT 22.955 152.68 54.145 153.08 ;
        RECT 23.355 153.08 54.145 153.48 ;
        RECT 23.755 153.48 54.145 153.88 ;
        RECT 24.155 153.88 54.145 154.28 ;
        RECT 24.555 154.28 54.145 154.68 ;
        RECT 24.955 154.68 54.145 155.08 ;
        RECT 25.355 155.08 54.145 155.48 ;
        RECT 25.755 155.48 54.145 155.88 ;
        RECT 26.155 155.88 54.145 156.28 ;
        RECT 26.555 156.28 54.145 156.68 ;
        RECT 26.955 156.68 54.145 157.08 ;
        RECT 27.355 157.08 54.145 157.48 ;
        RECT 27.755 157.48 54.145 157.88 ;
        RECT 28.155 157.88 54.145 158.28 ;
        RECT 28.555 158.28 54.145 158.68 ;
        RECT 28.955 158.68 54.145 159.08 ;
        RECT 29.26 159.08 54.145 159.385 ;
        RECT 29.26 159.385 54.145 197.6 ;
        RECT 29.26 197.6 54.145 198 ;
        RECT 29.26 198 54.545 198.4 ;
        RECT 29.26 198.4 54.945 198.8 ;
        RECT 29.26 198.8 55.345 199.2 ;
        RECT 29.26 199.2 55.745 199.6 ;
        RECT 29.26 199.6 56.145 200 ;
        RECT 29.26 200 56.545 200.4 ;
        RECT 29.26 200.4 56.945 200.8 ;
        RECT 29.26 200.8 57.345 201.2 ;
        RECT 29.26 201.2 57.745 201.6 ;
        RECT 29.26 201.6 58.145 202 ;
        RECT 29.26 202 58.545 202.4 ;
        RECT 29.26 202.4 58.945 202.8 ;
        RECT 29.26 202.8 59.345 203.2 ;
        RECT 29.26 203.2 59.745 203.6 ;
        RECT 29.26 203.6 60.145 204 ;
        RECT 29.26 204 60.545 204.4 ;
        RECT 29.26 204.4 60.945 204.49 ;
        RECT 29.26 204.49 422.295 204.89 ;
        RECT 29.26 204.89 421.895 205.29 ;
        RECT 29.26 205.29 421.495 205.69 ;
        RECT 29.26 205.69 421.095 206.09 ;
        RECT 29.26 206.09 420.695 206.49 ;
        RECT 29.26 206.49 420.295 206.89 ;
        RECT 29.26 206.89 419.895 207.29 ;
        RECT 29.26 207.29 419.86 207.325 ;
        RECT 29.66 207.325 419.46 207.725 ;
        RECT 30.06 207.725 419.06 208.125 ;
        RECT 30.46 208.125 418.66 208.525 ;
        RECT 30.86 208.525 418.26 208.925 ;
        RECT 31.26 208.925 417.86 209.325 ;
        RECT 31.66 209.325 417.46 209.725 ;
        RECT 32.06 209.725 417.06 210.125 ;
        RECT 32.46 210.125 416.66 210.525 ;
        RECT 32.86 210.525 416.26 210.925 ;
        RECT 33.26 210.925 415.86 211.325 ;
        RECT 33.66 211.325 415.46 211.725 ;
        RECT 34.06 211.725 415.06 212.125 ;
        RECT 34.46 212.125 414.66 212.525 ;
        RECT 34.86 212.525 414.26 212.925 ;
        RECT 35.26 212.925 413.86 213.325 ;
        RECT 35.66 213.325 413.46 213.725 ;
        RECT 36.06 213.725 413.06 214.125 ;
        RECT 36.46 214.125 412.66 214.525 ;
        RECT 36.86 214.525 412.26 214.925 ;
        RECT 37.26 214.925 411.86 215.325 ;
        RECT 37.66 215.325 411.46 215.725 ;
        RECT 38.06 215.725 411.06 216.125 ;
        RECT 38.46 216.125 410.66 216.525 ;
        RECT 38.86 216.525 410.26 216.925 ;
        RECT 39.26 216.925 409.86 217.325 ;
        RECT 39.66 217.325 409.46 217.725 ;
        RECT 40.06 217.725 409.06 218.125 ;
        RECT 40.46 218.125 408.66 218.525 ;
        RECT 40.86 218.525 408.26 218.925 ;
        RECT 41.26 218.925 407.86 219.325 ;
        RECT 41.66 219.325 407.46 219.725 ;
        RECT 42.06 219.725 407.06 220.125 ;
        RECT 42.46 220.125 406.66 220.525 ;
        RECT 42.86 220.525 406.26 220.925 ;
        RECT 43.26 220.925 405.86 221.325 ;
        RECT 43.66 221.325 405.46 221.725 ;
        RECT 44.06 221.725 405.06 222.125 ;
        RECT 44.46 222.125 404.66 222.525 ;
        RECT 44.86 222.525 404.26 222.925 ;
        RECT 45.26 222.925 403.86 223.325 ;
        RECT 45.66 223.325 403.46 223.725 ;
        RECT 46.06 223.725 403.06 224.125 ;
        RECT 46.46 224.125 402.66 224.525 ;
        RECT 46.86 224.525 402.26 224.925 ;
        RECT 47.26 224.925 401.86 225.325 ;
        RECT 47.66 225.325 401.46 225.725 ;
        RECT 48.06 225.725 401.06 226.125 ;
        RECT 48.46 226.125 400.66 226.525 ;
        RECT 48.86 226.525 400.26 226.925 ;
        RECT 49.26 226.925 399.86 227.325 ;
        RECT 49.66 227.325 399.46 227.725 ;
        RECT 49.835 227.725 399.285 227.9 ;
        RECT 0 145.925 50.99 146.325 ;
        RECT 0 146.325 51.39 146.725 ;
        RECT 0 146.725 51.79 147.125 ;
        RECT 0 147.125 52.19 147.525 ;
        RECT 0 147.525 52.59 147.925 ;
        RECT 0 147.925 52.99 148.325 ;
        RECT 0 148.325 53.39 148.715 ;
        RECT 0 145.905 50.99 145.925 ;
        RECT 0 133.35 38.48 133.415 ;
        RECT 388.29 204.17 422.695 204.49 ;
        RECT 388.69 203.77 423.015 204.17 ;
        RECT 389.09 203.37 423.415 203.77 ;
        RECT 389.49 202.97 423.815 203.37 ;
        RECT 389.89 202.57 424.215 202.97 ;
        RECT 390.29 202.17 424.615 202.57 ;
        RECT 390.69 201.77 425.015 202.17 ;
        RECT 391.09 201.37 425.415 201.77 ;
        RECT 391.49 200.97 425.815 201.37 ;
        RECT 391.89 200.57 426.215 200.97 ;
        RECT 392.29 200.17 426.615 200.57 ;
        RECT 392.69 199.77 427.015 200.17 ;
        RECT 393.09 199.37 427.415 199.77 ;
        RECT 393.49 198.97 427.815 199.37 ;
        RECT 393.89 198.57 428.215 198.97 ;
        RECT 394.29 198.17 428.615 198.57 ;
        RECT 394.69 197.77 429.015 198.17 ;
        RECT 395.09 197.37 429.415 197.77 ;
        RECT 395.49 196.97 429.815 197.37 ;
        RECT 395.89 196.57 430.215 196.97 ;
        RECT 396.29 196.17 430.615 196.57 ;
        RECT 396.69 195.77 431.015 196.17 ;
        RECT 397.09 195.37 431.415 195.77 ;
        RECT 397.49 194.97 431.815 195.37 ;
        RECT 397.89 194.57 432.215 194.97 ;
        RECT 398.29 194.17 432.615 194.57 ;
        RECT 398.69 193.77 433.015 194.17 ;
        RECT 399.09 193.37 433.415 193.77 ;
        RECT 399.49 192.97 433.815 193.37 ;
        RECT 399.89 192.57 434.215 192.97 ;
        RECT 400.29 192.17 434.615 192.57 ;
        RECT 400.69 191.77 435.015 192.17 ;
        RECT 401.09 191.37 435.415 191.77 ;
        RECT 401.49 190.97 435.815 191.37 ;
        RECT 401.89 190.57 436.215 190.97 ;
        RECT 402.29 190.17 436.615 190.57 ;
        RECT 402.69 189.77 437.015 190.17 ;
        RECT 403.09 189.37 437.415 189.77 ;
        RECT 403.49 188.97 437.815 189.37 ;
        RECT 403.89 188.57 438.215 188.97 ;
        RECT 404.29 188.17 438.615 188.57 ;
        RECT 404.69 187.77 439.015 188.17 ;
        RECT 405.09 187.37 439.415 187.77 ;
        RECT 405.49 186.97 439.815 187.37 ;
        RECT 405.89 186.57 440.215 186.97 ;
        RECT 406.29 186.17 440.615 186.57 ;
        RECT 406.69 185.77 441.015 186.17 ;
        RECT 407.09 185.37 441.415 185.77 ;
        RECT 407.49 184.97 441.815 185.37 ;
        RECT 407.89 184.57 442.215 184.97 ;
        RECT 408.29 184.17 442.615 184.57 ;
        RECT 408.69 183.77 443.015 184.17 ;
        RECT 409.09 183.37 443.415 183.77 ;
        RECT 409.49 182.97 443.815 183.37 ;
        RECT 409.89 182.57 444.215 182.97 ;
        RECT 410.29 182.17 444.615 182.57 ;
        RECT 410.69 181.77 445.015 182.17 ;
        RECT 411.09 181.37 445.415 181.77 ;
        RECT 411.49 180.97 445.815 181.37 ;
        RECT 411.89 180.57 446.215 180.97 ;
        RECT 412.29 180.17 446.615 180.57 ;
        RECT 412.69 179.77 447.015 180.17 ;
        RECT 413.09 179.37 447.415 179.77 ;
        RECT 413.49 178.97 447.815 179.37 ;
        RECT 413.89 178.57 448.215 178.97 ;
        RECT 414.29 178.17 448.615 178.57 ;
        RECT 414.69 177.77 449.015 178.17 ;
        RECT 415.09 177.37 449.415 177.77 ;
        RECT 415.49 176.97 449.815 177.37 ;
        RECT 415.89 176.57 450.215 176.97 ;
        RECT 416.29 176.17 450.615 176.57 ;
        RECT 416.69 175.77 451.015 176.17 ;
        RECT 417.09 175.37 451.415 175.77 ;
        RECT 417.49 174.97 451.815 175.37 ;
        RECT 417.89 174.57 452.215 174.97 ;
        RECT 418.29 174.17 452.615 174.57 ;
        RECT 418.69 173.77 453.015 174.17 ;
        RECT 419.09 173.37 453.415 173.77 ;
        RECT 419.49 172.97 453.815 173.37 ;
        RECT 419.89 172.57 454.215 172.97 ;
        RECT 420.29 172.17 454.615 172.57 ;
        RECT 420.69 171.77 455.015 172.17 ;
        RECT 421.09 171.37 455.415 171.77 ;
        RECT 421.49 170.97 455.815 171.37 ;
        RECT 421.89 170.57 456.215 170.97 ;
        RECT 422.29 170.17 456.615 170.57 ;
        RECT 422.69 169.77 457.015 170.17 ;
        RECT 423.09 169.37 457.415 169.77 ;
        RECT 423.49 168.97 457.815 169.37 ;
        RECT 423.89 168.57 458.215 168.97 ;
        RECT 424.29 168.17 458.615 168.57 ;
        RECT 424.69 167.77 459.015 168.17 ;
        RECT 425.09 167.37 459.415 167.77 ;
        RECT 425.49 166.97 459.815 167.37 ;
        RECT 425.89 166.57 460.215 166.97 ;
        RECT 426.29 166.17 460.615 166.57 ;
        RECT 426.69 165.77 461.015 166.17 ;
        RECT 427.09 165.37 461.415 165.77 ;
        RECT 427.49 164.97 461.815 165.37 ;
        RECT 427.89 164.57 462.215 164.97 ;
        RECT 428.29 164.17 462.615 164.57 ;
        RECT 428.69 163.77 463.015 164.17 ;
        RECT 429.09 163.37 463.415 163.77 ;
        RECT 429.49 162.97 463.815 163.37 ;
        RECT 429.89 162.57 464.215 162.97 ;
        RECT 430.29 162.17 464.615 162.57 ;
        RECT 430.69 161.77 465.015 162.17 ;
        RECT 431.09 161.37 465.415 161.77 ;
        RECT 431.49 160.97 465.815 161.37 ;
        RECT 431.89 160.57 466.215 160.97 ;
        RECT 432.29 160.17 466.615 160.57 ;
        RECT 432.69 159.77 467.015 160.17 ;
        RECT 433.09 159.37 467.415 159.77 ;
        RECT 433.49 158.97 467.815 159.37 ;
        RECT 433.89 158.57 468.215 158.97 ;
        RECT 434.29 158.17 468.615 158.57 ;
        RECT 434.69 157.77 469.015 158.17 ;
        RECT 435.09 157.37 469.415 157.77 ;
        RECT 435.49 156.97 469.815 157.37 ;
        RECT 435.89 156.57 470.215 156.97 ;
        RECT 436.29 156.17 470.615 156.57 ;
        RECT 436.69 155.77 471.015 156.17 ;
        RECT 437.09 155.37 471.415 155.77 ;
        RECT 437.49 154.97 471.815 155.37 ;
        RECT 437.89 154.57 472.215 154.97 ;
        RECT 438.29 154.17 472.615 154.57 ;
        RECT 438.69 153.77 473.015 154.17 ;
        RECT 439.09 153.37 473.415 153.77 ;
        RECT 439.49 152.97 473.815 153.37 ;
        RECT 439.89 152.57 474.215 152.97 ;
        RECT 440.29 152.17 474.615 152.57 ;
        RECT 440.69 151.77 475.015 152.17 ;
        RECT 440.69 151.75 475.425 151.76 ;
        RECT 440.69 151.76 475.415 151.77 ;
        RECT 443.76 148.7 478.085 149.1 ;
        RECT 443.36 149.1 477.685 149.5 ;
        RECT 442.96 149.5 477.285 149.9 ;
        RECT 442.56 149.9 476.885 150.3 ;
        RECT 442.16 150.3 476.485 150.7 ;
        RECT 441.76 150.7 476.085 151.1 ;
        RECT 441.36 151.1 475.685 151.5 ;
        RECT 440.96 151.5 475.435 151.75 ;
        RECT 446.89 145.51 480 145.57 ;
        RECT 446.89 145.57 480 145.97 ;
        RECT 446.49 145.97 480 146.37 ;
        RECT 446.09 146.37 480 146.77 ;
        RECT 445.69 146.77 480 147.17 ;
        RECT 445.29 147.17 480 147.57 ;
        RECT 444.89 147.57 480 147.97 ;
        RECT 444.49 147.97 480 148.37 ;
        RECT 444.09 148.37 480 148.7 ;
        RECT 468.71 123.75 480 124.15 ;
        RECT 468.31 124.15 480 124.55 ;
        RECT 467.91 124.55 480 124.95 ;
        RECT 467.51 124.95 480 125.35 ;
        RECT 467.11 125.35 480 125.75 ;
        RECT 466.71 125.75 480 126.15 ;
        RECT 466.31 126.15 480 126.55 ;
        RECT 465.91 126.55 480 126.95 ;
        RECT 465.51 126.95 480 127.35 ;
        RECT 465.11 127.35 480 127.75 ;
        RECT 464.71 127.75 480 128.15 ;
        RECT 464.31 128.15 480 128.55 ;
        RECT 463.91 128.55 480 128.95 ;
        RECT 463.51 128.95 480 129.35 ;
        RECT 463.11 129.35 480 129.75 ;
        RECT 462.71 129.75 480 130.15 ;
        RECT 462.31 130.15 480 130.55 ;
        RECT 461.91 130.55 480 130.95 ;
        RECT 461.51 130.95 480 131.35 ;
        RECT 461.11 131.35 480 131.75 ;
        RECT 460.71 131.75 480 132.15 ;
        RECT 460.31 132.15 480 132.55 ;
        RECT 459.91 132.55 480 132.95 ;
        RECT 459.51 132.95 480 133.35 ;
        RECT 459.11 133.35 480 133.75 ;
        RECT 458.71 133.75 480 134.15 ;
        RECT 458.31 134.15 480 134.55 ;
        RECT 457.91 134.55 480 134.95 ;
        RECT 457.51 134.95 480 135.35 ;
        RECT 457.11 135.35 480 135.75 ;
        RECT 456.71 135.75 480 136.15 ;
        RECT 456.31 136.15 480 136.55 ;
        RECT 455.91 136.55 480 136.95 ;
        RECT 455.51 136.95 480 137.35 ;
        RECT 455.11 137.35 480 137.75 ;
        RECT 454.71 137.75 480 138.15 ;
        RECT 454.31 138.15 480 138.55 ;
        RECT 453.91 138.55 480 138.95 ;
        RECT 453.51 138.95 480 139.35 ;
        RECT 453.11 139.35 480 139.75 ;
        RECT 452.71 139.75 480 140.15 ;
        RECT 452.31 140.15 480 140.55 ;
        RECT 451.91 140.55 480 140.95 ;
        RECT 451.51 140.95 480 141.35 ;
        RECT 451.11 141.35 480 141.75 ;
        RECT 450.71 141.75 480 142.15 ;
        RECT 450.31 142.15 480 142.55 ;
        RECT 449.91 142.55 480 142.95 ;
        RECT 449.51 142.95 480 143.35 ;
        RECT 449.11 143.35 480 143.75 ;
        RECT 448.71 143.75 480 144.15 ;
        RECT 448.31 144.15 480 144.55 ;
        RECT 447.91 144.55 480 144.95 ;
        RECT 447.51 144.95 480 145.35 ;
        RECT 447.11 145.35 480 145.51 ;
        RECT 0 133.415 38.48 133.815 ;
        RECT 0 133.815 38.88 134.215 ;
        RECT 0 134.215 39.28 134.615 ;
        RECT 0 134.615 39.68 135.015 ;
        RECT 0 135.015 40.08 135.415 ;
        RECT 0 135.415 40.48 135.815 ;
        RECT 0 135.815 40.88 136.215 ;
        RECT 0 136.215 41.28 136.615 ;
        RECT 0 136.615 41.68 137.015 ;
        RECT 0 137.015 42.08 137.415 ;
        RECT 0 137.415 42.48 137.815 ;
        RECT 0 137.815 42.88 138.215 ;
        RECT 0 138.215 43.28 138.615 ;
        RECT 0 138.615 43.68 139.015 ;
        RECT 0 139.015 44.08 139.415 ;
        RECT 0 139.415 44.48 139.815 ;
        RECT 0 139.815 44.88 140.215 ;
        RECT 0 140.215 45.28 140.615 ;
        RECT 0 140.615 45.68 141.015 ;
        RECT 0 141.015 46.08 141.415 ;
        RECT 0 141.415 46.48 141.815 ;
        RECT 0 141.815 46.88 142.215 ;
        RECT 0 142.215 47.28 142.615 ;
        RECT 0 142.615 47.68 143.015 ;
        RECT 0 143.015 48.08 143.415 ;
        RECT 0 143.415 48.48 143.815 ;
        RECT 0 143.815 48.88 144.215 ;
        RECT 0 144.215 49.28 144.615 ;
        RECT 0 144.615 49.68 145.015 ;
        RECT 0 145.015 50.08 145.415 ;
        RECT 0 145.415 50.48 145.815 ;
        RECT 0 145.815 50.88 145.905 ;
        RECT 0 123.75 28.815 124.15 ;
        RECT 0 124.15 29.215 124.55 ;
        RECT 0 124.55 29.615 124.95 ;
        RECT 0 124.95 30.015 125.35 ;
        RECT 0 125.35 30.415 125.75 ;
        RECT 0 125.75 30.815 126.15 ;
        RECT 0 126.15 31.215 126.55 ;
        RECT 0 126.55 31.615 126.95 ;
        RECT 0 126.95 32.015 127.35 ;
        RECT 0 127.35 32.415 127.75 ;
        RECT 0 127.75 32.815 128.15 ;
        RECT 0 128.15 33.215 128.55 ;
        RECT 0 128.55 33.615 128.95 ;
        RECT 0 128.95 34.015 129.35 ;
        RECT 0 129.35 34.415 129.75 ;
        RECT 0 129.75 34.815 130.15 ;
        RECT 0 130.15 35.215 130.55 ;
        RECT 0 130.55 35.615 130.95 ;
        RECT 0 130.95 36.015 131.35 ;
        RECT 0 131.35 36.415 131.75 ;
        RECT 0 131.75 36.815 132.15 ;
        RECT 0 132.15 37.215 132.55 ;
        RECT 0 132.55 37.615 132.95 ;
        RECT 0 132.95 38.015 133.35 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 73.5 480 78.15 ;
        RECT 9.665 73.415 457.925 73.455 ;
        RECT 9.625 73.455 457.965 73.495 ;
        RECT 9.585 73.495 458.005 73.5 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.835 227.875 399.285 227.9 ;
        RECT 49.81 227.725 399.31 227.875 ;
        RECT 49.66 227.575 399.46 227.725 ;
        RECT 49.51 227.425 399.61 227.575 ;
        RECT 49.36 227.275 399.76 227.425 ;
        RECT 49.21 227.125 399.91 227.275 ;
        RECT 49.06 226.975 400.06 227.125 ;
        RECT 48.91 226.825 400.21 226.975 ;
        RECT 48.76 226.675 400.36 226.825 ;
        RECT 48.61 226.525 400.51 226.675 ;
        RECT 48.46 226.375 400.66 226.525 ;
        RECT 48.31 226.225 400.81 226.375 ;
        RECT 48.16 226.075 400.96 226.225 ;
        RECT 48.01 225.925 401.11 226.075 ;
        RECT 47.86 225.775 401.26 225.925 ;
        RECT 47.71 225.625 401.41 225.775 ;
        RECT 47.56 225.475 401.56 225.625 ;
        RECT 47.41 225.325 401.71 225.475 ;
        RECT 47.26 225.175 401.86 225.325 ;
        RECT 47.11 225.025 402.01 225.175 ;
        RECT 46.96 224.875 402.16 225.025 ;
        RECT 46.81 224.725 402.31 224.875 ;
        RECT 46.66 224.575 402.46 224.725 ;
        RECT 46.51 224.425 402.61 224.575 ;
        RECT 46.36 224.275 402.76 224.425 ;
        RECT 46.21 224.125 402.91 224.275 ;
        RECT 46.06 223.975 403.06 224.125 ;
        RECT 45.91 223.825 403.21 223.975 ;
        RECT 45.76 223.675 403.36 223.825 ;
        RECT 45.61 223.525 403.51 223.675 ;
        RECT 45.46 223.375 403.66 223.525 ;
        RECT 45.31 223.225 403.81 223.375 ;
        RECT 45.16 223.075 403.96 223.225 ;
        RECT 45.01 222.925 404.11 223.075 ;
        RECT 44.86 222.775 404.26 222.925 ;
        RECT 44.71 222.625 404.41 222.775 ;
        RECT 44.56 222.475 404.56 222.625 ;
        RECT 44.41 222.325 404.71 222.475 ;
        RECT 44.26 222.175 404.86 222.325 ;
        RECT 44.11 222.025 405.01 222.175 ;
        RECT 43.96 221.875 405.16 222.025 ;
        RECT 43.81 221.725 405.31 221.875 ;
        RECT 43.66 221.575 405.46 221.725 ;
        RECT 43.51 221.425 405.61 221.575 ;
        RECT 43.36 221.275 405.76 221.425 ;
        RECT 43.21 221.125 405.91 221.275 ;
        RECT 43.06 220.975 406.06 221.125 ;
        RECT 42.91 220.825 406.21 220.975 ;
        RECT 42.76 220.675 406.36 220.825 ;
        RECT 42.61 220.525 406.51 220.675 ;
        RECT 42.46 220.375 406.66 220.525 ;
        RECT 42.31 220.225 406.81 220.375 ;
        RECT 42.16 220.075 406.96 220.225 ;
        RECT 42.01 219.925 407.11 220.075 ;
        RECT 41.86 219.775 407.26 219.925 ;
        RECT 41.71 219.625 407.41 219.775 ;
        RECT 41.56 219.475 407.56 219.625 ;
        RECT 41.41 219.325 407.71 219.475 ;
        RECT 41.26 219.175 407.86 219.325 ;
        RECT 41.11 219.025 408.01 219.175 ;
        RECT 40.96 218.875 408.16 219.025 ;
        RECT 40.81 218.725 408.31 218.875 ;
        RECT 40.66 218.575 408.46 218.725 ;
        RECT 40.51 218.425 408.61 218.575 ;
        RECT 40.36 218.275 408.76 218.425 ;
        RECT 40.21 218.125 408.91 218.275 ;
        RECT 40.06 217.975 409.06 218.125 ;
        RECT 39.91 217.825 409.21 217.975 ;
        RECT 39.76 217.675 409.36 217.825 ;
        RECT 39.61 217.525 409.51 217.675 ;
        RECT 39.46 217.375 409.66 217.525 ;
        RECT 39.31 217.225 409.81 217.375 ;
        RECT 39.16 217.075 409.96 217.225 ;
        RECT 39.01 216.925 410.11 217.075 ;
        RECT 38.86 216.775 410.26 216.925 ;
        RECT 38.71 216.625 410.41 216.775 ;
        RECT 38.56 216.475 410.56 216.625 ;
        RECT 38.41 216.325 410.71 216.475 ;
        RECT 38.26 216.175 410.86 216.325 ;
        RECT 38.11 216.025 411.01 216.175 ;
        RECT 37.96 215.875 411.16 216.025 ;
        RECT 37.81 215.725 411.31 215.875 ;
        RECT 37.66 215.575 411.46 215.725 ;
        RECT 37.51 215.425 411.61 215.575 ;
        RECT 37.36 215.275 411.76 215.425 ;
        RECT 37.21 215.125 411.91 215.275 ;
        RECT 37.06 214.975 412.06 215.125 ;
        RECT 36.91 214.825 412.21 214.975 ;
        RECT 36.76 214.675 412.36 214.825 ;
        RECT 36.61 214.525 412.51 214.675 ;
        RECT 36.46 214.375 412.66 214.525 ;
        RECT 36.31 214.225 412.81 214.375 ;
        RECT 36.16 214.075 412.96 214.225 ;
        RECT 36.01 213.925 413.11 214.075 ;
        RECT 35.86 213.775 413.26 213.925 ;
        RECT 35.71 213.625 413.41 213.775 ;
        RECT 35.56 213.475 413.56 213.625 ;
        RECT 35.41 213.325 413.71 213.475 ;
        RECT 35.26 213.175 413.86 213.325 ;
        RECT 35.11 213.025 414.01 213.175 ;
        RECT 34.96 212.875 414.16 213.025 ;
        RECT 34.81 212.725 414.31 212.875 ;
        RECT 34.66 212.575 414.46 212.725 ;
        RECT 34.51 212.425 414.61 212.575 ;
        RECT 34.36 212.275 414.76 212.425 ;
        RECT 34.21 212.125 414.91 212.275 ;
        RECT 34.06 211.975 415.06 212.125 ;
        RECT 33.91 211.825 415.21 211.975 ;
        RECT 33.76 211.675 415.36 211.825 ;
        RECT 33.61 211.525 415.51 211.675 ;
        RECT 33.46 211.375 415.66 211.525 ;
        RECT 33.31 211.225 415.81 211.375 ;
        RECT 33.16 211.075 415.96 211.225 ;
        RECT 33.01 210.925 416.11 211.075 ;
        RECT 32.86 210.775 416.26 210.925 ;
        RECT 32.71 210.625 416.41 210.775 ;
        RECT 32.56 210.475 416.56 210.625 ;
        RECT 32.41 210.325 416.71 210.475 ;
        RECT 32.26 210.175 416.86 210.325 ;
        RECT 32.11 210.025 417.01 210.175 ;
        RECT 31.96 209.875 417.16 210.025 ;
        RECT 31.81 209.725 417.31 209.875 ;
        RECT 31.66 209.575 417.46 209.725 ;
        RECT 31.51 209.425 417.61 209.575 ;
        RECT 31.36 209.275 417.76 209.425 ;
        RECT 31.21 209.125 417.91 209.275 ;
        RECT 31.06 208.975 418.06 209.125 ;
        RECT 30.91 208.825 418.21 208.975 ;
        RECT 30.76 208.675 418.36 208.825 ;
        RECT 30.61 208.525 418.51 208.675 ;
        RECT 30.46 208.375 418.66 208.525 ;
        RECT 30.31 208.225 418.81 208.375 ;
        RECT 30.16 208.075 418.96 208.225 ;
        RECT 30.01 207.925 419.11 208.075 ;
        RECT 29.86 207.775 419.26 207.925 ;
        RECT 29.71 207.625 419.41 207.775 ;
        RECT 29.56 207.475 419.56 207.625 ;
        RECT 29.41 207.325 419.71 207.475 ;
        RECT 29.26 204.505 422.53 204.655 ;
        RECT 29.26 204.655 422.38 204.805 ;
        RECT 29.26 204.805 422.23 204.955 ;
        RECT 29.26 204.955 422.08 205.105 ;
        RECT 29.26 205.105 421.93 205.255 ;
        RECT 29.26 205.255 421.78 205.405 ;
        RECT 29.26 205.405 421.63 205.555 ;
        RECT 29.26 205.555 421.48 205.705 ;
        RECT 29.26 205.705 421.33 205.855 ;
        RECT 29.26 205.855 421.18 206.005 ;
        RECT 29.26 206.005 421.03 206.155 ;
        RECT 29.26 206.155 420.88 206.305 ;
        RECT 29.26 206.305 420.73 206.455 ;
        RECT 29.26 206.455 420.58 206.605 ;
        RECT 29.26 206.605 420.43 206.755 ;
        RECT 29.26 206.755 420.28 206.905 ;
        RECT 29.26 206.905 420.13 207.055 ;
        RECT 29.26 207.055 419.98 207.205 ;
        RECT 29.26 207.205 419.86 207.325 ;
        RECT 29.26 197.6 54.145 197.75 ;
        RECT 29.26 197.75 54.295 197.9 ;
        RECT 29.26 197.9 54.445 198.05 ;
        RECT 29.26 198.05 54.595 198.2 ;
        RECT 29.26 198.2 54.745 198.35 ;
        RECT 29.26 198.35 54.895 198.5 ;
        RECT 29.26 198.5 55.045 198.65 ;
        RECT 29.26 198.65 55.195 198.8 ;
        RECT 29.26 198.8 55.345 198.95 ;
        RECT 29.26 198.95 55.495 199.1 ;
        RECT 29.26 199.1 55.645 199.25 ;
        RECT 29.26 199.25 55.795 199.4 ;
        RECT 29.26 199.4 55.945 199.55 ;
        RECT 29.26 199.55 56.095 199.7 ;
        RECT 29.26 199.7 56.245 199.85 ;
        RECT 29.26 199.85 56.395 200 ;
        RECT 29.26 200 56.545 200.15 ;
        RECT 29.26 200.15 56.695 200.3 ;
        RECT 29.26 200.3 56.845 200.45 ;
        RECT 29.26 200.45 56.995 200.6 ;
        RECT 29.26 200.6 57.145 200.75 ;
        RECT 29.26 200.75 57.295 200.9 ;
        RECT 29.26 200.9 57.445 201.05 ;
        RECT 29.26 201.05 57.595 201.2 ;
        RECT 29.26 201.2 57.745 201.35 ;
        RECT 29.26 201.35 57.895 201.5 ;
        RECT 29.26 201.5 58.045 201.65 ;
        RECT 29.26 201.65 58.195 201.8 ;
        RECT 29.26 201.8 58.345 201.95 ;
        RECT 29.26 201.95 58.495 202.1 ;
        RECT 29.26 202.1 58.645 202.25 ;
        RECT 29.26 202.25 58.795 202.4 ;
        RECT 29.26 202.4 58.945 202.55 ;
        RECT 29.26 202.55 59.095 202.7 ;
        RECT 29.26 202.7 59.245 202.85 ;
        RECT 29.26 202.85 59.395 203 ;
        RECT 29.26 203 59.545 203.15 ;
        RECT 29.26 203.15 59.695 203.3 ;
        RECT 29.26 203.3 59.845 203.45 ;
        RECT 29.26 203.45 59.995 203.6 ;
        RECT 29.26 203.6 60.145 203.75 ;
        RECT 29.26 203.75 60.295 203.9 ;
        RECT 29.26 203.9 60.445 204.05 ;
        RECT 29.26 204.05 60.595 204.2 ;
        RECT 29.26 204.2 60.745 204.35 ;
        RECT 29.26 204.35 60.895 204.5 ;
        RECT 29.26 204.5 61.045 204.505 ;
        RECT 29.26 159.385 54.145 197.6 ;
        RECT 29.26 159.28 54.145 159.385 ;
        RECT 29.155 159.13 54.145 159.28 ;
        RECT 29.005 158.98 54.145 159.13 ;
        RECT 28.855 158.83 54.145 158.98 ;
        RECT 28.705 158.68 54.145 158.83 ;
        RECT 28.555 158.53 54.145 158.68 ;
        RECT 28.405 158.38 54.145 158.53 ;
        RECT 28.255 158.23 54.145 158.38 ;
        RECT 28.105 158.08 54.145 158.23 ;
        RECT 27.955 157.93 54.145 158.08 ;
        RECT 27.805 157.78 54.145 157.93 ;
        RECT 27.655 157.63 54.145 157.78 ;
        RECT 27.505 157.48 54.145 157.63 ;
        RECT 27.355 157.33 54.145 157.48 ;
        RECT 27.205 157.18 54.145 157.33 ;
        RECT 27.055 157.03 54.145 157.18 ;
        RECT 26.905 156.88 54.145 157.03 ;
        RECT 26.755 156.73 54.145 156.88 ;
        RECT 26.605 156.58 54.145 156.73 ;
        RECT 26.455 156.43 54.145 156.58 ;
        RECT 26.305 156.28 54.145 156.43 ;
        RECT 26.155 156.13 54.145 156.28 ;
        RECT 26.005 155.98 54.145 156.13 ;
        RECT 25.855 155.83 54.145 155.98 ;
        RECT 25.705 155.68 54.145 155.83 ;
        RECT 25.555 155.53 54.145 155.68 ;
        RECT 25.405 155.38 54.145 155.53 ;
        RECT 25.255 155.23 54.145 155.38 ;
        RECT 25.105 155.08 54.145 155.23 ;
        RECT 24.955 154.93 54.145 155.08 ;
        RECT 24.805 154.78 54.145 154.93 ;
        RECT 24.655 154.63 54.145 154.78 ;
        RECT 24.505 154.48 54.145 154.63 ;
        RECT 24.355 154.33 54.145 154.48 ;
        RECT 24.205 154.18 54.145 154.33 ;
        RECT 24.055 154.03 54.145 154.18 ;
        RECT 23.905 153.88 54.145 154.03 ;
        RECT 23.755 153.73 54.145 153.88 ;
        RECT 23.605 153.58 54.145 153.73 ;
        RECT 23.455 153.43 54.145 153.58 ;
        RECT 23.305 153.28 54.145 153.43 ;
        RECT 23.155 153.13 54.145 153.28 ;
        RECT 23.005 152.98 54.145 153.13 ;
        RECT 22.855 152.83 54.145 152.98 ;
        RECT 22.705 152.68 54.145 152.83 ;
        RECT 22.555 152.53 54.145 152.68 ;
        RECT 22.405 152.38 54.145 152.53 ;
        RECT 22.255 152.23 54.145 152.38 ;
        RECT 22.105 152.08 54.145 152.23 ;
        RECT 21.955 151.93 54.145 152.08 ;
        RECT 21.805 151.78 54.145 151.93 ;
        RECT 21.655 151.63 54.145 151.78 ;
        RECT 21.505 151.48 54.145 151.63 ;
        RECT 21.355 151.33 54.145 151.48 ;
        RECT 21.205 151.18 54.145 151.33 ;
        RECT 21.055 151.03 54.145 151.18 ;
        RECT 20.905 150.88 54.145 151.03 ;
        RECT 20.755 150.73 54.145 150.88 ;
        RECT 20.605 150.58 54.145 150.73 ;
        RECT 20.455 150.43 54.145 150.58 ;
        RECT 20.305 150.28 54.145 150.43 ;
        RECT 20.155 150.13 54.145 150.28 ;
        RECT 20.005 149.98 54.145 150.13 ;
        RECT 19.855 149.83 54.145 149.98 ;
        RECT 19.705 149.68 54.145 149.83 ;
        RECT 19.555 149.53 54.145 149.68 ;
        RECT 19.405 149.38 54.145 149.53 ;
        RECT 19.255 149.23 54.145 149.38 ;
        RECT 19.105 149.08 54.145 149.23 ;
        RECT 388.11 204.365 422.68 204.505 ;
        RECT 388.26 204.215 422.82 204.365 ;
        RECT 388.41 204.065 422.97 204.215 ;
        RECT 388.56 203.915 423.12 204.065 ;
        RECT 388.71 203.765 423.27 203.915 ;
        RECT 388.86 203.615 423.42 203.765 ;
        RECT 389.01 203.465 423.57 203.615 ;
        RECT 389.16 203.315 423.72 203.465 ;
        RECT 389.31 203.165 423.87 203.315 ;
        RECT 389.46 203.015 424.02 203.165 ;
        RECT 389.61 202.865 424.17 203.015 ;
        RECT 389.76 202.715 424.32 202.865 ;
        RECT 389.91 202.565 424.47 202.715 ;
        RECT 390.06 202.415 424.62 202.565 ;
        RECT 390.21 202.265 424.77 202.415 ;
        RECT 390.36 202.115 424.92 202.265 ;
        RECT 390.51 201.965 425.07 202.115 ;
        RECT 390.66 201.815 425.22 201.965 ;
        RECT 390.81 201.665 425.37 201.815 ;
        RECT 390.96 201.515 425.52 201.665 ;
        RECT 391.11 201.365 425.67 201.515 ;
        RECT 391.26 201.215 425.82 201.365 ;
        RECT 391.41 201.065 425.97 201.215 ;
        RECT 391.56 200.915 426.12 201.065 ;
        RECT 391.71 200.765 426.27 200.915 ;
        RECT 391.86 200.615 426.42 200.765 ;
        RECT 392.01 200.465 426.57 200.615 ;
        RECT 392.16 200.315 426.72 200.465 ;
        RECT 392.31 200.165 426.87 200.315 ;
        RECT 392.46 200.015 427.02 200.165 ;
        RECT 392.61 199.865 427.17 200.015 ;
        RECT 392.76 199.715 427.32 199.865 ;
        RECT 392.91 199.565 427.47 199.715 ;
        RECT 393.06 199.415 427.62 199.565 ;
        RECT 393.21 199.265 427.77 199.415 ;
        RECT 393.36 199.115 427.92 199.265 ;
        RECT 393.51 198.965 428.07 199.115 ;
        RECT 393.66 198.815 428.22 198.965 ;
        RECT 393.81 198.665 428.37 198.815 ;
        RECT 393.96 198.515 428.52 198.665 ;
        RECT 394.11 198.365 428.67 198.515 ;
        RECT 394.26 198.215 428.82 198.365 ;
        RECT 394.41 198.065 428.97 198.215 ;
        RECT 394.56 197.915 429.12 198.065 ;
        RECT 394.71 197.765 429.27 197.915 ;
        RECT 394.86 197.615 429.42 197.765 ;
        RECT 395.01 197.465 429.57 197.615 ;
        RECT 395.16 197.315 429.72 197.465 ;
        RECT 395.31 197.165 429.87 197.315 ;
        RECT 395.46 197.015 430.02 197.165 ;
        RECT 395.61 196.865 430.17 197.015 ;
        RECT 395.76 196.715 430.32 196.865 ;
        RECT 395.91 196.565 430.47 196.715 ;
        RECT 396.06 196.415 430.62 196.565 ;
        RECT 396.21 196.265 430.77 196.415 ;
        RECT 396.36 196.115 430.92 196.265 ;
        RECT 396.51 195.965 431.07 196.115 ;
        RECT 396.66 195.815 431.22 195.965 ;
        RECT 396.81 195.665 431.37 195.815 ;
        RECT 396.96 195.515 431.52 195.665 ;
        RECT 397.11 195.365 431.67 195.515 ;
        RECT 397.26 195.215 431.82 195.365 ;
        RECT 397.41 195.065 431.97 195.215 ;
        RECT 397.56 194.915 432.12 195.065 ;
        RECT 397.71 194.765 432.27 194.915 ;
        RECT 397.86 194.615 432.42 194.765 ;
        RECT 398.01 194.465 432.57 194.615 ;
        RECT 398.16 194.315 432.72 194.465 ;
        RECT 398.31 194.165 432.87 194.315 ;
        RECT 398.46 194.015 433.02 194.165 ;
        RECT 398.61 193.865 433.17 194.015 ;
        RECT 398.76 193.715 433.32 193.865 ;
        RECT 398.91 193.565 433.47 193.715 ;
        RECT 399.06 193.415 433.62 193.565 ;
        RECT 399.21 193.265 433.77 193.415 ;
        RECT 399.36 193.115 433.92 193.265 ;
        RECT 399.51 192.965 434.07 193.115 ;
        RECT 399.66 192.815 434.22 192.965 ;
        RECT 399.81 192.665 434.37 192.815 ;
        RECT 399.96 192.515 434.52 192.665 ;
        RECT 400.11 192.365 434.67 192.515 ;
        RECT 400.26 192.215 434.82 192.365 ;
        RECT 400.41 192.065 434.97 192.215 ;
        RECT 400.56 191.915 435.12 192.065 ;
        RECT 400.71 191.765 435.27 191.915 ;
        RECT 400.86 191.615 435.42 191.765 ;
        RECT 401.01 191.465 435.57 191.615 ;
        RECT 401.16 191.315 435.72 191.465 ;
        RECT 401.31 191.165 435.87 191.315 ;
        RECT 401.46 191.015 436.02 191.165 ;
        RECT 401.61 190.865 436.17 191.015 ;
        RECT 401.76 190.715 436.32 190.865 ;
        RECT 401.91 190.565 436.47 190.715 ;
        RECT 402.06 190.415 436.62 190.565 ;
        RECT 402.21 190.265 436.77 190.415 ;
        RECT 402.36 190.115 436.92 190.265 ;
        RECT 402.51 189.965 437.07 190.115 ;
        RECT 402.66 189.815 437.22 189.965 ;
        RECT 402.81 189.665 437.37 189.815 ;
        RECT 402.96 189.515 437.52 189.665 ;
        RECT 403.11 189.365 437.67 189.515 ;
        RECT 403.26 189.215 437.82 189.365 ;
        RECT 403.41 189.065 437.97 189.215 ;
        RECT 403.56 188.915 438.12 189.065 ;
        RECT 403.71 188.765 438.27 188.915 ;
        RECT 403.86 188.615 438.42 188.765 ;
        RECT 404.01 188.465 438.57 188.615 ;
        RECT 404.16 188.315 438.72 188.465 ;
        RECT 404.31 188.165 438.87 188.315 ;
        RECT 404.46 188.015 439.02 188.165 ;
        RECT 404.61 187.865 439.17 188.015 ;
        RECT 404.76 187.715 439.32 187.865 ;
        RECT 404.91 187.565 439.47 187.715 ;
        RECT 405.06 187.415 439.62 187.565 ;
        RECT 405.21 187.265 439.77 187.415 ;
        RECT 405.36 187.115 439.92 187.265 ;
        RECT 405.51 186.965 440.07 187.115 ;
        RECT 405.66 186.815 440.22 186.965 ;
        RECT 405.81 186.665 440.37 186.815 ;
        RECT 405.96 186.515 440.52 186.665 ;
        RECT 406.11 186.365 440.67 186.515 ;
        RECT 406.26 186.215 440.82 186.365 ;
        RECT 406.41 186.065 440.97 186.215 ;
        RECT 406.56 185.915 441.12 186.065 ;
        RECT 406.71 185.765 441.27 185.915 ;
        RECT 406.86 185.615 441.42 185.765 ;
        RECT 407.01 185.465 441.57 185.615 ;
        RECT 407.16 185.315 441.72 185.465 ;
        RECT 407.31 185.165 441.87 185.315 ;
        RECT 407.46 185.015 442.02 185.165 ;
        RECT 407.61 184.865 442.17 185.015 ;
        RECT 407.76 184.715 442.32 184.865 ;
        RECT 407.91 184.565 442.47 184.715 ;
        RECT 408.06 184.415 442.62 184.565 ;
        RECT 408.21 184.265 442.77 184.415 ;
        RECT 408.36 184.115 442.92 184.265 ;
        RECT 408.51 183.965 443.07 184.115 ;
        RECT 408.66 183.815 443.22 183.965 ;
        RECT 408.81 183.665 443.37 183.815 ;
        RECT 408.96 183.515 443.52 183.665 ;
        RECT 409.11 183.365 443.67 183.515 ;
        RECT 409.26 183.215 443.82 183.365 ;
        RECT 409.41 183.065 443.97 183.215 ;
        RECT 409.56 182.915 444.12 183.065 ;
        RECT 409.71 182.765 444.27 182.915 ;
        RECT 409.86 182.615 444.42 182.765 ;
        RECT 410.01 182.465 444.57 182.615 ;
        RECT 410.16 182.315 444.72 182.465 ;
        RECT 410.31 182.165 444.87 182.315 ;
        RECT 410.46 182.015 445.02 182.165 ;
        RECT 410.61 181.865 445.17 182.015 ;
        RECT 410.76 181.715 445.32 181.865 ;
        RECT 410.91 181.565 445.47 181.715 ;
        RECT 411.06 181.415 445.62 181.565 ;
        RECT 411.21 181.265 445.77 181.415 ;
        RECT 411.36 181.115 445.92 181.265 ;
        RECT 411.51 180.965 446.07 181.115 ;
        RECT 411.66 180.815 446.22 180.965 ;
        RECT 411.81 180.665 446.37 180.815 ;
        RECT 411.96 180.515 446.52 180.665 ;
        RECT 412.11 180.365 446.67 180.515 ;
        RECT 412.26 180.215 446.82 180.365 ;
        RECT 412.41 180.065 446.97 180.215 ;
        RECT 412.56 179.915 447.12 180.065 ;
        RECT 412.71 179.765 447.27 179.915 ;
        RECT 412.86 179.615 447.42 179.765 ;
        RECT 413.01 179.465 447.57 179.615 ;
        RECT 413.16 179.315 447.72 179.465 ;
        RECT 413.31 179.165 447.87 179.315 ;
        RECT 413.46 179.015 448.02 179.165 ;
        RECT 413.61 178.865 448.17 179.015 ;
        RECT 413.76 178.715 448.32 178.865 ;
        RECT 413.91 178.565 448.47 178.715 ;
        RECT 414.06 178.415 448.62 178.565 ;
        RECT 414.21 178.265 448.77 178.415 ;
        RECT 414.36 178.115 448.92 178.265 ;
        RECT 414.51 177.965 449.07 178.115 ;
        RECT 414.66 177.815 449.22 177.965 ;
        RECT 414.81 177.665 449.37 177.815 ;
        RECT 414.96 177.515 449.52 177.665 ;
        RECT 415.11 177.365 449.67 177.515 ;
        RECT 415.26 177.215 449.82 177.365 ;
        RECT 415.41 177.065 449.97 177.215 ;
        RECT 415.56 176.915 450.12 177.065 ;
        RECT 415.71 176.765 450.27 176.915 ;
        RECT 415.86 176.615 450.42 176.765 ;
        RECT 416.01 176.465 450.57 176.615 ;
        RECT 416.16 176.315 450.72 176.465 ;
        RECT 416.31 176.165 450.87 176.315 ;
        RECT 416.46 176.015 451.02 176.165 ;
        RECT 416.61 175.865 451.17 176.015 ;
        RECT 416.76 175.715 451.32 175.865 ;
        RECT 416.91 175.565 451.47 175.715 ;
        RECT 417.06 175.415 451.62 175.565 ;
        RECT 417.21 175.265 451.77 175.415 ;
        RECT 417.36 175.115 451.92 175.265 ;
        RECT 417.51 174.965 452.07 175.115 ;
        RECT 417.66 174.815 452.22 174.965 ;
        RECT 417.81 174.665 452.37 174.815 ;
        RECT 417.96 174.515 452.52 174.665 ;
        RECT 418.11 174.365 452.67 174.515 ;
        RECT 418.26 174.215 452.82 174.365 ;
        RECT 418.41 174.065 452.97 174.215 ;
        RECT 418.56 173.915 453.12 174.065 ;
        RECT 418.71 173.765 453.27 173.915 ;
        RECT 418.86 173.615 453.42 173.765 ;
        RECT 419.01 173.465 453.57 173.615 ;
        RECT 419.16 173.315 453.72 173.465 ;
        RECT 419.31 173.165 453.87 173.315 ;
        RECT 419.46 173.015 454.02 173.165 ;
        RECT 419.61 172.865 454.17 173.015 ;
        RECT 419.76 172.715 454.32 172.865 ;
        RECT 419.91 172.565 454.47 172.715 ;
        RECT 420.06 172.415 454.62 172.565 ;
        RECT 420.21 172.265 454.77 172.415 ;
        RECT 420.36 172.115 454.92 172.265 ;
        RECT 420.51 171.965 455.07 172.115 ;
        RECT 420.66 171.815 455.22 171.965 ;
        RECT 420.81 171.665 455.37 171.815 ;
        RECT 420.96 171.515 455.52 171.665 ;
        RECT 421.11 171.365 455.67 171.515 ;
        RECT 421.26 171.215 455.82 171.365 ;
        RECT 421.41 171.065 455.97 171.215 ;
        RECT 421.56 170.915 456.12 171.065 ;
        RECT 421.71 170.765 456.27 170.915 ;
        RECT 421.86 170.615 456.42 170.765 ;
        RECT 422.01 170.465 456.57 170.615 ;
        RECT 422.16 170.315 456.72 170.465 ;
        RECT 422.31 170.165 456.87 170.315 ;
        RECT 422.46 170.015 457.02 170.165 ;
        RECT 422.61 169.865 457.17 170.015 ;
        RECT 422.76 169.715 457.32 169.865 ;
        RECT 422.91 169.565 457.47 169.715 ;
        RECT 423.06 169.415 457.62 169.565 ;
        RECT 423.21 169.265 457.77 169.415 ;
        RECT 423.36 169.115 457.92 169.265 ;
        RECT 423.51 168.965 458.07 169.115 ;
        RECT 423.66 168.815 458.22 168.965 ;
        RECT 423.81 168.665 458.37 168.815 ;
        RECT 423.96 168.515 458.52 168.665 ;
        RECT 424.11 168.365 458.67 168.515 ;
        RECT 424.26 168.215 458.82 168.365 ;
        RECT 424.41 168.065 458.97 168.215 ;
        RECT 424.56 167.915 459.12 168.065 ;
        RECT 424.71 167.765 459.27 167.915 ;
        RECT 424.86 167.615 459.42 167.765 ;
        RECT 425.01 167.465 459.57 167.615 ;
        RECT 425.16 167.315 459.72 167.465 ;
        RECT 425.31 167.165 459.87 167.315 ;
        RECT 425.46 167.015 460.02 167.165 ;
        RECT 425.61 166.865 460.17 167.015 ;
        RECT 425.76 166.715 460.32 166.865 ;
        RECT 425.91 166.565 460.47 166.715 ;
        RECT 426.06 166.415 460.62 166.565 ;
        RECT 426.21 166.265 460.77 166.415 ;
        RECT 426.36 166.115 460.92 166.265 ;
        RECT 426.51 165.965 461.07 166.115 ;
        RECT 426.66 165.815 461.22 165.965 ;
        RECT 426.81 165.665 461.37 165.815 ;
        RECT 426.96 165.515 461.52 165.665 ;
        RECT 427.11 165.365 461.67 165.515 ;
        RECT 427.26 165.215 461.82 165.365 ;
        RECT 427.41 165.065 461.97 165.215 ;
        RECT 427.56 164.915 462.12 165.065 ;
        RECT 427.71 164.765 462.27 164.915 ;
        RECT 427.86 164.615 462.42 164.765 ;
        RECT 428.01 164.465 462.57 164.615 ;
        RECT 428.16 164.315 462.72 164.465 ;
        RECT 428.31 164.165 462.87 164.315 ;
        RECT 428.46 164.015 463.02 164.165 ;
        RECT 428.61 163.865 463.17 164.015 ;
        RECT 428.76 163.715 463.32 163.865 ;
        RECT 428.91 163.565 463.47 163.715 ;
        RECT 429.06 163.415 463.62 163.565 ;
        RECT 429.21 163.265 463.77 163.415 ;
        RECT 429.36 163.115 463.92 163.265 ;
        RECT 429.51 162.965 464.07 163.115 ;
        RECT 429.66 162.815 464.22 162.965 ;
        RECT 429.81 162.665 464.37 162.815 ;
        RECT 429.96 162.515 464.52 162.665 ;
        RECT 430.11 162.365 464.67 162.515 ;
        RECT 430.26 162.215 464.82 162.365 ;
        RECT 430.41 162.065 464.97 162.215 ;
        RECT 430.56 161.915 465.12 162.065 ;
        RECT 430.71 161.765 465.27 161.915 ;
        RECT 430.86 161.615 465.42 161.765 ;
        RECT 431.01 161.465 465.57 161.615 ;
        RECT 431.16 161.315 465.72 161.465 ;
        RECT 431.31 161.165 465.87 161.315 ;
        RECT 431.46 161.015 466.02 161.165 ;
        RECT 431.61 160.865 466.17 161.015 ;
        RECT 431.76 160.715 466.32 160.865 ;
        RECT 431.91 160.565 466.47 160.715 ;
        RECT 432.06 160.415 466.62 160.565 ;
        RECT 432.21 160.265 466.77 160.415 ;
        RECT 432.36 160.115 466.92 160.265 ;
        RECT 432.51 159.965 467.07 160.115 ;
        RECT 432.66 159.815 467.22 159.965 ;
        RECT 432.81 159.665 467.37 159.815 ;
        RECT 432.96 159.515 467.52 159.665 ;
        RECT 433.11 159.365 467.67 159.515 ;
        RECT 433.26 159.215 467.82 159.365 ;
        RECT 433.41 159.065 467.97 159.215 ;
        RECT 433.56 158.915 468.12 159.065 ;
        RECT 433.71 158.765 468.27 158.915 ;
        RECT 433.86 158.615 468.42 158.765 ;
        RECT 434.01 158.465 468.57 158.615 ;
        RECT 434.16 158.315 468.72 158.465 ;
        RECT 434.31 158.165 468.87 158.315 ;
        RECT 434.46 158.015 469.02 158.165 ;
        RECT 434.61 157.865 469.17 158.015 ;
        RECT 434.76 157.715 469.32 157.865 ;
        RECT 434.91 157.565 469.47 157.715 ;
        RECT 435.06 157.415 469.62 157.565 ;
        RECT 435.21 157.265 469.77 157.415 ;
        RECT 435.36 157.115 469.92 157.265 ;
        RECT 435.51 156.965 470.07 157.115 ;
        RECT 435.66 156.815 470.22 156.965 ;
        RECT 435.81 156.665 470.37 156.815 ;
        RECT 435.96 156.515 470.52 156.665 ;
        RECT 436.11 156.365 470.67 156.515 ;
        RECT 436.26 156.215 470.82 156.365 ;
        RECT 436.41 156.065 470.97 156.215 ;
        RECT 436.56 155.915 471.12 156.065 ;
        RECT 436.71 155.765 471.27 155.915 ;
        RECT 436.86 155.615 471.42 155.765 ;
        RECT 437.01 155.465 471.57 155.615 ;
        RECT 437.16 155.315 471.72 155.465 ;
        RECT 437.31 155.165 471.87 155.315 ;
        RECT 437.46 155.015 472.02 155.165 ;
        RECT 437.61 154.865 472.17 155.015 ;
        RECT 437.76 154.715 472.32 154.865 ;
        RECT 437.91 154.565 472.47 154.715 ;
        RECT 438.06 154.415 472.62 154.565 ;
        RECT 438.21 154.265 472.77 154.415 ;
        RECT 438.36 154.115 472.92 154.265 ;
        RECT 438.51 153.965 473.07 154.115 ;
        RECT 438.66 153.815 473.22 153.965 ;
        RECT 438.81 153.665 473.37 153.815 ;
        RECT 438.96 153.515 473.52 153.665 ;
        RECT 439.11 153.365 473.67 153.515 ;
        RECT 439.26 153.215 473.82 153.365 ;
        RECT 439.41 153.065 473.97 153.215 ;
        RECT 439.56 152.915 474.12 153.065 ;
        RECT 439.71 152.765 474.27 152.915 ;
        RECT 439.86 152.615 474.42 152.765 ;
        RECT 440.01 152.465 474.57 152.615 ;
        RECT 440.16 152.315 474.72 152.465 ;
        RECT 440.31 152.165 474.87 152.315 ;
        RECT 440.46 152.015 475.02 152.165 ;
        RECT 440.61 151.865 475.17 152.015 ;
        RECT 440.76 151.715 475.32 151.865 ;
        RECT 440.91 151.565 475.47 151.715 ;
        RECT 441.06 151.415 475.62 151.565 ;
        RECT 441.21 151.265 475.77 151.415 ;
        RECT 441.36 151.115 475.92 151.265 ;
        RECT 441.51 150.965 476.07 151.115 ;
        RECT 441.66 150.815 476.22 150.965 ;
        RECT 441.81 150.665 476.37 150.815 ;
        RECT 441.96 150.515 476.52 150.665 ;
        RECT 442.11 150.365 476.67 150.515 ;
        RECT 442.26 150.215 476.82 150.365 ;
        RECT 442.41 150.065 476.97 150.215 ;
        RECT 442.56 149.915 477.12 150.065 ;
        RECT 442.71 149.765 477.27 149.915 ;
        RECT 442.86 149.615 477.42 149.765 ;
        RECT 443.01 149.465 477.57 149.615 ;
        RECT 443.16 149.315 477.72 149.465 ;
        RECT 443.31 149.165 477.87 149.315 ;
        RECT 443.46 149.015 478.02 149.165 ;
        RECT 443.61 148.865 478.17 149.015 ;
        RECT 443.76 148.715 478.32 148.865 ;
        RECT 18.74 148.715 53.78 148.865 ;
        RECT 18.89 148.865 53.93 149.015 ;
        RECT 18.955 149.015 54.08 149.08 ;
        RECT 0 148.615 53.68 148.715 ;
        RECT 0 148.465 53.53 148.615 ;
        RECT 0 148.315 53.38 148.465 ;
        RECT 0 148.165 53.23 148.315 ;
        RECT 0 148.015 53.08 148.165 ;
        RECT 0 147.865 52.93 148.015 ;
        RECT 0 147.715 52.78 147.865 ;
        RECT 0 147.565 52.63 147.715 ;
        RECT 0 147.415 52.48 147.565 ;
        RECT 0 147.265 52.33 147.415 ;
        RECT 0 147.115 52.18 147.265 ;
        RECT 0 146.965 52.03 147.115 ;
        RECT 0 146.815 51.88 146.965 ;
        RECT 0 146.665 51.73 146.815 ;
        RECT 0 146.515 51.58 146.665 ;
        RECT 0 146.365 51.43 146.515 ;
        RECT 0 146.215 51.28 146.365 ;
        RECT 0 146.065 51.13 146.215 ;
        RECT 0 145.915 50.98 146.065 ;
        RECT 0 145.765 50.83 145.915 ;
        RECT 0 145.615 50.68 145.765 ;
        RECT 0 145.465 50.53 145.615 ;
        RECT 0 145.315 50.38 145.465 ;
        RECT 0 145.165 50.23 145.315 ;
        RECT 0 145.015 50.08 145.165 ;
        RECT 0 144.865 49.93 145.015 ;
        RECT 0 144.715 49.78 144.865 ;
        RECT 0 144.565 49.63 144.715 ;
        RECT 0 144.415 49.48 144.565 ;
        RECT 0 144.265 49.33 144.415 ;
        RECT 0 144.115 49.18 144.265 ;
        RECT 0 143.965 49.03 144.115 ;
        RECT 0 143.815 48.88 143.965 ;
        RECT 0 143.665 48.73 143.815 ;
        RECT 0 143.515 48.58 143.665 ;
        RECT 0 143.365 48.43 143.515 ;
        RECT 0 143.215 48.28 143.365 ;
        RECT 0 143.065 48.13 143.215 ;
        RECT 0 142.915 47.98 143.065 ;
        RECT 0 142.765 47.83 142.915 ;
        RECT 0 142.615 47.68 142.765 ;
        RECT 0 142.465 47.53 142.615 ;
        RECT 0 142.315 47.38 142.465 ;
        RECT 0 142.165 47.23 142.315 ;
        RECT 0 142.015 47.08 142.165 ;
        RECT 0 141.865 46.93 142.015 ;
        RECT 0 141.715 46.78 141.865 ;
        RECT 0 141.565 46.63 141.715 ;
        RECT 0 141.415 46.48 141.565 ;
        RECT 0 141.265 46.33 141.415 ;
        RECT 0 141.115 46.18 141.265 ;
        RECT 0 140.965 46.03 141.115 ;
        RECT 0 140.815 45.88 140.965 ;
        RECT 0 140.665 45.73 140.815 ;
        RECT 0 140.515 45.58 140.665 ;
        RECT 0 140.365 45.43 140.515 ;
        RECT 0 140.215 45.28 140.365 ;
        RECT 0 140.065 45.13 140.215 ;
        RECT 0 139.915 44.98 140.065 ;
        RECT 0 139.765 44.83 139.915 ;
        RECT 0 139.615 44.68 139.765 ;
        RECT 0 139.465 44.53 139.615 ;
        RECT 0 139.315 44.38 139.465 ;
        RECT 0 139.165 44.23 139.315 ;
        RECT 0 139.015 44.08 139.165 ;
        RECT 0 138.865 43.93 139.015 ;
        RECT 0 138.715 43.78 138.865 ;
        RECT 0 138.565 43.63 138.715 ;
        RECT 0 138.415 43.48 138.565 ;
        RECT 0 138.265 43.33 138.415 ;
        RECT 0 138.115 43.18 138.265 ;
        RECT 0 137.965 43.03 138.115 ;
        RECT 0 137.815 42.88 137.965 ;
        RECT 0 137.665 42.73 137.815 ;
        RECT 0 137.515 42.58 137.665 ;
        RECT 0 137.365 42.43 137.515 ;
        RECT 0 137.215 42.28 137.365 ;
        RECT 0 137.065 42.13 137.215 ;
        RECT 0 136.915 41.98 137.065 ;
        RECT 0 136.765 41.83 136.915 ;
        RECT 0 136.615 41.68 136.765 ;
        RECT 0 136.465 41.53 136.615 ;
        RECT 0 136.315 41.38 136.465 ;
        RECT 0 136.165 41.23 136.315 ;
        RECT 0 136.015 41.08 136.165 ;
        RECT 0 135.865 40.93 136.015 ;
        RECT 0 135.715 40.78 135.865 ;
        RECT 0 135.565 40.63 135.715 ;
        RECT 0 135.415 40.48 135.565 ;
        RECT 0 135.265 40.33 135.415 ;
        RECT 0 135.115 40.18 135.265 ;
        RECT 0 134.965 40.03 135.115 ;
        RECT 0 134.815 39.88 134.965 ;
        RECT 0 134.665 39.73 134.815 ;
        RECT 0 134.515 39.58 134.665 ;
        RECT 0 134.365 39.43 134.515 ;
        RECT 0 134.215 39.28 134.365 ;
        RECT 0 134.065 39.13 134.215 ;
        RECT 0 133.915 38.98 134.065 ;
        RECT 0 133.765 38.83 133.915 ;
        RECT 0 133.615 38.68 133.765 ;
        RECT 0 133.465 38.53 133.615 ;
        RECT 0 133.315 38.38 133.465 ;
        RECT 0 133.165 38.23 133.315 ;
        RECT 0 133.015 38.08 133.165 ;
        RECT 0 132.865 37.93 133.015 ;
        RECT 0 132.715 37.78 132.865 ;
        RECT 0 132.565 37.63 132.715 ;
        RECT 0 132.415 37.48 132.565 ;
        RECT 0 132.265 37.33 132.415 ;
        RECT 0 132.115 37.18 132.265 ;
        RECT 0 131.965 37.03 132.115 ;
        RECT 0 131.815 36.88 131.965 ;
        RECT 0 131.665 36.73 131.815 ;
        RECT 0 131.515 36.58 131.665 ;
        RECT 0 131.365 36.43 131.515 ;
        RECT 0 131.215 36.28 131.365 ;
        RECT 0 131.065 36.13 131.215 ;
        RECT 0 130.915 35.98 131.065 ;
        RECT 0 130.765 35.83 130.915 ;
        RECT 0 130.615 35.68 130.765 ;
        RECT 0 130.465 35.53 130.615 ;
        RECT 0 130.315 35.38 130.465 ;
        RECT 0 130.165 35.23 130.315 ;
        RECT 0 130.015 35.08 130.165 ;
        RECT 0 129.865 34.93 130.015 ;
        RECT 0 129.715 34.78 129.865 ;
        RECT 0 129.565 34.63 129.715 ;
        RECT 0 129.415 34.48 129.565 ;
        RECT 0 129.265 34.33 129.415 ;
        RECT 0 129.115 34.18 129.265 ;
        RECT 0 128.965 34.03 129.115 ;
        RECT 0 128.815 33.88 128.965 ;
        RECT 0 128.665 33.73 128.815 ;
        RECT 0 128.515 33.58 128.665 ;
        RECT 0 128.365 33.43 128.515 ;
        RECT 0 128.215 33.28 128.365 ;
        RECT 0 128.065 33.13 128.215 ;
        RECT 0 127.915 32.98 128.065 ;
        RECT 0 127.765 32.83 127.915 ;
        RECT 0 127.615 32.68 127.765 ;
        RECT 0 127.465 32.53 127.615 ;
        RECT 0 127.315 32.38 127.465 ;
        RECT 0 127.165 32.23 127.315 ;
        RECT 0 127.015 32.08 127.165 ;
        RECT 0 126.865 31.93 127.015 ;
        RECT 0 126.715 31.78 126.865 ;
        RECT 0 126.565 31.63 126.715 ;
        RECT 0 126.415 31.48 126.565 ;
        RECT 0 126.265 31.33 126.415 ;
        RECT 0 126.115 31.18 126.265 ;
        RECT 0 125.965 31.03 126.115 ;
        RECT 0 125.815 30.88 125.965 ;
        RECT 0 125.665 30.73 125.815 ;
        RECT 0 125.515 30.58 125.665 ;
        RECT 0 125.365 30.43 125.515 ;
        RECT 0 125.215 30.28 125.365 ;
        RECT 0 125.065 30.13 125.215 ;
        RECT 0 124.915 29.98 125.065 ;
        RECT 0 124.765 29.83 124.915 ;
        RECT 0 124.615 29.68 124.765 ;
        RECT 0 124.465 29.53 124.615 ;
        RECT 0 124.315 29.38 124.465 ;
        RECT 0 124.165 29.23 124.315 ;
        RECT 0 124.015 29.08 124.165 ;
        RECT 0 123.865 28.93 124.015 ;
        RECT 443.825 148.65 480 148.715 ;
        RECT 443.975 148.5 480 148.65 ;
        RECT 444.125 148.35 480 148.5 ;
        RECT 444.275 148.2 480 148.35 ;
        RECT 444.425 148.05 480 148.2 ;
        RECT 444.575 147.9 480 148.05 ;
        RECT 444.725 147.75 480 147.9 ;
        RECT 444.875 147.6 480 147.75 ;
        RECT 445.025 147.45 480 147.6 ;
        RECT 445.175 147.3 480 147.45 ;
        RECT 445.325 147.15 480 147.3 ;
        RECT 445.475 147 480 147.15 ;
        RECT 445.625 146.85 480 147 ;
        RECT 445.775 146.7 480 146.85 ;
        RECT 445.925 146.55 480 146.7 ;
        RECT 446.075 146.4 480 146.55 ;
        RECT 446.225 146.25 480 146.4 ;
        RECT 446.375 146.1 480 146.25 ;
        RECT 446.525 145.95 480 146.1 ;
        RECT 446.675 145.8 480 145.95 ;
        RECT 446.825 145.65 480 145.8 ;
        RECT 446.975 145.5 480 145.65 ;
        RECT 447.125 145.35 480 145.5 ;
        RECT 447.275 145.2 480 145.35 ;
        RECT 447.425 145.05 480 145.2 ;
        RECT 447.575 144.9 480 145.05 ;
        RECT 447.725 144.75 480 144.9 ;
        RECT 447.875 144.6 480 144.75 ;
        RECT 448.025 144.45 480 144.6 ;
        RECT 448.175 144.3 480 144.45 ;
        RECT 448.325 144.15 480 144.3 ;
        RECT 448.475 144 480 144.15 ;
        RECT 448.625 143.85 480 144 ;
        RECT 448.775 143.7 480 143.85 ;
        RECT 448.925 143.55 480 143.7 ;
        RECT 449.075 143.4 480 143.55 ;
        RECT 449.225 143.25 480 143.4 ;
        RECT 449.375 143.1 480 143.25 ;
        RECT 449.525 142.95 480 143.1 ;
        RECT 449.675 142.8 480 142.95 ;
        RECT 449.825 142.65 480 142.8 ;
        RECT 449.975 142.5 480 142.65 ;
        RECT 450.125 142.35 480 142.5 ;
        RECT 450.275 142.2 480 142.35 ;
        RECT 450.425 142.05 480 142.2 ;
        RECT 450.575 141.9 480 142.05 ;
        RECT 450.725 141.75 480 141.9 ;
        RECT 450.875 141.6 480 141.75 ;
        RECT 451.025 141.45 480 141.6 ;
        RECT 451.175 141.3 480 141.45 ;
        RECT 451.325 141.15 480 141.3 ;
        RECT 451.475 141 480 141.15 ;
        RECT 451.625 140.85 480 141 ;
        RECT 451.775 140.7 480 140.85 ;
        RECT 451.925 140.55 480 140.7 ;
        RECT 452.075 140.4 480 140.55 ;
        RECT 452.225 140.25 480 140.4 ;
        RECT 452.375 140.1 480 140.25 ;
        RECT 452.525 139.95 480 140.1 ;
        RECT 452.675 139.8 480 139.95 ;
        RECT 452.825 139.65 480 139.8 ;
        RECT 452.975 139.5 480 139.65 ;
        RECT 453.125 139.35 480 139.5 ;
        RECT 453.275 139.2 480 139.35 ;
        RECT 453.425 139.05 480 139.2 ;
        RECT 453.575 138.9 480 139.05 ;
        RECT 453.725 138.75 480 138.9 ;
        RECT 453.875 138.6 480 138.75 ;
        RECT 454.025 138.45 480 138.6 ;
        RECT 454.175 138.3 480 138.45 ;
        RECT 454.325 138.15 480 138.3 ;
        RECT 454.475 138 480 138.15 ;
        RECT 454.625 137.85 480 138 ;
        RECT 454.775 137.7 480 137.85 ;
        RECT 454.925 137.55 480 137.7 ;
        RECT 455.075 137.4 480 137.55 ;
        RECT 455.225 137.25 480 137.4 ;
        RECT 455.375 137.1 480 137.25 ;
        RECT 455.525 136.95 480 137.1 ;
        RECT 455.675 136.8 480 136.95 ;
        RECT 455.825 136.65 480 136.8 ;
        RECT 455.975 136.5 480 136.65 ;
        RECT 456.125 136.35 480 136.5 ;
        RECT 456.275 136.2 480 136.35 ;
        RECT 456.425 136.05 480 136.2 ;
        RECT 456.575 135.9 480 136.05 ;
        RECT 456.725 135.75 480 135.9 ;
        RECT 456.875 135.6 480 135.75 ;
        RECT 457.025 135.45 480 135.6 ;
        RECT 457.175 135.3 480 135.45 ;
        RECT 457.325 135.15 480 135.3 ;
        RECT 457.475 135 480 135.15 ;
        RECT 457.625 134.85 480 135 ;
        RECT 457.775 134.7 480 134.85 ;
        RECT 457.925 134.55 480 134.7 ;
        RECT 458.075 134.4 480 134.55 ;
        RECT 458.225 134.25 480 134.4 ;
        RECT 458.375 134.1 480 134.25 ;
        RECT 458.525 133.95 480 134.1 ;
        RECT 458.675 133.8 480 133.95 ;
        RECT 458.825 133.65 480 133.8 ;
        RECT 458.975 133.5 480 133.65 ;
        RECT 459.125 133.35 480 133.5 ;
        RECT 459.275 133.2 480 133.35 ;
        RECT 459.425 133.05 480 133.2 ;
        RECT 459.575 132.9 480 133.05 ;
        RECT 459.725 132.75 480 132.9 ;
        RECT 459.875 132.6 480 132.75 ;
        RECT 460.025 132.45 480 132.6 ;
        RECT 460.175 132.3 480 132.45 ;
        RECT 460.325 132.15 480 132.3 ;
        RECT 460.475 132 480 132.15 ;
        RECT 460.625 131.85 480 132 ;
        RECT 460.775 131.7 480 131.85 ;
        RECT 460.925 131.55 480 131.7 ;
        RECT 461.075 131.4 480 131.55 ;
        RECT 461.225 131.25 480 131.4 ;
        RECT 461.375 131.1 480 131.25 ;
        RECT 461.525 130.95 480 131.1 ;
        RECT 461.675 130.8 480 130.95 ;
        RECT 461.825 130.65 480 130.8 ;
        RECT 461.975 130.5 480 130.65 ;
        RECT 462.125 130.35 480 130.5 ;
        RECT 462.275 130.2 480 130.35 ;
        RECT 462.425 130.05 480 130.2 ;
        RECT 462.575 129.9 480 130.05 ;
        RECT 462.725 129.75 480 129.9 ;
        RECT 462.875 129.6 480 129.75 ;
        RECT 463.025 129.45 480 129.6 ;
        RECT 463.175 129.3 480 129.45 ;
        RECT 463.325 129.15 480 129.3 ;
        RECT 463.475 129 480 129.15 ;
        RECT 463.625 128.85 480 129 ;
        RECT 463.775 128.7 480 128.85 ;
        RECT 463.925 128.55 480 128.7 ;
        RECT 464.075 128.4 480 128.55 ;
        RECT 464.225 128.25 480 128.4 ;
        RECT 464.375 128.1 480 128.25 ;
        RECT 464.525 127.95 480 128.1 ;
        RECT 464.675 127.8 480 127.95 ;
        RECT 464.825 127.65 480 127.8 ;
        RECT 464.975 127.5 480 127.65 ;
        RECT 465.125 127.35 480 127.5 ;
        RECT 465.275 127.2 480 127.35 ;
        RECT 465.425 127.05 480 127.2 ;
        RECT 465.575 126.9 480 127.05 ;
        RECT 465.725 126.75 480 126.9 ;
        RECT 465.875 126.6 480 126.75 ;
        RECT 466.025 126.45 480 126.6 ;
        RECT 466.175 126.3 480 126.45 ;
        RECT 466.325 126.15 480 126.3 ;
        RECT 466.475 126 480 126.15 ;
        RECT 466.625 125.85 480 126 ;
        RECT 466.775 125.7 480 125.85 ;
        RECT 466.925 125.55 480 125.7 ;
        RECT 467.075 125.4 480 125.55 ;
        RECT 467.225 125.25 480 125.4 ;
        RECT 467.375 125.1 480 125.25 ;
        RECT 467.525 124.95 480 125.1 ;
        RECT 467.675 124.8 480 124.95 ;
        RECT 467.825 124.65 480 124.8 ;
        RECT 467.975 124.5 480 124.65 ;
        RECT 468.125 124.35 480 124.5 ;
        RECT 468.275 124.2 480 124.35 ;
        RECT 468.425 124.05 480 124.2 ;
        RECT 468.575 123.9 480 124.05 ;
        RECT 468.725 123.75 480 123.9 ;
        RECT 0 123.75 28.815 123.8 ;
        RECT 0 123.8 28.865 123.85 ;
        RECT 0 123.85 28.93 123.865 ;
    END
  END vddio

  PIN vddio_q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 117.9 480 122.15 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 117.8 480 122.25 ;
    END
  END vddio_q

  PIN pad[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 218.815 132.205 284.215 194.545 ;
        RECT 219.215 194.545 283.815 194.945 ;
        RECT 219.615 194.945 283.415 195.345 ;
        RECT 220.015 195.345 283.015 195.745 ;
        RECT 220.415 195.745 282.615 196.145 ;
        RECT 220.815 196.145 282.215 196.545 ;
        RECT 221.215 196.545 281.815 196.945 ;
        RECT 221.615 196.945 281.415 197.345 ;
        RECT 222.015 197.345 281.015 197.745 ;
        RECT 222.415 197.745 280.615 198.145 ;
        RECT 222.815 198.145 280.215 198.545 ;
        RECT 223.215 198.545 279.815 198.945 ;
        RECT 223.615 198.945 279.415 199.345 ;
        RECT 224.015 199.345 279.015 199.745 ;
        RECT 224.415 199.745 278.615 200.145 ;
        RECT 224.815 200.145 278.215 200.545 ;
        RECT 225.215 200.545 277.815 200.945 ;
        RECT 225.345 200.945 277.685 201.075 ;
        RECT 225.345 125.675 277.685 126.075 ;
        RECT 224.945 126.075 278.085 126.475 ;
        RECT 224.545 126.475 278.485 126.875 ;
        RECT 224.145 126.875 278.885 127.275 ;
        RECT 223.745 127.275 279.285 127.675 ;
        RECT 223.345 127.675 279.685 128.075 ;
        RECT 222.945 128.075 280.085 128.475 ;
        RECT 222.545 128.475 280.485 128.875 ;
        RECT 222.145 128.875 280.885 129.275 ;
        RECT 221.745 129.275 281.285 129.675 ;
        RECT 221.345 129.675 281.685 130.075 ;
        RECT 220.945 130.075 282.085 130.475 ;
        RECT 220.545 130.475 282.485 130.875 ;
        RECT 220.145 130.875 282.885 131.275 ;
        RECT 219.745 131.275 283.285 131.675 ;
        RECT 219.345 131.675 283.685 132.075 ;
        RECT 218.945 132.075 284.085 132.205 ;
    END
    ANTENNADIFFAREA 3991.436 LAYER met1 ;
    ANTENNADIFFAREA 3991.436 LAYER met2 ;
    ANTENNADIFFAREA 3991.436 LAYER met3 ;
    ANTENNADIFFAREA 3991.436 LAYER met4 ;
    ANTENNADIFFAREA 3991.436 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 200.987 LAYER met5 ;
  END pad[1]

  PIN vssio_q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 112.05 480 116.3 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 111.95 480 116.4 ;
    END
  END vssio_q

  PIN pad[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 105.79 132.205 171.19 194.545 ;
        RECT 106.19 194.545 170.79 194.945 ;
        RECT 106.59 194.945 170.39 195.345 ;
        RECT 106.99 195.345 169.99 195.745 ;
        RECT 107.39 195.745 169.59 196.145 ;
        RECT 107.79 196.145 169.19 196.545 ;
        RECT 108.19 196.545 168.79 196.945 ;
        RECT 108.59 196.945 168.39 197.345 ;
        RECT 108.99 197.345 167.99 197.745 ;
        RECT 109.39 197.745 167.59 198.145 ;
        RECT 109.79 198.145 167.19 198.545 ;
        RECT 110.19 198.545 166.79 198.945 ;
        RECT 110.59 198.945 166.39 199.345 ;
        RECT 110.99 199.345 165.99 199.745 ;
        RECT 111.39 199.745 165.59 200.145 ;
        RECT 111.79 200.145 165.19 200.545 ;
        RECT 112.19 200.545 164.79 200.945 ;
        RECT 112.32 200.945 164.66 201.075 ;
        RECT 112.32 125.675 164.66 126.075 ;
        RECT 111.92 126.075 165.06 126.475 ;
        RECT 111.52 126.475 165.46 126.875 ;
        RECT 111.12 126.875 165.86 127.275 ;
        RECT 110.72 127.275 166.26 127.675 ;
        RECT 110.32 127.675 166.66 128.075 ;
        RECT 109.92 128.075 167.06 128.475 ;
        RECT 109.52 128.475 167.46 128.875 ;
        RECT 109.12 128.875 167.86 129.275 ;
        RECT 108.72 129.275 168.26 129.675 ;
        RECT 108.32 129.675 168.66 130.075 ;
        RECT 107.92 130.075 169.06 130.475 ;
        RECT 107.52 130.475 169.46 130.875 ;
        RECT 107.12 130.875 169.86 131.275 ;
        RECT 106.72 131.275 170.26 131.675 ;
        RECT 106.32 131.675 170.66 132.075 ;
        RECT 105.92 132.075 171.06 132.205 ;
    END
    ANTENNADIFFAREA 3991.436 LAYER met1 ;
    ANTENNADIFFAREA 3991.436 LAYER met2 ;
    ANTENNADIFFAREA 3991.436 LAYER met3 ;
    ANTENNADIFFAREA 3991.436 LAYER met4 ;
    ANTENNADIFFAREA 3991.436 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 200.987 LAYER met5 ;
  END pad[0]

  PIN vssio
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 79.65 480 84.1 ;
    END
    PORT
      LAYER met5 ;
        RECT 0 229.5 480 253.715 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 79.55 480 84.2 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 229.5 480 253.715 ;
    END
  END vssio

  PIN vswitch
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 85.7 480 88.95 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 85.6 480 89.05 ;
    END
  END vswitch

  PIN vssa
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 90.55 480 93.8 ;
    END
    PORT
      LAYER met5 ;
        RECT 0 101.45 480 110.45 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 90.45 480 93.9 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 101.45 480 101.78 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 105.36 480 106.54 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 110.12 480 110.45 ;
    END
  END vssa

  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 95.4 480 99.85 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 95.3 480 99.95 ;
    END
  END vssd
  OBS
    LAYER met2 ;
      RECT 248.14 1.935 248.23 2.025 ;
      RECT 141.685 1.935 141.865 2.025 ;
      RECT 280.055 1.895 282.18 17.295 ;
      RECT 107.825 1.895 109.95 17.295 ;
      RECT 248.945 1.82 254.03 2.025 ;
      RECT 135.975 1.82 140.855 2.025 ;
      RECT 304.885 0 402.7 23.28 ;
      RECT 403.24 0 404.855 14.71 ;
      RECT 405.395 0 419.305 5.175 ;
      RECT 419.845 0 422.55 5.175 ;
      RECT 453.555 0 453.765 237.35 ;
      RECT 452.805 0 453.015 237.03 ;
      RECT 452.055 0 452.265 236.71 ;
      RECT 451.305 0 451.515 236.39 ;
      RECT 450.555 0 450.765 236.07 ;
      RECT 449.805 0 450.015 83.685 ;
      RECT 448.305 0 448.515 83.5 ;
      RECT 449.055 0 449.265 83.455 ;
      RECT 454.305 0 464.39 60.435 ;
      RECT 465.31 0 465.89 60.435 ;
      RECT 466.81 0 480 60.435 ;
      RECT 423.09 0 444.7 23.155 ;
      RECT 445.24 0 447.765 22.245 ;
      RECT 240.34 0 241.99 28.31 ;
      RECT 268.69 0 279.515 17.525 ;
      RECT 242.93 0 247.2 10.73 ;
      RECT 254.97 0 261.48 10.235 ;
      RECT 262.02 0 268.15 10.005 ;
      RECT 283.435 1.41 302.77 2.125 ;
      RECT 248.14 0 248.32 1.935 ;
      RECT 280.055 1.18 282.18 1.895 ;
      RECT 248.945 0 254.03 1.82 ;
      RECT 283.435 0 302.77 1.41 ;
      RECT 280.055 0 282.895 1.18 ;
      RECT 110.49 0 121.315 17.525 ;
      RECT 179.13 0 210.875 24.37 ;
      RECT 234.165 0 235.795 33.975 ;
      RECT 213.155 0 233.225 24.37 ;
      RECT 236.735 0 239.8 2.13 ;
      RECT 154.21 0 155.84 33.975 ;
      RECT 148.015 0 149.665 28.31 ;
      RECT 156.78 0 176.85 24.37 ;
      RECT 142.805 0 147.075 10.73 ;
      RECT 128.525 0 135.035 10.235 ;
      RECT 121.855 0 127.985 10.005 ;
      RECT 150.205 0 153.27 2.155 ;
      RECT 141.685 0 141.865 1.935 ;
      RECT 135.975 0 141.06 1.82 ;
      RECT 0 0 85.12 30.685 ;
      RECT 87.235 1.41 107.285 2.125 ;
      RECT 107.11 1.18 109.95 1.895 ;
      RECT 87.235 0 106.57 1.41 ;
      RECT 107.11 0 109.95 1.18 ;
      RECT 268.69 36.24 279.77 36.26 ;
      RECT 110.215 36.24 121.315 36.26 ;
      RECT 236.335 35.085 239.8 42.155 ;
      RECT 150.205 35.085 153.67 42.155 ;
      RECT 154.21 33.975 235.795 41.925 ;
      RECT 280.33 33.375 447.765 36.47 ;
      RECT 0 33.375 109.675 36.47 ;
      RECT 156.38 33.235 233.625 33.975 ;
      RECT 236.735 31.7 239.8 35.085 ;
      RECT 150.205 31.7 153.27 35.085 ;
      RECT 240.34 31.205 241.99 46.275 ;
      RECT 148.015 31.205 149.665 46.275 ;
      RECT 236.735 31.16 239.8 31.7 ;
      RECT 150.745 31.16 153.27 31.7 ;
      RECT 303.9 30.685 447.765 33.375 ;
      RECT 0 30.685 86.105 33.375 ;
      RECT 239.8 30.665 241.99 31.205 ;
      RECT 148.015 30.665 149.665 31.205 ;
      RECT 256.01 30.43 261.745 42.465 ;
      RECT 254.57 30.43 255.47 36.505 ;
      RECT 128.26 30.43 133.995 42.465 ;
      RECT 134.535 30.43 135.435 36.505 ;
      RECT 254.57 30.385 255.47 30.43 ;
      RECT 256.055 30.385 261.745 30.43 ;
      RECT 128.26 30.385 133.995 30.43 ;
      RECT 134.58 30.385 135.435 30.43 ;
      RECT 254.57 30.025 255.315 30.385 ;
      RECT 135.045 30.025 135.435 30.385 ;
      RECT 256.39 29.845 261.745 30.385 ;
      RECT 128.26 29.845 133.615 30.385 ;
      RECT 255.5 29.8 261.745 29.845 ;
      RECT 128.26 29.8 134.46 29.845 ;
      RECT 254.57 29.54 254.96 30.025 ;
      RECT 135.045 29.54 135.435 30.025 ;
      RECT 255.5 29.31 261.745 29.8 ;
      RECT 254.57 29.15 254.96 29.54 ;
      RECT 128.26 29.31 134.505 29.8 ;
      RECT 239.8 28.845 241.99 30.665 ;
      RECT 148.015 28.845 150.205 30.665 ;
      RECT 254.97 28.78 261.745 29.31 ;
      RECT 128.26 28.78 134.505 29.31 ;
      RECT 242.53 28.56 243.97 46.275 ;
      RECT 146.035 28.56 147.475 46.275 ;
      RECT 150.745 28.355 153.27 31.16 ;
      RECT 236.735 28.355 239.26 31.16 ;
      RECT 244.51 28.33 254.03 37.09 ;
      RECT 135.975 28.33 145.495 37.09 ;
      RECT 240.34 28.31 241.99 28.845 ;
      RECT 148.015 28.31 150.205 28.845 ;
      RECT 242.53 27.115 243.97 28.56 ;
      RECT 236.735 27.815 239.26 28.355 ;
      RECT 150.205 27.815 153.27 28.355 ;
      RECT 242.93 26.75 254.03 28.33 ;
      RECT 135.975 26.75 145.495 28.33 ;
      RECT 262.285 24.435 268.15 43.05 ;
      RECT 121.855 24.435 127.72 43.05 ;
      RECT 156.78 24.37 233.225 33.235 ;
      RECT 254.97 24.205 261.745 28.78 ;
      RECT 128.26 24.205 135.035 28.78 ;
      RECT 262.885 23.83 268.15 24.435 ;
      RECT 121.855 23.83 127.72 24.435 ;
      RECT 254.97 23.605 261.745 24.205 ;
      RECT 127.66 23.605 135.035 24.205 ;
      RECT 304.885 23.28 447.765 30.685 ;
      RECT 423.09 23.155 447.765 23.28 ;
      RECT 445.31 22.315 447.765 23.155 ;
      RECT 445.24 22.245 447.765 22.315 ;
      RECT 280.33 18.295 302.77 33.375 ;
      RECT 87.235 18.295 109.675 33.375 ;
      RECT 268.69 17.795 279.79 36.24 ;
      RECT 110.215 17.795 121.315 36.24 ;
      RECT 280.33 17.57 282.18 18.295 ;
      RECT 107.825 17.57 109.675 18.295 ;
      RECT 268.69 17.525 279.79 17.795 ;
      RECT 110.49 17.525 121.315 17.795 ;
      RECT 280.055 17.295 282.18 17.57 ;
      RECT 107.825 17.295 109.675 17.57 ;
      RECT 403.24 15.21 422.55 23.28 ;
      RECT 403.24 14.75 404.815 15.21 ;
      RECT 403.24 14.71 404.815 14.75 ;
      RECT 405.735 14.67 422.55 15.21 ;
      RECT 405.395 14.625 422.55 14.67 ;
      RECT 254.97 11.1 262.345 23.605 ;
      RECT 127.66 11.1 135.035 23.605 ;
      RECT 262.885 10.87 268.15 23.83 ;
      RECT 121.855 10.87 127.12 23.83 ;
      RECT 242.93 10.73 254.03 26.75 ;
      RECT 135.975 10.73 147.075 26.75 ;
      RECT 254.97 10.235 262.345 11.1 ;
      RECT 128.525 10.235 135.035 11.1 ;
      RECT 262.02 10.005 268.15 10.87 ;
      RECT 121.855 10.005 127.12 10.87 ;
      RECT 247.74 7.72 254.03 10.73 ;
      RECT 135.975 7.72 142.265 10.73 ;
      RECT 405.395 5.175 422.55 14.625 ;
      RECT 236.735 3.11 239.8 27.815 ;
      RECT 150.205 3.085 153.27 27.815 ;
      RECT 236.78 3.065 239.8 3.11 ;
      RECT 150.205 3.065 153.27 3.085 ;
      RECT 248.14 2.485 254.03 7.72 ;
      RECT 135.975 2.485 141.865 7.72 ;
      RECT 236.78 2.175 239.8 3.065 ;
      RECT 150.205 2.175 153.25 3.065 ;
      RECT 150.205 2.155 153.25 2.175 ;
      RECT 236.735 2.13 239.8 2.175 ;
      RECT 282.72 2.125 302.77 18.295 ;
      RECT 87.235 2.125 107.285 18.295 ;
      RECT 249.15 2.025 254.03 2.485 ;
      RECT 248.14 2.025 248.23 2.485 ;
      RECT 141.775 2.025 141.865 2.485 ;
      RECT 135.975 2.025 140.855 2.485 ;
      RECT 297.84 111.66 446.945 111.9 ;
      RECT 0 111.66 92.405 111.9 ;
      RECT 93.485 111.36 296.52 112.28 ;
      RECT 92.735 111.315 297.225 111.36 ;
      RECT 92.735 103.125 297.27 111.315 ;
      RECT 297.84 102.925 446.945 111.66 ;
      RECT 0 102.925 92.165 111.66 ;
      RECT 100.755 95.1 297.27 103.125 ;
      RECT 289.475 94.56 446.945 102.925 ;
      RECT 0 94.56 92.165 102.925 ;
      RECT 106.235 94.31 284.56 95.1 ;
      RECT 284.335 94.105 446.945 94.56 ;
      RECT 0 94.105 105.215 94.56 ;
      RECT 106.235 89.625 283.77 94.31 ;
      RECT 284.335 89.42 446.945 94.105 ;
      RECT 0 89.42 105.67 94.105 ;
      RECT 108.15 87.71 283.77 89.625 ;
      RECT 282.395 87.48 446.945 89.42 ;
      RECT 0 87.48 105.67 89.42 ;
      RECT 447.485 86.005 450.015 235.84 ;
      RECT 282.395 85.775 446.945 87.48 ;
      RECT 449.805 83.685 450.015 86.005 ;
      RECT 282.395 83.5 446.945 85.775 ;
      RECT 449.055 83.455 449.22 83.5 ;
      RECT 108.15 76.675 281.855 87.71 ;
      RECT 0 76.45 107.61 87.48 ;
      RECT 282.395 76.45 447.765 83.5 ;
      RECT 109.78 75.05 281.855 76.675 ;
      RECT 280.765 74.82 447.765 76.45 ;
      RECT 0 74.82 107.61 76.45 ;
      RECT 454.305 60.435 480 237.67 ;
      RECT 109.78 58.665 280.225 75.05 ;
      RECT 150.585 58.125 239.42 58.665 ;
      RECT 150.205 58.08 239.755 58.125 ;
      RECT 280.765 57.435 447.765 74.82 ;
      RECT 0 57.435 109.24 74.82 ;
      RECT 240.34 57.205 280.225 58.665 ;
      RECT 109.78 57.205 149.665 58.665 ;
      RECT 281.575 56.625 447.765 57.435 ;
      RECT 0 56.625 109.24 57.435 ;
      RECT 240.34 56.395 280.225 57.205 ;
      RECT 108.97 56.395 149.665 57.205 ;
      RECT 240.34 51.985 281.035 56.395 ;
      RECT 108.97 51.985 149.665 56.395 ;
      RECT 240.34 49.755 263.81 51.985 ;
      RECT 126.195 49.755 149.665 51.985 ;
      RECT 244.89 49.215 263.81 49.755 ;
      RECT 126.195 49.215 145.115 49.755 ;
      RECT 244.51 49.17 263.81 49.215 ;
      RECT 126.195 49.17 145.45 49.215 ;
      RECT 264.795 48.91 281.035 51.985 ;
      RECT 244.51 48.91 263.81 49.17 ;
      RECT 108.97 48.91 125.21 51.985 ;
      RECT 126.195 48.91 145.495 49.17 ;
      RECT 244.51 48.77 263.81 48.91 ;
      RECT 126.055 48.77 145.495 48.91 ;
      RECT 264.49 48.605 281.035 48.91 ;
      RECT 108.97 48.605 125.21 48.91 ;
      RECT 264.49 47.63 281.035 48.605 ;
      RECT 108.97 47.63 125.515 48.605 ;
      RECT 264.49 47.53 281.035 47.63 ;
      RECT 109.07 47.53 125.515 47.63 ;
      RECT 281.575 47.4 447.765 56.625 ;
      RECT 0 47.4 108.43 56.625 ;
      RECT 244.51 47.3 263.95 48.77 ;
      RECT 126.055 47.3 145.495 48.77 ;
      RECT 265.285 46.735 280.935 47.53 ;
      RECT 109.865 46.735 125.515 47.53 ;
      RECT 280.68 46.505 447.765 47.4 ;
      RECT 0 46.505 108.43 47.4 ;
      RECT 265.6 46.42 280.14 46.735 ;
      RECT 109.865 46.42 124.72 46.735 ;
      RECT 240.34 46.275 243.97 49.755 ;
      RECT 146.035 46.275 149.665 49.755 ;
      RECT 268.69 46.02 280.14 46.42 ;
      RECT 109.865 46.02 121.315 46.42 ;
      RECT 244.51 45.88 263.95 47.3 ;
      RECT 124.63 45.88 145.495 47.3 ;
      RECT 280.68 45.79 447.765 46.505 ;
      RECT 0 45.79 109.325 46.505 ;
      RECT 244.51 45.78 268.05 45.88 ;
      RECT 121.855 45.78 145.495 45.88 ;
      RECT 268.69 45.65 280.14 46.02 ;
      RECT 110.235 45.65 121.315 46.02 ;
      RECT 280.31 45.42 447.765 45.79 ;
      RECT 0 45.42 109.325 45.79 ;
      RECT 244.51 43.05 268.15 45.78 ;
      RECT 150.205 43.05 239.8 58.08 ;
      RECT 121.855 43.05 145.495 45.78 ;
      RECT 244.51 42.88 260.985 43.05 ;
      RECT 129.02 42.88 145.495 43.05 ;
      RECT 256.01 42.51 260.985 42.88 ;
      RECT 129.02 42.51 133.995 42.88 ;
      RECT 256.01 42.465 261.7 42.51 ;
      RECT 128.26 42.465 133.995 42.51 ;
      RECT 236.325 42.165 239.8 43.05 ;
      RECT 150.205 42.165 153.68 43.05 ;
      RECT 236.335 42.155 239.8 42.165 ;
      RECT 150.205 42.155 153.68 42.165 ;
      RECT 154.22 41.935 235.785 43.05 ;
      RECT 154.21 41.925 235.785 41.935 ;
      RECT 244.51 37.09 255.47 42.88 ;
      RECT 134.535 37.09 145.495 42.88 ;
      RECT 254.95 36.55 255.47 37.09 ;
      RECT 134.535 36.55 135.055 37.09 ;
      RECT 254.57 36.505 255.47 36.55 ;
      RECT 134.535 36.505 135.39 36.55 ;
      RECT 280.31 36.49 447.765 45.42 ;
      RECT 0 36.49 109.695 45.42 ;
      RECT 280.33 36.47 447.765 36.49 ;
      RECT 0 36.47 109.695 36.49 ;
      RECT 268.69 36.26 279.77 45.65 ;
      RECT 110.235 36.26 121.315 45.65 ;
      RECT 0 245.955 480 253.715 ;
      RECT 0 245.555 449.105 245.955 ;
      RECT 0 245.155 448.355 245.555 ;
      RECT 0 244.755 447.605 245.155 ;
      RECT 0 244.295 446.78 244.755 ;
      RECT 0 244.13 446.78 244.295 ;
      RECT 447.485 244.11 447.605 244.215 ;
      RECT 449.645 242.365 480 245.955 ;
      RECT 449.645 241.925 450.975 242.365 ;
      RECT 451.145 241.7 451.23 241.825 ;
      RECT 449.645 240.855 450.605 241.925 ;
      RECT 451.895 240.08 480 242.365 ;
      RECT 451.145 239.85 451.355 241.7 ;
      RECT 451.145 239.76 451.355 239.85 ;
      RECT 450.395 239.53 450.605 240.855 ;
      RECT 450.395 239.44 450.605 239.53 ;
      RECT 449.645 239.21 449.855 240.855 ;
      RECT 449.645 239.12 449.855 239.21 ;
      RECT 448.895 238.89 449.105 245.555 ;
      RECT 448.895 238.8 449.105 238.89 ;
      RECT 448.145 238.57 448.355 245.155 ;
      RECT 448.145 238.48 448.355 238.57 ;
      RECT 447.485 238.25 447.605 244.11 ;
      RECT 454.305 237.67 480 240.08 ;
      RECT 453.555 237.35 453.765 237.44 ;
      RECT 452.805 237.03 453.015 237.12 ;
      RECT 452.055 236.71 452.265 236.8 ;
      RECT 451.305 236.39 451.515 236.48 ;
      RECT 450.555 236.07 450.765 236.16 ;
      RECT 447.485 235.84 447.605 238.25 ;
      RECT 0 112.28 446.945 244.13 ;
      RECT 297.06 111.96 446.945 112.28 ;
      RECT 0 111.96 92.945 112.28 ;
      RECT 297.12 111.9 446.945 111.96 ;
      RECT 0 111.9 92.945 111.96 ;
      RECT 449.455 84.23 449.875 84.3 ;
      RECT 449.525 84.16 449.875 84.23 ;
      RECT 449.595 84.09 449.875 84.16 ;
      RECT 449.665 84.02 449.875 84.09 ;
      RECT 449.735 83.95 449.875 84.02 ;
      RECT 449.805 83.88 449.875 83.95 ;
      RECT 447.625 235.785 449.805 235.855 ;
      RECT 447.625 235.855 449.735 235.925 ;
      RECT 447.625 235.925 449.665 235.995 ;
      RECT 447.625 235.995 449.595 236.065 ;
      RECT 447.625 236.065 449.525 236.135 ;
      RECT 447.625 236.135 449.455 236.205 ;
      RECT 447.625 236.205 449.385 236.275 ;
      RECT 447.625 236.275 449.315 236.345 ;
      RECT 447.625 236.345 449.245 236.415 ;
      RECT 447.625 236.415 449.175 236.485 ;
      RECT 447.625 236.485 449.105 236.555 ;
      RECT 447.625 236.555 449.035 236.625 ;
      RECT 447.625 236.625 448.965 236.695 ;
      RECT 447.625 236.695 448.895 236.765 ;
      RECT 447.625 236.765 448.825 236.835 ;
      RECT 447.625 236.835 448.755 236.905 ;
      RECT 447.625 236.905 448.685 236.975 ;
      RECT 447.625 236.975 448.615 237.045 ;
      RECT 447.625 237.045 448.545 237.115 ;
      RECT 447.625 237.115 448.475 237.185 ;
      RECT 447.625 237.185 448.405 237.255 ;
      RECT 447.625 237.255 448.335 237.325 ;
      RECT 447.625 237.325 448.265 237.395 ;
      RECT 447.625 237.395 448.195 237.465 ;
      RECT 447.625 237.465 448.125 237.535 ;
      RECT 447.625 237.535 448.055 237.605 ;
      RECT 447.625 237.605 447.985 237.675 ;
      RECT 447.625 237.675 447.915 237.745 ;
      RECT 447.625 237.745 447.845 237.815 ;
      RECT 447.625 237.815 447.775 237.885 ;
      RECT 447.625 237.885 447.705 237.955 ;
      RECT 447.625 237.955 447.635 238.025 ;
      RECT 94.935 101.12 295.07 101.19 ;
      RECT 95.005 101.05 295.0 101.12 ;
      RECT 95.075 100.98 294.93 101.05 ;
      RECT 95.145 100.91 294.86 100.98 ;
      RECT 95.215 100.84 294.79 100.91 ;
      RECT 95.285 100.77 294.72 100.84 ;
      RECT 95.355 100.7 294.65 100.77 ;
      RECT 95.425 100.63 294.58 100.7 ;
      RECT 95.495 100.56 294.51 100.63 ;
      RECT 95.565 100.49 294.44 100.56 ;
      RECT 95.635 100.42 294.37 100.49 ;
      RECT 95.705 100.35 294.3 100.42 ;
      RECT 95.775 100.28 294.23 100.35 ;
      RECT 95.845 100.21 294.16 100.28 ;
      RECT 95.915 100.14 294.09 100.21 ;
      RECT 95.985 100.07 294.02 100.14 ;
      RECT 96.055 100 293.95 100.07 ;
      RECT 96.125 99.93 293.88 100 ;
      RECT 96.195 99.86 293.81 99.93 ;
      RECT 96.265 99.79 293.74 99.86 ;
      RECT 96.335 99.72 293.67 99.79 ;
      RECT 96.405 99.65 293.6 99.72 ;
      RECT 96.475 99.58 293.53 99.65 ;
      RECT 96.545 99.51 293.46 99.58 ;
      RECT 96.615 99.44 293.39 99.51 ;
      RECT 96.685 99.37 293.32 99.44 ;
      RECT 96.755 99.3 293.25 99.37 ;
      RECT 96.825 99.23 293.18 99.3 ;
      RECT 96.895 99.16 293.11 99.23 ;
      RECT 96.965 99.09 293.04 99.16 ;
      RECT 97.035 99.02 292.97 99.09 ;
      RECT 97.105 98.95 292.9 99.02 ;
      RECT 97.175 98.88 292.83 98.95 ;
      RECT 97.245 98.81 292.76 98.88 ;
      RECT 97.315 98.74 292.69 98.81 ;
      RECT 97.385 98.67 292.62 98.74 ;
      RECT 97.455 98.6 292.55 98.67 ;
      RECT 97.525 98.53 292.48 98.6 ;
      RECT 97.595 98.46 292.41 98.53 ;
      RECT 97.665 98.39 292.34 98.46 ;
      RECT 97.735 98.32 292.27 98.39 ;
      RECT 97.805 98.25 292.2 98.32 ;
      RECT 97.875 98.18 292.13 98.25 ;
      RECT 97.945 98.11 292.06 98.18 ;
      RECT 98.015 98.04 291.99 98.11 ;
      RECT 98.085 97.97 291.92 98.04 ;
      RECT 98.155 97.9 291.85 97.97 ;
      RECT 98.225 97.83 291.78 97.9 ;
      RECT 98.295 97.76 291.71 97.83 ;
      RECT 98.365 97.69 291.64 97.76 ;
      RECT 98.435 97.62 291.57 97.69 ;
      RECT 98.505 97.55 291.5 97.62 ;
      RECT 98.575 97.48 291.43 97.55 ;
      RECT 98.645 97.41 291.36 97.48 ;
      RECT 98.715 97.34 291.29 97.41 ;
      RECT 98.785 97.27 291.22 97.34 ;
      RECT 98.855 97.2 291.15 97.27 ;
      RECT 98.925 97.13 291.08 97.2 ;
      RECT 98.995 97.06 291.01 97.13 ;
      RECT 99.065 96.99 290.94 97.06 ;
      RECT 99.135 96.92 290.87 96.99 ;
      RECT 99.205 96.85 290.8 96.92 ;
      RECT 99.275 96.78 290.73 96.85 ;
      RECT 99.345 96.71 290.66 96.78 ;
      RECT 99.415 96.64 290.59 96.71 ;
      RECT 99.485 96.57 290.52 96.64 ;
      RECT 99.555 96.5 290.45 96.57 ;
      RECT 99.625 96.43 290.38 96.5 ;
      RECT 99.695 96.36 290.31 96.43 ;
      RECT 99.765 96.29 290.24 96.36 ;
      RECT 99.835 96.22 290.17 96.29 ;
      RECT 99.905 96.15 290.1 96.22 ;
      RECT 99.975 96.08 290.03 96.15 ;
      RECT 100.045 96.01 289.96 96.08 ;
      RECT 100.115 95.94 289.89 96.01 ;
      RECT 100.185 95.87 289.82 95.94 ;
      RECT 100.255 95.8 289.75 95.87 ;
      RECT 100.325 95.73 289.68 95.8 ;
      RECT 100.395 95.66 289.61 95.73 ;
      RECT 100.465 95.59 289.54 95.66 ;
      RECT 100.535 95.52 289.47 95.59 ;
      RECT 100.605 95.45 289.4 95.52 ;
      RECT 100.675 95.38 289.33 95.45 ;
      RECT 100.745 95.31 289.26 95.38 ;
      RECT 100.815 95.24 289.19 95.31 ;
      RECT 0 244.075 446.735 244.145 ;
      RECT 0 244.145 446.665 244.215 ;
      RECT 0 244.215 446.64 244.24 ;
      RECT 297.655 112.04 446.805 112.11 ;
      RECT 297.585 112.11 446.805 112.18 ;
      RECT 297.515 112.18 446.805 112.25 ;
      RECT 297.445 112.25 446.805 112.32 ;
      RECT 297.375 112.32 446.805 112.39 ;
      RECT 297.305 112.39 446.805 112.42 ;
      RECT 297.98 111.715 446.805 111.785 ;
      RECT 297.91 111.785 446.805 111.855 ;
      RECT 297.84 111.855 446.805 111.925 ;
      RECT 297.77 111.925 446.805 111.995 ;
      RECT 297.7 111.995 446.805 112.04 ;
      RECT 447.625 86.06 449.875 235.785 ;
      RECT 447.635 86.05 449.875 86.06 ;
      RECT 447.705 85.98 449.875 86.05 ;
      RECT 447.775 85.91 449.875 85.98 ;
      RECT 447.845 85.84 449.875 85.91 ;
      RECT 447.915 85.77 449.875 85.84 ;
      RECT 447.985 85.7 449.875 85.77 ;
      RECT 448.055 85.63 449.875 85.7 ;
      RECT 448.125 85.56 449.875 85.63 ;
      RECT 448.195 85.49 449.875 85.56 ;
      RECT 448.265 85.42 449.875 85.49 ;
      RECT 448.335 85.35 449.875 85.42 ;
      RECT 448.405 85.28 449.875 85.35 ;
      RECT 448.475 85.21 449.875 85.28 ;
      RECT 448.545 85.14 449.875 85.21 ;
      RECT 448.615 85.07 449.875 85.14 ;
      RECT 448.685 85 449.875 85.07 ;
      RECT 448.755 84.93 449.875 85 ;
      RECT 448.825 84.86 449.875 84.93 ;
      RECT 448.895 84.79 449.875 84.86 ;
      RECT 448.965 84.72 449.875 84.79 ;
      RECT 449.035 84.65 449.875 84.72 ;
      RECT 449.105 84.58 449.875 84.65 ;
      RECT 449.175 84.51 449.875 84.58 ;
      RECT 449.245 84.44 449.875 84.51 ;
      RECT 449.315 84.37 449.875 84.44 ;
      RECT 449.385 84.3 449.875 84.37 ;
      RECT 296.32 101.14 446.805 101.21 ;
      RECT 296.25 101.07 446.805 101.14 ;
      RECT 296.18 101 446.805 101.07 ;
      RECT 296.11 100.93 446.805 101 ;
      RECT 296.04 100.86 446.805 100.93 ;
      RECT 295.97 100.79 446.805 100.86 ;
      RECT 295.9 100.72 446.805 100.79 ;
      RECT 295.83 100.65 446.805 100.72 ;
      RECT 295.76 100.58 446.805 100.65 ;
      RECT 295.69 100.51 446.805 100.58 ;
      RECT 295.62 100.44 446.805 100.51 ;
      RECT 295.55 100.37 446.805 100.44 ;
      RECT 295.48 100.3 446.805 100.37 ;
      RECT 295.41 100.23 446.805 100.3 ;
      RECT 295.34 100.16 446.805 100.23 ;
      RECT 295.27 100.09 446.805 100.16 ;
      RECT 295.2 100.02 446.805 100.09 ;
      RECT 295.13 99.95 446.805 100.02 ;
      RECT 295.06 99.88 446.805 99.95 ;
      RECT 294.99 99.81 446.805 99.88 ;
      RECT 294.92 99.74 446.805 99.81 ;
      RECT 294.85 99.67 446.805 99.74 ;
      RECT 294.78 99.6 446.805 99.67 ;
      RECT 294.71 99.53 446.805 99.6 ;
      RECT 294.64 99.46 446.805 99.53 ;
      RECT 294.57 99.39 446.805 99.46 ;
      RECT 294.5 99.32 446.805 99.39 ;
      RECT 294.43 99.25 446.805 99.32 ;
      RECT 294.36 99.18 446.805 99.25 ;
      RECT 294.29 99.11 446.805 99.18 ;
      RECT 294.22 99.04 446.805 99.11 ;
      RECT 294.15 98.97 446.805 99.04 ;
      RECT 294.08 98.9 446.805 98.97 ;
      RECT 294.01 98.83 446.805 98.9 ;
      RECT 293.94 98.76 446.805 98.83 ;
      RECT 293.87 98.69 446.805 98.76 ;
      RECT 293.8 98.62 446.805 98.69 ;
      RECT 293.73 98.55 446.805 98.62 ;
      RECT 293.66 98.48 446.805 98.55 ;
      RECT 293.59 98.41 446.805 98.48 ;
      RECT 293.52 98.34 446.805 98.41 ;
      RECT 293.45 98.27 446.805 98.34 ;
      RECT 293.38 98.2 446.805 98.27 ;
      RECT 293.31 98.13 446.805 98.2 ;
      RECT 293.24 98.06 446.805 98.13 ;
      RECT 293.17 97.99 446.805 98.06 ;
      RECT 293.1 97.92 446.805 97.99 ;
      RECT 293.03 97.85 446.805 97.92 ;
      RECT 292.96 97.78 446.805 97.85 ;
      RECT 292.89 97.71 446.805 97.78 ;
      RECT 292.82 97.64 446.805 97.71 ;
      RECT 292.75 97.57 446.805 97.64 ;
      RECT 292.68 97.5 446.805 97.57 ;
      RECT 292.61 97.43 446.805 97.5 ;
      RECT 292.54 97.36 446.805 97.43 ;
      RECT 292.47 97.29 446.805 97.36 ;
      RECT 292.4 97.22 446.805 97.29 ;
      RECT 292.33 97.15 446.805 97.22 ;
      RECT 292.26 97.08 446.805 97.15 ;
      RECT 292.19 97.01 446.805 97.08 ;
      RECT 292.12 96.94 446.805 97.01 ;
      RECT 292.05 96.87 446.805 96.94 ;
      RECT 291.98 96.8 446.805 96.87 ;
      RECT 291.91 96.73 446.805 96.8 ;
      RECT 291.84 96.66 446.805 96.73 ;
      RECT 291.77 96.59 446.805 96.66 ;
      RECT 291.7 96.52 446.805 96.59 ;
      RECT 291.63 96.45 446.805 96.52 ;
      RECT 291.56 96.38 446.805 96.45 ;
      RECT 291.49 96.31 446.805 96.38 ;
      RECT 291.42 96.24 446.805 96.31 ;
      RECT 291.35 96.17 446.805 96.24 ;
      RECT 291.28 96.1 446.805 96.17 ;
      RECT 291.21 96.03 446.805 96.1 ;
      RECT 291.14 95.96 446.805 96.03 ;
      RECT 291.07 95.89 446.805 95.96 ;
      RECT 291.0 95.82 446.805 95.89 ;
      RECT 290.93 95.75 446.805 95.82 ;
      RECT 290.86 95.68 446.805 95.75 ;
      RECT 290.79 95.61 446.805 95.68 ;
      RECT 290.72 95.54 446.805 95.61 ;
      RECT 290.65 95.47 446.805 95.54 ;
      RECT 290.58 95.4 446.805 95.47 ;
      RECT 290.51 95.33 446.805 95.4 ;
      RECT 290.44 95.26 446.805 95.33 ;
      RECT 290.37 95.19 446.805 95.26 ;
      RECT 290.3 95.12 446.805 95.19 ;
      RECT 290.23 95.05 446.805 95.12 ;
      RECT 290.16 94.98 446.805 95.05 ;
      RECT 290.09 94.91 446.805 94.98 ;
      RECT 290.02 94.84 446.805 94.91 ;
      RECT 289.95 94.77 446.805 94.84 ;
      RECT 289.88 94.7 446.805 94.77 ;
      RECT 289.81 94.63 446.805 94.7 ;
      RECT 289.74 94.56 446.805 94.63 ;
      RECT 289.67 94.49 446.805 94.56 ;
      RECT 289.6 94.42 446.805 94.49 ;
      RECT 92.905 103.15 297.1 103.18 ;
      RECT 92.975 103.08 297.03 103.15 ;
      RECT 93.045 103.01 296.96 103.08 ;
      RECT 93.115 102.94 296.89 103.01 ;
      RECT 93.185 102.87 296.82 102.94 ;
      RECT 93.255 102.8 296.75 102.87 ;
      RECT 93.325 102.73 296.68 102.8 ;
      RECT 93.395 102.66 296.61 102.73 ;
      RECT 93.465 102.59 296.54 102.66 ;
      RECT 93.535 102.52 296.47 102.59 ;
      RECT 93.605 102.45 296.4 102.52 ;
      RECT 93.675 102.38 296.33 102.45 ;
      RECT 93.745 102.31 296.26 102.38 ;
      RECT 93.815 102.24 296.19 102.31 ;
      RECT 93.885 102.17 296.12 102.24 ;
      RECT 93.955 102.1 296.05 102.17 ;
      RECT 94.025 102.03 295.98 102.1 ;
      RECT 94.095 101.96 295.91 102.03 ;
      RECT 94.165 101.89 295.84 101.96 ;
      RECT 94.235 101.82 295.77 101.89 ;
      RECT 94.305 101.75 295.7 101.82 ;
      RECT 94.375 101.68 295.63 101.75 ;
      RECT 94.445 101.61 295.56 101.68 ;
      RECT 94.515 101.54 295.49 101.61 ;
      RECT 94.585 101.47 295.42 101.54 ;
      RECT 94.655 101.4 295.35 101.47 ;
      RECT 94.725 101.33 295.28 101.4 ;
      RECT 94.795 101.26 295.21 101.33 ;
      RECT 94.865 101.19 295.14 101.26 ;
      RECT 0 57.31 108.92 57.38 ;
      RECT 0 57.38 108.99 57.45 ;
      RECT 0 57.45 109.06 57.49 ;
      RECT 0 46.45 109.115 46.52 ;
      RECT 0 46.52 109.045 46.59 ;
      RECT 0 46.59 108.975 46.66 ;
      RECT 0 46.66 108.905 46.73 ;
      RECT 0 46.73 108.835 46.8 ;
      RECT 0 46.8 108.765 46.87 ;
      RECT 0 46.87 108.695 46.94 ;
      RECT 0 46.94 108.625 47.01 ;
      RECT 0 47.01 108.555 47.08 ;
      RECT 0 47.08 108.485 47.15 ;
      RECT 0 47.15 108.415 47.22 ;
      RECT 0 47.22 108.345 47.29 ;
      RECT 0 47.29 108.29 47.345 ;
      RECT 0 45.365 109.485 45.435 ;
      RECT 0 45.435 109.415 45.505 ;
      RECT 0 45.505 109.345 45.575 ;
      RECT 0 45.575 109.275 45.645 ;
      RECT 0 45.645 109.205 45.715 ;
      RECT 0 45.715 109.185 45.735 ;
      RECT 0 36.525 109.535 36.535 ;
      RECT 0 36.535 109.545 36.545 ;
      RECT 126.265 48.715 145.355 48.785 ;
      RECT 126.335 48.785 145.355 48.855 ;
      RECT 268.83 45.705 279.63 45.775 ;
      RECT 268.83 45.775 279.7 45.845 ;
      RECT 268.83 45.845 279.77 45.915 ;
      RECT 268.83 45.915 279.84 45.985 ;
      RECT 268.83 45.985 279.91 46.055 ;
      RECT 268.83 46.055 279.98 46.075 ;
      RECT 268.83 36.185 279.64 36.195 ;
      RECT 268.83 36.195 279.63 36.205 ;
      RECT 244.65 48.715 263.74 48.785 ;
      RECT 244.65 48.785 263.67 48.855 ;
      RECT 244.65 45.74 265.245 45.81 ;
      RECT 244.65 45.81 265.175 45.88 ;
      RECT 244.65 45.88 265.105 45.95 ;
      RECT 244.65 45.95 265.035 46.02 ;
      RECT 244.65 46.02 264.965 46.09 ;
      RECT 244.65 46.09 264.895 46.16 ;
      RECT 244.65 46.16 264.825 46.23 ;
      RECT 244.65 46.23 264.755 46.3 ;
      RECT 244.65 46.3 264.685 46.37 ;
      RECT 244.65 46.37 264.615 46.44 ;
      RECT 244.65 46.44 264.545 46.51 ;
      RECT 244.65 46.51 264.475 46.58 ;
      RECT 244.65 46.58 264.405 46.65 ;
      RECT 244.65 46.65 264.335 46.72 ;
      RECT 244.65 46.72 264.265 46.79 ;
      RECT 244.65 46.79 264.195 46.86 ;
      RECT 244.65 46.86 264.125 46.93 ;
      RECT 244.65 46.93 264.055 47 ;
      RECT 244.65 47 263.985 47.07 ;
      RECT 244.65 47.07 263.915 47.14 ;
      RECT 244.65 47.14 263.845 47.21 ;
      RECT 244.65 47.21 263.81 47.245 ;
      RECT 264.7 48.55 280.895 48.62 ;
      RECT 264.77 48.62 280.895 48.69 ;
      RECT 264.84 48.69 280.895 48.76 ;
      RECT 264.91 48.76 280.895 48.83 ;
      RECT 264.935 48.83 280.895 48.855 ;
      RECT 264.63 47.68 280.885 47.685 ;
      RECT 280.52 45.365 447.625 45.435 ;
      RECT 280.59 45.435 447.625 45.505 ;
      RECT 280.66 45.505 447.625 45.575 ;
      RECT 280.73 45.575 447.625 45.645 ;
      RECT 280.8 45.645 447.625 45.715 ;
      RECT 280.82 45.715 447.625 45.735 ;
      RECT 280.47 36.525 447.625 36.535 ;
      RECT 280.46 36.535 447.625 36.545 ;
      RECT 280.89 46.45 447.625 46.52 ;
      RECT 280.96 46.52 447.625 46.59 ;
      RECT 281.03 46.59 447.625 46.66 ;
      RECT 281.1 46.66 447.625 46.73 ;
      RECT 281.17 46.73 447.625 46.8 ;
      RECT 281.24 46.8 447.625 46.87 ;
      RECT 281.31 46.87 447.625 46.94 ;
      RECT 281.38 46.94 447.625 47.01 ;
      RECT 281.45 47.01 447.625 47.08 ;
      RECT 281.52 47.08 447.625 47.15 ;
      RECT 281.59 47.15 447.625 47.22 ;
      RECT 281.66 47.22 447.625 47.29 ;
      RECT 281.715 47.29 447.625 47.345 ;
      RECT 281.715 56.68 447.625 56.75 ;
      RECT 281.645 56.75 447.625 56.82 ;
      RECT 281.575 56.82 447.625 56.89 ;
      RECT 281.505 56.89 447.625 56.96 ;
      RECT 281.435 56.96 447.625 57.03 ;
      RECT 281.365 57.03 447.625 57.1 ;
      RECT 281.295 57.1 447.625 57.17 ;
      RECT 281.225 57.17 447.625 57.24 ;
      RECT 281.155 57.24 447.625 57.31 ;
      RECT 281.085 57.31 447.625 57.38 ;
      RECT 281.015 57.38 447.625 57.45 ;
      RECT 280.945 57.45 447.625 57.49 ;
      RECT 297.98 102.82 446.805 102.87 ;
      RECT 297.93 102.75 446.805 102.82 ;
      RECT 297.86 102.68 446.805 102.75 ;
      RECT 297.79 102.61 446.805 102.68 ;
      RECT 297.72 102.54 446.805 102.61 ;
      RECT 297.65 102.47 446.805 102.54 ;
      RECT 297.58 102.4 446.805 102.47 ;
      RECT 297.51 102.33 446.805 102.4 ;
      RECT 297.44 102.26 446.805 102.33 ;
      RECT 297.37 102.19 446.805 102.26 ;
      RECT 297.3 102.12 446.805 102.19 ;
      RECT 297.23 102.05 446.805 102.12 ;
      RECT 297.16 101.98 446.805 102.05 ;
      RECT 297.09 101.91 446.805 101.98 ;
      RECT 297.02 101.84 446.805 101.91 ;
      RECT 296.95 101.77 446.805 101.84 ;
      RECT 296.88 101.7 446.805 101.77 ;
      RECT 296.81 101.63 446.805 101.7 ;
      RECT 296.74 101.56 446.805 101.63 ;
      RECT 296.67 101.49 446.805 101.56 ;
      RECT 296.6 101.42 446.805 101.49 ;
      RECT 296.53 101.35 446.805 101.42 ;
      RECT 296.46 101.28 446.805 101.35 ;
      RECT 296.39 101.21 446.805 101.28 ;
      RECT 0 101.63 93.195 101.7 ;
      RECT 0 101.56 93.265 101.63 ;
      RECT 0 101.49 93.335 101.56 ;
      RECT 0 101.42 93.405 101.49 ;
      RECT 0 101.35 93.475 101.42 ;
      RECT 0 101.28 93.545 101.35 ;
      RECT 0 101.21 93.615 101.28 ;
      RECT 0 101.14 93.685 101.21 ;
      RECT 0 101.07 93.755 101.14 ;
      RECT 0 101 93.825 101.07 ;
      RECT 0 100.93 93.895 101 ;
      RECT 0 100.86 93.965 100.93 ;
      RECT 0 100.79 94.035 100.86 ;
      RECT 0 100.72 94.105 100.79 ;
      RECT 0 100.65 94.175 100.72 ;
      RECT 0 100.58 94.245 100.65 ;
      RECT 0 100.51 94.315 100.58 ;
      RECT 0 100.44 94.385 100.51 ;
      RECT 0 100.37 94.455 100.44 ;
      RECT 0 100.3 94.525 100.37 ;
      RECT 0 100.23 94.595 100.3 ;
      RECT 0 100.16 94.665 100.23 ;
      RECT 0 100.09 94.735 100.16 ;
      RECT 0 100.02 94.805 100.09 ;
      RECT 0 99.95 94.875 100.02 ;
      RECT 0 99.88 94.945 99.95 ;
      RECT 0 99.81 95.015 99.88 ;
      RECT 0 99.74 95.085 99.81 ;
      RECT 0 99.67 95.155 99.74 ;
      RECT 0 99.6 95.225 99.67 ;
      RECT 0 99.53 95.295 99.6 ;
      RECT 0 99.46 95.365 99.53 ;
      RECT 0 99.39 95.435 99.46 ;
      RECT 0 99.32 95.505 99.39 ;
      RECT 0 99.25 95.575 99.32 ;
      RECT 0 99.18 95.645 99.25 ;
      RECT 0 99.11 95.715 99.18 ;
      RECT 0 99.04 95.785 99.11 ;
      RECT 0 98.97 95.855 99.04 ;
      RECT 0 98.9 95.925 98.97 ;
      RECT 0 98.83 95.995 98.9 ;
      RECT 0 98.76 96.065 98.83 ;
      RECT 0 98.69 96.135 98.76 ;
      RECT 0 98.62 96.205 98.69 ;
      RECT 0 98.55 96.275 98.62 ;
      RECT 0 98.48 96.345 98.55 ;
      RECT 0 98.41 96.415 98.48 ;
      RECT 0 98.34 96.485 98.41 ;
      RECT 0 98.27 96.555 98.34 ;
      RECT 0 98.2 96.625 98.27 ;
      RECT 0 98.13 96.695 98.2 ;
      RECT 0 98.06 96.765 98.13 ;
      RECT 0 97.99 96.835 98.06 ;
      RECT 0 97.92 96.905 97.99 ;
      RECT 0 97.85 96.975 97.92 ;
      RECT 0 97.78 97.045 97.85 ;
      RECT 0 97.71 97.115 97.78 ;
      RECT 0 97.64 97.185 97.71 ;
      RECT 0 97.57 97.255 97.64 ;
      RECT 0 97.5 97.325 97.57 ;
      RECT 0 97.43 97.395 97.5 ;
      RECT 0 97.36 97.465 97.43 ;
      RECT 0 97.29 97.535 97.36 ;
      RECT 0 97.22 97.605 97.29 ;
      RECT 0 97.15 97.675 97.22 ;
      RECT 0 97.08 97.745 97.15 ;
      RECT 0 97.01 97.815 97.08 ;
      RECT 0 96.94 97.885 97.01 ;
      RECT 0 96.87 97.955 96.94 ;
      RECT 0 96.8 98.025 96.87 ;
      RECT 0 96.73 98.095 96.8 ;
      RECT 0 96.66 98.165 96.73 ;
      RECT 0 96.59 98.235 96.66 ;
      RECT 0 96.52 98.305 96.59 ;
      RECT 0 96.45 98.375 96.52 ;
      RECT 0 96.38 98.445 96.45 ;
      RECT 0 96.31 98.515 96.38 ;
      RECT 0 96.24 98.585 96.31 ;
      RECT 0 96.17 98.655 96.24 ;
      RECT 0 96.1 98.725 96.17 ;
      RECT 0 96.03 98.795 96.1 ;
      RECT 0 95.96 98.865 96.03 ;
      RECT 0 95.89 98.935 95.96 ;
      RECT 0 95.82 99.005 95.89 ;
      RECT 0 95.75 99.075 95.82 ;
      RECT 0 95.68 99.145 95.75 ;
      RECT 0 95.61 99.215 95.68 ;
      RECT 0 95.54 99.285 95.61 ;
      RECT 0 95.47 99.355 95.54 ;
      RECT 0 95.4 99.425 95.47 ;
      RECT 0 95.33 99.495 95.4 ;
      RECT 0 95.26 99.565 95.33 ;
      RECT 0 95.19 99.635 95.26 ;
      RECT 0 95.12 99.705 95.19 ;
      RECT 0 95.05 99.775 95.12 ;
      RECT 0 94.98 99.845 95.05 ;
      RECT 0 94.91 99.915 94.98 ;
      RECT 0 94.84 99.985 94.91 ;
      RECT 0 94.77 100.055 94.84 ;
      RECT 0 94.7 100.125 94.77 ;
      RECT 0 94.63 100.195 94.7 ;
      RECT 0 94.56 100.265 94.63 ;
      RECT 0 94.49 100.335 94.56 ;
      RECT 0 94.42 100.405 94.49 ;
      RECT 0 111.715 92.025 111.785 ;
      RECT 0 111.785 92.095 111.855 ;
      RECT 0 111.855 92.165 111.925 ;
      RECT 0 111.925 92.235 111.995 ;
      RECT 0 111.995 92.305 112.04 ;
      RECT 110.375 45.705 121.175 45.775 ;
      RECT 110.305 45.775 121.175 45.845 ;
      RECT 110.235 45.845 121.175 45.915 ;
      RECT 110.165 45.915 121.175 45.985 ;
      RECT 110.095 45.985 121.175 46.055 ;
      RECT 110.025 46.055 121.175 46.075 ;
      RECT 110.365 36.185 121.175 36.195 ;
      RECT 110.375 36.195 121.175 36.205 ;
      RECT 0 56.68 108.29 56.75 ;
      RECT 0 56.75 108.36 56.82 ;
      RECT 0 56.82 108.43 56.89 ;
      RECT 0 56.89 108.5 56.96 ;
      RECT 0 56.96 108.57 57.03 ;
      RECT 0 57.03 108.64 57.1 ;
      RECT 0 57.1 108.71 57.17 ;
      RECT 0 57.17 108.78 57.24 ;
      RECT 0 57.24 108.85 57.31 ;
      RECT 283.015 2.025 302.63 2.095 ;
      RECT 282.945 2.095 302.63 2.165 ;
      RECT 282.875 2.165 302.63 2.18 ;
      RECT 280.975 74.765 447.625 74.835 ;
      RECT 281.045 74.835 447.625 74.905 ;
      RECT 281.115 74.905 447.625 74.975 ;
      RECT 281.185 74.975 447.625 75.045 ;
      RECT 281.255 75.045 447.625 75.115 ;
      RECT 281.325 75.115 447.625 75.185 ;
      RECT 281.395 75.185 447.625 75.255 ;
      RECT 281.465 75.255 447.625 75.325 ;
      RECT 281.535 75.325 447.625 75.395 ;
      RECT 281.605 75.395 447.625 75.465 ;
      RECT 281.675 75.465 447.625 75.535 ;
      RECT 281.745 75.535 447.625 75.605 ;
      RECT 281.815 75.605 447.625 75.675 ;
      RECT 281.885 75.675 447.625 75.745 ;
      RECT 281.955 75.745 447.625 75.815 ;
      RECT 282.025 75.815 447.625 75.885 ;
      RECT 282.095 75.885 447.625 75.955 ;
      RECT 282.165 75.955 447.625 76.025 ;
      RECT 282.235 76.025 447.625 76.095 ;
      RECT 282.305 76.095 447.625 76.165 ;
      RECT 282.375 76.165 447.625 76.235 ;
      RECT 282.445 76.235 447.625 76.305 ;
      RECT 282.515 76.305 447.625 76.375 ;
      RECT 282.535 76.375 447.625 76.395 ;
      RECT 282.605 87.425 446.805 87.495 ;
      RECT 282.675 87.495 446.805 87.565 ;
      RECT 282.745 87.565 446.805 87.635 ;
      RECT 282.815 87.635 446.805 87.705 ;
      RECT 282.885 87.705 446.805 87.775 ;
      RECT 282.955 87.775 446.805 87.845 ;
      RECT 283.025 87.845 446.805 87.915 ;
      RECT 283.095 87.915 446.805 87.985 ;
      RECT 283.165 87.985 446.805 88.055 ;
      RECT 283.235 88.055 446.805 88.125 ;
      RECT 283.305 88.125 446.805 88.195 ;
      RECT 283.375 88.195 446.805 88.265 ;
      RECT 283.445 88.265 446.805 88.335 ;
      RECT 283.515 88.335 446.805 88.405 ;
      RECT 283.585 88.405 446.805 88.475 ;
      RECT 283.655 88.475 446.805 88.545 ;
      RECT 283.725 88.545 446.805 88.615 ;
      RECT 283.795 88.615 446.805 88.685 ;
      RECT 283.865 88.685 446.805 88.755 ;
      RECT 283.935 88.755 446.805 88.825 ;
      RECT 284.005 88.825 446.805 88.895 ;
      RECT 284.075 88.895 446.805 88.965 ;
      RECT 284.145 88.965 446.805 89.035 ;
      RECT 284.215 89.035 446.805 89.105 ;
      RECT 284.285 89.105 446.805 89.175 ;
      RECT 284.355 89.175 446.805 89.245 ;
      RECT 284.425 89.245 446.805 89.315 ;
      RECT 284.475 89.315 446.805 89.365 ;
      RECT 282.535 84.9 447.555 84.97 ;
      RECT 282.535 84.97 447.485 85.04 ;
      RECT 282.535 85.04 447.415 85.11 ;
      RECT 282.535 85.11 447.345 85.18 ;
      RECT 282.535 85.18 447.275 85.25 ;
      RECT 282.535 85.25 447.205 85.32 ;
      RECT 282.535 85.32 447.135 85.39 ;
      RECT 282.535 85.39 447.065 85.46 ;
      RECT 282.535 85.46 446.995 85.53 ;
      RECT 282.535 85.53 446.925 85.6 ;
      RECT 282.535 85.6 446.855 85.67 ;
      RECT 282.535 85.67 446.805 85.72 ;
      RECT 284.545 94.05 446.805 94.12 ;
      RECT 284.615 94.12 446.805 94.19 ;
      RECT 284.685 94.19 446.805 94.26 ;
      RECT 284.755 94.26 446.805 94.33 ;
      RECT 284.825 94.33 446.805 94.4 ;
      RECT 284.845 94.4 446.805 94.42 ;
      RECT 452.065 240.105 480 240.135 ;
      RECT 452.135 240.035 480 240.105 ;
      RECT 452.205 239.965 480 240.035 ;
      RECT 452.275 239.895 480 239.965 ;
      RECT 452.345 239.825 480 239.895 ;
      RECT 452.415 239.755 480 239.825 ;
      RECT 452.485 239.685 480 239.755 ;
      RECT 452.555 239.615 480 239.685 ;
      RECT 452.625 239.545 480 239.615 ;
      RECT 452.695 239.475 480 239.545 ;
      RECT 452.765 239.405 480 239.475 ;
      RECT 452.835 239.335 480 239.405 ;
      RECT 452.905 239.265 480 239.335 ;
      RECT 452.975 239.195 480 239.265 ;
      RECT 453.045 239.125 480 239.195 ;
      RECT 453.115 239.055 480 239.125 ;
      RECT 453.185 238.985 480 239.055 ;
      RECT 453.255 238.915 480 238.985 ;
      RECT 453.325 238.845 480 238.915 ;
      RECT 453.395 238.775 480 238.845 ;
      RECT 453.465 238.705 480 238.775 ;
      RECT 453.535 238.635 480 238.705 ;
      RECT 453.605 238.565 480 238.635 ;
      RECT 453.675 238.495 480 238.565 ;
      RECT 453.745 238.425 480 238.495 ;
      RECT 453.815 238.355 480 238.425 ;
      RECT 453.885 238.285 480 238.355 ;
      RECT 453.955 238.215 480 238.285 ;
      RECT 454.025 238.145 480 238.215 ;
      RECT 454.095 238.075 480 238.145 ;
      RECT 454.165 238.005 480 238.075 ;
      RECT 454.235 237.935 480 238.005 ;
      RECT 454.305 237.865 480 237.935 ;
      RECT 454.375 237.795 480 237.865 ;
      RECT 454.445 237.725 480 237.795 ;
      RECT 0 102.82 92.025 102.87 ;
      RECT 0 102.75 92.075 102.82 ;
      RECT 0 102.68 92.145 102.75 ;
      RECT 0 102.61 92.215 102.68 ;
      RECT 0 102.54 92.285 102.61 ;
      RECT 0 102.47 92.355 102.54 ;
      RECT 0 102.4 92.425 102.47 ;
      RECT 0 102.33 92.495 102.4 ;
      RECT 0 102.26 92.565 102.33 ;
      RECT 0 102.19 92.635 102.26 ;
      RECT 0 102.12 92.705 102.19 ;
      RECT 0 102.05 92.775 102.12 ;
      RECT 0 101.98 92.845 102.05 ;
      RECT 0 101.91 92.915 101.98 ;
      RECT 0 101.84 92.985 101.91 ;
      RECT 0 101.77 93.055 101.84 ;
      RECT 0 101.7 93.125 101.77 ;
      RECT 108.73 76.295 281.275 76.365 ;
      RECT 108.66 76.365 281.345 76.435 ;
      RECT 108.59 76.435 281.415 76.505 ;
      RECT 108.52 76.505 281.485 76.575 ;
      RECT 108.45 76.575 281.555 76.645 ;
      RECT 108.38 76.645 281.625 76.715 ;
      RECT 108.31 76.715 281.695 76.735 ;
      RECT 243.14 26.695 253.89 26.765 ;
      RECT 243.21 26.765 253.89 26.835 ;
      RECT 243.28 26.835 253.89 26.905 ;
      RECT 243.35 26.905 253.89 26.975 ;
      RECT 243.42 26.975 253.89 27.045 ;
      RECT 243.49 27.045 253.89 27.115 ;
      RECT 243.56 27.115 253.89 27.185 ;
      RECT 243.63 27.185 253.89 27.255 ;
      RECT 243.7 27.255 253.89 27.325 ;
      RECT 243.77 27.325 253.89 27.395 ;
      RECT 243.84 27.395 253.89 27.465 ;
      RECT 243.91 27.465 253.89 27.535 ;
      RECT 243.98 27.535 253.89 27.605 ;
      RECT 244.05 27.605 253.89 27.675 ;
      RECT 244.12 27.675 253.89 27.745 ;
      RECT 244.19 27.745 253.89 27.815 ;
      RECT 244.26 27.815 253.89 27.885 ;
      RECT 244.33 27.885 253.89 27.955 ;
      RECT 244.4 27.955 253.89 28.025 ;
      RECT 244.47 28.025 253.89 28.095 ;
      RECT 244.54 28.095 253.89 28.165 ;
      RECT 244.61 28.165 253.89 28.235 ;
      RECT 244.65 28.235 253.89 28.275 ;
      RECT 255.11 10.29 261.34 10.36 ;
      RECT 255.11 10.36 261.41 10.43 ;
      RECT 255.11 10.43 261.48 10.5 ;
      RECT 255.11 10.5 261.55 10.57 ;
      RECT 255.11 10.57 261.62 10.64 ;
      RECT 255.11 10.64 261.69 10.71 ;
      RECT 255.11 10.71 261.76 10.78 ;
      RECT 255.11 10.78 261.83 10.85 ;
      RECT 255.11 10.85 261.9 10.92 ;
      RECT 255.11 10.92 261.97 10.99 ;
      RECT 255.11 10.99 262.04 11.06 ;
      RECT 255.11 11.06 262.11 11.13 ;
      RECT 255.11 11.13 262.18 11.155 ;
      RECT 255.18 28.725 261.605 28.795 ;
      RECT 255.25 28.795 261.605 28.865 ;
      RECT 255.32 28.865 261.605 28.935 ;
      RECT 255.39 28.935 261.605 29.005 ;
      RECT 255.46 29.005 261.605 29.075 ;
      RECT 255.53 29.075 261.605 29.145 ;
      RECT 255.6 29.145 261.605 29.215 ;
      RECT 255.64 29.215 261.605 29.255 ;
      RECT 255.11 23.55 262.135 23.62 ;
      RECT 255.11 23.62 262.065 23.69 ;
      RECT 255.11 23.69 261.995 23.76 ;
      RECT 255.11 23.76 261.925 23.83 ;
      RECT 255.11 23.83 261.855 23.9 ;
      RECT 255.11 23.9 261.785 23.97 ;
      RECT 255.11 23.97 261.715 24.04 ;
      RECT 255.11 24.04 261.645 24.11 ;
      RECT 255.11 24.11 261.605 24.15 ;
      RECT 255.71 29.255 261.605 29.325 ;
      RECT 255.78 29.325 261.605 29.395 ;
      RECT 255.85 29.395 261.605 29.465 ;
      RECT 255.92 29.465 261.605 29.535 ;
      RECT 255.99 29.535 261.605 29.605 ;
      RECT 256.06 29.605 261.605 29.675 ;
      RECT 256.09 29.675 261.605 29.705 ;
      RECT 262.23 9.95 268.01 10.02 ;
      RECT 262.3 10.02 268.01 10.09 ;
      RECT 262.37 10.09 268.01 10.16 ;
      RECT 262.44 10.16 268.01 10.23 ;
      RECT 262.51 10.23 268.01 10.3 ;
      RECT 262.58 10.3 268.01 10.37 ;
      RECT 262.65 10.37 268.01 10.44 ;
      RECT 262.72 10.44 268.01 10.51 ;
      RECT 262.79 10.51 268.01 10.58 ;
      RECT 262.86 10.58 268.01 10.65 ;
      RECT 262.93 10.65 268.01 10.72 ;
      RECT 263.0 10.72 268.01 10.79 ;
      RECT 263.025 10.79 268.01 10.815 ;
      RECT 263.025 23.89 268.01 23.96 ;
      RECT 262.955 23.96 268.01 24.03 ;
      RECT 262.885 24.03 268.01 24.1 ;
      RECT 262.815 24.1 268.01 24.17 ;
      RECT 262.745 24.17 268.01 24.24 ;
      RECT 262.675 24.24 268.01 24.31 ;
      RECT 262.605 24.31 268.01 24.38 ;
      RECT 262.535 24.38 268.01 24.45 ;
      RECT 262.465 24.45 268.01 24.49 ;
      RECT 240.48 56.34 280.825 56.41 ;
      RECT 240.48 56.41 280.755 56.48 ;
      RECT 240.48 56.48 280.685 56.55 ;
      RECT 240.48 56.55 280.615 56.62 ;
      RECT 240.48 56.62 280.545 56.69 ;
      RECT 240.48 56.69 280.475 56.76 ;
      RECT 240.48 56.76 280.405 56.83 ;
      RECT 240.48 56.83 280.335 56.9 ;
      RECT 240.48 56.9 280.265 56.97 ;
      RECT 240.48 56.97 280.195 57.04 ;
      RECT 240.48 57.04 280.125 57.11 ;
      RECT 240.48 57.11 280.085 57.15 ;
      RECT 268.83 17.58 279.375 17.65 ;
      RECT 268.83 17.65 279.445 17.72 ;
      RECT 268.83 17.72 279.515 17.79 ;
      RECT 268.83 17.79 279.585 17.855 ;
      RECT 265.425 46.79 280 46.86 ;
      RECT 265.355 46.86 280.07 46.93 ;
      RECT 265.285 46.93 280.14 47 ;
      RECT 265.215 47 280.21 47.035 ;
      RECT 265.655 46.56 280 46.63 ;
      RECT 265.585 46.63 280 46.7 ;
      RECT 265.515 46.7 280 46.77 ;
      RECT 265.445 46.77 280 46.79 ;
      RECT 283.575 1.465 302.63 1.535 ;
      RECT 283.505 1.535 302.63 1.605 ;
      RECT 283.435 1.605 302.63 1.675 ;
      RECT 283.365 1.675 302.63 1.745 ;
      RECT 283.295 1.745 302.63 1.815 ;
      RECT 283.225 1.815 302.63 1.885 ;
      RECT 283.155 1.885 302.63 1.955 ;
      RECT 283.085 1.955 302.63 2.025 ;
      RECT 121.995 10.37 127.355 10.44 ;
      RECT 121.995 10.44 127.285 10.51 ;
      RECT 121.995 10.51 127.215 10.58 ;
      RECT 121.995 10.58 127.145 10.65 ;
      RECT 121.995 10.65 127.075 10.72 ;
      RECT 121.995 10.72 127.005 10.79 ;
      RECT 121.995 10.79 126.98 10.815 ;
      RECT 124.76 45.74 145.355 45.81 ;
      RECT 124.83 45.81 145.355 45.88 ;
      RECT 124.9 45.88 145.355 45.95 ;
      RECT 124.97 45.95 145.355 46.02 ;
      RECT 125.04 46.02 145.355 46.09 ;
      RECT 125.11 46.09 145.355 46.16 ;
      RECT 125.18 46.16 145.355 46.23 ;
      RECT 125.25 46.23 145.355 46.3 ;
      RECT 125.32 46.3 145.355 46.37 ;
      RECT 125.39 46.37 145.355 46.44 ;
      RECT 125.46 46.44 145.355 46.51 ;
      RECT 125.53 46.51 145.355 46.58 ;
      RECT 125.6 46.58 145.355 46.65 ;
      RECT 125.67 46.65 145.355 46.72 ;
      RECT 125.74 46.72 145.355 46.79 ;
      RECT 125.81 46.79 145.355 46.86 ;
      RECT 125.88 46.86 145.355 46.93 ;
      RECT 125.95 46.93 145.355 47 ;
      RECT 126.02 47 145.355 47.07 ;
      RECT 126.09 47.07 145.355 47.14 ;
      RECT 126.16 47.14 145.355 47.21 ;
      RECT 126.195 47.21 145.355 47.245 ;
      RECT 127.87 23.55 134.895 23.62 ;
      RECT 127.94 23.62 134.895 23.69 ;
      RECT 128.01 23.69 134.895 23.76 ;
      RECT 128.08 23.76 134.895 23.83 ;
      RECT 128.15 23.83 134.895 23.9 ;
      RECT 128.22 23.9 134.895 23.97 ;
      RECT 128.29 23.97 134.895 24.04 ;
      RECT 128.36 24.04 134.895 24.11 ;
      RECT 128.4 24.11 134.895 24.15 ;
      RECT 128.4 29.255 134.295 29.325 ;
      RECT 128.4 29.325 134.225 29.395 ;
      RECT 128.4 29.395 134.155 29.465 ;
      RECT 128.4 29.465 134.085 29.535 ;
      RECT 128.4 29.535 134.015 29.605 ;
      RECT 128.4 29.605 133.945 29.675 ;
      RECT 128.4 29.675 133.915 29.705 ;
      RECT 128.4 28.725 134.825 28.795 ;
      RECT 128.4 28.795 134.755 28.865 ;
      RECT 128.4 28.865 134.685 28.935 ;
      RECT 128.4 28.935 134.615 29.005 ;
      RECT 128.4 29.005 134.545 29.075 ;
      RECT 128.4 29.075 134.475 29.145 ;
      RECT 128.4 29.145 134.405 29.215 ;
      RECT 128.4 29.215 134.365 29.255 ;
      RECT 128.665 10.29 134.895 10.36 ;
      RECT 128.595 10.36 134.895 10.43 ;
      RECT 128.525 10.43 134.895 10.5 ;
      RECT 128.455 10.5 134.895 10.57 ;
      RECT 128.385 10.57 134.895 10.64 ;
      RECT 128.315 10.64 134.895 10.71 ;
      RECT 128.245 10.71 134.895 10.78 ;
      RECT 128.175 10.78 134.895 10.85 ;
      RECT 128.105 10.85 134.895 10.92 ;
      RECT 128.035 10.92 134.895 10.99 ;
      RECT 127.965 10.99 134.895 11.06 ;
      RECT 127.895 11.06 134.895 11.13 ;
      RECT 127.825 11.13 134.895 11.155 ;
      RECT 136.115 26.695 146.865 26.765 ;
      RECT 136.115 26.765 146.795 26.835 ;
      RECT 136.115 26.835 146.725 26.905 ;
      RECT 136.115 26.905 146.655 26.975 ;
      RECT 136.115 26.975 146.585 27.045 ;
      RECT 136.115 27.045 146.515 27.115 ;
      RECT 136.115 27.115 146.445 27.185 ;
      RECT 136.115 27.185 146.375 27.255 ;
      RECT 136.115 27.255 146.305 27.325 ;
      RECT 136.115 27.325 146.235 27.395 ;
      RECT 136.115 27.395 146.165 27.465 ;
      RECT 136.115 27.465 146.095 27.535 ;
      RECT 136.115 27.535 146.025 27.605 ;
      RECT 136.115 27.605 145.955 27.675 ;
      RECT 136.115 27.675 145.885 27.745 ;
      RECT 136.115 27.745 145.815 27.815 ;
      RECT 136.115 27.815 145.745 27.885 ;
      RECT 136.115 27.885 145.675 27.955 ;
      RECT 136.115 27.955 145.605 28.025 ;
      RECT 136.115 28.025 145.535 28.095 ;
      RECT 136.115 28.095 145.465 28.165 ;
      RECT 136.115 28.165 145.395 28.235 ;
      RECT 136.115 28.235 145.355 28.275 ;
      RECT 109.18 56.34 149.525 56.41 ;
      RECT 109.25 56.41 149.525 56.48 ;
      RECT 109.32 56.48 149.525 56.55 ;
      RECT 109.39 56.55 149.525 56.62 ;
      RECT 109.46 56.62 149.525 56.69 ;
      RECT 109.53 56.69 149.525 56.76 ;
      RECT 109.6 56.76 149.525 56.83 ;
      RECT 109.67 56.83 149.525 56.9 ;
      RECT 109.74 56.9 149.525 56.97 ;
      RECT 109.81 56.97 149.525 57.04 ;
      RECT 109.88 57.04 149.525 57.11 ;
      RECT 109.92 57.11 149.525 57.15 ;
      RECT 150.345 42.21 153.53 42.215 ;
      RECT 150.345 42.215 153.535 42.22 ;
      RECT 154.355 41.87 235.65 41.875 ;
      RECT 154.36 41.875 235.645 41.88 ;
      RECT 236.475 42.21 239.66 42.215 ;
      RECT 236.47 42.215 239.66 42.22 ;
      RECT 109.92 75.105 280.085 75.175 ;
      RECT 109.85 75.175 280.155 75.245 ;
      RECT 109.78 75.245 280.225 75.315 ;
      RECT 109.71 75.315 280.295 75.385 ;
      RECT 109.64 75.385 280.365 75.455 ;
      RECT 109.57 75.455 280.435 75.525 ;
      RECT 109.5 75.525 280.505 75.595 ;
      RECT 109.43 75.595 280.575 75.665 ;
      RECT 109.36 75.665 280.645 75.735 ;
      RECT 109.29 75.735 280.715 75.805 ;
      RECT 109.22 75.805 280.785 75.875 ;
      RECT 109.15 75.875 280.855 75.945 ;
      RECT 109.08 75.945 280.925 76.015 ;
      RECT 109.01 76.015 280.995 76.085 ;
      RECT 108.94 76.085 281.065 76.155 ;
      RECT 108.87 76.155 281.135 76.225 ;
      RECT 108.8 76.225 281.205 76.295 ;
      RECT 0 89.245 105.58 89.315 ;
      RECT 0 89.315 105.53 89.365 ;
      RECT 0 74.765 109.03 74.835 ;
      RECT 0 74.835 108.96 74.905 ;
      RECT 0 74.905 108.89 74.975 ;
      RECT 0 74.975 108.82 75.045 ;
      RECT 0 75.045 108.75 75.115 ;
      RECT 0 75.115 108.68 75.185 ;
      RECT 0 75.185 108.61 75.255 ;
      RECT 0 75.255 108.54 75.325 ;
      RECT 0 75.325 108.47 75.395 ;
      RECT 0 75.395 108.4 75.465 ;
      RECT 0 75.465 108.33 75.535 ;
      RECT 0 75.535 108.26 75.605 ;
      RECT 0 75.605 108.19 75.675 ;
      RECT 0 75.675 108.12 75.745 ;
      RECT 0 75.745 108.05 75.815 ;
      RECT 0 75.815 107.98 75.885 ;
      RECT 0 75.885 107.91 75.955 ;
      RECT 0 75.955 107.84 76.025 ;
      RECT 0 76.025 107.77 76.095 ;
      RECT 0 76.095 107.7 76.165 ;
      RECT 0 76.165 107.63 76.235 ;
      RECT 0 76.235 107.56 76.305 ;
      RECT 0 76.305 107.49 76.375 ;
      RECT 0 76.375 107.47 76.395 ;
      RECT 87.375 1.465 106.43 1.535 ;
      RECT 87.375 1.535 106.5 1.605 ;
      RECT 87.375 1.605 106.57 1.675 ;
      RECT 87.375 1.675 106.64 1.745 ;
      RECT 87.375 1.745 106.71 1.815 ;
      RECT 87.375 1.815 106.78 1.885 ;
      RECT 87.375 1.885 106.85 1.955 ;
      RECT 87.375 1.955 106.92 2.025 ;
      RECT 87.375 2.025 106.99 2.095 ;
      RECT 87.375 2.095 107.06 2.165 ;
      RECT 87.375 2.165 107.13 2.18 ;
      RECT 106.375 94.365 283.63 94.435 ;
      RECT 106.305 94.435 283.7 94.505 ;
      RECT 106.235 94.505 283.77 94.575 ;
      RECT 106.165 94.575 283.84 94.645 ;
      RECT 106.095 94.645 283.91 94.715 ;
      RECT 106.025 94.715 283.98 94.785 ;
      RECT 105.955 94.785 284.05 94.855 ;
      RECT 105.885 94.855 284.12 94.925 ;
      RECT 105.815 94.925 284.19 94.995 ;
      RECT 105.745 94.995 284.26 95.065 ;
      RECT 105.675 95.065 284.33 95.135 ;
      RECT 105.605 95.135 284.4 95.205 ;
      RECT 105.535 95.205 284.47 95.24 ;
      RECT 108.29 87.765 281.715 87.835 ;
      RECT 108.22 87.835 281.785 87.905 ;
      RECT 108.15 87.905 281.855 87.975 ;
      RECT 108.08 87.975 281.925 88.045 ;
      RECT 108.01 88.045 281.995 88.115 ;
      RECT 107.94 88.115 282.065 88.185 ;
      RECT 107.87 88.185 282.135 88.255 ;
      RECT 107.8 88.255 282.205 88.325 ;
      RECT 107.73 88.325 282.275 88.395 ;
      RECT 107.66 88.395 282.345 88.465 ;
      RECT 107.59 88.465 282.415 88.535 ;
      RECT 107.52 88.535 282.485 88.605 ;
      RECT 107.45 88.605 282.555 88.675 ;
      RECT 107.38 88.675 282.625 88.745 ;
      RECT 107.31 88.745 282.695 88.815 ;
      RECT 107.24 88.815 282.765 88.885 ;
      RECT 107.17 88.885 282.835 88.955 ;
      RECT 107.1 88.955 282.905 89.025 ;
      RECT 107.03 89.025 282.975 89.095 ;
      RECT 106.96 89.095 283.045 89.165 ;
      RECT 106.89 89.165 283.115 89.235 ;
      RECT 106.82 89.235 283.185 89.305 ;
      RECT 106.75 89.305 283.255 89.375 ;
      RECT 106.68 89.375 283.325 89.445 ;
      RECT 106.61 89.445 283.395 89.515 ;
      RECT 106.54 89.515 283.465 89.585 ;
      RECT 106.47 89.585 283.535 89.655 ;
      RECT 106.4 89.655 283.605 89.68 ;
      RECT 109.21 47.585 125.375 47.635 ;
      RECT 109.16 47.635 125.375 47.685 ;
      RECT 109.11 48.55 125.305 48.62 ;
      RECT 109.11 48.62 125.235 48.69 ;
      RECT 109.11 48.69 125.165 48.76 ;
      RECT 109.11 48.76 125.095 48.83 ;
      RECT 109.11 48.83 125.07 48.855 ;
      RECT 110.005 46.79 124.58 46.86 ;
      RECT 109.935 46.86 124.65 46.93 ;
      RECT 109.865 46.93 124.72 47 ;
      RECT 109.795 47 124.79 47.07 ;
      RECT 109.725 47.07 124.86 47.14 ;
      RECT 109.655 47.14 124.93 47.21 ;
      RECT 109.585 47.21 125.0 47.28 ;
      RECT 109.515 47.28 125.07 47.35 ;
      RECT 109.445 47.35 125.14 47.42 ;
      RECT 109.375 47.42 125.21 47.49 ;
      RECT 109.305 47.49 125.28 47.56 ;
      RECT 109.235 47.56 125.35 47.585 ;
      RECT 110.005 46.56 124.35 46.63 ;
      RECT 110.005 46.63 124.42 46.7 ;
      RECT 110.005 46.7 124.49 46.77 ;
      RECT 110.005 46.77 124.56 46.79 ;
      RECT 110.63 17.58 121.175 17.65 ;
      RECT 110.56 17.65 121.175 17.72 ;
      RECT 110.49 17.72 121.175 17.79 ;
      RECT 110.42 17.79 121.175 17.855 ;
      RECT 121.995 23.89 126.98 23.96 ;
      RECT 121.995 23.96 127.05 24.03 ;
      RECT 121.995 24.03 127.12 24.1 ;
      RECT 121.995 24.1 127.19 24.17 ;
      RECT 121.995 24.17 127.26 24.24 ;
      RECT 121.995 24.24 127.33 24.31 ;
      RECT 121.995 24.31 127.4 24.38 ;
      RECT 121.995 24.38 127.47 24.45 ;
      RECT 121.995 24.45 127.54 24.49 ;
      RECT 121.995 9.95 127.775 10.02 ;
      RECT 121.995 10.02 127.705 10.09 ;
      RECT 121.995 10.09 127.635 10.16 ;
      RECT 121.995 10.16 127.565 10.23 ;
      RECT 121.995 10.23 127.495 10.3 ;
      RECT 121.995 10.3 127.425 10.37 ;
      RECT 292.05 96.87 446.805 96.94 ;
      RECT 291.98 96.8 446.805 96.87 ;
      RECT 291.91 96.73 446.805 96.8 ;
      RECT 291.84 96.66 446.805 96.73 ;
      RECT 291.77 96.59 446.805 96.66 ;
      RECT 291.7 96.52 446.805 96.59 ;
      RECT 291.63 96.45 446.805 96.52 ;
      RECT 291.56 96.38 446.805 96.45 ;
      RECT 291.49 96.31 446.805 96.38 ;
      RECT 291.42 96.24 446.805 96.31 ;
      RECT 291.35 96.17 446.805 96.24 ;
      RECT 291.28 96.1 446.805 96.17 ;
      RECT 291.21 96.03 446.805 96.1 ;
      RECT 291.14 95.96 446.805 96.03 ;
      RECT 291.07 95.89 446.805 95.96 ;
      RECT 291.0 95.82 446.805 95.89 ;
      RECT 290.93 95.75 446.805 95.82 ;
      RECT 290.86 95.68 446.805 95.75 ;
      RECT 290.79 95.61 446.805 95.68 ;
      RECT 290.72 95.54 446.805 95.61 ;
      RECT 290.65 95.47 446.805 95.54 ;
      RECT 290.58 95.4 446.805 95.47 ;
      RECT 290.51 95.33 446.805 95.4 ;
      RECT 290.44 95.26 446.805 95.33 ;
      RECT 290.37 95.19 446.805 95.26 ;
      RECT 290.3 95.12 446.805 95.19 ;
      RECT 290.23 95.05 446.805 95.12 ;
      RECT 290.16 94.98 446.805 95.05 ;
      RECT 290.09 94.91 446.805 94.98 ;
      RECT 290.02 94.84 446.805 94.91 ;
      RECT 289.95 94.77 446.805 94.84 ;
      RECT 289.88 94.7 446.805 94.77 ;
      RECT 289.81 94.63 446.805 94.7 ;
      RECT 289.74 94.56 446.805 94.63 ;
      RECT 289.67 94.49 446.805 94.56 ;
      RECT 289.6 94.42 446.805 94.49 ;
      RECT 297.655 112.04 446.805 112.11 ;
      RECT 297.585 112.11 446.805 112.18 ;
      RECT 297.515 112.18 446.805 112.25 ;
      RECT 297.445 112.25 446.805 112.32 ;
      RECT 297.375 112.32 446.805 112.39 ;
      RECT 297.305 112.39 446.805 112.42 ;
      RECT 297.98 111.715 446.805 111.785 ;
      RECT 297.91 111.785 446.805 111.855 ;
      RECT 297.84 111.855 446.805 111.925 ;
      RECT 297.77 111.925 446.805 111.995 ;
      RECT 297.7 111.995 446.805 112.04 ;
      RECT 452.065 240.105 480 240.135 ;
      RECT 452.135 240.035 480 240.105 ;
      RECT 452.205 239.965 480 240.035 ;
      RECT 452.275 239.895 480 239.965 ;
      RECT 452.345 239.825 480 239.895 ;
      RECT 452.415 239.755 480 239.825 ;
      RECT 452.485 239.685 480 239.755 ;
      RECT 452.555 239.615 480 239.685 ;
      RECT 452.625 239.545 480 239.615 ;
      RECT 452.695 239.475 480 239.545 ;
      RECT 452.765 239.405 480 239.475 ;
      RECT 452.835 239.335 480 239.405 ;
      RECT 452.905 239.265 480 239.335 ;
      RECT 452.975 239.195 480 239.265 ;
      RECT 453.045 239.125 480 239.195 ;
      RECT 453.115 239.055 480 239.125 ;
      RECT 453.185 238.985 480 239.055 ;
      RECT 453.255 238.915 480 238.985 ;
      RECT 453.325 238.845 480 238.915 ;
      RECT 453.395 238.775 480 238.845 ;
      RECT 453.465 238.705 480 238.775 ;
      RECT 453.535 238.635 480 238.705 ;
      RECT 453.605 238.565 480 238.635 ;
      RECT 453.675 238.495 480 238.565 ;
      RECT 453.745 238.425 480 238.495 ;
      RECT 453.815 238.355 480 238.425 ;
      RECT 453.885 238.285 480 238.355 ;
      RECT 453.955 238.215 480 238.285 ;
      RECT 454.025 238.145 480 238.215 ;
      RECT 454.095 238.075 480 238.145 ;
      RECT 454.165 238.005 480 238.075 ;
      RECT 454.235 237.935 480 238.005 ;
      RECT 454.305 237.865 480 237.935 ;
      RECT 454.375 237.795 480 237.865 ;
      RECT 454.445 237.725 480 237.795 ;
      RECT 264.71 47.585 280.795 47.63 ;
      RECT 264.67 47.63 280.84 47.675 ;
      RECT 264.635 47.675 280.885 47.68 ;
      RECT 265.18 47.035 280.245 47.105 ;
      RECT 265.12 47.105 280.315 47.175 ;
      RECT 265.06 47.175 280.385 47.245 ;
      RECT 265.0 47.245 280.455 47.315 ;
      RECT 264.94 47.315 280.525 47.385 ;
      RECT 264.88 47.385 280.595 47.455 ;
      RECT 264.82 47.455 280.665 47.525 ;
      RECT 264.76 47.525 280.735 47.585 ;
      RECT 0 94.05 105.46 94.12 ;
      RECT 0 94.12 105.39 94.19 ;
      RECT 0 94.19 105.32 94.26 ;
      RECT 0 94.26 105.25 94.33 ;
      RECT 0 94.33 105.18 94.4 ;
      RECT 0 94.4 105.16 94.42 ;
      RECT 0 87.425 107.4 87.495 ;
      RECT 0 87.495 107.33 87.565 ;
      RECT 0 87.565 107.26 87.635 ;
      RECT 0 87.635 107.19 87.705 ;
      RECT 0 87.705 107.12 87.775 ;
      RECT 0 87.775 107.05 87.845 ;
      RECT 0 87.845 106.98 87.915 ;
      RECT 0 87.915 106.91 87.985 ;
      RECT 0 87.985 106.84 88.055 ;
      RECT 0 88.055 106.77 88.125 ;
      RECT 0 88.125 106.7 88.195 ;
      RECT 0 88.195 106.63 88.265 ;
      RECT 0 88.265 106.56 88.335 ;
      RECT 0 88.335 106.49 88.405 ;
      RECT 0 88.405 106.42 88.475 ;
      RECT 0 88.475 106.35 88.545 ;
      RECT 0 88.545 106.28 88.615 ;
      RECT 0 88.615 106.21 88.685 ;
      RECT 0 88.685 106.14 88.755 ;
      RECT 0 88.755 106.07 88.825 ;
      RECT 0 88.825 106.0 88.895 ;
      RECT 0 88.895 105.93 88.965 ;
      RECT 0 88.965 105.86 89.035 ;
      RECT 0 89.035 105.79 89.105 ;
      RECT 0 89.105 105.72 89.175 ;
      RECT 0 89.175 105.65 89.245 ;
      RECT 283.725 88.545 446.805 88.615 ;
      RECT 283.795 88.615 446.805 88.685 ;
      RECT 283.865 88.685 446.805 88.755 ;
      RECT 283.935 88.755 446.805 88.825 ;
      RECT 284.005 88.825 446.805 88.895 ;
      RECT 284.075 88.895 446.805 88.965 ;
      RECT 284.145 88.965 446.805 89.035 ;
      RECT 284.215 89.035 446.805 89.105 ;
      RECT 284.285 89.105 446.805 89.175 ;
      RECT 284.355 89.175 446.805 89.245 ;
      RECT 284.425 89.245 446.805 89.315 ;
      RECT 284.475 89.315 446.805 89.365 ;
      RECT 282.535 84.9 447.555 84.97 ;
      RECT 282.535 84.97 447.485 85.04 ;
      RECT 282.535 85.04 447.415 85.11 ;
      RECT 282.535 85.11 447.345 85.18 ;
      RECT 282.535 85.18 447.275 85.25 ;
      RECT 282.535 85.25 447.205 85.32 ;
      RECT 282.535 85.32 447.135 85.39 ;
      RECT 282.535 85.39 447.065 85.46 ;
      RECT 282.535 85.46 446.995 85.53 ;
      RECT 282.535 85.53 446.925 85.6 ;
      RECT 282.535 85.6 446.855 85.67 ;
      RECT 282.535 85.67 446.805 85.72 ;
      RECT 283.575 1.465 302.63 1.535 ;
      RECT 283.505 1.535 302.63 1.605 ;
      RECT 283.435 1.605 302.63 1.675 ;
      RECT 283.365 1.675 302.63 1.745 ;
      RECT 283.295 1.745 302.63 1.815 ;
      RECT 283.225 1.815 302.63 1.885 ;
      RECT 283.155 1.885 302.63 1.955 ;
      RECT 283.085 1.955 302.63 2.025 ;
      RECT 283.015 2.025 302.63 2.095 ;
      RECT 282.945 2.095 302.63 2.165 ;
      RECT 282.875 2.165 302.63 2.18 ;
      RECT 284.545 94.05 446.805 94.12 ;
      RECT 284.615 94.12 446.805 94.19 ;
      RECT 284.685 94.19 446.805 94.26 ;
      RECT 284.755 94.26 446.805 94.33 ;
      RECT 284.825 94.33 446.805 94.4 ;
      RECT 284.845 94.4 446.805 94.42 ;
      RECT 297.98 102.82 446.805 102.87 ;
      RECT 297.93 102.75 446.805 102.82 ;
      RECT 297.86 102.68 446.805 102.75 ;
      RECT 297.79 102.61 446.805 102.68 ;
      RECT 297.72 102.54 446.805 102.61 ;
      RECT 297.65 102.47 446.805 102.54 ;
      RECT 297.58 102.4 446.805 102.47 ;
      RECT 297.51 102.33 446.805 102.4 ;
      RECT 297.44 102.26 446.805 102.33 ;
      RECT 297.37 102.19 446.805 102.26 ;
      RECT 297.3 102.12 446.805 102.19 ;
      RECT 297.23 102.05 446.805 102.12 ;
      RECT 297.16 101.98 446.805 102.05 ;
      RECT 297.09 101.91 446.805 101.98 ;
      RECT 297.02 101.84 446.805 101.91 ;
      RECT 296.95 101.77 446.805 101.84 ;
      RECT 296.88 101.7 446.805 101.77 ;
      RECT 296.81 101.63 446.805 101.7 ;
      RECT 296.74 101.56 446.805 101.63 ;
      RECT 296.67 101.49 446.805 101.56 ;
      RECT 296.6 101.42 446.805 101.49 ;
      RECT 296.53 101.35 446.805 101.42 ;
      RECT 296.46 101.28 446.805 101.35 ;
      RECT 296.39 101.21 446.805 101.28 ;
      RECT 296.32 101.14 446.805 101.21 ;
      RECT 296.25 101.07 446.805 101.14 ;
      RECT 296.18 101 446.805 101.07 ;
      RECT 296.11 100.93 446.805 101 ;
      RECT 296.04 100.86 446.805 100.93 ;
      RECT 295.97 100.79 446.805 100.86 ;
      RECT 295.9 100.72 446.805 100.79 ;
      RECT 295.83 100.65 446.805 100.72 ;
      RECT 295.76 100.58 446.805 100.65 ;
      RECT 295.69 100.51 446.805 100.58 ;
      RECT 295.62 100.44 446.805 100.51 ;
      RECT 295.55 100.37 446.805 100.44 ;
      RECT 295.48 100.3 446.805 100.37 ;
      RECT 295.41 100.23 446.805 100.3 ;
      RECT 295.34 100.16 446.805 100.23 ;
      RECT 295.27 100.09 446.805 100.16 ;
      RECT 295.2 100.02 446.805 100.09 ;
      RECT 295.13 99.95 446.805 100.02 ;
      RECT 295.06 99.88 446.805 99.95 ;
      RECT 294.99 99.81 446.805 99.88 ;
      RECT 294.92 99.74 446.805 99.81 ;
      RECT 294.85 99.67 446.805 99.74 ;
      RECT 294.78 99.6 446.805 99.67 ;
      RECT 294.71 99.53 446.805 99.6 ;
      RECT 294.64 99.46 446.805 99.53 ;
      RECT 294.57 99.39 446.805 99.46 ;
      RECT 294.5 99.32 446.805 99.39 ;
      RECT 294.43 99.25 446.805 99.32 ;
      RECT 294.36 99.18 446.805 99.25 ;
      RECT 294.29 99.11 446.805 99.18 ;
      RECT 294.22 99.04 446.805 99.11 ;
      RECT 294.15 98.97 446.805 99.04 ;
      RECT 294.08 98.9 446.805 98.97 ;
      RECT 294.01 98.83 446.805 98.9 ;
      RECT 293.94 98.76 446.805 98.83 ;
      RECT 293.87 98.69 446.805 98.76 ;
      RECT 293.8 98.62 446.805 98.69 ;
      RECT 293.73 98.55 446.805 98.62 ;
      RECT 293.66 98.48 446.805 98.55 ;
      RECT 293.59 98.41 446.805 98.48 ;
      RECT 293.52 98.34 446.805 98.41 ;
      RECT 293.45 98.27 446.805 98.34 ;
      RECT 293.38 98.2 446.805 98.27 ;
      RECT 293.31 98.13 446.805 98.2 ;
      RECT 293.24 98.06 446.805 98.13 ;
      RECT 293.17 97.99 446.805 98.06 ;
      RECT 293.1 97.92 446.805 97.99 ;
      RECT 293.03 97.85 446.805 97.92 ;
      RECT 292.96 97.78 446.805 97.85 ;
      RECT 292.89 97.71 446.805 97.78 ;
      RECT 292.82 97.64 446.805 97.71 ;
      RECT 292.75 97.57 446.805 97.64 ;
      RECT 292.68 97.5 446.805 97.57 ;
      RECT 292.61 97.43 446.805 97.5 ;
      RECT 292.54 97.36 446.805 97.43 ;
      RECT 292.47 97.29 446.805 97.36 ;
      RECT 292.4 97.22 446.805 97.29 ;
      RECT 292.33 97.15 446.805 97.22 ;
      RECT 292.26 97.08 446.805 97.15 ;
      RECT 292.19 97.01 446.805 97.08 ;
      RECT 292.12 96.94 446.805 97.01 ;
      RECT 262.955 23.96 268.01 24.03 ;
      RECT 262.885 24.03 268.01 24.1 ;
      RECT 262.815 24.1 268.01 24.17 ;
      RECT 262.745 24.17 268.01 24.24 ;
      RECT 262.675 24.24 268.01 24.31 ;
      RECT 262.605 24.31 268.01 24.38 ;
      RECT 262.535 24.38 268.01 24.45 ;
      RECT 262.465 24.45 268.01 24.49 ;
      RECT 264.71 47.585 280.795 47.63 ;
      RECT 264.67 47.63 280.84 47.675 ;
      RECT 264.635 47.675 280.885 47.68 ;
      RECT 264.63 47.68 280.885 47.685 ;
      RECT 264.7 48.55 280.895 48.62 ;
      RECT 264.77 48.62 280.895 48.69 ;
      RECT 264.84 48.69 280.895 48.76 ;
      RECT 264.91 48.76 280.895 48.83 ;
      RECT 264.935 48.83 280.895 48.855 ;
      RECT 265.18 47.035 280.245 47.105 ;
      RECT 265.12 47.105 280.315 47.175 ;
      RECT 265.06 47.175 280.385 47.245 ;
      RECT 265.0 47.245 280.455 47.315 ;
      RECT 264.94 47.315 280.525 47.385 ;
      RECT 264.88 47.385 280.595 47.455 ;
      RECT 264.82 47.455 280.665 47.525 ;
      RECT 264.76 47.525 280.735 47.585 ;
      RECT 265.425 46.79 280 46.86 ;
      RECT 265.355 46.86 280.07 46.93 ;
      RECT 265.285 46.93 280.14 47 ;
      RECT 265.215 47 280.21 47.035 ;
      RECT 265.655 46.56 280 46.63 ;
      RECT 265.585 46.63 280 46.7 ;
      RECT 265.515 46.7 280 46.77 ;
      RECT 265.445 46.77 280 46.79 ;
      RECT 268.83 36.185 279.64 36.195 ;
      RECT 268.83 36.195 279.63 36.205 ;
      RECT 268.83 45.705 279.63 45.775 ;
      RECT 268.83 45.775 279.7 45.845 ;
      RECT 268.83 45.845 279.77 45.915 ;
      RECT 268.83 45.915 279.84 45.985 ;
      RECT 268.83 45.985 279.91 46.055 ;
      RECT 268.83 46.055 279.98 46.075 ;
      RECT 268.83 17.58 279.375 17.65 ;
      RECT 268.83 17.65 279.445 17.72 ;
      RECT 268.83 17.72 279.515 17.79 ;
      RECT 268.83 17.79 279.585 17.855 ;
      RECT 280.52 45.365 447.625 45.435 ;
      RECT 280.59 45.435 447.625 45.505 ;
      RECT 280.66 45.505 447.625 45.575 ;
      RECT 280.73 45.575 447.625 45.645 ;
      RECT 280.8 45.645 447.625 45.715 ;
      RECT 280.82 45.715 447.625 45.735 ;
      RECT 280.47 36.525 447.625 36.535 ;
      RECT 280.46 36.535 447.625 36.545 ;
      RECT 280.89 46.45 447.625 46.52 ;
      RECT 280.96 46.52 447.625 46.59 ;
      RECT 281.03 46.59 447.625 46.66 ;
      RECT 281.1 46.66 447.625 46.73 ;
      RECT 281.17 46.73 447.625 46.8 ;
      RECT 281.24 46.8 447.625 46.87 ;
      RECT 281.31 46.87 447.625 46.94 ;
      RECT 281.38 46.94 447.625 47.01 ;
      RECT 281.45 47.01 447.625 47.08 ;
      RECT 281.52 47.08 447.625 47.15 ;
      RECT 281.59 47.15 447.625 47.22 ;
      RECT 281.66 47.22 447.625 47.29 ;
      RECT 281.715 47.29 447.625 47.345 ;
      RECT 280.975 74.765 447.625 74.835 ;
      RECT 281.045 74.835 447.625 74.905 ;
      RECT 281.115 74.905 447.625 74.975 ;
      RECT 281.185 74.975 447.625 75.045 ;
      RECT 281.255 75.045 447.625 75.115 ;
      RECT 281.325 75.115 447.625 75.185 ;
      RECT 281.395 75.185 447.625 75.255 ;
      RECT 281.465 75.255 447.625 75.325 ;
      RECT 281.535 75.325 447.625 75.395 ;
      RECT 281.605 75.395 447.625 75.465 ;
      RECT 281.675 75.465 447.625 75.535 ;
      RECT 281.745 75.535 447.625 75.605 ;
      RECT 281.815 75.605 447.625 75.675 ;
      RECT 281.885 75.675 447.625 75.745 ;
      RECT 281.955 75.745 447.625 75.815 ;
      RECT 282.025 75.815 447.625 75.885 ;
      RECT 282.095 75.885 447.625 75.955 ;
      RECT 282.165 75.955 447.625 76.025 ;
      RECT 282.235 76.025 447.625 76.095 ;
      RECT 282.305 76.095 447.625 76.165 ;
      RECT 282.375 76.165 447.625 76.235 ;
      RECT 282.445 76.235 447.625 76.305 ;
      RECT 282.515 76.305 447.625 76.375 ;
      RECT 282.535 76.375 447.625 76.395 ;
      RECT 281.715 56.68 447.625 56.75 ;
      RECT 281.645 56.75 447.625 56.82 ;
      RECT 281.575 56.82 447.625 56.89 ;
      RECT 281.505 56.89 447.625 56.96 ;
      RECT 281.435 56.96 447.625 57.03 ;
      RECT 281.365 57.03 447.625 57.1 ;
      RECT 281.295 57.1 447.625 57.17 ;
      RECT 281.225 57.17 447.625 57.24 ;
      RECT 281.155 57.24 447.625 57.31 ;
      RECT 281.085 57.31 447.625 57.38 ;
      RECT 281.015 57.38 447.625 57.45 ;
      RECT 280.945 57.45 447.625 57.49 ;
      RECT 282.605 87.425 446.805 87.495 ;
      RECT 282.675 87.495 446.805 87.565 ;
      RECT 282.745 87.565 446.805 87.635 ;
      RECT 282.815 87.635 446.805 87.705 ;
      RECT 282.885 87.705 446.805 87.775 ;
      RECT 282.955 87.775 446.805 87.845 ;
      RECT 283.025 87.845 446.805 87.915 ;
      RECT 283.095 87.915 446.805 87.985 ;
      RECT 283.165 87.985 446.805 88.055 ;
      RECT 283.235 88.055 446.805 88.125 ;
      RECT 283.305 88.125 446.805 88.195 ;
      RECT 283.375 88.195 446.805 88.265 ;
      RECT 283.445 88.265 446.805 88.335 ;
      RECT 283.515 88.335 446.805 88.405 ;
      RECT 283.585 88.405 446.805 88.475 ;
      RECT 283.655 88.475 446.805 88.545 ;
      RECT 136.115 27.745 145.815 27.815 ;
      RECT 136.115 27.815 145.745 27.885 ;
      RECT 136.115 27.885 145.675 27.955 ;
      RECT 136.115 27.955 145.605 28.025 ;
      RECT 136.115 28.025 145.535 28.095 ;
      RECT 136.115 28.095 145.465 28.165 ;
      RECT 136.115 28.165 145.395 28.235 ;
      RECT 136.115 28.235 145.355 28.275 ;
      RECT 150.345 42.21 153.53 42.215 ;
      RECT 150.345 42.215 153.535 42.22 ;
      RECT 154.355 41.87 235.65 41.875 ;
      RECT 154.36 41.875 235.645 41.88 ;
      RECT 236.475 42.21 239.66 42.215 ;
      RECT 236.47 42.215 239.66 42.22 ;
      RECT 240.48 56.34 280.825 56.41 ;
      RECT 240.48 56.41 280.755 56.48 ;
      RECT 240.48 56.48 280.685 56.55 ;
      RECT 240.48 56.55 280.615 56.62 ;
      RECT 240.48 56.62 280.545 56.69 ;
      RECT 240.48 56.69 280.475 56.76 ;
      RECT 240.48 56.76 280.405 56.83 ;
      RECT 240.48 56.83 280.335 56.9 ;
      RECT 240.48 56.9 280.265 56.97 ;
      RECT 240.48 56.97 280.195 57.04 ;
      RECT 240.48 57.04 280.125 57.11 ;
      RECT 240.48 57.11 280.085 57.15 ;
      RECT 243.14 26.695 253.89 26.765 ;
      RECT 243.21 26.765 253.89 26.835 ;
      RECT 243.28 26.835 253.89 26.905 ;
      RECT 243.35 26.905 253.89 26.975 ;
      RECT 243.42 26.975 253.89 27.045 ;
      RECT 243.49 27.045 253.89 27.115 ;
      RECT 243.56 27.115 253.89 27.185 ;
      RECT 243.63 27.185 253.89 27.255 ;
      RECT 243.7 27.255 253.89 27.325 ;
      RECT 243.77 27.325 253.89 27.395 ;
      RECT 243.84 27.395 253.89 27.465 ;
      RECT 243.91 27.465 253.89 27.535 ;
      RECT 243.98 27.535 253.89 27.605 ;
      RECT 244.05 27.605 253.89 27.675 ;
      RECT 244.12 27.675 253.89 27.745 ;
      RECT 244.19 27.745 253.89 27.815 ;
      RECT 244.26 27.815 253.89 27.885 ;
      RECT 244.33 27.885 253.89 27.955 ;
      RECT 244.4 27.955 253.89 28.025 ;
      RECT 244.47 28.025 253.89 28.095 ;
      RECT 244.54 28.095 253.89 28.165 ;
      RECT 244.61 28.165 253.89 28.235 ;
      RECT 244.65 28.235 253.89 28.275 ;
      RECT 244.65 48.715 263.74 48.785 ;
      RECT 244.65 48.785 263.67 48.855 ;
      RECT 244.65 45.74 265.245 45.81 ;
      RECT 244.65 45.81 265.175 45.88 ;
      RECT 244.65 45.88 265.105 45.95 ;
      RECT 244.65 45.95 265.035 46.02 ;
      RECT 244.65 46.02 264.965 46.09 ;
      RECT 244.65 46.09 264.895 46.16 ;
      RECT 244.65 46.16 264.825 46.23 ;
      RECT 244.65 46.23 264.755 46.3 ;
      RECT 244.65 46.3 264.685 46.37 ;
      RECT 244.65 46.37 264.615 46.44 ;
      RECT 244.65 46.44 264.545 46.51 ;
      RECT 244.65 46.51 264.475 46.58 ;
      RECT 244.65 46.58 264.405 46.65 ;
      RECT 244.65 46.65 264.335 46.72 ;
      RECT 244.65 46.72 264.265 46.79 ;
      RECT 244.65 46.79 264.195 46.86 ;
      RECT 244.65 46.86 264.125 46.93 ;
      RECT 244.65 46.93 264.055 47 ;
      RECT 244.65 47 263.985 47.07 ;
      RECT 244.65 47.07 263.915 47.14 ;
      RECT 244.65 47.14 263.845 47.21 ;
      RECT 244.65 47.21 263.81 47.245 ;
      RECT 255.11 23.55 262.135 23.62 ;
      RECT 255.11 23.62 262.065 23.69 ;
      RECT 255.11 23.69 261.995 23.76 ;
      RECT 255.11 23.76 261.925 23.83 ;
      RECT 255.11 23.83 261.855 23.9 ;
      RECT 255.11 23.9 261.785 23.97 ;
      RECT 255.11 23.97 261.715 24.04 ;
      RECT 255.11 24.04 261.645 24.11 ;
      RECT 255.11 24.11 261.605 24.15 ;
      RECT 255.11 10.29 261.34 10.36 ;
      RECT 255.11 10.36 261.41 10.43 ;
      RECT 255.11 10.43 261.48 10.5 ;
      RECT 255.11 10.5 261.55 10.57 ;
      RECT 255.11 10.57 261.62 10.64 ;
      RECT 255.11 10.64 261.69 10.71 ;
      RECT 255.11 10.71 261.76 10.78 ;
      RECT 255.11 10.78 261.83 10.85 ;
      RECT 255.11 10.85 261.9 10.92 ;
      RECT 255.11 10.92 261.97 10.99 ;
      RECT 255.11 10.99 262.04 11.06 ;
      RECT 255.11 11.06 262.11 11.13 ;
      RECT 255.11 11.13 262.18 11.155 ;
      RECT 255.18 28.725 261.605 28.795 ;
      RECT 255.25 28.795 261.605 28.865 ;
      RECT 255.32 28.865 261.605 28.935 ;
      RECT 255.39 28.935 261.605 29.005 ;
      RECT 255.46 29.005 261.605 29.075 ;
      RECT 255.53 29.075 261.605 29.145 ;
      RECT 255.6 29.145 261.605 29.215 ;
      RECT 255.64 29.215 261.605 29.255 ;
      RECT 255.71 29.255 261.605 29.325 ;
      RECT 255.78 29.325 261.605 29.395 ;
      RECT 255.85 29.395 261.605 29.465 ;
      RECT 255.92 29.465 261.605 29.535 ;
      RECT 255.99 29.535 261.605 29.605 ;
      RECT 256.06 29.605 261.605 29.675 ;
      RECT 256.09 29.675 261.605 29.705 ;
      RECT 262.23 9.95 268.01 10.02 ;
      RECT 262.3 10.02 268.01 10.09 ;
      RECT 262.37 10.09 268.01 10.16 ;
      RECT 262.44 10.16 268.01 10.23 ;
      RECT 262.51 10.23 268.01 10.3 ;
      RECT 262.58 10.3 268.01 10.37 ;
      RECT 262.65 10.37 268.01 10.44 ;
      RECT 262.72 10.44 268.01 10.51 ;
      RECT 262.79 10.51 268.01 10.58 ;
      RECT 262.86 10.58 268.01 10.65 ;
      RECT 262.93 10.65 268.01 10.72 ;
      RECT 263.0 10.72 268.01 10.79 ;
      RECT 263.025 10.79 268.01 10.815 ;
      RECT 263.025 23.89 268.01 23.96 ;
      RECT 109.655 47.14 124.93 47.21 ;
      RECT 109.585 47.21 125.0 47.28 ;
      RECT 109.515 47.28 125.07 47.35 ;
      RECT 109.445 47.35 125.14 47.42 ;
      RECT 109.375 47.42 125.21 47.49 ;
      RECT 109.305 47.49 125.28 47.56 ;
      RECT 109.235 47.56 125.35 47.585 ;
      RECT 110.375 45.705 121.175 45.775 ;
      RECT 110.305 45.775 121.175 45.845 ;
      RECT 110.235 45.845 121.175 45.915 ;
      RECT 110.165 45.915 121.175 45.985 ;
      RECT 110.095 45.985 121.175 46.055 ;
      RECT 110.025 46.055 121.175 46.075 ;
      RECT 110.005 46.56 124.35 46.63 ;
      RECT 110.005 46.63 124.42 46.7 ;
      RECT 110.005 46.7 124.49 46.77 ;
      RECT 110.005 46.77 124.56 46.79 ;
      RECT 110.365 36.185 121.175 36.195 ;
      RECT 110.375 36.195 121.175 36.205 ;
      RECT 110.63 17.58 121.175 17.65 ;
      RECT 110.56 17.65 121.175 17.72 ;
      RECT 110.49 17.72 121.175 17.79 ;
      RECT 110.42 17.79 121.175 17.855 ;
      RECT 121.995 23.89 126.98 23.96 ;
      RECT 121.995 23.96 127.05 24.03 ;
      RECT 121.995 24.03 127.12 24.1 ;
      RECT 121.995 24.1 127.19 24.17 ;
      RECT 121.995 24.17 127.26 24.24 ;
      RECT 121.995 24.24 127.33 24.31 ;
      RECT 121.995 24.31 127.4 24.38 ;
      RECT 121.995 24.38 127.47 24.45 ;
      RECT 121.995 24.45 127.54 24.49 ;
      RECT 121.995 9.95 127.775 10.02 ;
      RECT 121.995 10.02 127.705 10.09 ;
      RECT 121.995 10.09 127.635 10.16 ;
      RECT 121.995 10.16 127.565 10.23 ;
      RECT 121.995 10.23 127.495 10.3 ;
      RECT 121.995 10.3 127.425 10.37 ;
      RECT 121.995 10.37 127.355 10.44 ;
      RECT 121.995 10.44 127.285 10.51 ;
      RECT 121.995 10.51 127.215 10.58 ;
      RECT 121.995 10.58 127.145 10.65 ;
      RECT 121.995 10.65 127.075 10.72 ;
      RECT 121.995 10.72 127.005 10.79 ;
      RECT 121.995 10.79 126.98 10.815 ;
      RECT 124.76 45.74 145.355 45.81 ;
      RECT 124.83 45.81 145.355 45.88 ;
      RECT 124.9 45.88 145.355 45.95 ;
      RECT 124.97 45.95 145.355 46.02 ;
      RECT 125.04 46.02 145.355 46.09 ;
      RECT 125.11 46.09 145.355 46.16 ;
      RECT 125.18 46.16 145.355 46.23 ;
      RECT 125.25 46.23 145.355 46.3 ;
      RECT 125.32 46.3 145.355 46.37 ;
      RECT 125.39 46.37 145.355 46.44 ;
      RECT 125.46 46.44 145.355 46.51 ;
      RECT 125.53 46.51 145.355 46.58 ;
      RECT 125.6 46.58 145.355 46.65 ;
      RECT 125.67 46.65 145.355 46.72 ;
      RECT 125.74 46.72 145.355 46.79 ;
      RECT 125.81 46.79 145.355 46.86 ;
      RECT 125.88 46.86 145.355 46.93 ;
      RECT 125.95 46.93 145.355 47 ;
      RECT 126.02 47 145.355 47.07 ;
      RECT 126.09 47.07 145.355 47.14 ;
      RECT 126.16 47.14 145.355 47.21 ;
      RECT 126.195 47.21 145.355 47.245 ;
      RECT 126.265 48.715 145.355 48.785 ;
      RECT 126.335 48.785 145.355 48.855 ;
      RECT 127.87 23.55 134.895 23.62 ;
      RECT 127.94 23.62 134.895 23.69 ;
      RECT 128.01 23.69 134.895 23.76 ;
      RECT 128.08 23.76 134.895 23.83 ;
      RECT 128.15 23.83 134.895 23.9 ;
      RECT 128.22 23.9 134.895 23.97 ;
      RECT 128.29 23.97 134.895 24.04 ;
      RECT 128.36 24.04 134.895 24.11 ;
      RECT 128.4 24.11 134.895 24.15 ;
      RECT 128.665 10.29 134.895 10.36 ;
      RECT 128.595 10.36 134.895 10.43 ;
      RECT 128.525 10.43 134.895 10.5 ;
      RECT 128.455 10.5 134.895 10.57 ;
      RECT 128.385 10.57 134.895 10.64 ;
      RECT 128.315 10.64 134.895 10.71 ;
      RECT 128.245 10.71 134.895 10.78 ;
      RECT 128.175 10.78 134.895 10.85 ;
      RECT 128.105 10.85 134.895 10.92 ;
      RECT 128.035 10.92 134.895 10.99 ;
      RECT 127.965 10.99 134.895 11.06 ;
      RECT 127.895 11.06 134.895 11.13 ;
      RECT 127.825 11.13 134.895 11.155 ;
      RECT 128.4 29.255 134.295 29.325 ;
      RECT 128.4 29.325 134.225 29.395 ;
      RECT 128.4 29.395 134.155 29.465 ;
      RECT 128.4 29.465 134.085 29.535 ;
      RECT 128.4 29.535 134.015 29.605 ;
      RECT 128.4 29.605 133.945 29.675 ;
      RECT 128.4 29.675 133.915 29.705 ;
      RECT 128.4 28.725 134.825 28.795 ;
      RECT 128.4 28.795 134.755 28.865 ;
      RECT 128.4 28.865 134.685 28.935 ;
      RECT 128.4 28.935 134.615 29.005 ;
      RECT 128.4 29.005 134.545 29.075 ;
      RECT 128.4 29.075 134.475 29.145 ;
      RECT 128.4 29.145 134.405 29.215 ;
      RECT 128.4 29.215 134.365 29.255 ;
      RECT 136.115 26.695 146.865 26.765 ;
      RECT 136.115 26.765 146.795 26.835 ;
      RECT 136.115 26.835 146.725 26.905 ;
      RECT 136.115 26.905 146.655 26.975 ;
      RECT 136.115 26.975 146.585 27.045 ;
      RECT 136.115 27.045 146.515 27.115 ;
      RECT 136.115 27.115 146.445 27.185 ;
      RECT 136.115 27.185 146.375 27.255 ;
      RECT 136.115 27.255 146.305 27.325 ;
      RECT 136.115 27.325 146.235 27.395 ;
      RECT 136.115 27.395 146.165 27.465 ;
      RECT 136.115 27.465 146.095 27.535 ;
      RECT 136.115 27.535 146.025 27.605 ;
      RECT 136.115 27.605 145.955 27.675 ;
      RECT 136.115 27.675 145.885 27.745 ;
      RECT 98.435 97.62 291.57 97.69 ;
      RECT 98.505 97.55 291.5 97.62 ;
      RECT 98.575 97.48 291.43 97.55 ;
      RECT 98.645 97.41 291.36 97.48 ;
      RECT 98.715 97.34 291.29 97.41 ;
      RECT 98.785 97.27 291.22 97.34 ;
      RECT 98.855 97.2 291.15 97.27 ;
      RECT 98.925 97.13 291.08 97.2 ;
      RECT 98.995 97.06 291.01 97.13 ;
      RECT 99.065 96.99 290.94 97.06 ;
      RECT 99.135 96.92 290.87 96.99 ;
      RECT 99.205 96.85 290.8 96.92 ;
      RECT 99.275 96.78 290.73 96.85 ;
      RECT 99.345 96.71 290.66 96.78 ;
      RECT 99.415 96.64 290.59 96.71 ;
      RECT 99.485 96.57 290.52 96.64 ;
      RECT 99.555 96.5 290.45 96.57 ;
      RECT 99.625 96.43 290.38 96.5 ;
      RECT 99.695 96.36 290.31 96.43 ;
      RECT 99.765 96.29 290.24 96.36 ;
      RECT 99.835 96.22 290.17 96.29 ;
      RECT 99.905 96.15 290.1 96.22 ;
      RECT 99.975 96.08 290.03 96.15 ;
      RECT 100.045 96.01 289.96 96.08 ;
      RECT 100.115 95.94 289.89 96.01 ;
      RECT 100.185 95.87 289.82 95.94 ;
      RECT 100.255 95.8 289.75 95.87 ;
      RECT 100.325 95.73 289.68 95.8 ;
      RECT 100.395 95.66 289.61 95.73 ;
      RECT 100.465 95.59 289.54 95.66 ;
      RECT 100.535 95.52 289.47 95.59 ;
      RECT 100.605 95.45 289.4 95.52 ;
      RECT 100.675 95.38 289.33 95.45 ;
      RECT 100.745 95.31 289.26 95.38 ;
      RECT 100.815 95.24 289.19 95.31 ;
      RECT 106.375 94.365 283.63 94.435 ;
      RECT 106.305 94.435 283.7 94.505 ;
      RECT 106.235 94.505 283.77 94.575 ;
      RECT 106.165 94.575 283.84 94.645 ;
      RECT 106.095 94.645 283.91 94.715 ;
      RECT 106.025 94.715 283.98 94.785 ;
      RECT 105.955 94.785 284.05 94.855 ;
      RECT 105.885 94.855 284.12 94.925 ;
      RECT 105.815 94.925 284.19 94.995 ;
      RECT 105.745 94.995 284.26 95.065 ;
      RECT 105.675 95.065 284.33 95.135 ;
      RECT 105.605 95.135 284.4 95.205 ;
      RECT 105.535 95.205 284.47 95.24 ;
      RECT 108.29 87.765 281.715 87.835 ;
      RECT 108.22 87.835 281.785 87.905 ;
      RECT 108.15 87.905 281.855 87.975 ;
      RECT 108.08 87.975 281.925 88.045 ;
      RECT 108.01 88.045 281.995 88.115 ;
      RECT 107.94 88.115 282.065 88.185 ;
      RECT 107.87 88.185 282.135 88.255 ;
      RECT 107.8 88.255 282.205 88.325 ;
      RECT 107.73 88.325 282.275 88.395 ;
      RECT 107.66 88.395 282.345 88.465 ;
      RECT 107.59 88.465 282.415 88.535 ;
      RECT 107.52 88.535 282.485 88.605 ;
      RECT 107.45 88.605 282.555 88.675 ;
      RECT 107.38 88.675 282.625 88.745 ;
      RECT 107.31 88.745 282.695 88.815 ;
      RECT 107.24 88.815 282.765 88.885 ;
      RECT 107.17 88.885 282.835 88.955 ;
      RECT 107.1 88.955 282.905 89.025 ;
      RECT 107.03 89.025 282.975 89.095 ;
      RECT 106.96 89.095 283.045 89.165 ;
      RECT 106.89 89.165 283.115 89.235 ;
      RECT 106.82 89.235 283.185 89.305 ;
      RECT 106.75 89.305 283.255 89.375 ;
      RECT 106.68 89.375 283.325 89.445 ;
      RECT 106.61 89.445 283.395 89.515 ;
      RECT 106.54 89.515 283.465 89.585 ;
      RECT 106.47 89.585 283.535 89.655 ;
      RECT 106.4 89.655 283.605 89.68 ;
      RECT 109.92 75.105 280.085 75.175 ;
      RECT 109.85 75.175 280.155 75.245 ;
      RECT 109.78 75.245 280.225 75.315 ;
      RECT 109.71 75.315 280.295 75.385 ;
      RECT 109.64 75.385 280.365 75.455 ;
      RECT 109.57 75.455 280.435 75.525 ;
      RECT 109.5 75.525 280.505 75.595 ;
      RECT 109.43 75.595 280.575 75.665 ;
      RECT 109.36 75.665 280.645 75.735 ;
      RECT 109.29 75.735 280.715 75.805 ;
      RECT 109.22 75.805 280.785 75.875 ;
      RECT 109.15 75.875 280.855 75.945 ;
      RECT 109.08 75.945 280.925 76.015 ;
      RECT 109.01 76.015 280.995 76.085 ;
      RECT 108.94 76.085 281.065 76.155 ;
      RECT 108.87 76.155 281.135 76.225 ;
      RECT 108.8 76.225 281.205 76.295 ;
      RECT 108.73 76.295 281.275 76.365 ;
      RECT 108.66 76.365 281.345 76.435 ;
      RECT 108.59 76.435 281.415 76.505 ;
      RECT 108.52 76.505 281.485 76.575 ;
      RECT 108.45 76.575 281.555 76.645 ;
      RECT 108.38 76.645 281.625 76.715 ;
      RECT 108.31 76.715 281.695 76.735 ;
      RECT 109.21 47.585 125.375 47.635 ;
      RECT 109.16 47.635 125.375 47.685 ;
      RECT 109.18 56.34 149.525 56.41 ;
      RECT 109.25 56.41 149.525 56.48 ;
      RECT 109.32 56.48 149.525 56.55 ;
      RECT 109.39 56.55 149.525 56.62 ;
      RECT 109.46 56.62 149.525 56.69 ;
      RECT 109.53 56.69 149.525 56.76 ;
      RECT 109.6 56.76 149.525 56.83 ;
      RECT 109.67 56.83 149.525 56.9 ;
      RECT 109.74 56.9 149.525 56.97 ;
      RECT 109.81 56.97 149.525 57.04 ;
      RECT 109.88 57.04 149.525 57.11 ;
      RECT 109.92 57.11 149.525 57.15 ;
      RECT 109.11 48.55 125.305 48.62 ;
      RECT 109.11 48.62 125.235 48.69 ;
      RECT 109.11 48.69 125.165 48.76 ;
      RECT 109.11 48.76 125.095 48.83 ;
      RECT 109.11 48.83 125.07 48.855 ;
      RECT 110.005 46.79 124.58 46.86 ;
      RECT 109.935 46.86 124.65 46.93 ;
      RECT 109.865 46.93 124.72 47 ;
      RECT 109.795 47 124.79 47.07 ;
      RECT 109.725 47.07 124.86 47.14 ;
      RECT 0 94.77 100.055 94.84 ;
      RECT 0 94.7 100.125 94.77 ;
      RECT 0 94.63 100.195 94.7 ;
      RECT 0 94.56 100.265 94.63 ;
      RECT 0 94.49 100.335 94.56 ;
      RECT 0 94.42 100.405 94.49 ;
      RECT 0 111.715 92.025 111.785 ;
      RECT 0 111.785 92.095 111.855 ;
      RECT 0 111.855 92.165 111.925 ;
      RECT 0 111.925 92.235 111.995 ;
      RECT 0 111.995 92.305 112.04 ;
      RECT 0 74.765 109.03 74.835 ;
      RECT 0 74.835 108.96 74.905 ;
      RECT 0 74.905 108.89 74.975 ;
      RECT 0 74.975 108.82 75.045 ;
      RECT 0 75.045 108.75 75.115 ;
      RECT 0 75.115 108.68 75.185 ;
      RECT 0 75.185 108.61 75.255 ;
      RECT 0 75.255 108.54 75.325 ;
      RECT 0 75.325 108.47 75.395 ;
      RECT 0 75.395 108.4 75.465 ;
      RECT 0 75.465 108.33 75.535 ;
      RECT 0 75.535 108.26 75.605 ;
      RECT 0 75.605 108.19 75.675 ;
      RECT 0 75.675 108.12 75.745 ;
      RECT 0 75.745 108.05 75.815 ;
      RECT 0 75.815 107.98 75.885 ;
      RECT 0 75.885 107.91 75.955 ;
      RECT 0 75.955 107.84 76.025 ;
      RECT 0 76.025 107.77 76.095 ;
      RECT 0 76.095 107.7 76.165 ;
      RECT 0 76.165 107.63 76.235 ;
      RECT 0 76.235 107.56 76.305 ;
      RECT 0 76.305 107.49 76.375 ;
      RECT 0 76.375 107.47 76.395 ;
      RECT 87.375 1.465 106.43 1.535 ;
      RECT 87.375 1.535 106.5 1.605 ;
      RECT 87.375 1.605 106.57 1.675 ;
      RECT 87.375 1.675 106.64 1.745 ;
      RECT 87.375 1.745 106.71 1.815 ;
      RECT 87.375 1.815 106.78 1.885 ;
      RECT 87.375 1.885 106.85 1.955 ;
      RECT 87.375 1.955 106.92 2.025 ;
      RECT 87.375 2.025 106.99 2.095 ;
      RECT 87.375 2.095 107.06 2.165 ;
      RECT 87.375 2.165 107.13 2.18 ;
      RECT 92.905 103.15 297.1 103.18 ;
      RECT 92.975 103.08 297.03 103.15 ;
      RECT 93.045 103.01 296.96 103.08 ;
      RECT 93.115 102.94 296.89 103.01 ;
      RECT 93.185 102.87 296.82 102.94 ;
      RECT 93.255 102.8 296.75 102.87 ;
      RECT 93.325 102.73 296.68 102.8 ;
      RECT 93.395 102.66 296.61 102.73 ;
      RECT 93.465 102.59 296.54 102.66 ;
      RECT 93.535 102.52 296.47 102.59 ;
      RECT 93.605 102.45 296.4 102.52 ;
      RECT 93.675 102.38 296.33 102.45 ;
      RECT 93.745 102.31 296.26 102.38 ;
      RECT 93.815 102.24 296.19 102.31 ;
      RECT 93.885 102.17 296.12 102.24 ;
      RECT 93.955 102.1 296.05 102.17 ;
      RECT 94.025 102.03 295.98 102.1 ;
      RECT 94.095 101.96 295.91 102.03 ;
      RECT 94.165 101.89 295.84 101.96 ;
      RECT 94.235 101.82 295.77 101.89 ;
      RECT 94.305 101.75 295.7 101.82 ;
      RECT 94.375 101.68 295.63 101.75 ;
      RECT 94.445 101.61 295.56 101.68 ;
      RECT 94.515 101.54 295.49 101.61 ;
      RECT 94.585 101.47 295.42 101.54 ;
      RECT 94.655 101.4 295.35 101.47 ;
      RECT 94.725 101.33 295.28 101.4 ;
      RECT 94.795 101.26 295.21 101.33 ;
      RECT 94.865 101.19 295.14 101.26 ;
      RECT 94.935 101.12 295.07 101.19 ;
      RECT 95.005 101.05 295.0 101.12 ;
      RECT 95.075 100.98 294.93 101.05 ;
      RECT 95.145 100.91 294.86 100.98 ;
      RECT 95.215 100.84 294.79 100.91 ;
      RECT 95.285 100.77 294.72 100.84 ;
      RECT 95.355 100.7 294.65 100.77 ;
      RECT 95.425 100.63 294.58 100.7 ;
      RECT 95.495 100.56 294.51 100.63 ;
      RECT 95.565 100.49 294.44 100.56 ;
      RECT 95.635 100.42 294.37 100.49 ;
      RECT 95.705 100.35 294.3 100.42 ;
      RECT 95.775 100.28 294.23 100.35 ;
      RECT 95.845 100.21 294.16 100.28 ;
      RECT 95.915 100.14 294.09 100.21 ;
      RECT 95.985 100.07 294.02 100.14 ;
      RECT 96.055 100 293.95 100.07 ;
      RECT 96.125 99.93 293.88 100 ;
      RECT 96.195 99.86 293.81 99.93 ;
      RECT 96.265 99.79 293.74 99.86 ;
      RECT 96.335 99.72 293.67 99.79 ;
      RECT 96.405 99.65 293.6 99.72 ;
      RECT 96.475 99.58 293.53 99.65 ;
      RECT 96.545 99.51 293.46 99.58 ;
      RECT 96.615 99.44 293.39 99.51 ;
      RECT 96.685 99.37 293.32 99.44 ;
      RECT 96.755 99.3 293.25 99.37 ;
      RECT 96.825 99.23 293.18 99.3 ;
      RECT 96.895 99.16 293.11 99.23 ;
      RECT 96.965 99.09 293.04 99.16 ;
      RECT 97.035 99.02 292.97 99.09 ;
      RECT 97.105 98.95 292.9 99.02 ;
      RECT 97.175 98.88 292.83 98.95 ;
      RECT 97.245 98.81 292.76 98.88 ;
      RECT 97.315 98.74 292.69 98.81 ;
      RECT 97.385 98.67 292.62 98.74 ;
      RECT 97.455 98.6 292.55 98.67 ;
      RECT 97.525 98.53 292.48 98.6 ;
      RECT 97.595 98.46 292.41 98.53 ;
      RECT 97.665 98.39 292.34 98.46 ;
      RECT 97.735 98.32 292.27 98.39 ;
      RECT 97.805 98.25 292.2 98.32 ;
      RECT 97.875 98.18 292.13 98.25 ;
      RECT 97.945 98.11 292.06 98.18 ;
      RECT 98.015 98.04 291.99 98.11 ;
      RECT 98.085 97.97 291.92 98.04 ;
      RECT 98.155 97.9 291.85 97.97 ;
      RECT 98.225 97.83 291.78 97.9 ;
      RECT 98.295 97.76 291.71 97.83 ;
      RECT 98.365 97.69 291.64 97.76 ;
      RECT 0 88.965 105.86 89.035 ;
      RECT 0 89.035 105.79 89.105 ;
      RECT 0 89.105 105.72 89.175 ;
      RECT 0 89.175 105.65 89.245 ;
      RECT 0 89.245 105.58 89.315 ;
      RECT 0 89.315 105.53 89.365 ;
      RECT 0 94.05 105.46 94.12 ;
      RECT 0 94.12 105.39 94.19 ;
      RECT 0 94.19 105.32 94.26 ;
      RECT 0 94.26 105.25 94.33 ;
      RECT 0 94.33 105.18 94.4 ;
      RECT 0 94.4 105.16 94.42 ;
      RECT 0 102.82 92.025 102.87 ;
      RECT 0 102.75 92.075 102.82 ;
      RECT 0 102.68 92.145 102.75 ;
      RECT 0 102.61 92.215 102.68 ;
      RECT 0 102.54 92.285 102.61 ;
      RECT 0 102.47 92.355 102.54 ;
      RECT 0 102.4 92.425 102.47 ;
      RECT 0 102.33 92.495 102.4 ;
      RECT 0 102.26 92.565 102.33 ;
      RECT 0 102.19 92.635 102.26 ;
      RECT 0 102.12 92.705 102.19 ;
      RECT 0 102.05 92.775 102.12 ;
      RECT 0 101.98 92.845 102.05 ;
      RECT 0 101.91 92.915 101.98 ;
      RECT 0 101.84 92.985 101.91 ;
      RECT 0 101.77 93.055 101.84 ;
      RECT 0 101.7 93.125 101.77 ;
      RECT 0 101.63 93.195 101.7 ;
      RECT 0 101.56 93.265 101.63 ;
      RECT 0 101.49 93.335 101.56 ;
      RECT 0 101.42 93.405 101.49 ;
      RECT 0 101.35 93.475 101.42 ;
      RECT 0 101.28 93.545 101.35 ;
      RECT 0 101.21 93.615 101.28 ;
      RECT 0 101.14 93.685 101.21 ;
      RECT 0 101.07 93.755 101.14 ;
      RECT 0 101 93.825 101.07 ;
      RECT 0 100.93 93.895 101 ;
      RECT 0 100.86 93.965 100.93 ;
      RECT 0 100.79 94.035 100.86 ;
      RECT 0 100.72 94.105 100.79 ;
      RECT 0 100.65 94.175 100.72 ;
      RECT 0 100.58 94.245 100.65 ;
      RECT 0 100.51 94.315 100.58 ;
      RECT 0 100.44 94.385 100.51 ;
      RECT 0 100.37 94.455 100.44 ;
      RECT 0 100.3 94.525 100.37 ;
      RECT 0 100.23 94.595 100.3 ;
      RECT 0 100.16 94.665 100.23 ;
      RECT 0 100.09 94.735 100.16 ;
      RECT 0 100.02 94.805 100.09 ;
      RECT 0 99.95 94.875 100.02 ;
      RECT 0 99.88 94.945 99.95 ;
      RECT 0 99.81 95.015 99.88 ;
      RECT 0 99.74 95.085 99.81 ;
      RECT 0 99.67 95.155 99.74 ;
      RECT 0 99.6 95.225 99.67 ;
      RECT 0 99.53 95.295 99.6 ;
      RECT 0 99.46 95.365 99.53 ;
      RECT 0 99.39 95.435 99.46 ;
      RECT 0 99.32 95.505 99.39 ;
      RECT 0 99.25 95.575 99.32 ;
      RECT 0 99.18 95.645 99.25 ;
      RECT 0 99.11 95.715 99.18 ;
      RECT 0 99.04 95.785 99.11 ;
      RECT 0 98.97 95.855 99.04 ;
      RECT 0 98.9 95.925 98.97 ;
      RECT 0 98.83 95.995 98.9 ;
      RECT 0 98.76 96.065 98.83 ;
      RECT 0 98.69 96.135 98.76 ;
      RECT 0 98.62 96.205 98.69 ;
      RECT 0 98.55 96.275 98.62 ;
      RECT 0 98.48 96.345 98.55 ;
      RECT 0 98.41 96.415 98.48 ;
      RECT 0 98.34 96.485 98.41 ;
      RECT 0 98.27 96.555 98.34 ;
      RECT 0 98.2 96.625 98.27 ;
      RECT 0 98.13 96.695 98.2 ;
      RECT 0 98.06 96.765 98.13 ;
      RECT 0 97.99 96.835 98.06 ;
      RECT 0 97.92 96.905 97.99 ;
      RECT 0 97.85 96.975 97.92 ;
      RECT 0 97.78 97.045 97.85 ;
      RECT 0 97.71 97.115 97.78 ;
      RECT 0 97.64 97.185 97.71 ;
      RECT 0 97.57 97.255 97.64 ;
      RECT 0 97.5 97.325 97.57 ;
      RECT 0 97.43 97.395 97.5 ;
      RECT 0 97.36 97.465 97.43 ;
      RECT 0 97.29 97.535 97.36 ;
      RECT 0 97.22 97.605 97.29 ;
      RECT 0 97.15 97.675 97.22 ;
      RECT 0 97.08 97.745 97.15 ;
      RECT 0 97.01 97.815 97.08 ;
      RECT 0 96.94 97.885 97.01 ;
      RECT 0 96.87 97.955 96.94 ;
      RECT 0 96.8 98.025 96.87 ;
      RECT 0 96.73 98.095 96.8 ;
      RECT 0 96.66 98.165 96.73 ;
      RECT 0 96.59 98.235 96.66 ;
      RECT 0 96.52 98.305 96.59 ;
      RECT 0 96.45 98.375 96.52 ;
      RECT 0 96.38 98.445 96.45 ;
      RECT 0 96.31 98.515 96.38 ;
      RECT 0 96.24 98.585 96.31 ;
      RECT 0 96.17 98.655 96.24 ;
      RECT 0 96.1 98.725 96.17 ;
      RECT 0 96.03 98.795 96.1 ;
      RECT 0 95.96 98.865 96.03 ;
      RECT 0 95.89 98.935 95.96 ;
      RECT 0 95.82 99.005 95.89 ;
      RECT 0 95.75 99.075 95.82 ;
      RECT 0 95.68 99.145 95.75 ;
      RECT 0 95.61 99.215 95.68 ;
      RECT 0 95.54 99.285 95.61 ;
      RECT 0 95.47 99.355 95.54 ;
      RECT 0 95.4 99.425 95.47 ;
      RECT 0 95.33 99.495 95.4 ;
      RECT 0 95.26 99.565 95.33 ;
      RECT 0 95.19 99.635 95.26 ;
      RECT 0 95.12 99.705 95.19 ;
      RECT 0 95.05 99.775 95.12 ;
      RECT 0 94.98 99.845 95.05 ;
      RECT 0 94.91 99.915 94.98 ;
      RECT 0 94.84 99.985 94.91 ;
      RECT 254.71 30.395 255.13 30.465 ;
      RECT 254.71 30.465 255.2 30.525 ;
      RECT 264.63 47.585 280.795 47.635 ;
      RECT 264.63 47.635 280.845 47.685 ;
      RECT 265.425 46.79 280 46.86 ;
      RECT 265.355 46.86 280.07 46.93 ;
      RECT 265.285 46.93 280.14 47 ;
      RECT 265.215 47 280.21 47.07 ;
      RECT 265.145 47.07 280.28 47.14 ;
      RECT 265.075 47.14 280.35 47.21 ;
      RECT 265.005 47.21 280.42 47.28 ;
      RECT 264.935 47.28 280.49 47.35 ;
      RECT 264.865 47.35 280.56 47.42 ;
      RECT 264.795 47.42 280.63 47.49 ;
      RECT 264.725 47.49 280.7 47.56 ;
      RECT 264.655 47.56 280.77 47.585 ;
      RECT 280.265 17.24 282.04 17.31 ;
      RECT 280.335 17.31 282.04 17.38 ;
      RECT 280.405 17.38 282.04 17.45 ;
      RECT 280.47 17.45 282.04 17.515 ;
      RECT 280.195 1.125 282.685 1.195 ;
      RECT 280.195 1.195 282.615 1.265 ;
      RECT 280.195 1.265 282.545 1.335 ;
      RECT 280.195 1.335 282.475 1.405 ;
      RECT 280.195 1.405 282.405 1.475 ;
      RECT 280.195 1.475 282.335 1.545 ;
      RECT 280.195 1.545 282.265 1.615 ;
      RECT 280.195 1.615 282.195 1.685 ;
      RECT 280.195 1.685 282.125 1.755 ;
      RECT 280.195 1.755 282.055 1.825 ;
      RECT 280.195 1.825 282.04 1.84 ;
      RECT 282.535 83.64 448.815 83.71 ;
      RECT 282.535 83.71 448.745 83.78 ;
      RECT 282.535 83.78 448.675 83.85 ;
      RECT 282.535 83.85 448.605 83.92 ;
      RECT 282.535 83.92 448.535 83.99 ;
      RECT 282.535 83.99 448.465 84.06 ;
      RECT 282.535 84.06 448.395 84.13 ;
      RECT 282.535 84.13 448.325 84.2 ;
      RECT 282.535 84.2 448.255 84.27 ;
      RECT 282.535 84.27 448.185 84.34 ;
      RECT 282.535 84.34 448.115 84.41 ;
      RECT 282.535 84.41 448.045 84.48 ;
      RECT 282.535 84.48 447.975 84.55 ;
      RECT 282.535 84.55 447.905 84.62 ;
      RECT 282.535 84.62 447.835 84.69 ;
      RECT 282.535 84.69 447.765 84.76 ;
      RECT 282.535 84.76 447.695 84.83 ;
      RECT 282.535 84.83 447.625 84.9 ;
      RECT 282.535 84.9 447.555 84.97 ;
      RECT 282.535 84.97 447.485 85.04 ;
      RECT 282.535 85.04 447.415 85.11 ;
      RECT 282.535 85.11 447.345 85.18 ;
      RECT 282.535 85.18 447.275 85.25 ;
      RECT 282.535 85.25 447.205 85.32 ;
      RECT 282.535 85.32 447.135 85.39 ;
      RECT 282.535 85.39 447.065 85.46 ;
      RECT 282.535 85.46 446.995 85.53 ;
      RECT 282.535 85.53 446.925 85.6 ;
      RECT 282.535 85.6 446.855 85.67 ;
      RECT 282.535 85.67 446.805 85.72 ;
      RECT 403.38 14.655 404.695 14.675 ;
      RECT 403.38 14.675 404.675 14.695 ;
      RECT 445.415 22.19 447.625 22.225 ;
      RECT 445.45 22.225 447.625 22.26 ;
      RECT 0 46.45 109.115 46.52 ;
      RECT 0 46.52 109.045 46.59 ;
      RECT 0 46.59 108.975 46.66 ;
      RECT 0 46.66 108.905 46.73 ;
      RECT 0 46.73 108.835 46.8 ;
      RECT 0 46.8 108.765 46.87 ;
      RECT 0 46.87 108.695 46.94 ;
      RECT 0 46.94 108.625 47.01 ;
      RECT 0 47.01 108.555 47.08 ;
      RECT 0 47.08 108.485 47.15 ;
      RECT 0 47.15 108.415 47.22 ;
      RECT 0 47.22 108.345 47.29 ;
      RECT 0 47.29 108.29 47.345 ;
      RECT 0 56.68 108.29 56.75 ;
      RECT 0 56.75 108.36 56.82 ;
      RECT 0 56.82 108.43 56.89 ;
      RECT 0 56.89 108.5 56.96 ;
      RECT 0 56.96 108.57 57.03 ;
      RECT 0 57.03 108.64 57.1 ;
      RECT 0 57.1 108.71 57.17 ;
      RECT 0 57.17 108.78 57.24 ;
      RECT 0 57.24 108.85 57.31 ;
      RECT 0 57.31 108.92 57.38 ;
      RECT 0 57.38 108.99 57.45 ;
      RECT 0 57.45 109.06 57.49 ;
      RECT 0 36.525 109.535 36.535 ;
      RECT 0 36.535 109.545 36.545 ;
      RECT 0 45.365 109.485 45.435 ;
      RECT 0 45.435 109.415 45.505 ;
      RECT 0 45.505 109.345 45.575 ;
      RECT 0 45.575 109.275 45.645 ;
      RECT 0 45.645 109.205 45.715 ;
      RECT 0 45.715 109.185 45.735 ;
      RECT 0 244.075 446.735 244.145 ;
      RECT 0 244.145 446.665 244.215 ;
      RECT 0 244.215 446.64 244.24 ;
      RECT 0 87.425 107.4 87.495 ;
      RECT 0 87.495 107.33 87.565 ;
      RECT 0 87.565 107.26 87.635 ;
      RECT 0 87.635 107.19 87.705 ;
      RECT 0 87.705 107.12 87.775 ;
      RECT 0 87.775 107.05 87.845 ;
      RECT 0 87.845 106.98 87.915 ;
      RECT 0 87.915 106.91 87.985 ;
      RECT 0 87.985 106.84 88.055 ;
      RECT 0 88.055 106.77 88.125 ;
      RECT 0 88.125 106.7 88.195 ;
      RECT 0 88.195 106.63 88.265 ;
      RECT 0 88.265 106.56 88.335 ;
      RECT 0 88.335 106.49 88.405 ;
      RECT 0 88.405 106.42 88.475 ;
      RECT 0 88.475 106.35 88.545 ;
      RECT 0 88.545 106.28 88.615 ;
      RECT 0 88.615 106.21 88.685 ;
      RECT 0 88.685 106.14 88.755 ;
      RECT 0 88.755 106.07 88.825 ;
      RECT 0 88.825 106.0 88.895 ;
      RECT 0 88.895 105.93 88.965 ;
      RECT 135.975 1.765 140.85 1.835 ;
      RECT 135.975 1.835 140.78 1.905 ;
      RECT 135.975 1.905 140.715 1.97 ;
      RECT 147.265 27.525 147.335 27.595 ;
      RECT 147.195 27.595 147.335 27.665 ;
      RECT 147.125 27.665 147.335 27.735 ;
      RECT 147.055 27.735 147.335 27.805 ;
      RECT 146.985 27.805 147.335 27.875 ;
      RECT 146.915 27.875 147.335 27.945 ;
      RECT 146.845 27.945 147.335 28.015 ;
      RECT 146.775 28.015 147.335 28.085 ;
      RECT 146.705 28.085 147.335 28.155 ;
      RECT 146.635 28.155 147.335 28.225 ;
      RECT 146.565 28.225 147.335 28.295 ;
      RECT 146.495 28.295 147.335 28.365 ;
      RECT 146.425 28.365 147.335 28.435 ;
      RECT 146.355 28.435 147.335 28.505 ;
      RECT 146.285 28.505 147.335 28.575 ;
      RECT 146.215 28.575 147.335 28.615 ;
      RECT 148.155 30.61 149.995 30.68 ;
      RECT 148.155 30.68 149.925 30.75 ;
      RECT 148.155 30.75 149.855 30.82 ;
      RECT 148.155 30.82 149.785 30.89 ;
      RECT 148.155 30.89 149.715 30.96 ;
      RECT 148.155 30.96 149.645 31.03 ;
      RECT 148.155 31.03 149.575 31.1 ;
      RECT 148.155 31.1 149.525 31.15 ;
      RECT 148.155 28.365 149.525 28.435 ;
      RECT 148.155 28.435 149.595 28.505 ;
      RECT 148.155 28.505 149.665 28.575 ;
      RECT 148.155 28.575 149.735 28.645 ;
      RECT 148.155 28.645 149.805 28.715 ;
      RECT 148.155 28.715 149.875 28.785 ;
      RECT 148.155 28.785 149.945 28.855 ;
      RECT 148.155 28.855 150.015 28.905 ;
      RECT 150.345 2.1 153.12 2.11 ;
      RECT 150.345 2.11 153.11 2.12 ;
      RECT 150.885 31.215 153.13 31.285 ;
      RECT 150.815 31.285 153.13 31.355 ;
      RECT 150.745 31.355 153.13 31.425 ;
      RECT 150.675 31.425 153.13 31.495 ;
      RECT 150.605 31.495 153.13 31.565 ;
      RECT 150.535 31.565 153.13 31.635 ;
      RECT 150.465 31.635 153.13 31.705 ;
      RECT 150.395 31.705 153.13 31.755 ;
      RECT 150.345 3.12 153.11 3.13 ;
      RECT 150.345 3.13 153.12 3.14 ;
      RECT 150.415 27.76 153.13 27.83 ;
      RECT 150.485 27.83 153.13 27.9 ;
      RECT 150.555 27.9 153.13 27.97 ;
      RECT 150.625 27.97 153.13 28.04 ;
      RECT 150.695 28.04 153.13 28.11 ;
      RECT 150.765 28.11 153.13 28.18 ;
      RECT 150.835 28.18 153.13 28.25 ;
      RECT 150.885 28.25 153.13 28.3 ;
      RECT 236.92 3.12 239.66 3.145 ;
      RECT 236.895 3.145 239.66 3.165 ;
      RECT 236.875 31.215 239.12 31.285 ;
      RECT 236.875 31.285 239.19 31.355 ;
      RECT 236.875 31.355 239.26 31.425 ;
      RECT 236.875 31.425 239.33 31.495 ;
      RECT 236.875 31.495 239.4 31.565 ;
      RECT 236.875 31.565 239.47 31.635 ;
      RECT 236.875 31.635 239.54 31.705 ;
      RECT 236.875 31.705 239.61 31.755 ;
      RECT 236.895 2.075 239.66 2.095 ;
      RECT 236.915 2.095 239.66 2.115 ;
      RECT 236.92 2.115 239.66 2.12 ;
      RECT 236.875 27.76 239.59 27.83 ;
      RECT 236.875 27.83 239.52 27.9 ;
      RECT 236.875 27.9 239.45 27.97 ;
      RECT 236.875 27.97 239.38 28.04 ;
      RECT 236.875 28.04 239.31 28.11 ;
      RECT 236.875 28.11 239.24 28.18 ;
      RECT 236.875 28.18 239.17 28.25 ;
      RECT 236.875 28.25 239.12 28.3 ;
      RECT 240.48 28.365 241.85 28.435 ;
      RECT 240.41 28.435 241.85 28.505 ;
      RECT 240.34 28.505 241.85 28.575 ;
      RECT 240.27 28.575 241.85 28.645 ;
      RECT 240.2 28.645 241.85 28.715 ;
      RECT 240.13 28.715 241.85 28.785 ;
      RECT 240.06 28.785 241.85 28.855 ;
      RECT 239.99 28.855 241.85 28.905 ;
      RECT 240.01 30.61 241.85 30.68 ;
      RECT 240.08 30.68 241.85 30.75 ;
      RECT 240.15 30.75 241.85 30.82 ;
      RECT 240.22 30.82 241.85 30.89 ;
      RECT 240.29 30.89 241.85 30.96 ;
      RECT 240.36 30.96 241.85 31.03 ;
      RECT 240.43 31.03 241.85 31.1 ;
      RECT 240.48 31.1 241.85 31.15 ;
      RECT 242.67 27.525 242.74 27.595 ;
      RECT 242.67 27.595 242.81 27.665 ;
      RECT 242.67 27.665 242.88 27.735 ;
      RECT 242.67 27.735 242.95 27.805 ;
      RECT 242.67 27.805 243.02 27.875 ;
      RECT 242.67 27.875 243.09 27.945 ;
      RECT 242.67 27.945 243.16 28.015 ;
      RECT 242.67 28.015 243.23 28.085 ;
      RECT 242.67 28.085 243.3 28.155 ;
      RECT 242.67 28.155 243.37 28.225 ;
      RECT 242.67 28.225 243.44 28.295 ;
      RECT 242.67 28.295 243.51 28.365 ;
      RECT 242.67 28.365 243.58 28.435 ;
      RECT 242.67 28.435 243.65 28.505 ;
      RECT 242.67 28.505 243.72 28.575 ;
      RECT 242.67 28.575 243.79 28.615 ;
      RECT 249.155 1.765 254.03 1.835 ;
      RECT 249.225 1.835 254.03 1.905 ;
      RECT 249.29 1.905 254.03 1.97 ;
      RECT 254.71 30.045 254.78 30.115 ;
      RECT 254.71 30.115 254.85 30.185 ;
      RECT 254.71 30.185 254.92 30.255 ;
      RECT 254.71 30.255 254.99 30.325 ;
      RECT 254.71 30.325 255.06 30.395 ;
      RECT 283.575 0 302.63 18.435 ;
      RECT 283.575 0 302.63 18.435 ;
      RECT 283.575 0 302.63 1.465 ;
      RECT 282.535 85.72 446.805 87.425 ;
      RECT 282.535 83.64 447.625 84.9 ;
      RECT 282.535 76.395 447.625 83.64 ;
      RECT 284.475 89.365 446.805 94.05 ;
      RECT 284.475 76.395 446.805 94.05 ;
      RECT 280.47 33.515 447.625 36.525 ;
      RECT 305.025 0 402.56 23.42 ;
      RECT 405.535 0 419.165 5.315 ;
      RECT 403.38 15.35 422.41 30.825 ;
      RECT 403.38 15.35 422.41 23.42 ;
      RECT 405.535 5.315 422.41 14.53 ;
      RECT 405.875 14.53 422.41 15.35 ;
      RECT 405.875 5.315 422.41 15.35 ;
      RECT 304.04 30.825 447.625 33.515 ;
      RECT 305.025 23.42 447.625 33.515 ;
      RECT 305.025 23.42 447.625 30.825 ;
      RECT 423.23 0 444.56 30.825 ;
      RECT 423.23 23.295 447.625 30.825 ;
      RECT 423.23 23.295 447.625 23.42 ;
      RECT 423.23 0 444.56 23.295 ;
      RECT 0 246.095 480 253.715 ;
      RECT 449.785 242.505 480 253.715 ;
      RECT 449.785 242.505 480 253.715 ;
      RECT 449.785 242.505 480 253.715 ;
      RECT 449.785 242.505 480 246.095 ;
      RECT 452.035 240.135 480 242.505 ;
      RECT 454.445 0 464.25 60.575 ;
      RECT 454.445 60.575 480 242.505 ;
      RECT 454.445 60.575 480 237.725 ;
      RECT 466.95 0 480 60.575 ;
      RECT 0 102.87 92.025 112.42 ;
      RECT 110.005 46.075 121.175 46.56 ;
      RECT 110.375 36.205 121.175 46.79 ;
      RECT 0 47.345 108.29 74.765 ;
      RECT 0 45.735 109.185 46.45 ;
      RECT 0 30.825 85.965 45.365 ;
      RECT 0 36.545 109.555 45.365 ;
      RECT 0 33.515 109.535 45.365 ;
      RECT 87.375 18.435 109.535 45.365 ;
      RECT 109.11 52.125 149.525 56.34 ;
      RECT 109.92 52.125 149.525 75.105 ;
      RECT 109.92 52.125 149.525 75.105 ;
      RECT 126.195 47.245 145.355 48.715 ;
      RECT 126.335 48.715 144.975 56.34 ;
      RECT 126.335 48.715 144.975 56.34 ;
      RECT 126.335 48.715 144.975 56.34 ;
      RECT 126.335 49.895 149.525 56.34 ;
      RECT 126.335 49.895 149.525 56.34 ;
      RECT 126.335 49.895 149.525 56.34 ;
      RECT 126.335 49.895 149.525 52.125 ;
      RECT 126.335 48.855 145.355 49.075 ;
      RECT 135.975 2.625 141.725 6.1 ;
      RECT 135.975 1.57 140.715 1.765 ;
      RECT 136.115 2.625 141.725 10.87 ;
      RECT 136.115 2.625 141.725 10.87 ;
      RECT 136.115 6.1 141.725 7.86 ;
      RECT 128.665 2.61 134.895 11.155 ;
      RECT 128.665 2.61 134.895 11.155 ;
      RECT 128.665 2.61 134.895 11.155 ;
      RECT 128.665 7.81 134.895 10.29 ;
      RECT 128.665 2.61 135.035 7.81 ;
      RECT 254.97 2.61 261.34 7.81 ;
      RECT 255.11 2.61 261.34 11.155 ;
      RECT 255.11 2.61 261.34 11.155 ;
      RECT 255.11 2.61 261.34 11.155 ;
      RECT 255.11 7.81 261.34 10.29 ;
      RECT 268.83 36.205 279.63 46.79 ;
      RECT 268.83 36.205 279.63 46.79 ;
      RECT 268.83 46.075 280 46.56 ;
      RECT 240.48 49.895 263.67 56.34 ;
      RECT 240.48 49.895 263.67 56.34 ;
      RECT 240.48 49.895 263.67 56.34 ;
      RECT 240.48 49.895 263.67 52.125 ;
      RECT 244.65 47.245 263.81 48.715 ;
      RECT 244.65 43.19 268.01 45.74 ;
      RECT 245.03 48.715 263.67 56.34 ;
      RECT 245.03 48.715 263.67 56.34 ;
      RECT 245.03 48.715 263.67 56.34 ;
      RECT 262.425 24.49 268.01 45.74 ;
      RECT 262.425 24.49 268.01 45.74 ;
      RECT 262.425 24.49 268.01 45.74 ;
      RECT 262.425 24.49 268.01 45.74 ;
      RECT 240.48 52.125 280.085 75.105 ;
      RECT 240.48 52.125 280.085 75.105 ;
      RECT 240.48 52.125 280.895 56.34 ;
      RECT 264.63 48.145 280.895 48.55 ;
      RECT 264.63 47.685 280.895 48.145 ;
      RECT 264.935 47.685 280.895 56.34 ;
      RECT 264.935 47.685 280.895 56.34 ;
      RECT 264.935 47.685 280.895 56.34 ;
      RECT 280.45 36.545 447.625 45.365 ;
      RECT 280.47 33.515 447.625 45.365 ;
      RECT 280.82 45.735 447.625 46.45 ;
      RECT 281.715 47.345 447.625 74.765 ;
      RECT 304.04 30.825 447.625 45.365 ;
      RECT 92.875 103.18 297.13 111.22 ;
      RECT 0 244.075 446.64 253.715 ;
      RECT 0 244.075 446.64 253.715 ;
      RECT 0 244.075 446.64 253.715 ;
      RECT 0 112.42 446.64 253.715 ;
      RECT 0 112.42 446.805 244.075 ;
      RECT 107.32 1.125 109.81 1.195 ;
      RECT 107.39 1.195 109.81 1.265 ;
      RECT 107.46 1.265 109.81 1.335 ;
      RECT 107.53 1.335 109.81 1.405 ;
      RECT 107.6 1.405 109.81 1.475 ;
      RECT 107.67 1.475 109.81 1.545 ;
      RECT 107.74 1.545 109.81 1.615 ;
      RECT 107.81 1.615 109.81 1.685 ;
      RECT 107.88 1.685 109.81 1.755 ;
      RECT 107.95 1.755 109.81 1.825 ;
      RECT 107.965 1.825 109.81 1.84 ;
      RECT 107.965 17.24 109.74 17.31 ;
      RECT 107.965 17.31 109.67 17.38 ;
      RECT 107.965 17.38 109.6 17.45 ;
      RECT 107.965 17.45 109.535 17.515 ;
      RECT 135.225 30.045 135.295 30.115 ;
      RECT 135.155 30.115 135.295 30.185 ;
      RECT 135.085 30.185 135.295 30.255 ;
      RECT 135.015 30.255 135.295 30.325 ;
      RECT 134.945 30.325 135.295 30.395 ;
      RECT 134.875 30.395 135.295 30.465 ;
      RECT 134.805 30.465 135.295 30.525 ;
      RECT 109.11 48.855 125.07 52.125 ;
      RECT 109.11 48.55 125.07 52.125 ;
      RECT 109.11 48.55 125.07 52.125 ;
      RECT 109.11 48.55 125.07 52.125 ;
      RECT 109.11 48.55 125.07 52.125 ;
      RECT 109.92 57.15 149.525 58.805 ;
      RECT 110.355 17.855 121.175 36.185 ;
      RECT 110.63 0 121.175 17.58 ;
      RECT 121.995 10.815 126.98 23.89 ;
      RECT 121.995 9.95 126.98 23.89 ;
      RECT 121.995 9.95 126.98 23.89 ;
      RECT 121.995 7.81 127.845 9.95 ;
      RECT 121.995 0 127.845 7.81 ;
      RECT 121.995 2.61 127.98 7.81 ;
      RECT 121.995 0 127.845 7.81 ;
      RECT 121.995 0 127.845 2.61 ;
      RECT 121.995 24.49 127.58 45.74 ;
      RECT 121.995 24.49 127.58 45.74 ;
      RECT 121.995 24.49 127.58 45.74 ;
      RECT 121.995 24.49 127.58 45.74 ;
      RECT 121.995 24.49 127.58 43.19 ;
      RECT 128.4 24.15 134.895 28.725 ;
      RECT 127.8 11.155 134.895 23.55 ;
      RECT 128.4 30.525 133.855 42.37 ;
      RECT 128.4 28.725 133.475 42.37 ;
      RECT 128.4 29.705 133.475 30.525 ;
      RECT 129.16 30.525 133.855 43.19 ;
      RECT 129.16 30.525 133.855 43.19 ;
      RECT 129.16 30.525 133.855 43.19 ;
      RECT 129.16 42.37 133.855 43.02 ;
      RECT 121.995 43.19 145.355 45.74 ;
      RECT 129.16 43.02 145.355 43.19 ;
      RECT 136.115 0 140.715 1.57 ;
      RECT 136.115 7.86 142.125 26.695 ;
      RECT 136.115 7.86 142.125 26.695 ;
      RECT 136.115 7.86 142.125 10.87 ;
      RECT 134.675 37.23 145.355 43.19 ;
      RECT 134.675 37.23 145.355 43.19 ;
      RECT 134.675 37.23 145.355 43.19 ;
      RECT 134.675 37.23 145.355 43.02 ;
      RECT 136.115 28.275 145.355 37.23 ;
      RECT 136.115 26.695 145.355 37.23 ;
      RECT 136.115 10.87 146.935 26.695 ;
      RECT 142.945 0 146.935 26.695 ;
      RECT 142.945 0 146.935 10.87 ;
      RECT 146.175 46.415 149.525 56.34 ;
      RECT 146.175 46.415 149.525 56.34 ;
      RECT 146.175 46.415 149.525 56.34 ;
      RECT 146.175 46.415 149.525 52.125 ;
      RECT 146.175 46.415 149.525 49.895 ;
      RECT 150.345 35.225 153.53 42.21 ;
      RECT 150.345 35.225 153.53 57.985 ;
      RECT 150.345 35.225 153.53 57.985 ;
      RECT 150.345 42.22 153.54 43.19 ;
      RECT 154.36 41.88 235.645 43.19 ;
      RECT 154.35 34.115 235.655 41.87 ;
      RECT 154.36 41.87 235.645 57.985 ;
      RECT 154.36 41.87 235.645 57.985 ;
      RECT 156.52 33.375 233.485 41.87 ;
      RECT 156.52 33.375 233.485 34.115 ;
      RECT 156.92 0 176.71 24.51 ;
      RECT 179.27 0 210.735 24.51 ;
      RECT 156.92 24.51 233.085 41.87 ;
      RECT 156.92 24.51 233.085 33.375 ;
      RECT 213.295 0 233.085 24.51 ;
      RECT 150.725 57.985 239.28 58.805 ;
      RECT 150.345 43.19 239.66 57.985 ;
      RECT 150.725 43.19 239.28 58.805 ;
      RECT 150.725 43.19 239.28 58.805 ;
      RECT 150.725 43.19 239.28 58.805 ;
      RECT 236.465 42.22 239.66 57.985 ;
      RECT 236.465 42.22 239.66 57.985 ;
      RECT 236.465 42.22 239.66 43.19 ;
      RECT 236.475 35.225 239.66 42.22 ;
      RECT 236.475 35.225 239.66 42.22 ;
      RECT 236.475 35.225 239.66 42.21 ;
      RECT 109.92 58.805 280.085 75.105 ;
      RECT 240.48 57.15 280.085 58.805 ;
      RECT 240.48 46.415 243.83 56.34 ;
      RECT 240.48 46.415 243.83 56.34 ;
      RECT 240.48 46.415 243.83 56.34 ;
      RECT 240.48 46.415 243.83 52.125 ;
      RECT 240.48 46.415 243.83 49.895 ;
      RECT 243.07 0 247.06 26.695 ;
      RECT 243.07 0 247.06 10.87 ;
      RECT 244.65 28.275 253.89 37.23 ;
      RECT 244.65 37.23 255.33 43.19 ;
      RECT 244.65 37.23 255.33 43.19 ;
      RECT 244.65 37.23 255.33 43.19 ;
      RECT 244.65 37.23 255.33 43.02 ;
      RECT 243.07 10.87 253.89 26.695 ;
      RECT 244.65 10.87 253.89 37.23 ;
      RECT 247.88 7.86 253.89 26.695 ;
      RECT 247.88 7.86 253.89 26.695 ;
      RECT 247.88 7.86 253.89 10.87 ;
      RECT 248.28 6.1 253.89 7.86 ;
      RECT 249.29 0 253.89 1.57 ;
      RECT 249.29 1.57 254.03 1.765 ;
      RECT 248.28 2.625 253.89 10.87 ;
      RECT 248.28 2.625 253.89 10.87 ;
      RECT 248.28 2.625 254.03 6.1 ;
      RECT 249.29 1.97 254.03 2.625 ;
      RECT 249.29 1.765 254.03 1.97 ;
      RECT 255.11 11.155 262.205 23.55 ;
      RECT 244.65 43.02 260.845 43.19 ;
      RECT 255.11 24.15 261.605 28.725 ;
      RECT 255.64 24.15 261.605 29.705 ;
      RECT 256.15 42.37 260.845 43.02 ;
      RECT 256.15 30.525 261.605 42.37 ;
      RECT 256.53 24.15 261.605 42.37 ;
      RECT 256.53 29.705 261.605 30.525 ;
      RECT 262.025 2.61 268.01 7.81 ;
      RECT 262.16 0 268.01 7.81 ;
      RECT 262.16 0 268.01 7.81 ;
      RECT 262.16 0 268.01 2.61 ;
      RECT 262.425 24.49 268.01 43.19 ;
      RECT 262.16 7.81 268.01 9.95 ;
      RECT 263.025 10.815 268.01 23.89 ;
      RECT 263.025 9.95 268.01 23.89 ;
      RECT 263.025 9.95 268.01 23.89 ;
      RECT 268.83 0 279.375 17.58 ;
      RECT 268.83 17.855 279.65 36.185 ;
      RECT 280.905 57.49 447.625 74.765 ;
      RECT 280.47 18.435 302.63 36.525 ;
      RECT 280.47 18.435 302.63 33.515 ;
      RECT 282.805 2.28 302.63 18.435 ;
      RECT 282.86 2.18 302.63 2.28 ;
      RECT 107.965 1.84 109.81 2.68 ;
      RECT 107.965 17.515 109.535 18.435 ;
      RECT 134.675 36.41 134.915 37.23 ;
      RECT 148.155 28.905 150.065 30.61 ;
      RECT 239.94 28.905 241.85 30.61 ;
      RECT 255.09 36.41 255.33 37.23 ;
      RECT 280.195 1.84 282.04 2.68 ;
      RECT 280.47 17.515 282.04 18.435 ;
      RECT 403.38 14.695 404.675 15.35 ;
      RECT 449.785 242.065 450.835 242.505 ;
      RECT 449.785 240.995 450.465 242.065 ;
      RECT 89.8 112.04 92.805 112.42 ;
      RECT 93.625 111.22 296.38 112.42 ;
      RECT 107.25 0 109.81 1.125 ;
      RECT 107.935 2.68 109.81 7.155 ;
      RECT 107.965 7.155 109.81 17.24 ;
      RECT 128.665 0 134.895 3.005 ;
      RECT 134.675 30.525 135.295 36.41 ;
      RECT 135.975 1.765 140.715 4.77 ;
      RECT 140.715 0 140.92 1.765 ;
      RECT 146.175 28.615 147.335 46.415 ;
      RECT 148.155 31.15 149.525 46.415 ;
      RECT 148.155 0 149.525 28.365 ;
      RECT 150.345 2.12 153.11 3.12 ;
      RECT 150.345 0 153.13 2.1 ;
      RECT 150.345 31.755 153.13 35.225 ;
      RECT 150.345 3.14 153.13 27.76 ;
      RECT 150.885 28.3 153.13 31.215 ;
      RECT 154.35 0 155.7 34.115 ;
      RECT 234.305 0 235.655 34.115 ;
      RECT 236.875 0 239.66 2.075 ;
      RECT 236.875 28.3 239.12 31.215 ;
      RECT 236.875 3.165 239.66 27.76 ;
      RECT 236.875 31.755 239.66 35.225 ;
      RECT 236.92 2.12 239.66 3.12 ;
      RECT 240.48 0 241.85 28.365 ;
      RECT 240.48 31.15 241.85 46.415 ;
      RECT 242.67 28.615 243.83 46.415 ;
      RECT 244.65 48.855 247.655 49.075 ;
      RECT 249.085 0 249.29 1.765 ;
      RECT 254.71 30.525 255.33 36.41 ;
      RECT 255.11 0 261.34 3.005 ;
      RECT 280.195 2.68 282.07 7.155 ;
      RECT 280.195 0 282.755 1.125 ;
      RECT 280.195 7.155 282.04 17.24 ;
      RECT 297.2 112.04 300.205 112.42 ;
      RECT 297.98 102.87 446.805 111.715 ;
      RECT 403.38 0 404.715 14.655 ;
      RECT 419.985 0 422.41 5.315 ;
      RECT 445.38 0 447.625 22.19 ;
      RECT 445.45 22.26 447.625 23.295 ;
      RECT 465.45 0 465.75 60.575 ;
      RECT 0 57.49 109.1 74.765 ;
      RECT 0 30.825 85.965 33.515 ;
      RECT 0 0 84.98 33.515 ;
      RECT 0 0 84.98 30.825 ;
      RECT 0 89.365 105.53 94.05 ;
      RECT 0 244.24 446.64 244.895 ;
      RECT 0 76.395 107.47 87.425 ;
      RECT 0 245.695 448.965 253.715 ;
      RECT 0 245.695 448.965 253.715 ;
      RECT 0 245.695 448.965 253.715 ;
      RECT 0 245.695 448.965 253.715 ;
      RECT 0 245.295 448.215 253.715 ;
      RECT 0 245.295 448.215 253.715 ;
      RECT 0 245.295 448.215 253.715 ;
      RECT 0 245.295 448.215 253.715 ;
      RECT 0 244.895 447.465 253.715 ;
      RECT 0 244.895 447.465 253.715 ;
      RECT 0 244.895 447.465 253.715 ;
      RECT 0 244.895 447.465 253.715 ;
      RECT 0 245.695 448.965 246.095 ;
      RECT 0 245.295 448.215 245.695 ;
      RECT 0 244.895 447.465 245.295 ;
      RECT 87.375 0 106.43 1.465 ;
      RECT 87.375 2.18 107.145 2.28 ;
      RECT 0 33.515 109.535 36.525 ;
      RECT 87.375 18.435 109.535 33.515 ;
      RECT 87.375 2.28 107.2 18.435 ;
      RECT 106.375 89.68 283.63 94.365 ;
      RECT 108.29 76.735 281.715 94.365 ;
      RECT 108.29 76.735 281.715 89.68 ;
      RECT 108.29 76.735 281.715 87.765 ;
      RECT 109.11 48.855 125.07 48.855 ;
      RECT 109.11 48.07 125.375 48.55 ;
      RECT 109.11 47.685 125.375 48.07 ;
    LAYER li1 ;
      RECT 208.065 113.91 211.065 164.9 ;
      RECT 169.92 113.91 172.92 164.9 ;
      RECT 217.085 113.91 220.085 164.9 ;
      RECT 160.9 113.91 163.9 164.9 ;
      RECT 174.43 113.91 177.43 164.9 ;
      RECT 212.575 113.91 215.575 164.9 ;
      RECT 165.41 113.91 168.41 164.9 ;
      RECT 183.45 113.91 186.45 164.9 ;
      RECT 203.555 113.91 206.555 164.9 ;
      RECT 226.105 113.91 229.105 164.9 ;
      RECT 221.595 113.91 224.595 164.9 ;
      RECT 230.615 113.91 233.615 164.9 ;
      RECT 239.635 113.91 242.635 164.9 ;
      RECT 248.655 113.91 251.655 164.9 ;
      RECT 257.675 113.91 260.675 164.9 ;
      RECT 266.695 113.91 269.695 164.9 ;
      RECT 275.715 113.91 278.715 164.9 ;
      RECT 284.735 113.91 287.735 164.9 ;
      RECT 235.125 113.91 238.125 164.9 ;
      RECT 244.145 113.91 247.145 164.9 ;
      RECT 253.165 113.91 256.165 164.9 ;
      RECT 262.185 113.91 265.185 164.9 ;
      RECT 271.205 113.91 274.205 164.9 ;
      RECT 280.225 113.91 283.225 164.9 ;
      RECT 293.755 113.91 296.755 164.9 ;
      RECT 289.245 113.91 292.245 164.9 ;
      RECT 37.485 230.175 37.655 245.125 ;
      RECT 34.965 230.175 35.135 245.125 ;
      RECT 32.445 230.175 32.615 245.125 ;
      RECT 29.925 230.175 30.095 245.125 ;
      RECT 52.09 224.125 62.09 226.445 ;
      RECT 66.16 225.16 76.16 227.48 ;
      RECT 52.09 228.735 62.09 230.645 ;
      RECT 66.16 230.445 76.16 232.185 ;
      RECT 90.025 229.425 100.025 232.185 ;
      RECT 90.025 224.125 100.025 226.46 ;
      RECT 78.08 229.425 88.08 232.185 ;
      RECT 78.08 224.125 88.08 226.46 ;
      RECT 101.735 229.425 111.735 232.185 ;
      RECT 101.735 224.125 111.735 226.46 ;
      RECT 113.445 229.425 123.445 232.185 ;
      RECT 113.445 224.125 123.445 226.46 ;
      RECT 125.155 229.425 135.155 232.185 ;
      RECT 125.155 224.125 135.155 226.46 ;
      RECT 142.24 221.465 161.95 222.075 ;
      RECT 142.24 225.365 161.95 225.975 ;
      RECT 142.24 226.925 161.95 227.535 ;
      RECT 142.24 228.485 161.95 229.095 ;
      RECT 142.24 230.045 161.95 230.655 ;
      RECT 228.055 221.465 247.765 222.075 ;
      RECT 228.055 225.365 247.765 225.975 ;
      RECT 228.055 226.925 247.765 227.535 ;
      RECT 228.055 228.485 247.765 229.095 ;
      RECT 228.055 230.045 247.765 230.655 ;
      RECT 254.85 229.425 264.85 232.185 ;
      RECT 254.85 224.125 264.85 226.46 ;
      RECT 278.27 229.425 288.27 232.185 ;
      RECT 266.56 229.425 276.56 232.185 ;
      RECT 278.27 224.125 288.27 226.46 ;
      RECT 266.56 224.125 276.56 226.46 ;
      RECT 289.98 229.425 299.98 232.185 ;
      RECT 289.98 224.125 299.98 226.46 ;
      RECT 301.925 229.425 311.925 232.185 ;
      RECT 301.925 224.125 311.925 226.46 ;
      RECT 313.845 225.16 323.845 227.48 ;
      RECT 313.845 230.445 323.845 232.185 ;
      RECT 327.915 224.125 337.915 226.445 ;
      RECT 327.915 228.735 337.915 230.645 ;
      RECT 349.52 228.345 350.27 246.62 ;
      RECT 349.52 246.62 362.855 247.375 ;
      RECT 362.105 228.345 362.855 246.62 ;
      RECT 349.52 227.595 362.855 228.345 ;
      RECT 359.13 230.095 359.3 245.125 ;
      RECT 353.13 230.095 353.3 245.125 ;
      RECT 351.57 230.095 351.74 245.125 ;
      RECT 355.65 230.095 355.82 245.125 ;
      RECT 354.09 230.095 354.26 245.125 ;
      RECT 358.17 230.095 358.34 245.125 ;
      RECT 356.61 230.095 356.78 245.125 ;
      RECT 352.35 230.175 352.52 245.125 ;
      RECT 354.87 230.175 355.04 245.125 ;
      RECT 357.39 230.175 357.56 245.125 ;
      RECT 359.91 230.175 360.08 245.125 ;
      RECT 360.69 230.095 360.86 245.125 ;
      RECT 450.77 222.01 465.61 222.18 ;
      RECT 450.77 210.765 465.61 210.935 ;
      RECT 52.09 232.935 62.09 235.255 ;
      RECT 52.09 236.415 62.09 238.735 ;
      RECT 66.16 235.15 76.16 237.91 ;
      RECT 52.09 241.7 62.09 242.935 ;
      RECT 66.16 240.875 76.16 242.11 ;
      RECT 90.025 235.15 100.025 237.91 ;
      RECT 90.025 240.875 100.025 243.21 ;
      RECT 78.08 235.15 88.08 237.91 ;
      RECT 78.08 240.875 88.08 242.11 ;
      RECT 101.735 235.15 111.735 237.91 ;
      RECT 113.445 235.15 123.445 237.91 ;
      RECT 101.735 240.875 111.735 243.21 ;
      RECT 113.445 240.875 123.445 243.21 ;
      RECT 125.155 235.15 135.155 237.91 ;
      RECT 125.155 240.875 135.155 243.21 ;
      RECT 142.24 233.665 161.95 234.16 ;
      RECT 142.24 234.33 161.95 234.825 ;
      RECT 142.24 235.775 161.95 236.27 ;
      RECT 142.24 236.465 161.95 236.96 ;
      RECT 142.24 237.91 161.95 238.405 ;
      RECT 142.24 232.22 161.95 232.715 ;
      RECT 142.24 232.885 161.965 233.495 ;
      RECT 142.24 234.995 161.95 235.605 ;
      RECT 228.055 234.33 247.765 234.825 ;
      RECT 228.055 235.775 247.765 236.27 ;
      RECT 228.055 236.465 247.765 236.96 ;
      RECT 228.055 237.91 247.765 238.405 ;
      RECT 228.055 232.22 247.765 232.715 ;
      RECT 228.055 233.665 247.765 234.16 ;
      RECT 228.04 232.885 247.765 233.495 ;
      RECT 228.055 234.995 247.765 235.605 ;
      RECT 254.85 235.15 264.85 237.91 ;
      RECT 254.85 240.875 264.85 243.21 ;
      RECT 278.27 235.15 288.27 237.91 ;
      RECT 266.56 235.15 276.56 237.91 ;
      RECT 278.27 240.875 288.27 243.21 ;
      RECT 266.56 240.875 276.56 243.21 ;
      RECT 289.98 235.15 299.98 237.91 ;
      RECT 289.98 240.875 299.98 243.21 ;
      RECT 301.925 235.15 311.925 237.91 ;
      RECT 301.925 240.875 311.925 242.11 ;
      RECT 313.845 235.15 323.845 237.91 ;
      RECT 313.845 240.875 323.845 242.11 ;
      RECT 327.915 232.935 337.915 235.255 ;
      RECT 327.915 236.415 337.915 238.735 ;
      RECT 327.915 241.7 337.915 242.935 ;
      RECT 450.77 233.27 465.61 233.44 ;
      RECT 37.01 54.98 62.41 55.15 ;
      RECT 327.595 54.98 352.995 55.15 ;
      RECT 448.34 146.92 448.51 181.625 ;
      RECT 420.815 236.82 449.625 237.07 ;
      RECT 93.25 113.91 96.25 164.9 ;
      RECT 156.39 113.91 159.39 164.9 ;
      RECT 147.37 113.91 150.37 164.9 ;
      RECT 138.35 113.91 141.35 164.9 ;
      RECT 129.33 113.91 132.33 164.9 ;
      RECT 120.31 113.91 123.31 164.9 ;
      RECT 111.29 113.91 114.29 164.9 ;
      RECT 102.27 113.91 105.27 164.9 ;
      RECT 151.88 113.91 154.88 164.9 ;
      RECT 142.86 113.91 145.86 164.9 ;
      RECT 133.84 113.91 136.84 164.9 ;
      RECT 124.82 113.91 127.82 164.9 ;
      RECT 115.8 113.91 118.8 164.9 ;
      RECT 106.78 113.91 109.78 164.9 ;
      RECT 97.76 113.91 100.76 164.9 ;
      RECT 178.94 113.91 181.94 164.9 ;
      RECT 310.63 186.19 325.66 186.36 ;
      RECT 310.63 186.97 325.66 187.14 ;
      RECT 326.425 186.19 341.375 186.36 ;
      RECT 326.425 186.97 341.375 187.14 ;
      RECT 314.925 172.105 324.925 174.82 ;
      RECT 20.865 193.48 28.865 193.65 ;
      RECT 48.63 189.67 63.58 189.84 ;
      RECT 48.63 190.45 63.58 190.62 ;
      RECT 48.63 187.93 63.58 188.1 ;
      RECT 48.63 188.71 63.58 188.88 ;
      RECT 48.63 191.41 63.58 191.58 ;
      RECT 48.63 192.19 63.58 192.36 ;
      RECT 64.345 192.19 79.375 192.36 ;
      RECT 64.345 187.93 79.295 188.1 ;
      RECT 64.345 188.71 79.375 188.88 ;
      RECT 64.345 189.67 79.295 189.84 ;
      RECT 64.345 190.45 79.375 190.62 ;
      RECT 64.345 191.41 79.295 191.58 ;
      RECT 86.46 200.495 86.99 215.995 ;
      RECT 90.58 200.495 91.11 215.995 ;
      RECT 82.04 217.365 157.33 218.215 ;
      RECT 82.04 198.275 157.33 199.125 ;
      RECT 82.04 199.125 85.95 217.365 ;
      RECT 153.42 199.125 157.33 217.365 ;
      RECT 88.52 200.495 89.05 215.995 ;
      RECT 94.7 200.495 95.23 215.995 ;
      RECT 98.82 200.495 99.35 215.995 ;
      RECT 92.64 200.495 93.17 215.995 ;
      RECT 96.76 200.495 97.29 215.995 ;
      RECT 100.88 200.495 101.41 215.995 ;
      RECT 105 200.495 105.53 215.995 ;
      RECT 109.12 200.495 109.65 215.995 ;
      RECT 113.24 200.495 113.77 215.995 ;
      RECT 102.94 200.495 103.47 215.995 ;
      RECT 107.06 200.495 107.59 215.995 ;
      RECT 111.18 200.495 111.71 215.995 ;
      RECT 117.36 200.495 117.89 215.995 ;
      RECT 121.48 200.495 122.01 215.995 ;
      RECT 125.6 200.495 126.13 215.995 ;
      RECT 129.72 200.495 130.25 215.995 ;
      RECT 133.84 200.495 134.37 215.995 ;
      RECT 115.3 200.495 115.83 215.995 ;
      RECT 119.42 200.495 119.95 215.995 ;
      RECT 123.54 200.495 124.07 215.995 ;
      RECT 127.66 200.495 128.19 215.995 ;
      RECT 131.78 200.495 132.31 215.995 ;
      RECT 146.2 200.495 146.73 215.995 ;
      RECT 150.32 200.495 150.85 215.995 ;
      RECT 137.96 200.495 138.49 215.995 ;
      RECT 142.08 200.495 142.61 215.995 ;
      RECT 152.38 200.495 152.91 215.995 ;
      RECT 135.9 200.495 136.43 215.995 ;
      RECT 140.02 200.495 140.55 215.995 ;
      RECT 144.14 200.495 144.67 215.995 ;
      RECT 148.26 200.495 148.79 215.995 ;
      RECT 165.55 207.38 165.72 217.23 ;
      RECT 168.67 207.38 168.84 217.23 ;
      RECT 166.33 207.38 166.5 217.23 ;
      RECT 167.11 207.38 167.28 217.23 ;
      RECT 167.89 207.38 168.06 217.23 ;
      RECT 224.285 207.38 224.455 217.23 ;
      RECT 221.165 207.38 221.335 217.23 ;
      RECT 239.155 200.495 239.685 215.995 ;
      RECT 232.675 217.365 307.965 218.215 ;
      RECT 232.675 198.275 307.965 199.125 ;
      RECT 232.675 199.125 236.585 217.365 ;
      RECT 304.055 199.125 307.965 217.365 ;
      RECT 237.095 200.495 237.625 215.995 ;
      RECT 241.215 200.495 241.745 215.995 ;
      RECT 223.505 207.38 223.675 217.23 ;
      RECT 222.725 207.38 222.895 217.23 ;
      RECT 221.945 207.38 222.115 217.23 ;
      RECT 243.275 200.495 243.805 215.995 ;
      RECT 259.755 200.495 260.285 215.995 ;
      RECT 255.635 200.495 256.165 215.995 ;
      RECT 251.515 200.495 252.045 215.995 ;
      RECT 247.395 200.495 247.925 215.995 ;
      RECT 261.815 200.495 262.345 215.995 ;
      RECT 257.695 200.495 258.225 215.995 ;
      RECT 253.575 200.495 254.105 215.995 ;
      RECT 249.455 200.495 249.985 215.995 ;
      RECT 245.335 200.495 245.865 215.995 ;
      RECT 284.475 200.495 285.005 215.995 ;
      RECT 280.355 200.495 280.885 215.995 ;
      RECT 276.235 200.495 276.765 215.995 ;
      RECT 272.115 200.495 272.645 215.995 ;
      RECT 267.995 200.495 268.525 215.995 ;
      RECT 263.875 200.495 264.405 215.995 ;
      RECT 282.415 200.495 282.945 215.995 ;
      RECT 278.295 200.495 278.825 215.995 ;
      RECT 274.175 200.495 274.705 215.995 ;
      RECT 270.055 200.495 270.585 215.995 ;
      RECT 265.935 200.495 266.465 215.995 ;
      RECT 303.015 200.495 303.545 215.995 ;
      RECT 298.895 200.495 299.425 215.995 ;
      RECT 294.775 200.495 295.305 215.995 ;
      RECT 290.655 200.495 291.185 215.995 ;
      RECT 300.955 200.495 301.485 215.995 ;
      RECT 296.835 200.495 297.365 215.995 ;
      RECT 292.715 200.495 293.245 215.995 ;
      RECT 288.595 200.495 289.125 215.995 ;
      RECT 286.535 200.495 287.065 215.995 ;
      RECT 326.425 191.41 341.375 191.58 ;
      RECT 326.425 192.19 341.375 192.36 ;
      RECT 310.71 189.67 325.66 189.84 ;
      RECT 310.63 190.45 325.66 190.62 ;
      RECT 310.71 191.41 325.66 191.58 ;
      RECT 310.63 192.19 325.66 192.36 ;
      RECT 310.71 187.93 325.66 188.1 ;
      RECT 310.63 188.71 325.66 188.88 ;
      RECT 326.425 189.67 341.375 189.84 ;
      RECT 326.425 190.45 341.375 190.62 ;
      RECT 326.425 187.93 341.375 188.1 ;
      RECT 326.425 188.71 341.375 188.88 ;
      RECT 361.14 193.48 369.14 193.65 ;
      RECT 27.15 246.62 40.485 247.375 ;
      RECT 39.735 228.345 40.485 246.62 ;
      RECT 27.15 227.595 40.485 228.345 ;
      RECT 27.15 228.345 27.9 246.62 ;
      RECT 29.145 230.095 29.315 245.125 ;
      RECT 30.705 230.095 30.875 245.125 ;
      RECT 36.705 230.095 36.875 245.125 ;
      RECT 38.265 230.095 38.435 245.125 ;
      RECT 34.185 230.095 34.355 245.125 ;
      RECT 35.745 230.095 35.915 245.125 ;
      RECT 31.665 230.095 31.835 245.125 ;
      RECT 33.225 230.095 33.395 245.125 ;
      RECT 298.63 64.425 305.885 64.435 ;
      RECT 319.73 58.795 319.9 68.685 ;
      RECT 318.55 58.795 318.72 68.685 ;
      RECT 316.19 58.795 316.36 68.685 ;
      RECT 315.01 58.795 315.18 68.685 ;
      RECT 317.37 58.795 317.54 68.685 ;
      RECT 346.18 59.435 354.46 59.605 ;
      RECT 346.315 59.39 354.4 59.435 ;
      RECT 398.74 64.77 398.91 74.66 ;
      RECT 407.3 64.77 407.47 74.66 ;
      RECT 398.74 75.84 398.91 85.73 ;
      RECT 407.3 75.84 407.47 85.73 ;
      RECT 412.9 75.84 413.07 85.73 ;
      RECT 412.9 64.77 413.07 74.66 ;
      RECT 411.58 64.77 411.75 74.66 ;
      RECT 411.58 75.84 411.75 85.73 ;
      RECT 403.02 64.77 403.19 74.66 ;
      RECT 403.02 75.84 403.19 85.73 ;
      RECT 417.18 75.84 417.35 85.73 ;
      RECT 417.18 64.77 417.35 74.66 ;
      RECT 424.02 75.84 424.19 85.73 ;
      RECT 424.02 64.77 424.19 74.66 ;
      RECT 421.74 75.84 421.91 85.73 ;
      RECT 419.46 75.84 419.63 85.73 ;
      RECT 421.74 64.77 421.91 74.66 ;
      RECT 419.46 64.77 419.63 74.66 ;
      RECT 19.555 87.175 27.555 87.345 ;
      RECT 19.555 94.825 27.555 94.995 ;
      RECT 19.7 87.345 27.44 94.825 ;
      RECT 362.45 87.175 370.45 87.345 ;
      RECT 362.45 94.825 370.45 94.995 ;
      RECT 362.565 87.345 370.305 94.825 ;
      RECT 398.74 98.035 398.91 107.925 ;
      RECT 407.3 98.035 407.47 107.925 ;
      RECT 398.74 86.965 398.91 96.855 ;
      RECT 407.3 86.965 407.47 96.855 ;
      RECT 412.9 98.035 413.07 107.925 ;
      RECT 411.58 86.965 411.75 96.855 ;
      RECT 412.9 86.965 413.07 96.855 ;
      RECT 411.58 98.035 411.75 107.925 ;
      RECT 403.02 98.035 403.19 107.925 ;
      RECT 403.02 86.965 403.19 96.855 ;
      RECT 417.18 98.035 417.35 107.925 ;
      RECT 417.18 86.965 417.35 96.855 ;
      RECT 424.02 86.965 424.19 96.855 ;
      RECT 424.02 98.035 424.19 107.925 ;
      RECT 421.74 86.965 421.91 96.855 ;
      RECT 419.46 86.965 419.63 96.855 ;
      RECT 421.74 98.035 421.91 107.925 ;
      RECT 419.46 98.035 419.63 107.925 ;
      RECT 19.555 117.195 27.555 117.365 ;
      RECT 19.555 124.845 27.555 125.015 ;
      RECT 19.7 117.365 27.44 124.845 ;
      RECT 362.45 117.195 370.45 117.365 ;
      RECT 362.45 124.845 370.45 125.015 ;
      RECT 362.565 117.365 370.305 124.845 ;
      RECT 401.71 110.765 401.88 120.655 ;
      RECT 399.35 110.765 399.52 120.655 ;
      RECT 406.43 110.765 406.6 120.655 ;
      RECT 404.07 110.765 404.24 120.655 ;
      RECT 409.49 110.765 409.66 120.655 ;
      RECT 411.85 110.765 412.02 120.655 ;
      RECT 408.9 109.66 417.33 109.84 ;
      RECT 398.765 109.66 407.19 109.84 ;
      RECT 408.9 110.605 409.08 120.97 ;
      RECT 407.01 110.605 407.19 120.97 ;
      RECT 407.015 110.405 407.185 110.605 ;
      RECT 398.76 110.605 398.94 120.97 ;
      RECT 398.765 110.405 398.935 110.605 ;
      RECT 414.21 110.765 414.38 120.655 ;
      RECT 416.57 110.765 416.74 120.655 ;
      RECT 417.15 110.605 417.33 120.97 ;
      RECT 19.915 133.415 26.675 133.585 ;
      RECT 19.915 133.405 26.615 133.415 ;
      RECT 34.25 142.27 47.84 142.44 ;
      RECT 38.585 132.01 38.755 141.97 ;
      RECT 36.305 132.01 36.475 141.86 ;
      RECT 40.865 132.01 41.035 141.86 ;
      RECT 43.145 132.01 43.315 141.97 ;
      RECT 47.705 132.01 47.875 141.97 ;
      RECT 45.425 132.01 45.595 141.86 ;
      RECT 34.025 132.01 34.195 141.97 ;
      RECT 342.165 142.27 355.755 142.44 ;
      RECT 348.97 132.01 349.14 141.86 ;
      RECT 346.69 132.01 346.86 141.97 ;
      RECT 342.13 132.01 342.3 141.97 ;
      RECT 344.41 132.01 344.58 141.86 ;
      RECT 351.25 132.01 351.42 141.97 ;
      RECT 353.53 132.01 353.7 141.86 ;
      RECT 355.81 132.01 355.98 141.97 ;
      RECT 363.33 133.415 370.09 133.585 ;
      RECT 363.39 133.405 370.09 133.415 ;
      RECT 22.62 148.07 34.85 148.24 ;
      RECT 28.885 155.27 34.995 155.44 ;
      RECT 64.375 146.75 64.545 156.6 ;
      RECT 54.445 147.505 54.615 157.355 ;
      RECT 53.265 147.505 53.435 157.355 ;
      RECT 52.715 147.505 52.885 157.355 ;
      RECT 51.535 147.505 51.705 157.355 ;
      RECT 68.655 146.75 68.825 156.6 ;
      RECT 65.08 162.48 75.08 165.195 ;
      RECT 77.215 146.75 77.385 156.6 ;
      RECT 81.495 146.75 81.665 156.6 ;
      RECT 72.935 146.75 73.105 156.6 ;
      RECT 85.775 146.75 85.945 156.6 ;
      RECT 76.72 162.48 86.72 165.195 ;
      RECT 304.06 146.75 304.23 156.6 ;
      RECT 303.285 162.48 313.285 165.195 ;
      RECT 325.46 146.75 325.63 156.6 ;
      RECT 312.62 146.75 312.79 156.6 ;
      RECT 308.34 146.75 308.51 156.6 ;
      RECT 321.18 146.75 321.35 156.6 ;
      RECT 316.9 146.75 317.07 156.6 ;
      RECT 314.925 162.48 324.925 165.195 ;
      RECT 335.39 147.505 335.56 157.355 ;
      RECT 336.57 147.505 336.74 157.355 ;
      RECT 337.12 147.505 337.29 157.355 ;
      RECT 338.3 147.505 338.47 157.355 ;
      RECT 355.01 155.27 361.12 155.44 ;
      RECT 355.155 148.07 367.385 148.24 ;
      RECT 48.63 186.19 63.58 186.36 ;
      RECT 48.63 186.97 63.58 187.14 ;
      RECT 64.345 186.19 79.375 186.36 ;
      RECT 64.345 186.97 79.375 187.14 ;
      RECT 65.08 172.105 75.08 174.82 ;
      RECT 76.72 172.105 86.72 174.82 ;
      RECT 303.285 172.105 313.285 174.82 ;
      RECT 458.9 249.43 459.07 252.14 ;
      RECT 462.4 248.71 464.085 248.88 ;
      RECT 461.47 249.25 461.72 249.37 ;
      RECT 460.66 249.37 462.55 252.14 ;
      RECT 463.26 249.43 463.43 252.14 ;
      RECT 464.14 249.43 464.31 252.14 ;
      RECT 420.63 252.495 465.16 253.385 ;
      RECT 420.63 250.89 454.055 252.495 ;
      RECT 464.72 247.445 465.16 252.495 ;
      RECT 449.985 244.735 467.055 246.035 ;
      RECT 466.045 246.035 467.055 253.445 ;
      RECT 13.59 4.675 13.76 14.525 ;
      RECT 12.41 4.675 12.58 14.565 ;
      RECT 48.5 11.525 58.39 11.695 ;
      RECT 59.84 11.525 69.73 11.695 ;
      RECT 320.275 11.525 330.165 11.695 ;
      RECT 331.615 11.525 341.505 11.695 ;
      RECT 376.245 4.675 376.415 14.525 ;
      RECT 377.425 4.675 377.595 14.565 ;
      RECT 45.385 17.34 45.555 27.19 ;
      RECT 46.565 17.34 46.735 27.19 ;
      RECT 44.205 17.34 44.375 27.19 ;
      RECT 48.5 19.295 58.39 19.465 ;
      RECT 48.5 20.475 58.39 20.645 ;
      RECT 48.5 17.495 58.39 17.665 ;
      RECT 48.5 18.675 58.39 18.845 ;
      RECT 48.5 14.505 58.39 14.675 ;
      RECT 48.5 13.325 58.39 13.495 ;
      RECT 48.5 15.685 58.39 15.855 ;
      RECT 48.5 16.315 58.39 16.485 ;
      RECT 48.5 12.705 58.39 12.875 ;
      RECT 28.52 32.335 38.41 32.505 ;
      RECT 28.52 31.155 38.41 31.325 ;
      RECT 40.11 32.335 50 32.505 ;
      RECT 40.11 31.155 50 31.325 ;
      RECT 28.52 33.515 38.41 33.685 ;
      RECT 40.11 33.515 50 33.685 ;
      RECT 59.84 12.705 69.73 12.875 ;
      RECT 59.84 19.295 69.73 19.465 ;
      RECT 59.84 20.475 69.73 20.645 ;
      RECT 59.84 17.495 69.73 17.665 ;
      RECT 59.84 16.315 69.73 16.485 ;
      RECT 59.84 14.505 69.73 14.675 ;
      RECT 59.84 15.685 69.73 15.855 ;
      RECT 59.84 18.675 69.73 18.845 ;
      RECT 59.84 13.325 69.73 13.495 ;
      RECT 137.165 26.945 144.19 27.115 ;
      RECT 245.815 26.945 252.84 27.115 ;
      RECT 320.275 12.705 330.165 12.875 ;
      RECT 320.275 19.295 330.165 19.465 ;
      RECT 320.275 20.475 330.165 20.645 ;
      RECT 320.275 17.495 330.165 17.665 ;
      RECT 320.275 16.315 330.165 16.485 ;
      RECT 320.275 14.505 330.165 14.675 ;
      RECT 320.275 15.685 330.165 15.855 ;
      RECT 320.275 18.675 330.165 18.845 ;
      RECT 320.275 13.325 330.165 13.495 ;
      RECT 344.45 17.34 344.62 27.19 ;
      RECT 343.27 17.34 343.44 27.19 ;
      RECT 345.63 17.34 345.8 27.19 ;
      RECT 331.615 12.705 341.505 12.875 ;
      RECT 331.615 19.295 341.505 19.465 ;
      RECT 331.615 20.475 341.505 20.645 ;
      RECT 331.615 17.495 341.505 17.665 ;
      RECT 331.615 18.675 341.505 18.845 ;
      RECT 331.615 14.505 341.505 14.675 ;
      RECT 331.615 13.325 341.505 13.495 ;
      RECT 331.615 15.685 341.505 15.855 ;
      RECT 331.615 16.315 341.505 16.485 ;
      RECT 340.005 32.335 349.895 32.505 ;
      RECT 340.005 31.155 349.895 31.325 ;
      RECT 340.005 33.515 349.895 33.685 ;
      RECT 351.595 32.335 361.485 32.505 ;
      RECT 351.595 31.155 361.485 31.325 ;
      RECT 351.595 33.515 361.485 33.685 ;
      RECT 21.07 42.415 21.24 52.305 ;
      RECT 23.43 42.415 23.6 52.305 ;
      RECT 16.43 42.415 16.6 52.305 ;
      RECT 45.59 50.56 62.41 50.73 ;
      RECT 45.63 50.53 62.355 50.56 ;
      RECT 28.52 35.875 38.41 36.045 ;
      RECT 28.52 34.695 38.41 34.865 ;
      RECT 40.11 35.875 50 36.045 ;
      RECT 40.11 34.695 50 34.865 ;
      RECT 81.015 50.44 89 50.61 ;
      RECT 81.225 50.61 88.955 50.665 ;
      RECT 72.48 50.44 79.05 50.61 ;
      RECT 72.62 50.61 78.91 50.665 ;
      RECT 144.795 50.33 153.885 59.67 ;
      RECT 236.12 50.33 245.21 59.67 ;
      RECT 301.005 50.44 308.99 50.61 ;
      RECT 301.05 50.61 308.78 50.665 ;
      RECT 310.955 50.44 317.525 50.61 ;
      RECT 311.095 50.61 317.385 50.665 ;
      RECT 327.595 50.56 344.415 50.73 ;
      RECT 327.65 50.53 344.375 50.56 ;
      RECT 340.005 35.875 349.895 36.045 ;
      RECT 340.005 34.695 349.895 34.865 ;
      RECT 351.595 35.875 361.485 36.045 ;
      RECT 351.595 34.695 361.485 34.865 ;
      RECT 368.765 42.415 368.935 52.305 ;
      RECT 366.405 42.415 366.575 52.305 ;
      RECT 373.405 42.415 373.575 52.305 ;
      RECT 408.62 51.38 408.79 61.23 ;
      RECT 408.62 40.92 408.79 50.77 ;
      RECT 398.74 40.92 398.91 50.77 ;
      RECT 407.3 40.92 407.47 50.77 ;
      RECT 398.74 51.38 398.91 61.23 ;
      RECT 407.3 51.38 407.47 61.23 ;
      RECT 412.9 51.38 413.07 61.23 ;
      RECT 403.02 40.92 403.19 50.77 ;
      RECT 412.9 40.92 413.07 50.77 ;
      RECT 403.02 51.38 403.19 61.23 ;
      RECT 417.18 51.38 417.35 61.23 ;
      RECT 417.18 40.92 417.35 50.77 ;
      RECT 35.545 59.435 43.825 59.605 ;
      RECT 35.605 59.39 43.69 59.435 ;
      RECT 70.105 58.795 70.275 68.685 ;
      RECT 71.285 58.795 71.455 68.685 ;
      RECT 73.645 58.795 73.815 68.685 ;
      RECT 74.825 58.795 74.995 68.685 ;
      RECT 72.465 58.795 72.635 68.685 ;
      RECT 82.175 64.435 92.135 64.605 ;
      RECT 84.12 64.425 91.375 64.435 ;
      RECT 160.59 74.745 168.4 74.915 ;
      RECT 221.605 74.745 229.415 74.915 ;
      RECT 297.87 64.435 307.83 64.605 ;
      RECT 407.94 249.475 408.55 252.915 ;
      RECT 412.615 249.475 413.225 252.915 ;
      RECT 390.24 249.565 391.17 252.425 ;
      RECT 387.345 248.775 387.735 252.275 ;
      RECT 387.345 248.605 387.875 248.775 ;
      RECT 389.245 248.605 389.775 248.775 ;
      RECT 389.365 247.065 389.645 248.605 ;
      RECT 389.83 246.775 390.095 248.075 ;
      RECT 388.785 246.265 391.15 246.775 ;
      RECT 388.92 246.775 389.185 248.075 ;
      RECT 390.745 246.775 391.01 248.075 ;
      RECT 390.34 247.065 390.51 248.075 ;
      RECT 387.41 245.925 388.08 248.415 ;
      RECT 388.905 248.995 390.285 249.165 ;
      RECT 393.46 246.265 395.825 246.775 ;
      RECT 394.505 246.775 394.77 248.075 ;
      RECT 393.595 246.775 393.86 248.075 ;
      RECT 395.42 246.775 395.685 248.075 ;
      RECT 390.735 248.605 391.405 248.775 ;
      RECT 391.585 247.405 391.84 249.565 ;
      RECT 391.46 249.565 391.84 252.275 ;
      RECT 392.02 248.775 392.41 252.275 ;
      RECT 392.02 248.605 392.55 248.775 ;
      RECT 392.595 249.565 393.525 252.425 ;
      RECT 393.92 248.605 394.45 248.775 ;
      RECT 394.04 247.065 394.32 248.605 ;
      RECT 393.58 248.995 394.96 249.165 ;
      RECT 394.915 249.565 395.845 252.425 ;
      RECT 396.26 247.405 396.515 249.565 ;
      RECT 396.135 249.565 396.515 252.275 ;
      RECT 395.015 247.065 395.185 248.075 ;
      RECT 395.41 248.605 396.08 248.775 ;
      RECT 398.135 246.265 400.5 246.775 ;
      RECT 398.27 246.775 398.535 248.075 ;
      RECT 399.18 246.775 399.445 248.075 ;
      RECT 400.095 246.775 400.36 248.075 ;
      RECT 396.695 248.775 397.085 252.275 ;
      RECT 396.695 248.605 397.225 248.775 ;
      RECT 397.27 249.565 398.2 252.425 ;
      RECT 398.595 248.605 399.125 248.775 ;
      RECT 398.715 247.065 398.995 248.605 ;
      RECT 398.255 248.995 399.635 249.165 ;
      RECT 399.59 249.565 400.52 252.425 ;
      RECT 400.935 247.405 401.19 249.565 ;
      RECT 400.81 249.565 401.19 252.275 ;
      RECT 399.69 247.065 399.86 248.075 ;
      RECT 400.085 248.605 400.755 248.775 ;
      RECT 401.37 248.775 401.76 252.275 ;
      RECT 401.37 248.605 401.9 248.775 ;
      RECT 401.945 249.565 402.875 252.425 ;
      RECT 402.81 246.265 405.175 246.775 ;
      RECT 402.945 246.775 403.21 248.075 ;
      RECT 403.855 246.775 404.12 248.075 ;
      RECT 404.77 246.775 405.035 248.075 ;
      RECT 407.485 246.265 409.85 246.775 ;
      RECT 407.62 246.775 407.885 248.075 ;
      RECT 408.53 246.775 408.795 248.075 ;
      RECT 409.445 246.775 409.71 248.075 ;
      RECT 402.93 248.995 404.31 249.165 ;
      RECT 403.27 248.605 403.8 248.775 ;
      RECT 403.39 247.065 403.67 248.605 ;
      RECT 404.265 249.565 405.195 252.425 ;
      RECT 405.61 247.405 405.865 249.565 ;
      RECT 405.485 249.565 405.865 252.275 ;
      RECT 404.365 247.065 404.535 248.075 ;
      RECT 404.76 248.605 405.43 248.775 ;
      RECT 406.62 249.565 407.55 252.425 ;
      RECT 406.045 248.775 406.435 252.275 ;
      RECT 406.045 248.605 406.575 248.775 ;
      RECT 407.605 248.995 408.985 249.165 ;
      RECT 407.945 248.605 408.475 248.775 ;
      RECT 408.065 247.065 408.345 248.605 ;
      RECT 412.16 246.265 414.525 246.775 ;
      RECT 412.295 246.775 412.56 248.075 ;
      RECT 413.205 246.775 413.47 248.075 ;
      RECT 414.12 246.775 414.385 248.075 ;
      RECT 408.94 249.565 409.87 252.425 ;
      RECT 410.285 247.405 410.54 249.565 ;
      RECT 410.16 249.565 410.54 252.275 ;
      RECT 409.04 247.065 409.21 248.075 ;
      RECT 409.435 248.605 410.105 248.775 ;
      RECT 410.72 248.775 411.11 252.275 ;
      RECT 410.72 248.605 411.25 248.775 ;
      RECT 411.295 249.565 412.225 252.425 ;
      RECT 412.62 248.605 413.15 248.775 ;
      RECT 412.74 247.065 413.02 248.605 ;
      RECT 412.28 248.995 413.66 249.165 ;
      RECT 413.615 249.565 414.545 252.425 ;
      RECT 413.715 247.065 413.885 248.075 ;
      RECT 414.96 247.405 415.215 249.565 ;
      RECT 414.835 249.565 415.215 252.275 ;
      RECT 414.11 248.605 414.78 248.775 ;
      RECT 422.25 247.19 422.42 249.9 ;
      RECT 420.75 247.19 420.92 249.9 ;
      RECT 423.75 247.19 423.92 249.9 ;
      RECT 426.13 247.19 426.3 249.9 ;
      RECT 430.01 247.19 430.18 249.9 ;
      RECT 429.39 247.19 429.56 249.9 ;
      RECT 425.51 247.19 425.68 249.9 ;
      RECT 427.63 247.19 427.8 249.9 ;
      RECT 435.39 247.19 435.56 249.9 ;
      RECT 433.01 247.19 433.18 249.9 ;
      RECT 434.77 247.19 434.94 249.9 ;
      RECT 436.89 247.19 437.06 249.9 ;
      RECT 439.27 247.19 439.44 249.9 ;
      RECT 438.65 247.19 438.82 249.9 ;
      RECT 442.275 247.19 442.445 249.9 ;
      RECT 448.535 247.19 448.705 249.9 ;
      RECT 447.915 247.19 448.085 249.9 ;
      RECT 446.155 247.19 446.325 249.9 ;
      RECT 444.655 247.19 444.825 249.9 ;
      RECT 444.035 247.19 444.205 249.9 ;
      RECT 443.155 238.04 443.325 250.205 ;
      RECT 452.085 247.25 452.255 250.23 ;
      RECT 450.325 247.25 450.495 250.23 ;
      RECT 452.965 247.52 453.135 250.23 ;
      RECT 450.55 246.265 461.585 246.97 ;
      RECT 453.845 247.25 454.015 250.23 ;
      RECT 451.205 247.52 451.375 250.23 ;
      RECT 456.325 250.7 456.86 251.38 ;
      RECT 454.91 251.38 456.86 251.73 ;
      RECT 455.635 250.665 455.805 251.195 ;
      RECT 454.6 250.48 455.055 251.03 ;
      RECT 454.6 250.31 456.53 250.48 ;
      RECT 458.905 248.71 460.605 248.88 ;
      RECT 457.085 250.78 458.5 251.08 ;
      RECT 459.78 249.43 459.95 252.14 ;
      RECT 247.945 244.345 248.695 246.365 ;
      RECT 388.42 241.395 388.59 244.105 ;
      RECT 389.3 241.335 390.62 244.105 ;
      RECT 388.615 244.325 389.285 244.495 ;
      RECT 392.18 243.835 392.85 244.495 ;
      RECT 392.18 241.215 392.85 241.295 ;
      RECT 390.825 241.215 391.13 243.905 ;
      RECT 390.65 240.675 392.85 240.845 ;
      RECT 390.825 240.845 392.85 241.215 ;
      RECT 391.33 241.395 391.5 244.105 ;
      RECT 392.18 241.905 392.91 243.225 ;
      RECT 394.9 243.845 395.57 245.095 ;
      RECT 392.085 245.095 395.57 245.765 ;
      RECT 392.085 245.765 392.755 248.415 ;
      RECT 393.19 243.59 393.36 243.86 ;
      RECT 392.76 243.42 393.36 243.59 ;
      RECT 393.19 243.19 393.36 243.42 ;
      RECT 396.86 241.765 397.03 241.93 ;
      RECT 396.01 241.595 397.03 241.765 ;
      RECT 396.86 241.26 397.03 241.595 ;
      RECT 396.01 241.765 396.66 244.495 ;
      RECT 393.19 241.765 393.36 241.93 ;
      RECT 393.19 241.595 394.21 241.765 ;
      RECT 393.19 241.26 393.36 241.595 ;
      RECT 393.56 241.765 394.21 244.495 ;
      RECT 397.37 243.835 398.04 244.495 ;
      RECT 397.37 241.215 398.04 241.295 ;
      RECT 399.09 241.215 399.395 243.905 ;
      RECT 397.37 240.675 399.57 240.845 ;
      RECT 397.37 240.845 399.395 241.215 ;
      RECT 398.72 241.395 398.89 244.105 ;
      RECT 401.63 241.395 401.8 244.105 ;
      RECT 397.31 241.905 398.04 243.225 ;
      RECT 399.6 241.335 400.92 244.105 ;
      RECT 401.435 244.695 402.105 248.415 ;
      RECT 396.76 244.71 397.43 248.415 ;
      RECT 396.86 243.59 397.03 243.86 ;
      RECT 396.86 243.42 397.46 243.59 ;
      RECT 396.86 243.19 397.03 243.42 ;
      RECT 400.935 244.325 401.605 244.495 ;
      RECT 406.33 241.395 406.5 244.105 ;
      RECT 407.21 241.335 408.53 244.105 ;
      RECT 406.11 245.11 406.78 248.415 ;
      RECT 406.525 244.325 407.195 244.495 ;
      RECT 410.09 243.835 410.76 244.495 ;
      RECT 410.09 241.215 410.76 241.295 ;
      RECT 408.735 241.215 409.04 243.905 ;
      RECT 408.56 240.675 410.76 240.845 ;
      RECT 408.735 240.845 410.76 241.215 ;
      RECT 409.24 241.395 409.41 244.105 ;
      RECT 410.09 241.905 410.82 243.225 ;
      RECT 410.785 245.51 411.455 248.415 ;
      RECT 412.98 241.695 418.055 244.245 ;
      RECT 416.4 244.245 418.055 244.73 ;
      RECT 416.4 244.77 420.665 245.98 ;
      RECT 416.4 245.98 419.855 246.265 ;
      RECT 416.4 244.73 419.855 244.77 ;
      RECT 416.965 246.265 419.855 253.125 ;
      RECT 411.1 243.59 411.27 243.86 ;
      RECT 410.67 243.42 411.27 243.59 ;
      RECT 411.1 243.19 411.27 243.42 ;
      RECT 411.1 241.765 411.27 241.93 ;
      RECT 411.1 241.595 412.12 241.765 ;
      RECT 411.1 241.26 411.27 241.595 ;
      RECT 411.47 241.765 412.12 244.495 ;
      RECT 420.75 237.915 420.92 238.965 ;
      RECT 422.25 237.915 422.42 238.965 ;
      RECT 423.75 237.915 423.92 238.98 ;
      RECT 424.63 238.04 424.8 250.205 ;
      RECT 426.13 237.915 426.3 238.965 ;
      RECT 427.63 237.915 427.8 238.98 ;
      RECT 430.01 237.915 430.18 238.965 ;
      RECT 427.01 237.915 427.18 250.22 ;
      RECT 428.51 238.04 428.68 250.205 ;
      RECT 435.39 237.915 435.56 238.965 ;
      RECT 436.89 237.915 437.06 238.98 ;
      RECT 433.01 237.915 433.18 238.98 ;
      RECT 436.27 237.915 436.44 250.205 ;
      RECT 433.89 238.04 434.06 250.205 ;
      RECT 439.27 237.915 439.44 238.965 ;
      RECT 442.275 237.915 442.445 238.98 ;
      RECT 437.77 238.04 437.94 250.205 ;
      RECT 448.535 237.915 448.705 238.965 ;
      RECT 445.535 239.235 446.065 239.405 ;
      RECT 445.535 239.405 445.705 250.205 ;
      RECT 445.535 237.915 445.705 239.235 ;
      RECT 444.655 237.915 444.825 238.965 ;
      RECT 446.155 237.915 446.325 238.98 ;
      RECT 447.035 238.04 447.205 250.205 ;
      RECT 449.415 237.915 449.585 250.205 ;
      RECT 451.06 240.3 452.66 240.47 ;
      RECT 451.835 240.72 452.005 241.73 ;
      RECT 451.835 237.935 452.005 239.21 ;
      RECT 451.15 237.965 451.32 238.975 ;
      RECT 450.27 238.075 450.445 238.965 ;
      RECT 450.27 238.965 450.44 238.975 ;
      RECT 450.27 237.965 450.44 238.075 ;
      RECT 459.275 239.45 459.945 239.62 ;
      RECT 457.06 241.45 463.32 241.62 ;
      RECT 457.24 239.45 457.91 239.62 ;
      RECT 456.965 241.81 465.08 241.995 ;
      RECT 456.965 241.995 457.495 242.085 ;
      RECT 463.6 241.45 465.08 241.81 ;
      RECT 454.42 240.3 456.14 240.47 ;
      RECT 456.03 237.935 456.2 238.945 ;
      RECT 455.315 240.72 455.485 241.73 ;
      RECT 169.25 246.125 171.96 246.295 ;
      RECT 169.25 247.685 171.96 247.855 ;
      RECT 169.25 248.235 171.96 248.405 ;
      RECT 169.25 249.795 171.96 249.965 ;
      RECT 169.25 249.015 171.96 249.185 ;
      RECT 169.25 246.905 171.96 247.075 ;
      RECT 172.15 246.35 172.32 249.82 ;
      RECT 218.045 246.125 220.755 246.295 ;
      RECT 218.045 247.685 220.755 247.855 ;
      RECT 218.045 248.235 220.755 248.405 ;
      RECT 218.045 249.795 220.755 249.965 ;
      RECT 217.685 246.35 217.855 249.82 ;
      RECT 218.045 249.015 220.755 249.185 ;
      RECT 218.045 246.905 220.755 247.075 ;
      RECT 387.92 249.565 388.85 252.425 ;
      RECT 389.24 249.475 389.85 252.915 ;
      RECT 386.44 252.915 415.045 253.535 ;
      RECT 386.44 246.7 387.06 252.915 ;
      RECT 393.915 249.475 394.525 252.915 ;
      RECT 398.59 249.475 399.2 252.915 ;
      RECT 403.265 249.475 403.875 252.915 ;
      RECT 440.12 230.315 440.29 235.935 ;
      RECT 439.24 234.995 439.41 236.06 ;
      RECT 438.62 234.57 438.79 236.06 ;
      RECT 437.74 230.315 437.91 235.935 ;
      RECT 438.62 230.62 438.79 233.33 ;
      RECT 438.04 237.415 438.55 237.745 ;
      RECT 438.11 237.745 438.48 250.37 ;
      RECT 438.04 250.37 438.55 250.7 ;
      RECT 439.54 237.415 440.05 237.745 ;
      RECT 439.54 250.37 440.05 250.7 ;
      RECT 438.65 239.24 439.98 239.75 ;
      RECT 439.61 239.75 439.98 250.37 ;
      RECT 439.61 237.745 439.98 239.24 ;
      RECT 438.65 237.915 438.82 239.24 ;
      RECT 441.62 235.01 441.79 236.06 ;
      RECT 441.62 230.62 441.79 233.33 ;
      RECT 441 230.62 441.17 233.33 ;
      RECT 442.545 237.415 443.055 237.745 ;
      RECT 442.545 250.37 443.055 250.7 ;
      RECT 442.615 239.75 442.985 250.37 ;
      RECT 442.615 237.745 442.985 239.24 ;
      RECT 440.15 239.24 442.985 239.75 ;
      RECT 440.15 239.75 440.32 250.205 ;
      RECT 440.15 237.915 440.32 239.24 ;
      RECT 446.495 237.745 446.865 250.37 ;
      RECT 446.425 250.37 446.935 250.7 ;
      RECT 446.425 237.665 446.935 237.745 ;
      RECT 446.345 237.495 446.935 237.665 ;
      RECT 446.425 237.415 446.935 237.495 ;
      RECT 443.415 237.495 443.945 237.665 ;
      RECT 443.495 237.745 443.865 250.37 ;
      RECT 443.425 250.37 443.935 250.7 ;
      RECT 443.425 237.665 443.935 237.745 ;
      RECT 443.425 237.415 443.935 237.495 ;
      RECT 447.295 237.495 447.825 237.665 ;
      RECT 447.305 250.37 447.815 250.7 ;
      RECT 447.375 246.105 447.905 246.275 ;
      RECT 447.305 237.665 447.815 237.745 ;
      RECT 447.305 237.415 447.815 237.495 ;
      RECT 447.375 246.275 447.745 250.37 ;
      RECT 447.375 237.745 447.745 246.105 ;
      RECT 444.925 237.415 445.435 237.745 ;
      RECT 444.925 250.37 445.435 250.7 ;
      RECT 444.035 239.24 445.365 239.75 ;
      RECT 444.995 239.75 445.365 250.37 ;
      RECT 444.995 237.745 445.365 239.24 ;
      RECT 444.035 237.915 444.205 239.24 ;
      RECT 446.49 233.27 450.49 233.44 ;
      RECT 450.46 237.545 451.13 237.715 ;
      RECT 448.805 237.415 449.315 237.745 ;
      RECT 448.805 250.37 449.315 250.7 ;
      RECT 447.915 239.24 449.245 239.75 ;
      RECT 448.875 239.75 449.245 250.37 ;
      RECT 448.875 237.745 449.245 239.24 ;
      RECT 447.915 237.915 448.085 239.24 ;
      RECT 452.715 236.365 455.32 238.945 ;
      RECT 459.955 236.19 460.125 238.9 ;
      RECT 457.045 236.19 457.215 238.9 ;
      RECT 458.735 236.19 459.245 236.395 ;
      RECT 457.925 236.19 458.435 236.395 ;
      RECT 457.925 236.395 459.245 238.96 ;
      RECT 463.38 236.19 463.55 240.94 ;
      RECT 461.62 236.19 461.79 240.94 ;
      RECT 465.14 236.19 465.65 241 ;
      RECT 462.5 236.19 462.67 240.94 ;
      RECT 464.26 236.19 464.43 240.94 ;
      RECT 141.23 242.025 146.425 243.72 ;
      RECT 141.23 239.55 146.095 241.24 ;
      RECT 141.31 244.175 141.68 244.345 ;
      RECT 141.31 243.89 143.665 244.175 ;
      RECT 141.31 244.345 142.06 246.365 ;
      RECT 142.23 244.175 143.665 246.535 ;
      RECT 141.31 246.365 141.68 246.535 ;
      RECT 141.31 246.535 143.665 246.935 ;
      RECT 146.615 239.55 152.28 241.24 ;
      RECT 146.955 242.03 152.18 243.72 ;
      RECT 152.94 243.7 158.99 243.72 ;
      RECT 152.82 242.09 158.99 243.7 ;
      RECT 152.94 242.03 158.99 242.09 ;
      RECT 152.8 239.55 161.42 241.24 ;
      RECT 149.545 244.175 151.72 246.535 ;
      RECT 149.545 243.89 152.64 244.175 ;
      RECT 149.545 246.535 152.64 246.935 ;
      RECT 152.27 244.175 152.64 244.345 ;
      RECT 152.27 246.365 152.64 246.535 ;
      RECT 151.89 244.345 152.64 246.365 ;
      RECT 161.965 239.55 163.79 241.16 ;
      RECT 162.135 241.16 163.79 241.24 ;
      RECT 161.385 242.03 163.79 243.72 ;
      RECT 165.72 238.05 170.47 238.545 ;
      RECT 165.72 239.495 170.47 239.99 ;
      RECT 167.66 245.655 168.51 250.435 ;
      RECT 167.66 244.805 173.41 245.655 ;
      RECT 167.66 250.435 173.41 251.715 ;
      RECT 167.85 251.715 173.22 251.845 ;
      RECT 172.56 245.655 173.41 250.435 ;
      RECT 165.72 238.715 170.47 239.325 ;
      RECT 216.595 244.805 222.345 245.655 ;
      RECT 221.495 245.655 222.345 250.435 ;
      RECT 216.595 250.435 222.345 251.715 ;
      RECT 216.785 251.715 222.155 251.845 ;
      RECT 216.595 245.655 217.445 250.435 ;
      RECT 219.535 238.05 224.285 238.545 ;
      RECT 219.535 239.495 224.285 239.99 ;
      RECT 219.535 238.715 224.285 239.325 ;
      RECT 226.215 242.03 228.62 243.72 ;
      RECT 226.215 239.55 228.04 241.16 ;
      RECT 226.215 241.16 227.87 241.24 ;
      RECT 231.015 242.09 237.185 243.7 ;
      RECT 231.015 243.7 237.065 243.72 ;
      RECT 231.015 242.03 237.065 242.09 ;
      RECT 228.585 239.55 237.205 241.24 ;
      RECT 237.825 242.03 243.05 243.72 ;
      RECT 237.725 239.55 243.39 241.24 ;
      RECT 237.365 244.175 237.735 244.345 ;
      RECT 237.365 243.89 240.46 244.175 ;
      RECT 237.365 244.345 238.115 246.365 ;
      RECT 238.285 244.175 240.46 246.535 ;
      RECT 237.365 246.365 237.735 246.535 ;
      RECT 237.365 246.535 240.46 246.935 ;
      RECT 243.91 239.55 248.775 241.24 ;
      RECT 243.58 242.025 248.775 243.72 ;
      RECT 246.34 244.175 247.775 246.535 ;
      RECT 246.34 243.89 248.695 244.175 ;
      RECT 246.34 246.535 248.695 246.935 ;
      RECT 248.325 244.175 248.695 244.345 ;
      RECT 248.325 246.365 248.695 246.535 ;
      RECT 412.155 231.76 412.325 234.47 ;
      RECT 411.095 237.24 412.555 237.91 ;
      RECT 409.9 237.24 410.07 238.26 ;
      RECT 408.795 236.07 409.325 236.24 ;
      RECT 409.155 235.47 409.325 236.07 ;
      RECT 411.01 235.47 411.18 236.48 ;
      RECT 408.13 233.22 408.66 234.23 ;
      RECT 408.13 231.54 408.66 232.55 ;
      RECT 408.535 238.53 409.125 238.7 ;
      RECT 408.58 236.9 409.125 238.53 ;
      RECT 408.075 236.9 408.245 238.26 ;
      RECT 409.325 236.42 410.3 236.54 ;
      RECT 409.325 236.54 409.935 237.04 ;
      RECT 409.325 238.53 409.915 238.7 ;
      RECT 409.325 237.04 409.7 238.53 ;
      RECT 409.58 235.47 410.3 236.42 ;
      RECT 409.96 231.04 412.1 231.21 ;
      RECT 408.265 236.48 408.935 236.65 ;
      RECT 410.125 236.73 411.125 236.9 ;
      RECT 419.55 230.115 419.72 233 ;
      RECT 417.79 230.115 417.96 233 ;
      RECT 418.52 236.31 419.05 236.48 ;
      RECT 418.45 234.66 419.12 234.83 ;
      RECT 417.135 233.55 420.375 233.72 ;
      RECT 418.63 234.83 418.97 236.31 ;
      RECT 418.63 233.72 418.97 234.66 ;
      RECT 416.91 230.29 417.08 233.27 ;
      RECT 419.15 235.01 419.32 236.09 ;
      RECT 418.27 235.01 418.44 236.09 ;
      RECT 418.67 230.29 418.84 233.27 ;
      RECT 421.34 230.62 421.51 233.33 ;
      RECT 421.34 235.01 421.51 236.06 ;
      RECT 422.84 230.62 423.01 233.33 ;
      RECT 424.895 237.495 425.425 237.665 ;
      RECT 424.97 237.745 425.34 250.37 ;
      RECT 424.9 250.37 425.41 250.7 ;
      RECT 424.9 237.665 425.41 237.745 ;
      RECT 424.9 237.415 425.41 237.495 ;
      RECT 425.22 230.3 425.39 235.935 ;
      RECT 422.84 235.01 423.01 236.06 ;
      RECT 424.34 234.995 424.51 236.06 ;
      RECT 424.34 230.62 424.51 233.33 ;
      RECT 424.02 237.415 424.53 237.745 ;
      RECT 424.02 250.37 424.53 250.7 ;
      RECT 424.09 239.75 424.46 250.37 ;
      RECT 424.09 237.745 424.46 239.24 ;
      RECT 423.13 239.24 424.46 239.75 ;
      RECT 423.13 239.75 423.3 250.205 ;
      RECT 423.13 237.915 423.3 239.24 ;
      RECT 421.02 237.415 421.53 237.745 ;
      RECT 420.93 239.235 421.46 239.405 ;
      RECT 421.02 250.37 421.53 250.7 ;
      RECT 421.09 239.405 421.46 250.37 ;
      RECT 421.09 237.745 421.46 239.235 ;
      RECT 422.52 237.415 423.03 237.745 ;
      RECT 422.52 250.37 423.03 250.7 ;
      RECT 422.59 239.75 422.96 250.37 ;
      RECT 422.59 237.745 422.96 239.24 ;
      RECT 421.63 239.24 422.96 239.75 ;
      RECT 421.63 239.75 421.8 250.205 ;
      RECT 421.63 237.915 421.8 239.24 ;
      RECT 420.43 230.29 420.6 233.27 ;
      RECT 426.1 230.62 426.27 233.33 ;
      RECT 426.72 234.995 426.89 236.06 ;
      RECT 427.6 230.315 427.77 235.935 ;
      RECT 426.72 230.62 426.89 233.33 ;
      RECT 428.48 230.62 428.65 233.33 ;
      RECT 426.1 234.57 426.27 236.06 ;
      RECT 427.9 237.415 428.41 237.745 ;
      RECT 427.81 239.795 428.34 239.965 ;
      RECT 427.9 250.37 428.41 250.7 ;
      RECT 427.97 239.965 428.34 250.37 ;
      RECT 427.97 237.745 428.34 239.795 ;
      RECT 426.4 237.415 426.91 237.745 ;
      RECT 426.4 250.37 426.91 250.7 ;
      RECT 425.51 239.24 426.84 239.75 ;
      RECT 426.47 239.75 426.84 250.37 ;
      RECT 426.47 237.745 426.84 239.24 ;
      RECT 425.51 237.915 425.68 239.24 ;
      RECT 429.1 235.01 429.27 236.06 ;
      RECT 430.6 234.995 430.77 236.06 ;
      RECT 430.6 230.62 430.77 233.33 ;
      RECT 429.1 230.62 429.27 233.33 ;
      RECT 428.78 237.415 429.29 237.745 ;
      RECT 428.85 237.745 429.22 250.37 ;
      RECT 428.78 250.37 429.29 250.7 ;
      RECT 430.28 237.415 430.79 237.745 ;
      RECT 430.28 250.37 430.79 250.7 ;
      RECT 429.39 239.24 430.72 239.75 ;
      RECT 430.35 239.75 430.72 250.37 ;
      RECT 430.35 237.745 430.72 239.24 ;
      RECT 429.39 237.915 429.56 239.24 ;
      RECT 431.48 230.315 431.65 235.935 ;
      RECT 434.145 237.495 434.675 237.665 ;
      RECT 434.23 237.745 434.6 250.37 ;
      RECT 434.16 250.37 434.67 250.7 ;
      RECT 434.16 237.665 434.67 237.745 ;
      RECT 434.16 237.415 434.67 237.495 ;
      RECT 432.36 234.57 432.53 236.06 ;
      RECT 432.36 230.62 432.53 233.33 ;
      RECT 432.98 234.995 433.15 236.06 ;
      RECT 433.86 230.315 434.03 235.935 ;
      RECT 432.98 230.62 433.15 233.33 ;
      RECT 433.28 237.415 433.79 237.745 ;
      RECT 433.28 250.37 433.79 250.7 ;
      RECT 430.89 239.24 433.72 239.75 ;
      RECT 433.35 239.75 433.72 250.37 ;
      RECT 433.35 237.745 433.72 239.24 ;
      RECT 430.89 239.75 431.06 250.205 ;
      RECT 430.89 237.915 431.06 239.24 ;
      RECT 434.74 230.62 434.91 233.33 ;
      RECT 435.36 230.62 435.53 233.33 ;
      RECT 435.36 235.01 435.53 236.06 ;
      RECT 436.86 234.995 437.03 236.06 ;
      RECT 436.86 230.62 437.03 233.33 ;
      RECT 435.66 237.415 436.17 237.745 ;
      RECT 435.66 250.37 436.17 250.7 ;
      RECT 434.77 239.24 436.1 239.75 ;
      RECT 435.73 239.75 436.1 250.37 ;
      RECT 435.73 237.745 436.1 239.24 ;
      RECT 434.77 237.915 434.94 239.24 ;
      RECT 437.16 237.415 437.67 237.745 ;
      RECT 437.07 239.795 437.6 239.965 ;
      RECT 437.16 250.37 437.67 250.7 ;
      RECT 437.23 239.965 437.6 250.37 ;
      RECT 437.23 237.745 437.6 239.795 ;
      RECT 439.24 230.62 439.41 233.33 ;
      RECT 165.72 237.385 170.47 237.88 ;
      RECT 170.64 234.695 170.885 236.485 ;
      RECT 165.33 236.485 170.885 236.655 ;
      RECT 165.33 236.655 165.5 239.66 ;
      RECT 165.33 236.27 165.5 236.485 ;
      RECT 167.18 234.495 170.155 234.99 ;
      RECT 165.72 236.825 170.47 237.215 ;
      RECT 167.18 230.595 169.89 231.205 ;
      RECT 167.18 231.375 170.155 231.985 ;
      RECT 167.18 232.155 169.89 232.765 ;
      RECT 167.18 232.935 170.155 233.545 ;
      RECT 167.18 233.715 169.89 234.325 ;
      RECT 219.535 235.94 224.285 236.215 ;
      RECT 219.63 236.215 224.12 236.315 ;
      RECT 219.535 237.385 224.285 237.88 ;
      RECT 219.85 234.495 222.825 234.99 ;
      RECT 219.12 234.695 219.365 236.485 ;
      RECT 224.505 236.655 224.675 239.66 ;
      RECT 219.12 236.485 224.675 236.655 ;
      RECT 224.505 236.27 224.675 236.485 ;
      RECT 219.535 236.825 224.285 237.215 ;
      RECT 220.115 230.595 222.825 231.205 ;
      RECT 219.85 231.375 222.825 231.985 ;
      RECT 220.115 232.155 222.825 232.765 ;
      RECT 219.85 232.935 222.825 233.545 ;
      RECT 220.115 233.715 222.825 234.325 ;
      RECT 227.24 232.55 227.605 238.03 ;
      RECT 227.335 238.03 227.505 238.05 ;
      RECT 228.055 237.13 247.765 237.74 ;
      RECT 228.055 230.825 247.765 231.435 ;
      RECT 312.695 237.1 313.675 239.845 ;
      RECT 312.695 239.845 323.78 240.135 ;
      RECT 312.695 240.135 324.48 240.705 ;
      RECT 324.015 234.66 324.645 235.96 ;
      RECT 324.015 233.17 324.545 234.66 ;
      RECT 323.95 239.795 324.48 239.965 ;
      RECT 324.31 237.1 324.645 238.4 ;
      RECT 324.31 238.4 324.48 239.795 ;
      RECT 388.345 235.7 388.515 238.41 ;
      RECT 387.465 235.7 387.635 238.41 ;
      RECT 389.855 235.64 390.385 235.81 ;
      RECT 389.965 235.81 390.135 236.14 ;
      RECT 389.965 235.47 390.135 235.64 ;
      RECT 390.22 233.22 390.75 234.23 ;
      RECT 386.68 233.22 387.535 234.23 ;
      RECT 390.22 231.54 390.75 232.55 ;
      RECT 390.165 236.9 390.335 238.26 ;
      RECT 387.085 232.8 390.345 232.97 ;
      RECT 390.355 236.48 391.025 236.65 ;
      RECT 387.875 231.54 388.405 232.55 ;
      RECT 388.035 234.95 388.565 234.98 ;
      RECT 387.665 235.12 388.335 235.15 ;
      RECT 387.665 234.98 388.565 235.12 ;
      RECT 389.04 233.22 389.57 234.23 ;
      RECT 387.875 233.22 388.405 234.23 ;
      RECT 395.805 231.76 395.975 234.47 ;
      RECT 391.825 231.76 391.995 234.47 ;
      RECT 392.345 234.32 392.875 234.49 ;
      RECT 392.705 231.76 392.875 234.32 ;
      RECT 393.365 231.76 393.535 234.47 ;
      RECT 394.245 231.76 394.415 234.47 ;
      RECT 393.185 237.24 394.645 237.91 ;
      RECT 391.99 237.24 392.16 238.26 ;
      RECT 390.885 236.07 391.415 236.24 ;
      RECT 391.245 235.47 391.415 236.07 ;
      RECT 390.625 238.53 391.215 238.7 ;
      RECT 390.67 236.9 391.215 238.53 ;
      RECT 391.415 236.42 392.39 236.54 ;
      RECT 391.415 236.54 392.025 237.04 ;
      RECT 391.415 238.53 392.005 238.7 ;
      RECT 391.415 237.04 391.79 238.53 ;
      RECT 391.67 235.47 392.39 236.42 ;
      RECT 393.1 235.47 393.27 236.48 ;
      RECT 396.03 231.04 398.17 231.21 ;
      RECT 392.05 231.04 394.19 231.21 ;
      RECT 395.575 237.24 397.035 237.91 ;
      RECT 392.215 236.73 393.215 236.9 ;
      RECT 398.225 231.76 398.395 234.47 ;
      RECT 397.345 234.32 397.875 234.49 ;
      RECT 397.345 231.76 397.515 234.32 ;
      RECT 396.685 231.76 396.855 234.47 ;
      RECT 399.47 233.22 400 234.23 ;
      RECT 399.47 231.54 400 232.55 ;
      RECT 399.875 232.8 403.135 232.97 ;
      RECT 401.815 231.54 402.345 232.55 ;
      RECT 400.65 233.22 401.18 234.23 ;
      RECT 401.815 233.22 402.345 234.23 ;
      RECT 398.06 237.24 398.23 238.26 ;
      RECT 398.805 236.07 399.335 236.24 ;
      RECT 398.805 235.47 398.975 236.07 ;
      RECT 399.005 238.53 399.595 238.7 ;
      RECT 399.005 236.9 399.55 238.53 ;
      RECT 397.83 236.42 398.805 236.54 ;
      RECT 398.195 236.54 398.805 237.04 ;
      RECT 398.215 238.53 398.805 238.7 ;
      RECT 398.43 237.04 398.805 238.53 ;
      RECT 397.83 235.47 398.55 236.42 ;
      RECT 396.95 235.47 397.12 236.48 ;
      RECT 399.195 236.48 399.865 236.65 ;
      RECT 397.005 236.73 398.005 236.9 ;
      RECT 401.705 235.7 401.875 238.41 ;
      RECT 399.835 235.64 400.365 235.81 ;
      RECT 400.085 235.81 400.255 236.14 ;
      RECT 400.085 235.47 400.255 235.64 ;
      RECT 399.885 236.9 400.055 238.26 ;
      RECT 401.655 234.95 402.185 234.98 ;
      RECT 401.885 235.12 402.555 235.15 ;
      RECT 401.655 234.98 402.555 235.12 ;
      RECT 406.255 235.7 406.425 238.41 ;
      RECT 405.375 235.7 405.545 238.41 ;
      RECT 402.585 235.7 402.755 238.41 ;
      RECT 407.765 235.64 408.295 235.81 ;
      RECT 407.875 235.81 408.045 236.14 ;
      RECT 407.875 235.47 408.045 235.64 ;
      RECT 402.685 233.22 403.54 234.23 ;
      RECT 404.59 233.22 405.445 234.23 ;
      RECT 404.995 232.8 408.255 232.97 ;
      RECT 405.785 231.54 406.315 232.55 ;
      RECT 405.945 234.95 406.475 234.98 ;
      RECT 405.575 235.12 406.245 235.15 ;
      RECT 405.575 234.98 406.475 235.12 ;
      RECT 406.95 233.22 407.48 234.23 ;
      RECT 405.785 233.22 406.315 234.23 ;
      RECT 409.735 231.76 409.905 234.47 ;
      RECT 410.255 234.32 410.785 234.49 ;
      RECT 410.615 231.76 410.785 234.32 ;
      RECT 411.275 231.76 411.445 234.47 ;
      RECT 429.37 236.23 429.88 236.56 ;
      RECT 428.48 234.225 429.81 234.735 ;
      RECT 429.44 234.735 429.81 236.23 ;
      RECT 429.44 230.07 429.81 234.225 ;
      RECT 428.48 234.735 428.65 236.06 ;
      RECT 430.79 229.9 431.46 230.07 ;
      RECT 430.87 236.23 431.38 236.56 ;
      RECT 429.98 234.225 431.31 234.735 ;
      RECT 430.94 234.735 431.31 236.23 ;
      RECT 430.94 230.07 431.31 234.225 ;
      RECT 429.98 234.735 430.15 236.06 ;
      RECT 429.98 230.315 430.15 234.225 ;
      RECT 427.645 222.65 427.815 225.36 ;
      RECT 428.165 222.63 428.695 222.8 ;
      RECT 428.525 222.8 428.695 225.36 ;
      RECT 429.185 222.65 429.355 225.36 ;
      RECT 430.065 222.65 430.235 225.36 ;
      RECT 426.04 222.89 426.57 223.9 ;
      RECT 426.04 224.57 426.57 225.58 ;
      RECT 428.775 226.57 429.285 227.58 ;
      RECT 426.715 226.57 427.225 227.58 ;
      RECT 427.915 226.57 428.085 227.6 ;
      RECT 427.485 226.27 427.655 227.58 ;
      RECT 428.345 226.27 428.515 227.58 ;
      RECT 427.87 225.91 430.01 226.08 ;
      RECT 427.28 227.83 428.72 228 ;
      RECT 431.67 229.9 432.34 230.07 ;
      RECT 431.82 230.07 432.19 236.23 ;
      RECT 431.735 236.31 432.265 236.48 ;
      RECT 431.75 236.48 432.26 236.56 ;
      RECT 431.75 236.23 432.26 236.31 ;
      RECT 433.17 229.9 433.84 230.07 ;
      RECT 433.16 234.01 433.69 234.18 ;
      RECT 433.25 236.23 433.76 236.56 ;
      RECT 433.32 234.18 433.69 236.23 ;
      RECT 433.32 230.07 433.69 234.01 ;
      RECT 434.05 229.9 434.72 230.07 ;
      RECT 434.2 230.07 434.57 236.23 ;
      RECT 434.13 236.23 434.64 236.56 ;
      RECT 435.55 229.9 436.22 230.07 ;
      RECT 435.63 236.23 436.14 236.56 ;
      RECT 434.74 234.225 436.07 234.735 ;
      RECT 435.7 234.735 436.07 236.23 ;
      RECT 435.7 230.07 436.07 234.225 ;
      RECT 434.74 234.735 434.91 236.06 ;
      RECT 434.045 222.65 434.215 225.36 ;
      RECT 433.165 222.63 433.695 222.8 ;
      RECT 433.165 222.8 433.335 225.36 ;
      RECT 432.505 222.65 432.675 225.36 ;
      RECT 431.625 222.65 431.795 225.36 ;
      RECT 435.29 222.89 435.82 223.9 ;
      RECT 435.29 224.57 435.82 225.58 ;
      RECT 436.42 226.57 436.93 227.58 ;
      RECT 432.575 226.57 433.085 227.58 ;
      RECT 434.635 226.57 435.145 227.58 ;
      RECT 433.775 226.57 433.945 227.6 ;
      RECT 434.205 226.27 434.375 227.58 ;
      RECT 433.345 226.27 433.515 227.58 ;
      RECT 435.695 224.15 438.955 224.32 ;
      RECT 436.595 224.56 436.875 225.77 ;
      RECT 436.595 225.77 439.22 226.02 ;
      RECT 437.995 226.02 438.275 227.59 ;
      RECT 437.135 226.02 437.415 227.59 ;
      RECT 438.955 224.56 439.22 225.77 ;
      RECT 436.47 222.89 437 223.9 ;
      RECT 431.85 225.91 433.99 226.08 ;
      RECT 433.14 227.83 434.58 228 ;
      RECT 441.81 229.9 442.48 230.07 ;
      RECT 441.89 236.23 442.4 236.56 ;
      RECT 441 234.225 442.33 234.735 ;
      RECT 441.96 234.735 442.33 236.23 ;
      RECT 441.96 230.07 442.33 234.225 ;
      RECT 441 234.735 441.17 236.06 ;
      RECT 440.31 229.9 440.98 230.07 ;
      RECT 440.39 236.23 440.9 236.56 ;
      RECT 440.46 233.875 441.06 234.045 ;
      RECT 440.46 234.045 440.83 236.23 ;
      RECT 440.46 230.07 440.83 233.875 ;
      RECT 439.43 229.9 440.1 230.07 ;
      RECT 439.58 230.07 439.95 236.23 ;
      RECT 439.475 236.31 440.02 236.48 ;
      RECT 439.51 236.48 440.02 236.56 ;
      RECT 439.51 236.23 440.02 236.31 ;
      RECT 437.05 229.9 437.72 230.07 ;
      RECT 437.13 236.23 437.64 236.56 ;
      RECT 436.24 234.225 437.57 234.735 ;
      RECT 437.2 234.735 437.57 236.23 ;
      RECT 437.2 230.07 437.57 234.225 ;
      RECT 436.24 234.735 436.41 236.06 ;
      RECT 436.24 230.315 436.41 234.225 ;
      RECT 437.93 229.9 438.6 230.07 ;
      RECT 438.08 230.07 438.45 236.23 ;
      RECT 438 236.31 438.53 236.48 ;
      RECT 438.01 236.48 438.52 236.56 ;
      RECT 438.01 236.23 438.52 236.31 ;
      RECT 438.505 222.89 439.36 223.9 ;
      RECT 438.48 226.57 438.99 227.58 ;
      RECT 444.665 218.755 444.835 223.505 ;
      RECT 442.385 218.755 442.555 223.505 ;
      RECT 442.385 223.505 444.835 228.605 ;
      RECT 437.62 226.57 437.79 227.58 ;
      RECT 442.655 230.005 443.185 230.175 ;
      RECT 442.5 230.315 443.005 236.06 ;
      RECT 442.655 230.175 443.005 230.315 ;
      RECT 437.635 224.57 438.165 225.58 ;
      RECT 437.635 222.89 438.165 223.9 ;
      RECT 436.985 227.83 438.425 228 ;
      RECT 446.265 223.2 446.435 233.05 ;
      RECT 450.545 223.2 450.715 233.05 ;
      RECT 459.105 223.2 459.275 233.05 ;
      RECT 454.825 223.2 454.995 233.05 ;
      RECT 463.385 223.2 463.555 233.05 ;
      RECT 465.665 223.2 465.835 233.05 ;
      RECT 65.36 234.66 65.99 235.96 ;
      RECT 65.46 233.17 65.99 234.66 ;
      RECT 65.525 239.795 66.055 239.965 ;
      RECT 65.36 237.1 65.695 238.4 ;
      RECT 65.525 238.4 65.695 239.795 ;
      RECT 76.33 237.1 77.31 239.845 ;
      RECT 66.225 239.845 77.31 240.135 ;
      RECT 65.525 240.135 77.31 240.705 ;
      RECT 142.24 237.13 161.95 237.74 ;
      RECT 142.24 230.825 161.95 231.435 ;
      RECT 162.4 232.55 162.765 238.03 ;
      RECT 162.5 238.03 162.67 238.05 ;
      RECT 165.72 235.94 170.47 236.215 ;
      RECT 165.885 236.215 170.375 236.315 ;
      RECT 402.175 229.53 402.455 231.1 ;
      RECT 400.775 231.35 401.055 232.56 ;
      RECT 403.135 231.35 403.4 232.56 ;
      RECT 401.8 229.54 401.97 230.55 ;
      RECT 401.165 229.12 402.605 229.29 ;
      RECT 401.165 227.83 402.605 228 ;
      RECT 402.685 222.89 403.54 223.9 ;
      RECT 404.59 222.89 405.445 223.9 ;
      RECT 405.785 222.89 406.315 223.9 ;
      RECT 406.95 222.89 407.48 223.9 ;
      RECT 402.66 226.57 403.17 227.58 ;
      RECT 404.73 225.77 407.355 226.02 ;
      RECT 404.73 224.56 404.995 225.77 ;
      RECT 406.535 226.02 406.815 227.59 ;
      RECT 407.075 224.56 407.355 225.77 ;
      RECT 405.675 226.02 405.955 227.59 ;
      RECT 407.02 226.57 407.53 227.58 ;
      RECT 404.96 226.57 405.47 227.58 ;
      RECT 406.16 226.57 406.33 227.58 ;
      RECT 405.785 224.57 406.315 225.58 ;
      RECT 404.995 224.15 408.255 224.32 ;
      RECT 402.66 229.54 403.17 230.55 ;
      RECT 407.02 229.54 407.53 230.55 ;
      RECT 404.96 229.54 405.47 230.55 ;
      RECT 406.535 229.53 406.815 231.1 ;
      RECT 404.73 231.1 407.355 231.35 ;
      RECT 405.675 229.53 405.955 231.1 ;
      RECT 407.075 231.35 407.355 232.56 ;
      RECT 404.73 231.35 404.995 232.56 ;
      RECT 406.16 229.54 406.33 230.55 ;
      RECT 405.525 229.12 406.965 229.29 ;
      RECT 405.525 227.83 406.965 228 ;
      RECT 413.715 222.65 413.885 225.36 ;
      RECT 409.735 222.65 409.905 225.36 ;
      RECT 410.255 222.63 410.785 222.8 ;
      RECT 410.615 222.8 410.785 225.36 ;
      RECT 411.275 222.65 411.445 225.36 ;
      RECT 412.155 222.65 412.325 225.36 ;
      RECT 408.13 222.89 408.66 223.9 ;
      RECT 408.13 224.57 408.66 225.58 ;
      RECT 410.865 226.57 411.375 227.58 ;
      RECT 408.805 226.57 409.315 227.58 ;
      RECT 410.865 229.54 411.375 230.55 ;
      RECT 408.805 229.54 409.315 230.55 ;
      RECT 410.435 226.27 410.605 227.58 ;
      RECT 410.435 229.54 410.605 230.85 ;
      RECT 410.005 226.57 410.175 227.6 ;
      RECT 410.005 229.52 410.175 230.55 ;
      RECT 409.575 226.27 409.745 227.58 ;
      RECT 409.575 229.54 409.745 230.85 ;
      RECT 409.37 229.12 410.81 229.29 ;
      RECT 409.96 225.91 412.1 226.08 ;
      RECT 409.37 227.83 410.81 228 ;
      RECT 416.135 222.65 416.305 225.36 ;
      RECT 415.255 222.63 415.785 222.8 ;
      RECT 415.255 222.8 415.425 225.36 ;
      RECT 414.595 222.65 414.765 225.36 ;
      RECT 417.38 222.89 417.91 223.9 ;
      RECT 417.38 224.57 417.91 225.58 ;
      RECT 418.51 226.57 419.02 227.58 ;
      RECT 414.665 226.57 415.175 227.58 ;
      RECT 416.725 226.57 417.235 227.58 ;
      RECT 415.865 226.57 416.035 227.6 ;
      RECT 416.295 226.27 416.465 227.58 ;
      RECT 419.225 226.02 419.505 227.59 ;
      RECT 418.685 225.77 421.31 226.02 ;
      RECT 418.685 224.56 418.965 225.77 ;
      RECT 420.085 226.02 420.365 227.59 ;
      RECT 421.045 224.56 421.31 225.77 ;
      RECT 415.435 226.27 415.605 227.58 ;
      RECT 417.785 224.15 421.045 224.32 ;
      RECT 418.56 222.89 419.09 223.9 ;
      RECT 419.075 227.83 420.515 228 ;
      RECT 413.94 225.91 416.08 226.08 ;
      RECT 415.23 227.83 416.67 228 ;
      RECT 420.595 222.89 421.45 223.9 ;
      RECT 419.725 222.89 420.255 223.9 ;
      RECT 422.5 222.89 423.355 223.9 ;
      RECT 423.695 222.89 424.225 223.9 ;
      RECT 424.86 222.89 425.39 223.9 ;
      RECT 419.725 224.57 420.255 225.58 ;
      RECT 422.64 224.56 422.905 225.77 ;
      RECT 422.64 225.77 425.265 226.02 ;
      RECT 424.985 224.56 425.265 225.77 ;
      RECT 423.585 226.02 423.865 227.59 ;
      RECT 424.445 226.02 424.725 227.59 ;
      RECT 423.695 224.57 424.225 225.58 ;
      RECT 422.905 224.15 426.165 224.32 ;
      RECT 421.53 229.9 422.2 230.07 ;
      RECT 421.52 234.57 422.05 234.74 ;
      RECT 421.61 236.23 422.12 236.56 ;
      RECT 421.68 234.74 422.05 236.23 ;
      RECT 421.68 230.07 422.05 234.57 ;
      RECT 420.57 226.57 421.08 227.58 ;
      RECT 419.71 226.57 419.88 227.58 ;
      RECT 423.03 229.9 423.7 230.07 ;
      RECT 423.11 236.23 423.62 236.56 ;
      RECT 423.18 234.735 423.55 236.23 ;
      RECT 423.18 230.07 423.55 234.225 ;
      RECT 422.22 234.225 423.55 234.735 ;
      RECT 422.22 234.735 422.39 236.06 ;
      RECT 422.22 230.315 422.39 234.225 ;
      RECT 424.53 229.9 425.2 230.07 ;
      RECT 424.61 236.23 425.12 236.56 ;
      RECT 424.68 234.735 425.05 236.23 ;
      RECT 424.68 230.07 425.05 234.225 ;
      RECT 423.72 234.225 425.05 234.735 ;
      RECT 423.72 234.735 423.89 236.06 ;
      RECT 423.72 230.315 423.89 234.225 ;
      RECT 424.93 226.57 425.44 227.58 ;
      RECT 422.87 226.57 423.38 227.58 ;
      RECT 424.07 226.57 424.24 227.58 ;
      RECT 423.435 227.83 424.875 228 ;
      RECT 425.41 229.9 426.08 230.07 ;
      RECT 425.56 230.07 425.93 236.23 ;
      RECT 425.485 236.31 426.015 236.48 ;
      RECT 425.49 236.48 426 236.56 ;
      RECT 425.49 236.23 426 236.31 ;
      RECT 426.91 229.9 427.58 230.07 ;
      RECT 426.9 234.01 427.43 234.18 ;
      RECT 426.99 236.23 427.5 236.56 ;
      RECT 427.06 234.18 427.43 236.23 ;
      RECT 427.06 230.07 427.43 234.01 ;
      RECT 427.79 229.9 428.46 230.07 ;
      RECT 427.94 230.07 428.31 236.23 ;
      RECT 427.87 236.23 428.38 236.56 ;
      RECT 429.29 229.9 429.96 230.07 ;
      RECT 265.28 229.255 266.13 232.355 ;
      RECT 276.99 229.255 277.84 232.355 ;
      RECT 253.91 232.355 313.205 233.39 ;
      RECT 288.7 229.255 289.55 232.355 ;
      RECT 300.41 229.255 301.26 232.355 ;
      RECT 312.355 229.255 313.205 232.355 ;
      RECT 253.91 228.22 313.205 229.255 ;
      RECT 314.02 224.26 323.75 224.59 ;
      RECT 324.72 224.26 325.25 224.59 ;
      RECT 324.815 224.59 325.145 240.725 ;
      RECT 325.315 224.76 325.845 230.315 ;
      RECT 325.31 223.865 325.845 224.035 ;
      RECT 325.42 224.035 325.845 224.76 ;
      RECT 323.95 224.34 324.48 224.51 ;
      RECT 324.015 226.75 324.645 228.05 ;
      RECT 324.015 224.51 324.48 226.75 ;
      RECT 326.04 223.865 326.6 224.205 ;
      RECT 326.04 224.205 327.03 224.735 ;
      RECT 326.5 224.735 327.03 237.925 ;
      RECT 326.5 237.925 327.465 239.225 ;
      RECT 327.2 224.035 327.565 233.745 ;
      RECT 326.77 223.865 327.565 224.035 ;
      RECT 351.085 229.105 361.38 229.275 ;
      RECT 351.085 245.69 361.38 245.865 ;
      RECT 353.61 229.275 353.78 245.69 ;
      RECT 356.13 229.275 356.3 245.69 ;
      RECT 358.65 229.275 358.82 245.69 ;
      RECT 361.17 229.275 361.38 245.69 ;
      RECT 351.085 229.275 351.26 245.69 ;
      RECT 354.23 229.695 355.68 229.865 ;
      RECT 351.71 229.695 353.16 229.865 ;
      RECT 359.27 229.695 360.72 229.865 ;
      RECT 356.75 229.695 358.2 229.865 ;
      RECT 386.68 222.89 387.535 223.9 ;
      RECT 390.22 222.89 390.75 223.9 ;
      RECT 387.875 222.89 388.405 223.9 ;
      RECT 389.04 222.89 389.57 223.9 ;
      RECT 386.82 224.56 387.085 225.77 ;
      RECT 386.82 225.77 389.445 226.02 ;
      RECT 388.625 226.02 388.905 227.59 ;
      RECT 389.165 224.56 389.445 225.77 ;
      RECT 387.765 226.02 388.045 227.59 ;
      RECT 387.05 226.57 387.56 227.58 ;
      RECT 387.085 224.15 390.345 224.32 ;
      RECT 390.22 224.57 390.75 225.58 ;
      RECT 389.11 226.57 389.62 227.58 ;
      RECT 388.25 226.57 388.42 227.58 ;
      RECT 387.875 224.57 388.405 225.58 ;
      RECT 387.05 229.54 387.56 230.55 ;
      RECT 386.07 239.055 413.105 239.06 ;
      RECT 413.28 239.055 420.055 239.06 ;
      RECT 386.07 238.89 420.055 239.055 ;
      RECT 412.935 237.3 420.055 238.89 ;
      RECT 386.07 228.645 386.24 238.89 ;
      RECT 395.025 228.645 395.195 238.89 ;
      RECT 403.98 228.645 404.15 238.89 ;
      RECT 412.935 228.645 415.84 237.3 ;
      RECT 386.07 228.475 439.97 228.645 ;
      RECT 386.07 218.34 386.24 228.475 ;
      RECT 395.025 218.34 395.195 228.475 ;
      RECT 403.98 218.34 404.15 228.475 ;
      RECT 412.935 218.34 413.105 228.475 ;
      RECT 421.89 218.34 422.06 228.475 ;
      RECT 430.845 218.34 431.015 228.475 ;
      RECT 439.8 218.34 439.97 228.475 ;
      RECT 386.07 218.17 439.97 218.34 ;
      RECT 389.11 229.54 389.62 230.55 ;
      RECT 388.625 229.53 388.905 231.1 ;
      RECT 386.82 231.1 389.445 231.35 ;
      RECT 387.765 229.53 388.045 231.1 ;
      RECT 389.165 231.35 389.445 232.56 ;
      RECT 386.82 231.35 387.085 232.56 ;
      RECT 388.25 229.54 388.42 230.55 ;
      RECT 387.615 229.12 389.055 229.29 ;
      RECT 387.615 227.83 389.055 228 ;
      RECT 395.805 222.65 395.975 225.36 ;
      RECT 391.825 222.65 391.995 225.36 ;
      RECT 392.345 222.63 392.875 222.8 ;
      RECT 392.705 222.8 392.875 225.36 ;
      RECT 393.365 222.65 393.535 225.36 ;
      RECT 394.245 222.65 394.415 225.36 ;
      RECT 392.955 229.54 393.465 230.55 ;
      RECT 390.895 229.54 391.405 230.55 ;
      RECT 392.955 226.57 393.465 227.58 ;
      RECT 390.895 226.57 391.405 227.58 ;
      RECT 392.525 226.27 392.695 227.58 ;
      RECT 392.525 229.54 392.695 230.85 ;
      RECT 392.095 226.57 392.265 227.6 ;
      RECT 392.095 229.52 392.265 230.55 ;
      RECT 391.665 226.27 391.835 227.58 ;
      RECT 391.665 229.54 391.835 230.85 ;
      RECT 391.46 229.12 392.9 229.29 ;
      RECT 396.03 225.91 398.17 226.08 ;
      RECT 392.05 225.91 394.19 226.08 ;
      RECT 391.46 227.83 392.9 228 ;
      RECT 398.225 222.65 398.395 225.36 ;
      RECT 397.345 222.63 397.875 222.8 ;
      RECT 397.345 222.8 397.515 225.36 ;
      RECT 396.685 222.65 396.855 225.36 ;
      RECT 399.47 222.89 400 223.9 ;
      RECT 401.815 222.89 402.345 223.9 ;
      RECT 400.65 222.89 401.18 223.9 ;
      RECT 399.47 224.57 400 225.58 ;
      RECT 396.755 226.57 397.265 227.58 ;
      RECT 398.815 226.57 399.325 227.58 ;
      RECT 397.525 226.27 397.695 227.58 ;
      RECT 397.955 226.57 398.125 227.6 ;
      RECT 398.385 226.27 398.555 227.58 ;
      RECT 400.6 226.57 401.11 227.58 ;
      RECT 401.315 226.02 401.595 227.59 ;
      RECT 400.775 225.77 403.4 226.02 ;
      RECT 400.775 224.56 401.055 225.77 ;
      RECT 402.175 226.02 402.455 227.59 ;
      RECT 403.135 224.56 403.4 225.77 ;
      RECT 401.8 226.57 401.97 227.58 ;
      RECT 401.815 224.57 402.345 225.58 ;
      RECT 399.875 224.15 403.135 224.32 ;
      RECT 396.755 229.54 397.265 230.55 ;
      RECT 398.815 229.54 399.325 230.55 ;
      RECT 397.525 229.54 397.695 230.85 ;
      RECT 397.955 229.52 398.125 230.55 ;
      RECT 398.385 229.54 398.555 230.85 ;
      RECT 397.32 229.12 398.76 229.29 ;
      RECT 397.32 227.83 398.76 228 ;
      RECT 400.6 229.54 401.11 230.55 ;
      RECT 401.315 229.53 401.595 231.1 ;
      RECT 400.775 231.1 403.4 231.35 ;
      RECT 62.44 223.865 63.235 224.035 ;
      RECT 66.255 224.26 75.985 224.59 ;
      RECT 65.46 229.68 65.99 232.355 ;
      RECT 65.46 228.83 76.63 229.68 ;
      RECT 65.46 232.355 76.63 232.985 ;
      RECT 75.78 228.05 76.63 228.83 ;
      RECT 66.315 232.985 76.63 233.56 ;
      RECT 76.33 225.65 77.31 226.63 ;
      RECT 77.14 234.98 77.31 235.96 ;
      RECT 89.085 225.65 89.255 226.63 ;
      RECT 88.25 234.98 89.855 235.745 ;
      RECT 100.795 225.65 100.965 226.63 ;
      RECT 88.875 235.745 89.855 238.08 ;
      RECT 100.795 234.98 100.965 235.96 ;
      RECT 112.505 225.65 112.675 226.63 ;
      RECT 124.215 225.65 124.385 226.63 ;
      RECT 100.795 237.1 100.965 238.08 ;
      RECT 112.505 234.98 112.675 235.96 ;
      RECT 135.925 225.65 136.095 226.63 ;
      RECT 112.505 237.1 112.675 238.08 ;
      RECT 124.215 234.98 124.385 235.96 ;
      RECT 124.215 237.1 124.385 238.08 ;
      RECT 135.925 234.98 136.095 235.96 ;
      RECT 135.925 237.1 136.095 238.08 ;
      RECT 75.78 227.73 136.095 228.05 ;
      RECT 66.315 233.56 136.095 234.41 ;
      RECT 76.33 226.63 136.095 227.73 ;
      RECT 76.33 234.41 136.095 234.98 ;
      RECT 88.875 238.08 136.095 239.5 ;
      RECT 123.875 229.255 124.725 232.355 ;
      RECT 76.8 229.255 77.65 232.355 ;
      RECT 88.745 229.255 89.595 232.355 ;
      RECT 76.8 228.22 136.095 229.255 ;
      RECT 100.455 229.255 101.305 232.355 ;
      RECT 112.165 229.255 113.015 232.355 ;
      RECT 76.8 232.355 136.095 233.39 ;
      RECT 142.24 222.245 161.95 222.855 ;
      RECT 142.24 223.805 161.95 224.415 ;
      RECT 142.24 226.145 161.95 226.755 ;
      RECT 142.24 227.705 161.95 228.315 ;
      RECT 142.24 229.265 161.95 229.875 ;
      RECT 142.24 224.585 161.95 225.195 ;
      RECT 142.24 223.025 161.95 223.635 ;
      RECT 165.72 227.705 170.47 228.2 ;
      RECT 164.99 231.315 166.52 235.42 ;
      RECT 165.67 228.585 166.52 231.315 ;
      RECT 166.69 228.7 167.01 235.275 ;
      RECT 166.69 235.275 170.155 235.77 ;
      RECT 165.72 222.245 170.47 222.855 ;
      RECT 165.72 223.025 170.47 223.635 ;
      RECT 165.72 223.805 170.47 224.415 ;
      RECT 165.72 224.585 170.47 225.195 ;
      RECT 165.72 225.365 170.47 225.975 ;
      RECT 165.72 226.145 170.47 226.755 ;
      RECT 165.72 226.925 170.47 227.535 ;
      RECT 167.18 228.37 170.155 228.865 ;
      RECT 167.18 229.035 169.89 229.645 ;
      RECT 167.18 229.815 170.155 230.425 ;
      RECT 219.535 227.705 224.285 228.2 ;
      RECT 219.535 222.245 224.285 222.855 ;
      RECT 219.535 223.025 224.285 223.635 ;
      RECT 219.535 223.805 224.285 224.415 ;
      RECT 219.535 224.585 224.285 225.195 ;
      RECT 219.535 225.365 224.285 225.975 ;
      RECT 219.535 226.145 224.285 226.755 ;
      RECT 219.535 226.925 224.285 227.535 ;
      RECT 219.85 228.37 222.825 228.865 ;
      RECT 220.115 229.035 222.825 229.645 ;
      RECT 219.85 229.815 222.825 230.425 ;
      RECT 223.485 231.315 225.015 235.42 ;
      RECT 223.485 228.585 224.335 231.315 ;
      RECT 222.995 228.7 223.315 235.275 ;
      RECT 219.85 235.275 223.315 235.77 ;
      RECT 228.055 222.245 247.765 222.855 ;
      RECT 228.055 223.805 247.765 224.415 ;
      RECT 228.055 226.145 247.765 226.755 ;
      RECT 228.055 227.705 247.765 228.315 ;
      RECT 228.055 229.265 247.765 229.875 ;
      RECT 228.055 224.585 247.765 225.195 ;
      RECT 228.055 223.025 247.765 223.635 ;
      RECT 313.375 228.05 314.225 228.83 ;
      RECT 313.375 228.83 324.545 229.68 ;
      RECT 324.015 229.68 324.545 232.355 ;
      RECT 313.375 232.355 324.545 232.985 ;
      RECT 313.375 232.985 323.69 233.56 ;
      RECT 253.91 225.65 254.08 226.63 ;
      RECT 265.62 225.65 265.79 226.63 ;
      RECT 277.33 225.65 277.5 226.63 ;
      RECT 289.04 225.65 289.21 226.63 ;
      RECT 300.75 225.65 300.92 226.63 ;
      RECT 312.695 225.65 313.675 226.63 ;
      RECT 312.695 234.98 312.865 235.96 ;
      RECT 300.15 234.98 301.755 235.745 ;
      RECT 300.15 235.745 301.13 238.08 ;
      RECT 289.04 234.98 289.21 235.96 ;
      RECT 289.04 237.1 289.21 238.08 ;
      RECT 277.33 234.98 277.5 235.96 ;
      RECT 277.33 237.1 277.5 238.08 ;
      RECT 265.62 234.98 265.79 235.96 ;
      RECT 265.62 237.1 265.79 238.08 ;
      RECT 253.91 234.98 254.08 235.96 ;
      RECT 253.91 237.1 254.08 238.08 ;
      RECT 253.91 227.73 314.225 228.05 ;
      RECT 253.91 226.63 313.675 227.73 ;
      RECT 253.91 233.56 323.69 234.41 ;
      RECT 253.91 234.41 313.675 234.98 ;
      RECT 253.91 238.08 301.13 239.5 ;
      RECT 253.81 223.695 254.42 225.35 ;
      RECT 300.41 223.695 301.02 225.35 ;
      RECT 252.335 223.695 253.185 243.64 ;
      RECT 252.335 243.64 339.535 244.49 ;
      RECT 265.28 223.695 266.13 225.35 ;
      RECT 276.99 223.695 277.84 225.35 ;
      RECT 288.7 223.695 289.55 225.35 ;
      RECT 252.495 244.49 331.14 244.52 ;
      RECT 326.085 224.905 326.255 230.57 ;
      RECT 338.685 223.695 339.535 243.64 ;
      RECT 300.41 240.705 301.26 242.54 ;
      RECT 300.41 242.54 327.275 243.46 ;
      RECT 325.405 239.805 327.275 242.54 ;
      RECT 325.405 230.57 326.255 239.805 ;
      RECT 253.91 239.67 301.26 240.705 ;
      RECT 265.28 240.705 266.13 243.64 ;
      RECT 276.99 240.705 277.84 243.64 ;
      RECT 288.7 240.705 289.55 243.64 ;
      RECT 300.41 243.46 327.245 243.64 ;
      RECT 252.335 222.845 339.535 223.695 ;
      RECT 405.93 222 406.83 222.14 ;
      RECT 411.095 219.21 412.555 219.88 ;
      RECT 409.9 219.185 410.43 219.88 ;
      RECT 409.155 220.98 409.325 221.65 ;
      RECT 408.535 218.52 409.125 218.69 ;
      RECT 408.58 218.69 409.125 220.22 ;
      RECT 409.325 220.58 410.3 220.79 ;
      RECT 409.325 220.08 409.935 220.58 ;
      RECT 409.58 220.79 410.3 221.65 ;
      RECT 409.325 218.52 409.915 218.69 ;
      RECT 409.325 218.69 409.7 220.08 ;
      RECT 411.01 220.64 411.18 221.65 ;
      RECT 408.265 220.47 408.935 220.64 ;
      RECT 410.125 220.22 411.125 220.39 ;
      RECT 413.485 219.21 414.945 219.88 ;
      RECT 419.26 218.71 419.43 221.42 ;
      RECT 415.61 219.185 416.14 219.88 ;
      RECT 416.715 220.98 416.885 221.65 ;
      RECT 417.995 220.98 418.165 221.87 ;
      RECT 416.915 218.52 417.505 218.69 ;
      RECT 416.915 218.69 417.46 220.22 ;
      RECT 417.795 219.125 418.325 220.22 ;
      RECT 415.74 220.58 416.715 220.79 ;
      RECT 416.105 220.08 416.715 220.58 ;
      RECT 415.74 220.79 416.46 221.65 ;
      RECT 416.125 218.52 416.715 218.69 ;
      RECT 416.34 218.69 416.715 220.08 ;
      RECT 414.86 220.64 415.03 221.65 ;
      RECT 417.105 220.47 417.775 220.64 ;
      RECT 414.915 220.22 415.915 220.39 ;
      RECT 419.44 221.97 420.11 222 ;
      RECT 419.21 222.14 419.74 222.17 ;
      RECT 419.21 222 420.11 222.14 ;
      RECT 424.52 218.71 424.69 221.42 ;
      RECT 423.64 218.71 423.81 221.42 ;
      RECT 420.14 218.71 420.31 221.42 ;
      RECT 423.84 221.97 424.51 222 ;
      RECT 424.21 222.14 424.74 222.17 ;
      RECT 423.84 222 424.74 222.14 ;
      RECT 429.005 219.21 430.465 219.88 ;
      RECT 427.81 219.185 428.34 219.88 ;
      RECT 427.065 220.98 427.235 221.65 ;
      RECT 425.785 220.98 425.955 221.87 ;
      RECT 426.445 218.52 427.035 218.69 ;
      RECT 426.49 218.69 427.035 220.22 ;
      RECT 425.625 219.125 426.155 220.22 ;
      RECT 427.235 220.58 428.21 220.79 ;
      RECT 427.235 220.08 427.845 220.58 ;
      RECT 427.49 220.79 428.21 221.65 ;
      RECT 427.235 218.52 427.825 218.69 ;
      RECT 427.235 218.69 427.61 220.08 ;
      RECT 428.92 220.64 429.09 221.65 ;
      RECT 426.175 220.47 426.845 220.64 ;
      RECT 428.035 220.22 429.035 220.39 ;
      RECT 431.395 219.21 432.855 219.88 ;
      RECT 433.52 219.185 434.05 219.88 ;
      RECT 434.625 220.98 434.795 221.65 ;
      RECT 435.905 220.98 436.075 221.87 ;
      RECT 434.825 218.52 435.415 218.69 ;
      RECT 434.825 218.69 435.37 220.22 ;
      RECT 435.705 219.125 436.235 220.22 ;
      RECT 433.65 220.58 434.625 220.79 ;
      RECT 434.015 220.08 434.625 220.58 ;
      RECT 433.65 220.79 434.37 221.65 ;
      RECT 434.035 218.52 434.625 218.69 ;
      RECT 434.25 218.69 434.625 220.08 ;
      RECT 432.77 220.64 432.94 221.65 ;
      RECT 435.015 220.47 435.685 220.64 ;
      RECT 432.825 220.22 433.825 220.39 ;
      RECT 437.17 218.71 437.34 221.42 ;
      RECT 438.05 218.71 438.22 221.42 ;
      RECT 442.61 218.175 444.61 218.345 ;
      RECT 443.125 218.345 444.065 222.18 ;
      RECT 437.35 221.97 438.02 222 ;
      RECT 437.12 222.14 437.65 222.17 ;
      RECT 437.12 222 438.02 222.14 ;
      RECT 446.265 211.94 446.435 221.79 ;
      RECT 446.49 222.01 450.49 222.18 ;
      RECT 450.545 211.94 450.715 221.79 ;
      RECT 454.825 211.94 454.995 221.79 ;
      RECT 459.105 211.94 459.275 221.79 ;
      RECT 463.385 211.94 463.555 221.79 ;
      RECT 465.665 211.94 465.835 221.79 ;
      RECT 28.625 229.105 38.92 229.275 ;
      RECT 28.625 245.69 38.92 245.865 ;
      RECT 31.185 229.275 31.355 245.69 ;
      RECT 36.225 229.275 36.395 245.69 ;
      RECT 33.705 229.275 33.875 245.69 ;
      RECT 28.625 229.275 28.835 245.69 ;
      RECT 38.745 229.275 38.92 245.69 ;
      RECT 29.285 229.695 30.735 229.865 ;
      RECT 34.325 229.695 35.775 229.865 ;
      RECT 36.845 229.695 38.295 229.865 ;
      RECT 31.805 229.695 33.255 229.865 ;
      RECT 50.47 243.64 137.67 244.49 ;
      RECT 88.985 223.695 89.595 225.35 ;
      RECT 135.585 223.695 136.195 225.35 ;
      RECT 136.82 223.695 137.67 243.64 ;
      RECT 58.865 244.49 137.51 244.52 ;
      RECT 100.455 223.695 101.305 225.35 ;
      RECT 112.165 223.695 113.015 225.35 ;
      RECT 123.875 223.695 124.725 225.35 ;
      RECT 63.75 224.905 63.92 230.57 ;
      RECT 63.75 230.57 64.6 239.805 ;
      RECT 50.47 223.695 51.32 243.64 ;
      RECT 62.73 239.805 64.6 242.54 ;
      RECT 62.73 242.54 89.595 243.46 ;
      RECT 88.745 240.705 89.595 242.54 ;
      RECT 88.745 239.67 136.095 240.705 ;
      RECT 100.455 240.705 101.305 243.64 ;
      RECT 112.165 240.705 113.015 243.64 ;
      RECT 123.875 240.705 124.725 243.64 ;
      RECT 62.76 243.46 89.595 243.64 ;
      RECT 50.47 222.845 137.67 223.695 ;
      RECT 64.755 224.26 65.285 224.59 ;
      RECT 64.86 224.59 65.19 240.725 ;
      RECT 64.16 224.76 64.69 230.315 ;
      RECT 64.16 223.865 64.695 224.035 ;
      RECT 64.16 224.035 64.585 224.76 ;
      RECT 65.525 224.34 66.055 224.51 ;
      RECT 65.36 226.75 65.99 228.05 ;
      RECT 65.525 224.51 65.99 226.75 ;
      RECT 63.405 223.865 63.965 224.205 ;
      RECT 62.975 224.205 63.965 224.735 ;
      RECT 62.975 224.735 63.505 237.925 ;
      RECT 62.54 237.925 63.505 239.225 ;
      RECT 62.44 224.035 62.805 233.745 ;
      RECT 145.1 216.235 145.77 216.405 ;
      RECT 147.16 216.235 147.83 216.405 ;
      RECT 143.04 216.235 143.71 216.405 ;
      RECT 151.28 216.235 151.95 216.405 ;
      RECT 149.22 216.235 149.89 216.405 ;
      RECT 165.72 221.465 170.47 222.075 ;
      RECT 169.26 220.235 171 220.765 ;
      RECT 170.64 220.765 171 222.01 ;
      RECT 165.195 221.91 165.5 230.71 ;
      RECT 162.5 230.71 165.5 230.99 ;
      RECT 162.5 221.91 162.755 230.71 ;
      RECT 163.93 230.99 164.82 238.295 ;
      RECT 219.535 221.465 224.285 222.075 ;
      RECT 219.005 220.765 219.365 222.01 ;
      RECT 219.005 220.235 220.745 220.765 ;
      RECT 219.535 221.045 248.345 221.215 ;
      RECT 225.455 238.575 248.345 239.105 ;
      RECT 226.245 232.05 227.07 238.575 ;
      RECT 230.885 239.105 239.335 239.275 ;
      RECT 226.245 231.16 227.07 231.605 ;
      RECT 248.175 232.05 248.345 238.575 ;
      RECT 226.245 231.605 248.345 232.05 ;
      RECT 218.665 221.045 218.835 240.355 ;
      RECT 225.455 239.105 225.625 240.355 ;
      RECT 218.665 240.355 225.625 240.525 ;
      RECT 224.98 221.215 227.08 230.235 ;
      RECT 248.175 221.215 248.345 231.605 ;
      RECT 224.505 221.91 224.81 230.71 ;
      RECT 224.505 230.71 227.505 230.99 ;
      RECT 227.25 221.91 227.505 230.71 ;
      RECT 225.185 230.99 226.075 238.295 ;
      RECT 238.055 216.235 238.725 216.405 ;
      RECT 240.115 216.235 240.785 216.405 ;
      RECT 244.235 216.235 244.905 216.405 ;
      RECT 242.175 216.235 242.845 216.405 ;
      RECT 250.415 216.235 251.085 216.405 ;
      RECT 248.355 216.235 249.025 216.405 ;
      RECT 246.295 216.235 246.965 216.405 ;
      RECT 250.72 221.23 341.15 222.08 ;
      RECT 250.72 245.255 341.15 246.105 ;
      RECT 340.3 222.08 341.15 245.255 ;
      RECT 250.72 222.08 251.57 245.255 ;
      RECT 252.475 216.235 253.145 216.405 ;
      RECT 256.595 216.235 257.265 216.405 ;
      RECT 254.535 216.235 255.205 216.405 ;
      RECT 262.775 216.235 263.445 216.405 ;
      RECT 258.655 216.235 259.325 216.405 ;
      RECT 260.715 216.235 261.385 216.405 ;
      RECT 264.835 216.235 265.505 216.405 ;
      RECT 268.955 216.235 269.625 216.405 ;
      RECT 266.895 216.235 267.565 216.405 ;
      RECT 273.075 216.235 273.745 216.405 ;
      RECT 271.015 216.235 271.685 216.405 ;
      RECT 279.255 216.235 279.925 216.405 ;
      RECT 275.135 216.235 275.805 216.405 ;
      RECT 277.195 216.235 277.865 216.405 ;
      RECT 281.315 216.235 281.985 216.405 ;
      RECT 285.435 216.235 286.105 216.405 ;
      RECT 283.375 216.235 284.045 216.405 ;
      RECT 287.495 216.235 288.165 216.405 ;
      RECT 312.4 215.155 315.24 215.385 ;
      RECT 316.54 215.155 319.38 215.385 ;
      RECT 328.955 215.155 331.8 215.385 ;
      RECT 333.1 215.155 335.94 215.385 ;
      RECT 354.925 214.38 355.095 217.34 ;
      RECT 355.15 217.56 357.43 217.73 ;
      RECT 356.375 217.73 357.37 217.735 ;
      RECT 357.71 217.56 359.99 217.73 ;
      RECT 358.05 217.73 358.815 217.735 ;
      RECT 360.045 214.38 360.215 217.34 ;
      RECT 358.765 214.63 358.935 217.34 ;
      RECT 360.27 217.56 362.55 217.73 ;
      RECT 360.33 217.73 361.325 217.735 ;
      RECT 361.325 214.63 361.495 217.34 ;
      RECT 356.205 214.63 356.375 217.34 ;
      RECT 357.485 214.38 357.655 217.34 ;
      RECT 365.165 214.38 365.335 217.34 ;
      RECT 362.83 217.56 365.11 217.73 ;
      RECT 363.235 217.73 364.23 217.735 ;
      RECT 363.885 214.63 364.055 217.34 ;
      RECT 362.605 214.38 362.775 217.34 ;
      RECT 388.7 218.71 388.87 221.42 ;
      RECT 387.82 218.71 387.99 221.42 ;
      RECT 389.965 220.98 390.135 221.87 ;
      RECT 389.805 219.125 390.335 220.22 ;
      RECT 390.355 220.47 391.025 220.64 ;
      RECT 388.02 221.97 388.69 222 ;
      RECT 388.39 222.14 388.92 222.17 ;
      RECT 388.02 222 388.92 222.14 ;
      RECT 390.67 218.69 391.215 220.22 ;
      RECT 390.625 218.52 391.215 218.69 ;
      RECT 393.185 219.21 394.645 219.88 ;
      RECT 391.99 219.185 392.52 219.88 ;
      RECT 391.245 220.98 391.415 221.65 ;
      RECT 391.415 220.58 392.39 220.79 ;
      RECT 391.415 220.08 392.025 220.58 ;
      RECT 391.67 220.79 392.39 221.65 ;
      RECT 391.415 218.52 392.005 218.69 ;
      RECT 391.415 218.69 391.79 220.08 ;
      RECT 393.1 220.64 393.27 221.65 ;
      RECT 392.215 220.22 393.215 220.39 ;
      RECT 395.575 219.21 397.035 219.88 ;
      RECT 401.35 218.71 401.52 221.42 ;
      RECT 397.7 219.185 398.23 219.88 ;
      RECT 398.805 220.98 398.975 221.65 ;
      RECT 400.085 220.98 400.255 221.87 ;
      RECT 399.005 218.52 399.595 218.69 ;
      RECT 399.005 218.69 399.55 220.22 ;
      RECT 399.885 219.125 400.415 220.22 ;
      RECT 397.83 220.58 398.805 220.79 ;
      RECT 398.195 220.08 398.805 220.58 ;
      RECT 397.83 220.79 398.55 221.65 ;
      RECT 398.215 218.52 398.805 218.69 ;
      RECT 398.43 218.69 398.805 220.08 ;
      RECT 396.95 220.64 397.12 221.65 ;
      RECT 399.195 220.47 399.865 220.64 ;
      RECT 397.005 220.22 398.005 220.39 ;
      RECT 401.53 221.97 402.2 222 ;
      RECT 401.3 222.14 401.83 222.17 ;
      RECT 401.3 222 402.2 222.14 ;
      RECT 406.61 218.71 406.78 221.42 ;
      RECT 405.73 218.71 405.9 221.42 ;
      RECT 402.23 218.71 402.4 221.42 ;
      RECT 407.875 220.98 408.045 221.87 ;
      RECT 407.715 219.125 408.245 220.22 ;
      RECT 405.93 221.97 406.6 222 ;
      RECT 406.3 222.14 406.83 222.17 ;
      RECT 399.6 207.34 400.92 210.11 ;
      RECT 400.935 206.95 401.605 207.12 ;
      RECT 396.86 207.855 397.46 208.025 ;
      RECT 396.86 208.025 397.03 208.255 ;
      RECT 396.86 207.585 397.03 207.855 ;
      RECT 406.33 207.34 406.5 210.05 ;
      RECT 407.21 207.34 408.53 210.11 ;
      RECT 406.525 206.95 407.195 207.12 ;
      RECT 410.09 207.44 410.76 207.61 ;
      RECT 408.56 210.325 410.76 210.995 ;
      RECT 410.09 210.15 410.76 210.325 ;
      RECT 408.735 207.54 409.04 210.325 ;
      RECT 409.24 207.34 409.41 210.05 ;
      RECT 410.09 208.22 410.82 209.54 ;
      RECT 410.67 207.855 411.27 208.025 ;
      RECT 411.1 208.025 411.27 208.255 ;
      RECT 411.1 207.585 411.27 207.855 ;
      RECT 411.1 209.68 412.12 209.85 ;
      RECT 411.1 209.85 411.27 210.185 ;
      RECT 411.1 209.515 411.27 209.68 ;
      RECT 411.47 207.41 412.12 209.68 ;
      RECT 415.28 207.44 415.95 207.61 ;
      RECT 415.28 210.325 417.48 210.995 ;
      RECT 415.28 210.15 415.95 210.325 ;
      RECT 417 207.54 417.305 210.325 ;
      RECT 416.63 207.34 416.8 210.05 ;
      RECT 419.54 207.34 419.71 210.05 ;
      RECT 415.22 208.22 415.95 209.54 ;
      RECT 417.51 207.34 418.83 210.11 ;
      RECT 418.845 206.95 419.515 207.12 ;
      RECT 414.77 207.855 415.37 208.025 ;
      RECT 414.77 208.025 414.94 208.255 ;
      RECT 414.77 207.585 414.94 207.855 ;
      RECT 413.92 209.68 414.94 209.85 ;
      RECT 414.77 209.85 414.94 210.185 ;
      RECT 414.77 209.515 414.94 209.68 ;
      RECT 413.92 207.41 414.57 209.68 ;
      RECT 424.24 207.34 424.41 210.05 ;
      RECT 425.12 207.34 426.44 210.11 ;
      RECT 424.435 206.95 425.105 207.12 ;
      RECT 428 207.44 428.67 207.61 ;
      RECT 426.47 210.325 428.67 210.995 ;
      RECT 428 210.15 428.67 210.325 ;
      RECT 426.645 207.54 426.95 210.325 ;
      RECT 427.15 207.34 427.32 210.05 ;
      RECT 428 208.22 428.73 209.54 ;
      RECT 428.58 207.855 429.18 208.025 ;
      RECT 429.01 208.025 429.18 208.255 ;
      RECT 429.01 207.585 429.18 207.855 ;
      RECT 429.01 209.68 430.03 209.85 ;
      RECT 429.01 209.85 429.18 210.185 ;
      RECT 429.01 209.515 429.18 209.68 ;
      RECT 429.38 207.41 430.03 209.68 ;
      RECT 433.19 207.44 433.86 207.61 ;
      RECT 433.19 210.325 435.39 210.995 ;
      RECT 433.19 210.15 433.86 210.325 ;
      RECT 434.91 207.54 435.215 210.325 ;
      RECT 434.54 207.34 434.71 210.05 ;
      RECT 433.13 208.22 433.86 209.54 ;
      RECT 435.42 207.34 436.74 210.11 ;
      RECT 436.755 206.95 437.425 207.12 ;
      RECT 432.68 207.855 433.28 208.025 ;
      RECT 432.68 208.025 432.85 208.255 ;
      RECT 432.68 207.585 432.85 207.855 ;
      RECT 431.83 209.68 432.85 209.85 ;
      RECT 432.68 209.85 432.85 210.185 ;
      RECT 432.68 209.515 432.85 209.68 ;
      RECT 431.83 207.41 432.48 209.68 ;
      RECT 437.45 207.34 437.62 210.05 ;
      RECT 446.49 210.765 450.49 210.935 ;
      RECT 24.67 214.38 24.84 217.34 ;
      RECT 24.895 217.56 27.175 217.73 ;
      RECT 25.775 217.73 26.77 217.735 ;
      RECT 30.015 217.56 32.295 217.73 ;
      RECT 31.19 217.73 31.955 217.735 ;
      RECT 29.79 214.38 29.96 217.34 ;
      RECT 31.07 214.63 31.24 217.34 ;
      RECT 25.95 214.63 26.12 217.34 ;
      RECT 27.455 217.56 29.735 217.73 ;
      RECT 28.68 217.73 29.675 217.735 ;
      RECT 28.51 214.63 28.68 217.34 ;
      RECT 27.23 214.38 27.4 217.34 ;
      RECT 34.91 214.38 35.08 217.34 ;
      RECT 33.63 214.63 33.8 217.34 ;
      RECT 32.575 217.56 34.855 217.73 ;
      RECT 32.635 217.73 33.63 217.735 ;
      RECT 32.35 214.38 32.52 217.34 ;
      RECT 54.065 215.155 56.905 215.385 ;
      RECT 58.205 215.155 61.05 215.385 ;
      RECT 70.625 215.155 73.465 215.385 ;
      RECT 74.765 215.155 77.605 215.385 ;
      RECT 103.9 216.235 104.57 216.405 ;
      RECT 105.96 216.235 106.63 216.405 ;
      RECT 101.84 216.235 102.51 216.405 ;
      RECT 110.08 216.235 110.75 216.405 ;
      RECT 108.02 216.235 108.69 216.405 ;
      RECT 112.14 216.235 112.81 216.405 ;
      RECT 114.2 216.235 114.87 216.405 ;
      RECT 116.26 216.235 116.93 216.405 ;
      RECT 118.32 216.235 118.99 216.405 ;
      RECT 120.38 216.235 121.05 216.405 ;
      RECT 122.44 216.235 123.11 216.405 ;
      RECT 126.56 216.235 127.23 216.405 ;
      RECT 124.5 216.235 125.17 216.405 ;
      RECT 128.62 216.235 129.29 216.405 ;
      RECT 130.68 216.235 131.35 216.405 ;
      RECT 132.74 216.235 133.41 216.405 ;
      RECT 134.8 216.235 135.47 216.405 ;
      RECT 138.92 216.235 139.59 216.405 ;
      RECT 136.86 216.235 137.53 216.405 ;
      RECT 140.98 216.235 141.65 216.405 ;
      RECT 48.855 221.23 139.285 222.08 ;
      RECT 48.855 245.255 139.285 246.105 ;
      RECT 48.855 222.08 49.705 245.255 ;
      RECT 138.435 222.08 139.285 245.255 ;
      RECT 141.66 221.045 170.47 221.215 ;
      RECT 141.66 238.575 164.55 239.105 ;
      RECT 162.935 232.05 163.76 238.575 ;
      RECT 150.67 239.105 159.12 239.275 ;
      RECT 162.935 231.16 163.76 231.605 ;
      RECT 141.66 232.05 141.83 238.575 ;
      RECT 141.66 231.605 163.76 232.05 ;
      RECT 171.17 221.045 171.34 240.355 ;
      RECT 164.38 239.105 164.55 240.355 ;
      RECT 164.38 240.355 171.34 240.525 ;
      RECT 162.925 221.215 165.025 230.235 ;
      RECT 141.66 221.215 141.83 231.605 ;
      RECT 445.655 229.45 445.825 232.32 ;
      RECT 466.22 222.67 466.45 233.7 ;
      RECT 445.625 211.185 466.45 211.415 ;
      RECT 445.625 222.44 466.45 222.67 ;
      RECT 446.265 200.695 446.435 210.545 ;
      RECT 450.545 200.695 450.715 210.545 ;
      RECT 454.825 200.695 454.995 210.545 ;
      RECT 459.105 200.695 459.275 210.545 ;
      RECT 463.385 200.695 463.555 210.545 ;
      RECT 465.665 200.695 465.835 210.545 ;
      RECT 25.6 209.8 25.77 212.51 ;
      RECT 22.45 208.335 36.68 209.185 ;
      RECT 22.45 209.185 25 213.44 ;
      RECT 22.48 219.39 32.945 219.455 ;
      RECT 29.785 209.185 30.295 213.44 ;
      RECT 35.49 209.185 36.68 213.44 ;
      RECT 22.64 207.86 36.68 208.335 ;
      RECT 35.49 213.95 36.68 218.195 ;
      RECT 35.3 218.195 36.68 218.2 ;
      RECT 22.48 219.33 36.68 219.39 ;
      RECT 22.45 218.2 36.68 219.33 ;
      RECT 22.45 213.44 36.68 213.95 ;
      RECT 22.45 213.95 24.145 218.2 ;
      RECT 30.92 209.68 31.09 210.69 ;
      RECT 30.92 212.245 31.09 213.115 ;
      RECT 26.48 209.8 26.65 212.51 ;
      RECT 28.24 209.8 28.41 212.51 ;
      RECT 27.36 209.8 27.53 212.51 ;
      RECT 25.755 212.73 26.425 212.9 ;
      RECT 31.145 210.91 32.625 211.08 ;
      RECT 26.705 212.73 28.185 212.9 ;
      RECT 31.075 211.785 31.745 211.955 ;
      RECT 32.68 209.68 32.85 210.69 ;
      RECT 32.68 212.185 32.85 212.915 ;
      RECT 31.8 209.68 31.97 210.69 ;
      RECT 31.8 212.245 31.97 213.115 ;
      RECT 32.025 211.785 32.695 211.955 ;
      RECT 55.4 199.985 55.57 214.985 ;
      RECT 59.54 199.985 59.71 214.985 ;
      RECT 63.68 199.985 63.85 214.985 ;
      RECT 67.82 199.985 67.99 214.985 ;
      RECT 71.96 199.985 72.13 214.985 ;
      RECT 76.1 199.985 76.27 214.985 ;
      RECT 164.39 206.465 164.56 213.315 ;
      RECT 161.27 206.465 161.44 213.255 ;
      RECT 159.35 208.205 160.075 208.735 ;
      RECT 162.05 206.465 162.22 213.255 ;
      RECT 163.61 206.465 163.78 213.255 ;
      RECT 162.83 206.465 163 213.255 ;
      RECT 165.84 206.8 168.55 206.98 ;
      RECT 165.84 217.44 168.55 217.62 ;
      RECT 168.23 206.98 168.5 217.44 ;
      RECT 167.45 206.98 167.72 217.44 ;
      RECT 166.67 206.98 166.94 217.44 ;
      RECT 165.89 206.98 166.16 217.44 ;
      RECT 221.455 206.8 224.165 206.98 ;
      RECT 221.455 217.44 224.165 217.62 ;
      RECT 221.505 206.98 221.775 217.44 ;
      RECT 222.285 206.98 222.555 217.44 ;
      RECT 223.065 206.98 223.335 217.44 ;
      RECT 223.845 206.98 224.115 217.44 ;
      RECT 225.445 206.465 225.615 213.315 ;
      RECT 227.785 206.465 227.955 213.255 ;
      RECT 226.225 206.465 226.395 213.255 ;
      RECT 227.005 206.465 227.175 213.255 ;
      RECT 228.565 206.465 228.735 213.255 ;
      RECT 229.93 208.205 230.655 208.735 ;
      RECT 313.735 199.985 313.905 214.985 ;
      RECT 317.875 199.985 318.045 214.985 ;
      RECT 322.015 199.985 322.185 214.985 ;
      RECT 326.155 199.985 326.325 214.985 ;
      RECT 330.295 199.985 330.465 214.985 ;
      RECT 334.435 199.985 334.605 214.985 ;
      RECT 353.325 208.335 367.555 209.185 ;
      RECT 365.005 209.185 367.555 213.44 ;
      RECT 357.06 219.39 367.525 219.455 ;
      RECT 353.325 207.86 367.365 208.335 ;
      RECT 353.325 218.195 354.705 218.2 ;
      RECT 353.325 213.95 354.515 218.195 ;
      RECT 359.71 209.185 360.22 213.44 ;
      RECT 353.325 209.185 354.515 213.44 ;
      RECT 353.325 219.33 367.525 219.39 ;
      RECT 353.325 213.44 367.555 213.95 ;
      RECT 365.86 213.95 367.555 218.2 ;
      RECT 353.325 218.2 367.555 219.33 ;
      RECT 357.155 209.68 357.325 210.69 ;
      RECT 358.915 209.68 359.085 210.69 ;
      RECT 357.155 212.185 357.325 212.915 ;
      RECT 358.915 212.245 359.085 213.115 ;
      RECT 361.595 209.8 361.765 212.51 ;
      RECT 358.26 211.785 358.93 211.955 ;
      RECT 358.035 209.68 358.205 210.69 ;
      RECT 357.38 210.91 358.86 211.08 ;
      RECT 358.035 212.245 358.205 213.115 ;
      RECT 357.31 211.785 357.98 211.955 ;
      RECT 363.355 209.8 363.525 212.51 ;
      RECT 364.235 209.8 364.405 212.51 ;
      RECT 362.475 209.8 362.645 212.51 ;
      RECT 363.58 212.73 364.25 212.9 ;
      RECT 361.82 212.73 363.3 212.9 ;
      RECT 388.42 207.34 388.59 210.05 ;
      RECT 389.3 207.34 390.62 210.11 ;
      RECT 388.615 206.95 389.285 207.12 ;
      RECT 392.18 207.44 392.85 207.61 ;
      RECT 390.65 210.325 392.85 210.995 ;
      RECT 392.18 210.15 392.85 210.325 ;
      RECT 390.825 207.54 391.13 210.325 ;
      RECT 391.33 207.34 391.5 210.05 ;
      RECT 392.18 208.22 392.91 209.54 ;
      RECT 392.76 207.855 393.36 208.025 ;
      RECT 393.19 208.025 393.36 208.255 ;
      RECT 393.19 207.585 393.36 207.855 ;
      RECT 393.19 209.68 394.21 209.85 ;
      RECT 393.19 209.85 393.36 210.185 ;
      RECT 393.19 209.515 393.36 209.68 ;
      RECT 393.56 207.41 394.21 209.68 ;
      RECT 396.01 207.41 396.66 209.68 ;
      RECT 396.86 209.85 397.03 210.185 ;
      RECT 396.01 209.68 397.03 209.85 ;
      RECT 396.86 209.515 397.03 209.68 ;
      RECT 397.37 207.44 398.04 207.61 ;
      RECT 397.37 210.325 399.57 210.995 ;
      RECT 397.37 210.15 398.04 210.325 ;
      RECT 399.09 207.54 399.395 210.325 ;
      RECT 398.72 207.34 398.89 210.05 ;
      RECT 401.63 207.34 401.8 210.05 ;
      RECT 397.31 208.22 398.04 209.54 ;
      RECT 226.225 198.815 226.395 205.605 ;
      RECT 228.565 198.815 228.735 205.605 ;
      RECT 238.055 200.085 238.725 200.255 ;
      RECT 238.055 199.685 238.715 200.085 ;
      RECT 240.115 200.085 240.785 200.255 ;
      RECT 244.235 200.085 244.905 200.255 ;
      RECT 242.175 200.085 242.845 200.255 ;
      RECT 250.415 200.085 251.085 200.255 ;
      RECT 248.355 200.085 249.025 200.255 ;
      RECT 246.295 200.085 246.965 200.255 ;
      RECT 254.535 200.085 255.205 200.255 ;
      RECT 252.475 200.085 253.145 200.255 ;
      RECT 256.595 200.085 257.265 200.255 ;
      RECT 260.715 200.085 261.385 200.255 ;
      RECT 262.775 200.085 263.445 200.255 ;
      RECT 258.655 200.085 259.325 200.255 ;
      RECT 268.955 200.085 269.625 200.255 ;
      RECT 266.895 200.085 267.565 200.255 ;
      RECT 264.835 200.085 265.505 200.255 ;
      RECT 273.075 200.085 273.745 200.255 ;
      RECT 271.015 200.085 271.685 200.255 ;
      RECT 271.085 199.3 271.615 200.085 ;
      RECT 272.295 199.685 272.825 200.255 ;
      RECT 274.175 199.3 274.705 200.255 ;
      RECT 277.195 200.085 277.865 200.255 ;
      RECT 279.255 200.085 279.925 200.255 ;
      RECT 275.135 200.085 275.805 200.255 ;
      RECT 280.355 199.685 280.885 200.255 ;
      RECT 278.295 199.3 278.825 200.255 ;
      RECT 276.235 199.685 276.765 200.255 ;
      RECT 283.375 200.085 284.045 200.255 ;
      RECT 281.315 200.085 281.985 200.255 ;
      RECT 285.435 200.085 286.105 200.255 ;
      RECT 284.475 199.685 285.005 200.255 ;
      RECT 282.415 199.3 282.945 200.255 ;
      RECT 291.615 200.085 292.285 200.255 ;
      RECT 289.035 216.18 290.225 216.405 ;
      RECT 289.355 200.085 290.225 200.255 ;
      RECT 289.555 200.255 290.225 216.18 ;
      RECT 287.495 200.085 288.165 200.255 ;
      RECT 288.415 199.685 288.945 200.255 ;
      RECT 286.535 199.3 287.065 200.255 ;
      RECT 293.675 200.085 294.345 200.255 ;
      RECT 295.735 200.085 296.405 200.255 ;
      RECT 297.795 200.085 298.465 200.255 ;
      RECT 301.65 200.085 302.585 200.255 ;
      RECT 299.855 200.085 300.525 200.255 ;
      RECT 312.955 199.965 313.125 214.935 ;
      RECT 314.515 199.965 314.685 214.935 ;
      RECT 310.815 198.455 337.525 199.305 ;
      RECT 315.41 199.305 316.37 199.985 ;
      RECT 319.55 199.305 320.51 199.985 ;
      RECT 323.69 199.305 324.65 199.985 ;
      RECT 327.83 199.305 328.79 199.985 ;
      RECT 331.97 199.305 332.93 199.985 ;
      RECT 315.295 199.985 316.485 214.935 ;
      RECT 319.435 199.985 320.625 214.935 ;
      RECT 323.575 199.985 324.765 214.935 ;
      RECT 327.715 199.985 328.905 214.935 ;
      RECT 331.855 199.985 333.045 214.935 ;
      RECT 315.41 214.935 316.37 215.605 ;
      RECT 319.55 214.935 320.51 215.605 ;
      RECT 323.69 214.935 324.65 215.605 ;
      RECT 327.83 214.935 328.785 215.605 ;
      RECT 331.97 214.935 332.93 215.605 ;
      RECT 310.815 199.305 312.125 199.985 ;
      RECT 310.815 214.935 312.125 215.605 ;
      RECT 335.995 199.985 337.525 214.935 ;
      RECT 336.215 214.935 337.525 215.605 ;
      RECT 336.215 199.305 337.525 199.985 ;
      RECT 310.815 215.605 337.525 218.285 ;
      RECT 310.815 199.985 312.345 214.935 ;
      RECT 312.4 199.505 315.24 199.675 ;
      RECT 317.095 199.965 317.265 214.935 ;
      RECT 318.655 199.965 318.825 214.935 ;
      RECT 320.68 199.505 323.52 199.675 ;
      RECT 320.68 215.155 323.52 215.385 ;
      RECT 323.135 199.675 323.405 215.155 ;
      RECT 316.54 199.505 319.38 199.675 ;
      RECT 325.375 199.965 325.545 214.935 ;
      RECT 322.795 199.965 322.965 214.935 ;
      RECT 321.235 199.965 321.405 214.935 ;
      RECT 324.82 199.505 327.66 199.675 ;
      RECT 324.82 215.155 327.66 215.385 ;
      RECT 324.935 199.675 325.205 215.155 ;
      RECT 326.935 199.965 327.105 214.935 ;
      RECT 329.515 199.965 329.685 214.935 ;
      RECT 331.075 199.965 331.245 214.935 ;
      RECT 328.96 199.505 331.8 199.675 ;
      RECT 335.215 199.965 335.385 214.935 ;
      RECT 333.655 199.965 333.825 214.935 ;
      RECT 333.1 199.505 335.94 199.675 ;
      RECT 349.185 205.1 369.515 205.12 ;
      RECT 349.185 217.345 352.475 223.55 ;
      RECT 368.315 223.34 369.515 223.55 ;
      RECT 368.315 206.33 369.52 223.34 ;
      RECT 349.44 205.07 352.875 205.1 ;
      RECT 349.185 205.12 369.52 206.33 ;
      RECT 349.185 223.55 369.515 224.82 ;
      RECT 349.185 206.33 352.875 217.345 ;
      RECT 430.95 198.725 431.28 199.375 ;
      RECT 435 198.725 435.33 199.375 ;
      RECT 434.19 198.725 434.52 199.375 ;
      RECT 436.62 198.725 436.95 199.375 ;
      RECT 432.57 198.725 432.9 199.375 ;
      RECT 431.76 198.725 432.09 199.375 ;
      RECT 435.81 198.725 436.14 199.375 ;
      RECT 433.38 198.725 433.71 199.375 ;
      RECT 438.24 198.725 438.57 199.375 ;
      RECT 437.43 198.725 437.76 199.375 ;
      RECT 439.86 198.725 440.19 199.375 ;
      RECT 439.05 198.725 439.38 199.375 ;
      RECT 440.67 198.725 441 199.375 ;
      RECT 445.625 201.28 445.855 206.125 ;
      RECT 445.625 215.23 445.855 219.275 ;
      RECT 445.625 232.32 445.855 233.7 ;
      RECT 445.625 199.915 466.45 200.145 ;
      RECT 445.625 233.7 466.45 233.93 ;
      RECT 445.655 200.145 445.825 201.28 ;
      RECT 466.22 200.145 466.45 211.185 ;
      RECT 445.655 211.91 445.825 215.23 ;
      RECT 445.625 211.415 445.855 211.91 ;
      RECT 445.655 206.125 445.825 209.62 ;
      RECT 445.625 209.62 445.855 211.185 ;
      RECT 445.625 222.67 445.855 229.45 ;
      RECT 445.655 219.275 445.825 222.44 ;
      RECT 466.22 211.415 466.45 222.44 ;
      RECT 69.495 199.305 70.455 199.985 ;
      RECT 73.635 199.305 74.595 199.985 ;
      RECT 65.24 199.985 66.43 214.935 ;
      RECT 61.1 199.985 62.29 214.935 ;
      RECT 69.38 199.985 70.57 214.935 ;
      RECT 73.52 199.985 74.71 214.935 ;
      RECT 57.075 214.935 58.035 215.605 ;
      RECT 65.355 214.935 66.315 215.605 ;
      RECT 61.22 214.935 62.175 215.605 ;
      RECT 69.495 214.935 70.455 215.605 ;
      RECT 73.635 214.935 74.595 215.605 ;
      RECT 52.48 199.985 54.01 214.935 ;
      RECT 77.88 199.305 79.19 199.985 ;
      RECT 52.48 214.935 53.79 215.605 ;
      RECT 52.48 199.305 53.79 199.985 ;
      RECT 77.88 214.935 79.19 215.605 ;
      RECT 52.48 215.605 79.19 218.285 ;
      RECT 77.66 199.985 79.19 214.935 ;
      RECT 64.46 199.965 64.63 214.935 ;
      RECT 62.9 199.965 63.07 214.935 ;
      RECT 62.345 199.505 65.185 199.675 ;
      RECT 62.345 215.155 65.185 215.385 ;
      RECT 64.8 199.675 65.07 215.155 ;
      RECT 67.04 199.965 67.21 214.935 ;
      RECT 68.6 199.965 68.77 214.935 ;
      RECT 71.18 199.965 71.35 214.935 ;
      RECT 70.625 199.505 73.465 199.675 ;
      RECT 66.485 199.505 69.325 199.675 ;
      RECT 66.485 215.155 69.325 215.385 ;
      RECT 66.6 199.675 66.87 215.155 ;
      RECT 76.88 199.965 77.05 214.935 ;
      RECT 75.32 199.965 75.49 214.935 ;
      RECT 72.74 199.965 72.91 214.935 ;
      RECT 74.765 199.505 77.605 199.675 ;
      RECT 87.42 200.085 88.355 200.255 ;
      RECT 93.6 200.085 94.27 200.255 ;
      RECT 89.48 200.085 90.15 200.255 ;
      RECT 91.54 200.085 92.21 200.255 ;
      RECT 97.72 200.085 98.39 200.255 ;
      RECT 95.66 200.085 96.33 200.255 ;
      RECT 99.78 216.18 100.97 216.405 ;
      RECT 99.78 200.085 100.65 200.255 ;
      RECT 99.78 200.255 100.45 216.18 ;
      RECT 105.96 200.085 106.63 200.255 ;
      RECT 101.84 200.085 102.51 200.255 ;
      RECT 103.9 200.085 104.57 200.255 ;
      RECT 101.06 199.685 101.59 200.255 ;
      RECT 102.94 199.3 103.47 200.255 ;
      RECT 105 199.685 105.53 200.255 ;
      RECT 112.14 200.085 112.81 200.255 ;
      RECT 110.08 200.085 110.75 200.255 ;
      RECT 108.02 200.085 108.69 200.255 ;
      RECT 107.06 199.3 107.59 200.255 ;
      RECT 109.12 199.685 109.65 200.255 ;
      RECT 111.18 199.3 111.71 200.255 ;
      RECT 116.26 200.085 116.93 200.255 ;
      RECT 114.2 200.085 114.87 200.255 ;
      RECT 118.32 200.085 118.99 200.255 ;
      RECT 118.39 199.3 118.92 200.085 ;
      RECT 117.18 199.685 117.71 200.255 ;
      RECT 113.24 199.685 113.77 200.255 ;
      RECT 115.3 199.3 115.83 200.255 ;
      RECT 122.44 200.085 123.11 200.255 ;
      RECT 120.38 200.085 121.05 200.255 ;
      RECT 128.62 200.085 129.29 200.255 ;
      RECT 126.56 200.085 127.23 200.255 ;
      RECT 124.5 200.085 125.17 200.255 ;
      RECT 132.74 200.085 133.41 200.255 ;
      RECT 130.68 200.085 131.35 200.255 ;
      RECT 134.8 200.085 135.47 200.255 ;
      RECT 138.92 200.085 139.59 200.255 ;
      RECT 136.86 200.085 137.53 200.255 ;
      RECT 140.98 200.085 141.65 200.255 ;
      RECT 145.1 200.085 145.77 200.255 ;
      RECT 147.16 200.085 147.83 200.255 ;
      RECT 143.04 200.085 143.71 200.255 ;
      RECT 149.22 200.085 149.89 200.255 ;
      RECT 151.28 200.085 151.95 200.255 ;
      RECT 151.29 199.685 151.95 200.085 ;
      RECT 164.39 198.815 164.56 205.605 ;
      RECT 161.27 198.815 161.44 205.605 ;
      RECT 162.83 198.815 163 205.605 ;
      RECT 162.05 198.815 162.22 205.605 ;
      RECT 163.61 198.815 163.78 205.605 ;
      RECT 165.55 204.255 170.42 204.425 ;
      RECT 165.55 203.705 170.425 203.875 ;
      RECT 165.55 202.925 170.425 203.095 ;
      RECT 165.55 198.705 170.425 198.875 ;
      RECT 165.55 200.265 170.425 200.435 ;
      RECT 165.55 202.375 170.425 202.545 ;
      RECT 165.55 200.815 170.425 200.985 ;
      RECT 165.55 205.815 170.42 205.985 ;
      RECT 165.55 205.035 170.425 205.205 ;
      RECT 165.55 199.485 170.425 199.655 ;
      RECT 165.55 201.595 170.425 201.765 ;
      RECT 170.685 199.005 170.98 200.255 ;
      RECT 170.81 200.255 170.98 200.28 ;
      RECT 170.81 198.93 170.98 199.005 ;
      RECT 170.685 201.02 170.98 202.27 ;
      RECT 170.81 202.27 170.98 202.32 ;
      RECT 170.81 200.97 170.98 201.02 ;
      RECT 170.675 204.48 170.98 205.76 ;
      RECT 170.705 204.205 170.875 204.48 ;
      RECT 170.675 203.15 170.98 203.82 ;
      RECT 219.025 199.005 219.32 200.255 ;
      RECT 219.025 200.255 219.195 200.28 ;
      RECT 219.025 198.93 219.195 199.005 ;
      RECT 219.025 201.02 219.32 202.27 ;
      RECT 219.025 202.27 219.195 202.32 ;
      RECT 219.025 200.97 219.195 201.02 ;
      RECT 219.58 203.705 224.455 203.875 ;
      RECT 219.58 202.925 224.455 203.095 ;
      RECT 219.58 198.705 224.455 198.875 ;
      RECT 219.58 200.265 224.455 200.435 ;
      RECT 219.58 202.375 224.455 202.545 ;
      RECT 219.58 200.815 224.455 200.985 ;
      RECT 219.585 205.815 224.455 205.985 ;
      RECT 219.585 204.255 224.455 204.425 ;
      RECT 219.025 204.48 219.33 205.76 ;
      RECT 219.13 204.205 219.3 204.48 ;
      RECT 219.025 203.15 219.33 203.82 ;
      RECT 219.58 205.035 224.455 205.205 ;
      RECT 219.58 199.485 224.455 199.655 ;
      RECT 219.58 201.595 224.455 201.765 ;
      RECT 225.445 198.815 225.615 205.605 ;
      RECT 227.005 198.815 227.175 205.605 ;
      RECT 227.785 198.815 227.955 205.605 ;
      RECT 144.02 192.7 144.56 192.87 ;
      RECT 144.05 192.87 144.56 192.95 ;
      RECT 144.05 192.62 144.56 192.7 ;
      RECT 144.34 190.925 153.64 191.365 ;
      RECT 140.19 191.365 155.14 191.535 ;
      RECT 161.56 198.425 164.27 198.595 ;
      RECT 161.56 205.815 164.27 206.245 ;
      RECT 161.61 198.595 161.88 205.815 ;
      RECT 162.39 198.595 162.66 205.815 ;
      RECT 163.17 198.595 163.44 205.815 ;
      RECT 163.95 198.595 164.22 205.815 ;
      RECT 163.435 192.285 164.105 193.605 ;
      RECT 163.435 193.605 169.14 194.135 ;
      RECT 159.745 197.515 160.075 198.485 ;
      RECT 164.97 217.81 169.42 217.98 ;
      RECT 159.745 198.485 160.86 198.655 ;
      RECT 160.69 198.655 160.86 213.855 ;
      RECT 160.69 198.235 160.86 198.485 ;
      RECT 164.97 198.235 165.14 206.44 ;
      RECT 160.69 198.065 171.34 198.235 ;
      RECT 160.69 213.855 165.14 214.025 ;
      RECT 164.97 206.44 171.34 206.61 ;
      RECT 169.25 206.61 169.42 217.81 ;
      RECT 164.97 214.025 165.14 217.81 ;
      RECT 164.97 206.61 165.14 213.855 ;
      RECT 171.17 198.235 171.34 206.44 ;
      RECT 167.275 192.395 167.945 192.875 ;
      RECT 167.275 192.875 169.14 193.405 ;
      RECT 171.125 192.395 171.795 192.565 ;
      RECT 172.405 192.395 173.075 192.565 ;
      RECT 222.06 192.395 222.73 192.875 ;
      RECT 220.865 192.875 222.73 193.405 ;
      RECT 218.21 192.395 218.88 192.565 ;
      RECT 216.93 192.395 217.6 192.565 ;
      RECT 220.585 217.81 225.035 217.98 ;
      RECT 229.93 197.515 230.26 198.485 ;
      RECT 218.665 198.065 229.315 198.235 ;
      RECT 229.145 198.655 229.315 213.855 ;
      RECT 229.145 198.235 229.315 198.485 ;
      RECT 224.865 214.025 225.035 217.81 ;
      RECT 229.145 198.485 230.26 198.655 ;
      RECT 218.665 198.235 218.835 206.44 ;
      RECT 218.665 206.44 225.035 206.61 ;
      RECT 220.585 206.61 220.755 217.81 ;
      RECT 224.865 206.61 225.035 213.855 ;
      RECT 224.865 213.855 229.315 214.025 ;
      RECT 224.865 198.235 225.035 206.44 ;
      RECT 220.865 193.605 226.57 194.135 ;
      RECT 225.9 192.285 226.57 193.605 ;
      RECT 225.735 198.425 228.445 198.595 ;
      RECT 225.735 205.815 228.445 206.245 ;
      RECT 225.785 198.595 226.055 205.815 ;
      RECT 226.565 198.595 226.835 205.815 ;
      RECT 227.345 198.595 227.615 205.815 ;
      RECT 228.125 198.595 228.395 205.815 ;
      RECT 245.445 192.7 245.985 192.87 ;
      RECT 245.445 192.87 245.955 192.95 ;
      RECT 245.445 192.62 245.955 192.7 ;
      RECT 250.035 191.195 250.545 191.225 ;
      RECT 245.835 190.925 250.545 191.195 ;
      RECT 250.035 190.895 250.545 190.925 ;
      RECT 236.365 190.925 245.665 191.365 ;
      RECT 234.865 191.365 249.815 191.535 ;
      RECT 267.405 191.195 267.915 191.225 ;
      RECT 263.205 190.925 267.915 191.195 ;
      RECT 267.405 190.895 267.915 190.925 ;
      RECT 253.735 190.925 263.035 191.365 ;
      RECT 252.235 191.365 267.185 191.535 ;
      RECT 284.145 192.96 288.165 193.71 ;
      RECT 308.58 193.74 308.75 193.855 ;
      RECT 308.58 192.845 308.75 192.97 ;
      RECT 304.85 192.97 308.75 193.74 ;
      RECT 304.85 193.74 305.18 193.775 ;
      RECT 304.85 192.925 305.18 192.97 ;
      RECT 305.32 192.63 308.105 192.8 ;
      RECT 310.59 193.68 311.125 193.85 ;
      RECT 310.595 193.85 311.125 193.965 ;
      RECT 310.595 193.605 311.125 193.68 ;
      RECT 310.23 191.55 310.4 192.22 ;
      RECT 321.315 193.685 321.875 193.855 ;
      RECT 321.315 193.855 321.825 193.935 ;
      RECT 321.315 193.605 321.825 193.685 ;
      RECT 341.595 192.15 341.765 192.22 ;
      RECT 341.58 191.62 341.765 192.15 ;
      RECT 341.595 191.55 341.765 191.62 ;
      RECT 360.915 192.22 361.085 193.23 ;
      RECT 356.635 192.22 356.805 193.23 ;
      RECT 356.86 191.62 360.86 191.79 ;
      RECT 361.14 191.62 369.14 191.79 ;
      RECT 356.86 193.48 360.86 193.65 ;
      RECT 368.37 194.885 369.38 195.055 ;
      RECT 368.37 194.005 369.38 194.175 ;
      RECT 368.48 194.175 369.325 194.18 ;
      RECT 369.195 192.22 369.365 193.23 ;
      RECT 367.98 194.23 368.15 194.9 ;
      RECT 387.7 197.84 388.03 198.49 ;
      RECT 389.59 197.84 389.92 198.49 ;
      RECT 388.33 197.84 388.66 198.49 ;
      RECT 388.96 197.84 389.29 198.49 ;
      RECT 390.22 197.84 390.55 198.49 ;
      RECT 395.03 194.52 395.365 198.25 ;
      RECT 390.85 197.84 391.18 198.49 ;
      RECT 405.63 194.52 405.8 198.25 ;
      RECT 416.28 194.52 416.45 198.25 ;
      RECT 426.725 194.52 427.05 198.25 ;
      RECT 445.98 194.525 446.15 198.525 ;
      RECT 446.56 194.3 456.41 194.47 ;
      RECT 446.56 198.58 456.41 198.75 ;
      RECT 20.49 205.1 40.82 205.12 ;
      RECT 20.49 223.55 40.82 224.82 ;
      RECT 37.13 205.07 40.565 205.1 ;
      RECT 20.49 223.34 21.69 223.55 ;
      RECT 20.485 206.33 21.69 223.34 ;
      RECT 37.53 217.345 40.82 223.55 ;
      RECT 20.485 205.12 40.82 206.33 ;
      RECT 37.13 206.33 40.82 217.345 ;
      RECT 54.62 199.965 54.79 214.935 ;
      RECT 54.065 199.505 56.905 199.675 ;
      RECT 56.18 199.965 56.35 214.935 ;
      RECT 60.32 199.965 60.49 214.935 ;
      RECT 58.76 199.965 58.93 214.935 ;
      RECT 58.205 199.505 61.045 199.675 ;
      RECT 57.075 199.305 58.035 199.985 ;
      RECT 56.96 199.985 58.15 214.935 ;
      RECT 52.48 198.455 79.19 199.305 ;
      RECT 65.355 199.305 66.315 199.985 ;
      RECT 61.215 199.305 62.175 199.985 ;
      RECT 365.315 187.325 365.885 187.495 ;
      RECT 365.315 187.495 365.485 187.55 ;
      RECT 365.315 187.22 365.485 187.325 ;
      RECT 366.015 183.955 366.185 185.625 ;
      RECT 365.655 183.785 366.185 183.955 ;
      RECT 364.665 184.125 365.635 184.375 ;
      RECT 364.665 184.375 364.975 185.455 ;
      RECT 363.925 185.455 364.975 185.625 ;
      RECT 367.3 186.95 367.83 187.12 ;
      RECT 367.54 187.12 367.82 187.555 ;
      RECT 365.48 187.77 369.63 187.94 ;
      RECT 365.79 189.63 367.79 189.8 ;
      RECT 365.85 189.8 367.72 189.81 ;
      RECT 368.805 187.22 370.045 187.55 ;
      RECT 367.68 189.16 368.21 189.33 ;
      RECT 367.845 189.33 368.015 189.41 ;
      RECT 367.845 189.08 368.015 189.16 ;
      RECT 369.195 190.36 369.365 191.37 ;
      RECT 376.275 182.95 376.605 183.55 ;
      RECT 377.085 182.95 377.415 183.55 ;
      RECT 375.465 182.95 375.795 183.555 ;
      RECT 377.895 182.95 378.225 183.55 ;
      RECT 378.705 182.95 379.035 183.55 ;
      RECT 379.515 182.95 379.845 183.54 ;
      RECT 389.59 188.795 389.92 189.445 ;
      RECT 388.33 188.795 388.66 189.445 ;
      RECT 388.96 188.795 389.29 189.445 ;
      RECT 390.22 188.795 390.55 189.445 ;
      RECT 387.7 187.765 388.03 188.415 ;
      RECT 389.59 187.765 389.92 188.415 ;
      RECT 390.22 187.765 390.55 188.415 ;
      RECT 388.96 187.765 389.29 188.415 ;
      RECT 388.33 187.765 388.66 188.415 ;
      RECT 387.7 188.795 388.03 189.445 ;
      RECT 395.03 190.24 395.365 193.97 ;
      RECT 394.98 183.61 395.15 188.37 ;
      RECT 395.86 183.61 396.03 188.36 ;
      RECT 395.205 188.87 396.685 189.04 ;
      RECT 395.69 188.53 396.22 188.87 ;
      RECT 390.85 188.795 391.18 189.445 ;
      RECT 390.85 187.765 391.18 188.415 ;
      RECT 394.61 199.02 427.47 199.2 ;
      RECT 427.29 183.135 427.47 189.29 ;
      RECT 427.29 189.47 427.47 199.02 ;
      RECT 395.56 198.44 426.71 199.02 ;
      RECT 394.39 189.29 427.47 189.47 ;
      RECT 394.39 183.135 394.57 189.29 ;
      RECT 395.56 190.05 415.82 194.16 ;
      RECT 406.28 194.33 415.82 198.44 ;
      RECT 416.88 190.05 426.12 194.16 ;
      RECT 395.56 194.16 426.71 194.33 ;
      RECT 416.88 194.33 426.12 198.44 ;
      RECT 395.56 189.47 426.71 190.05 ;
      RECT 395.56 194.33 405.395 198.44 ;
      RECT 394.61 189.47 394.79 199.02 ;
      RECT 413.37 188.87 414.04 189.29 ;
      RECT 394.39 182.955 427.47 183.135 ;
      RECT 399.3 183.61 399.47 188.37 ;
      RECT 396.74 183.61 396.91 188.37 ;
      RECT 401.86 183.61 402.03 188.37 ;
      RECT 397.03 188.87 406.76 189.04 ;
      RECT 398.02 183.61 398.19 188.36 ;
      RECT 400.58 183.61 400.75 188.36 ;
      RECT 407.86 183.61 408.03 188.36 ;
      RECT 406.98 183.61 407.15 188.37 ;
      RECT 404.42 183.61 404.59 188.37 ;
      RECT 407.34 188.87 407.67 189.04 ;
      RECT 407.42 188.11 407.59 188.87 ;
      RECT 405.7 183.61 405.87 188.36 ;
      RECT 403.14 183.61 403.31 188.36 ;
      RECT 412.98 183.61 413.15 188.37 ;
      RECT 410.42 183.61 410.59 188.37 ;
      RECT 408.25 188.87 412.905 189.04 ;
      RECT 409.14 183.61 409.31 188.36 ;
      RECT 411.7 183.61 411.87 188.36 ;
      RECT 416.28 190.24 416.45 193.97 ;
      RECT 418.1 183.61 418.27 188.475 ;
      RECT 415.54 183.61 415.71 188.37 ;
      RECT 418.44 188.87 425.56 189.04 ;
      RECT 414.5 188.87 417.88 189.04 ;
      RECT 419.38 183.61 419.55 188.36 ;
      RECT 416.82 183.61 416.99 188.36 ;
      RECT 414.26 183.61 414.43 188.36 ;
      RECT 423.22 183.61 423.39 188.475 ;
      RECT 420.66 183.61 420.83 188.475 ;
      RECT 421.94 183.61 422.11 188.36 ;
      RECT 424.5 183.61 424.67 188.36 ;
      RECT 426.725 190.24 427.05 193.97 ;
      RECT 425.78 183.61 425.95 188.475 ;
      RECT 426.56 183.61 426.73 188.475 ;
      RECT 426.93 188.11 427.1 188.87 ;
      RECT 426.005 188.87 427.1 189.04 ;
      RECT 20.625 194.885 21.635 195.055 ;
      RECT 20.625 194.005 21.635 194.175 ;
      RECT 20.68 194.175 21.525 194.18 ;
      RECT 20.64 192.22 20.81 193.23 ;
      RECT 20.865 191.62 28.865 191.79 ;
      RECT 21.855 194.23 22.025 194.9 ;
      RECT 28.92 192.22 29.09 193.23 ;
      RECT 29.145 191.62 33.145 191.79 ;
      RECT 29.145 193.48 33.145 193.65 ;
      RECT 33.2 192.22 33.37 193.23 ;
      RECT 48.24 192.15 48.41 192.22 ;
      RECT 48.24 191.62 48.425 192.15 ;
      RECT 48.24 191.55 48.41 191.62 ;
      RECT 68.13 193.685 68.69 193.855 ;
      RECT 68.18 193.855 68.69 193.935 ;
      RECT 68.18 193.605 68.69 193.685 ;
      RECT 78.88 193.68 79.415 193.85 ;
      RECT 78.88 193.85 79.41 193.965 ;
      RECT 78.88 193.605 79.41 193.68 ;
      RECT 81.255 193.74 81.425 193.855 ;
      RECT 81.255 192.845 81.425 192.97 ;
      RECT 81.255 192.97 85.155 193.74 ;
      RECT 84.825 193.74 85.155 193.775 ;
      RECT 84.825 192.925 85.155 192.97 ;
      RECT 79.605 191.55 79.775 192.22 ;
      RECT 81.9 192.63 84.685 192.8 ;
      RECT 101.84 192.96 105.86 193.71 ;
      RECT 122.09 190.925 126.8 191.195 ;
      RECT 122.09 191.195 122.6 191.225 ;
      RECT 122.09 190.895 122.6 190.925 ;
      RECT 126.97 190.925 136.27 191.365 ;
      RECT 122.82 191.365 137.77 191.535 ;
      RECT 139.46 190.925 144.17 191.195 ;
      RECT 139.46 191.195 139.97 191.225 ;
      RECT 139.46 190.895 139.97 190.925 ;
      RECT 26.255 189.005 28.965 189.175 ;
      RECT 26.04 187.245 28.965 187.415 ;
      RECT 28.92 190.36 29.09 191.37 ;
      RECT 29.185 188.35 29.355 189.02 ;
      RECT 29.185 187.4 29.355 188.07 ;
      RECT 35.605 183.62 42.115 183.79 ;
      RECT 33.2 190.94 33.785 191.11 ;
      RECT 33.2 191.11 33.37 191.37 ;
      RECT 33.2 190.36 33.37 190.94 ;
      RECT 48.24 190.41 48.41 190.48 ;
      RECT 48.24 189.88 48.425 190.41 ;
      RECT 48.24 189.81 48.41 189.88 ;
      RECT 48.24 186.33 48.41 186.475 ;
      RECT 48.255 187 48.425 187.005 ;
      RECT 48.24 186.475 48.425 187 ;
      RECT 48.24 188.14 48.425 188.67 ;
      RECT 48.24 188.67 48.41 188.74 ;
      RECT 48.24 188.07 48.41 188.14 ;
      RECT 79.605 188.07 79.775 188.74 ;
      RECT 79.605 189.805 79.775 190.475 ;
      RECT 79.605 186.33 79.775 187 ;
      RECT 101.84 186.39 105.86 187.365 ;
      RECT 122.09 190.145 124.65 190.415 ;
      RECT 122.09 190.415 122.6 190.445 ;
      RECT 122.09 190.115 122.6 190.145 ;
      RECT 122.91 186.175 137.86 186.345 ;
      RECT 126.97 189.975 136.27 190.415 ;
      RECT 122.82 189.805 137.77 189.975 ;
      RECT 122.82 190.585 137.77 190.755 ;
      RECT 138.08 186.005 138.59 186.035 ;
      RECT 133.88 185.735 138.59 186.005 ;
      RECT 138.08 185.705 138.59 185.735 ;
      RECT 124.41 185.565 133.71 186.005 ;
      RECT 122.91 185.395 137.86 185.565 ;
      RECT 124.41 186.515 133.71 186.955 ;
      RECT 122.91 186.955 137.86 187.125 ;
      RECT 139.46 190.145 142.02 190.415 ;
      RECT 139.46 190.415 139.97 190.445 ;
      RECT 139.46 190.115 139.97 190.145 ;
      RECT 139.46 185.735 144.17 186.005 ;
      RECT 139.46 186.005 139.97 186.035 ;
      RECT 139.46 185.705 139.97 185.735 ;
      RECT 139.46 186.515 142.02 186.785 ;
      RECT 139.46 186.785 139.97 186.815 ;
      RECT 139.46 186.485 139.97 186.515 ;
      RECT 136.03 186.515 138.59 186.785 ;
      RECT 138.08 186.785 138.59 186.815 ;
      RECT 138.08 186.485 138.59 186.515 ;
      RECT 144.34 185.565 153.64 186.005 ;
      RECT 140.19 185.395 155.14 185.565 ;
      RECT 144.34 189.975 153.64 190.415 ;
      RECT 140.19 189.805 155.14 189.975 ;
      RECT 144.34 186.515 153.64 186.955 ;
      RECT 140.19 186.955 155.14 187.125 ;
      RECT 140.19 190.585 155.14 190.755 ;
      RECT 140.19 186.175 155.14 186.345 ;
      RECT 169.845 186.225 170.515 188.785 ;
      RECT 169.76 184.235 171.78 184.985 ;
      RECT 168.555 189.915 169.225 192.565 ;
      RECT 169.845 189.915 170.515 192.565 ;
      RECT 219.49 186.225 220.16 188.785 ;
      RECT 218.225 184.235 220.245 184.985 ;
      RECT 220.78 189.915 221.45 192.565 ;
      RECT 219.49 189.915 220.16 192.565 ;
      RECT 234.865 190.585 249.815 190.755 ;
      RECT 234.865 186.175 249.815 186.345 ;
      RECT 236.365 186.515 245.665 186.955 ;
      RECT 234.865 186.955 249.815 187.125 ;
      RECT 250.035 186.005 250.545 186.035 ;
      RECT 245.835 185.735 250.545 186.005 ;
      RECT 250.035 185.705 250.545 185.735 ;
      RECT 236.365 185.565 245.665 186.005 ;
      RECT 234.865 185.395 249.815 185.565 ;
      RECT 236.365 189.975 245.665 190.415 ;
      RECT 234.865 189.805 249.815 189.975 ;
      RECT 247.985 190.145 250.545 190.415 ;
      RECT 250.035 190.415 250.545 190.445 ;
      RECT 250.035 190.115 250.545 190.145 ;
      RECT 247.985 186.515 250.545 186.785 ;
      RECT 250.035 186.785 250.545 186.815 ;
      RECT 250.035 186.485 250.545 186.515 ;
      RECT 251.415 185.735 256.125 186.005 ;
      RECT 251.415 186.005 251.925 186.035 ;
      RECT 251.415 185.705 251.925 185.735 ;
      RECT 251.415 186.515 253.975 186.785 ;
      RECT 251.415 186.785 251.925 186.815 ;
      RECT 251.415 186.485 251.925 186.515 ;
      RECT 252.235 190.585 267.185 190.755 ;
      RECT 256.295 186.515 265.595 186.955 ;
      RECT 252.145 186.955 267.095 187.125 ;
      RECT 252.145 186.175 267.095 186.345 ;
      RECT 256.295 185.565 265.595 186.005 ;
      RECT 252.145 185.395 267.095 185.565 ;
      RECT 253.735 189.975 263.035 190.415 ;
      RECT 252.235 189.805 267.185 189.975 ;
      RECT 265.355 190.145 267.915 190.415 ;
      RECT 267.405 190.415 267.915 190.445 ;
      RECT 267.405 190.115 267.915 190.145 ;
      RECT 284.145 186.39 288.165 187.365 ;
      RECT 310.23 186.33 310.4 187 ;
      RECT 310.23 188.07 310.4 188.74 ;
      RECT 310.23 189.805 310.4 190.475 ;
      RECT 341.595 190.41 341.765 190.48 ;
      RECT 341.58 189.88 341.765 190.41 ;
      RECT 341.595 189.81 341.765 189.88 ;
      RECT 341.595 186.33 341.765 186.475 ;
      RECT 341.58 187 341.75 187.005 ;
      RECT 341.58 186.475 341.765 187 ;
      RECT 341.58 188.14 341.765 188.67 ;
      RECT 341.595 188.67 341.765 188.74 ;
      RECT 341.595 188.07 341.765 188.14 ;
      RECT 347.89 183.62 354.4 183.79 ;
      RECT 361.04 188.125 364 188.295 ;
      RECT 361.04 189.005 363.75 189.175 ;
      RECT 361.04 187.245 363.965 187.415 ;
      RECT 360.915 190.36 361.085 191.37 ;
      RECT 356.22 190.94 356.805 191.11 ;
      RECT 356.635 191.11 356.805 191.37 ;
      RECT 356.635 190.36 356.805 190.94 ;
      RECT 360.65 188.35 360.82 189.02 ;
      RECT 360.65 187.4 360.82 188.07 ;
      RECT 365.175 184.645 365.705 185.655 ;
      RECT 365.345 184.635 365.515 184.645 ;
      RECT 362.9 183.725 363.07 185.625 ;
      RECT 362.725 183.145 363.255 183.725 ;
      RECT 362.465 184.635 362.635 185.685 ;
      RECT 365.565 188.455 365.735 189.41 ;
      RECT 367.715 179.455 367.885 179.895 ;
      RECT 367.135 180.36 367.885 180.975 ;
      RECT 363.555 182.795 363.725 183.275 ;
      RECT 363.555 183.945 363.725 184.675 ;
      RECT 363.555 182.465 363.915 182.795 ;
      RECT 363.555 183.275 364.085 183.945 ;
      RECT 363.345 184.675 363.725 185.685 ;
      RECT 362.465 182.265 363.3 182.795 ;
      RECT 362.465 181.885 363.885 182.265 ;
      RECT 362.54 179.575 362.71 179.625 ;
      RECT 362.51 179.625 362.71 180.825 ;
      RECT 362.51 180.825 362.68 180.975 ;
      RECT 363.29 181.145 365.02 181.315 ;
      RECT 363.29 179.625 363.46 181.145 ;
      RECT 364.85 179.625 365.02 181.145 ;
      RECT 365.175 182.265 366.225 182.895 ;
      RECT 365.175 181.885 366.935 182.265 ;
      RECT 363.895 184.585 364.465 184.915 ;
      RECT 364.295 181.885 364.465 183.385 ;
      RECT 364.295 183.385 366.34 183.555 ;
      RECT 364.295 183.555 364.915 183.725 ;
      RECT 364.295 183.725 364.465 184.585 ;
      RECT 363.895 184.915 364.065 184.975 ;
      RECT 366.58 182.465 367.005 182.795 ;
      RECT 366.58 182.795 366.75 183.275 ;
      RECT 366.58 183.275 366.865 183.945 ;
      RECT 366.58 183.945 366.75 184.645 ;
      RECT 366.395 184.645 366.75 185.655 ;
      RECT 387.7 178.72 388.03 179.37 ;
      RECT 389.59 178.72 389.92 179.37 ;
      RECT 390.22 178.72 390.55 179.37 ;
      RECT 388.96 178.72 389.29 179.37 ;
      RECT 388.33 178.72 388.66 179.37 ;
      RECT 387.7 177.69 388.03 178.34 ;
      RECT 388.96 177.69 389.29 178.34 ;
      RECT 388.33 177.69 388.66 178.34 ;
      RECT 389.59 177.69 389.92 178.34 ;
      RECT 390.22 177.69 390.55 178.34 ;
      RECT 396.2 180.455 399.77 180.785 ;
      RECT 395.76 175.275 395.93 180.125 ;
      RECT 390.85 178.72 391.18 179.37 ;
      RECT 390.85 177.69 391.18 178.34 ;
      RECT 400.48 180.455 404.05 180.785 ;
      RECT 400.04 175.275 400.21 180.125 ;
      RECT 404.32 175.275 404.49 180.125 ;
      RECT 413.66 180.455 417.23 180.785 ;
      RECT 409.38 180.455 412.95 180.785 ;
      RECT 408.94 175.275 409.11 180.125 ;
      RECT 413.22 175.275 413.39 180.125 ;
      RECT 417.5 175.275 417.67 180.125 ;
      RECT 425.28 179.535 425.61 180.185 ;
      RECT 423.66 179.535 423.99 180.185 ;
      RECT 424.47 179.535 424.8 180.185 ;
      RECT 422.85 179.535 423.18 180.185 ;
      RECT 422.04 179.535 422.37 180.185 ;
      RECT 421.18 181.095 423.525 181.84 ;
      RECT 430.14 179.535 430.47 180.185 ;
      RECT 430.95 179.535 431.28 180.185 ;
      RECT 429.33 179.535 429.66 180.185 ;
      RECT 428.52 179.535 428.85 180.185 ;
      RECT 427.71 179.535 428.04 180.185 ;
      RECT 426.9 179.535 427.23 180.185 ;
      RECT 426.09 179.535 426.42 180.185 ;
      RECT 431.76 179.535 432.09 180.185 ;
      RECT 432.57 179.535 432.9 180.185 ;
      RECT 435 179.535 435.33 180.185 ;
      RECT 433.38 179.535 433.71 180.185 ;
      RECT 434.19 179.535 434.52 180.185 ;
      RECT 436.62 179.535 436.95 180.185 ;
      RECT 435.81 179.535 436.14 180.185 ;
      RECT 438.24 179.535 438.57 180.185 ;
      RECT 437.43 179.535 437.76 180.185 ;
      RECT 439.86 179.535 440.19 180.185 ;
      RECT 439.05 179.535 439.38 180.185 ;
      RECT 440.67 179.535 441 180.185 ;
      RECT 450.32 176.255 456.455 176.785 ;
      RECT 450.32 180.685 456.455 181.215 ;
      RECT 450.32 175.545 456.025 176.075 ;
      RECT 450.32 179.975 456.025 180.505 ;
      RECT 450.32 179.07 455.595 179.6 ;
      RECT 448.865 176.14 449.875 176.31 ;
      RECT 448.865 175.26 449.875 175.43 ;
      RECT 448.865 176.965 458.585 177.23 ;
      RECT 448.865 180.57 449.875 180.74 ;
      RECT 448.865 179.69 449.875 179.86 ;
      RECT 448.865 177.89 458.585 178.155 ;
      RECT 448.865 178.81 449.875 178.98 ;
      RECT 448.865 181.395 458.585 181.66 ;
      RECT 456.695 175.205 458.575 175.485 ;
      RECT 457.565 178.755 459.345 179.035 ;
      RECT 459.095 177.74 459.345 178.755 ;
      RECT 459.095 180.795 459.345 181.81 ;
      RECT 457.565 180.515 459.345 180.795 ;
      RECT 459.095 179.035 459.345 180.515 ;
      RECT 456.695 179.635 458.575 179.915 ;
      RECT 456.675 178.37 457.345 178.54 ;
      RECT 13.4 182.95 13.73 183.55 ;
      RECT 12.59 182.95 12.92 183.55 ;
      RECT 11.78 182.95 12.11 183.55 ;
      RECT 10.97 182.95 11.3 183.55 ;
      RECT 10.16 182.95 10.49 183.54 ;
      RECT 14.21 182.95 14.54 183.555 ;
      RECT 24.3 184.645 24.83 185.655 ;
      RECT 24.49 184.635 24.66 184.645 ;
      RECT 24.27 188.455 24.44 189.41 ;
      RECT 21.795 189.16 22.325 189.33 ;
      RECT 21.99 189.33 22.16 189.41 ;
      RECT 21.99 189.08 22.16 189.16 ;
      RECT 24.12 187.325 24.69 187.495 ;
      RECT 24.52 187.495 24.69 187.55 ;
      RECT 24.52 187.22 24.69 187.325 ;
      RECT 19.96 187.22 21.2 187.55 ;
      RECT 23.82 183.955 23.99 185.625 ;
      RECT 23.82 183.785 24.35 183.955 ;
      RECT 24.37 184.125 25.34 184.375 ;
      RECT 25.03 184.375 25.34 185.455 ;
      RECT 25.03 185.455 26.08 185.625 ;
      RECT 20.64 190.36 20.81 191.37 ;
      RECT 22.175 186.95 22.705 187.12 ;
      RECT 22.185 187.12 22.465 187.555 ;
      RECT 20.375 187.77 24.525 187.94 ;
      RECT 22.215 189.63 24.215 189.8 ;
      RECT 22.285 189.8 24.155 189.81 ;
      RECT 26.935 183.725 27.105 185.625 ;
      RECT 26.75 183.145 27.28 183.725 ;
      RECT 27.37 184.635 27.54 185.685 ;
      RECT 26.005 188.125 28.965 188.295 ;
      RECT 231.155 183.525 249.755 184.375 ;
      RECT 268.94 180.515 293.52 183.71 ;
      RECT 267.665 180.175 293.52 180.515 ;
      RECT 231.155 179.155 293.52 180.175 ;
      RECT 231.155 180.175 234.11 183.525 ;
      RECT 225.85 251.735 346.52 251.76 ;
      RECT 224.715 247.105 346.52 251.735 ;
      RECT 224.715 244.355 236.945 247.105 ;
      RECT 224.715 242.435 225.565 244.355 ;
      RECT 217.055 241.585 225.565 242.435 ;
      RECT 342.15 220.085 346.52 247.105 ;
      RECT 249.105 220.085 249.955 247.105 ;
      RECT 217.055 220.065 217.905 241.585 ;
      RECT 249.105 220.065 346.52 220.085 ;
      RECT 217.055 219.215 346.52 220.065 ;
      RECT 217.055 218.74 231.675 219.215 ;
      RECT 338.705 216.295 346.52 219.215 ;
      RECT 225.795 214.785 231.675 218.74 ;
      RECT 217.055 207.37 219.825 218.74 ;
      RECT 230.075 209.275 231.675 214.785 ;
      RECT 338.705 199.885 343.725 216.295 ;
      RECT 308.965 197.275 309.815 219.215 ;
      RECT 230.825 197.275 231.675 209.275 ;
      RECT 217.055 197.275 217.905 207.37 ;
      RECT 338.705 197.275 344.705 199.885 ;
      RECT 217.055 196.425 344.705 197.275 ;
      RECT 343.565 182.95 344.705 196.425 ;
      RECT 229.205 178.905 230.055 196.425 ;
      RECT 294.365 178.905 344.705 182.95 ;
      RECT 229.205 178.21 344.705 178.905 ;
      RECT 229.205 176.905 298.85 178.21 ;
      RECT 347.665 180.74 347.835 183.45 ;
      RECT 347.665 177.27 347.835 179.98 ;
      RECT 349.225 180.74 349.395 183.45 ;
      RECT 348.445 180.15 351.735 180.57 ;
      RECT 350.005 180.57 350.175 183.45 ;
      RECT 348.445 180.57 348.615 183.45 ;
      RECT 351.565 180.57 351.735 183.45 ;
      RECT 348.445 177.27 348.615 180.15 ;
      RECT 350.005 177.27 350.175 180.15 ;
      RECT 351.565 177.27 351.735 180.15 ;
      RECT 349.225 177.27 349.395 179.98 ;
      RECT 347.89 176.6 354.4 176.77 ;
      RECT 347.89 176.77 352.93 176.8 ;
      RECT 354.455 177.27 354.625 179.98 ;
      RECT 352.895 177.27 353.065 179.98 ;
      RECT 354.455 180.74 354.625 183.45 ;
      RECT 352.895 180.74 353.065 183.45 ;
      RECT 352.345 180.74 352.515 183.45 ;
      RECT 352.345 177.27 352.515 179.98 ;
      RECT 350.785 180.74 350.955 183.45 ;
      RECT 353.675 177.27 353.845 183.45 ;
      RECT 350.785 177.27 350.955 179.98 ;
      RECT 356.965 177.155 357.135 182.9 ;
      RECT 358.725 177.155 358.895 182.9 ;
      RECT 356.355 176.655 356.865 176.985 ;
      RECT 356.355 183.065 356.865 183.395 ;
      RECT 356.425 176.985 356.795 183.065 ;
      RECT 357.235 183.065 358.625 183.395 ;
      RECT 357.235 176.655 358.625 176.985 ;
      RECT 357.305 176.985 357.675 183.065 ;
      RECT 358.185 176.985 358.555 183.065 ;
      RECT 358.995 176.655 359.505 176.985 ;
      RECT 358.995 183.065 359.505 183.395 ;
      RECT 359.065 176.985 359.435 183.065 ;
      RECT 360.155 177.155 360.325 182.9 ;
      RECT 361.375 176.985 361.745 183.065 ;
      RECT 361.305 183.065 361.815 183.395 ;
      RECT 361.285 176.69 361.815 176.86 ;
      RECT 361.305 176.86 361.815 176.985 ;
      RECT 361.305 176.655 361.815 176.69 ;
      RECT 360.495 176.985 360.865 183.065 ;
      RECT 360.425 176.655 360.935 176.985 ;
      RECT 360.425 183.065 360.935 183.395 ;
      RECT 356.085 177.155 356.255 178.205 ;
      RECT 356.085 178.435 356.255 178.765 ;
      RECT 357.845 178.435 358.015 178.765 ;
      RECT 357.845 177.155 358.015 178.205 ;
      RECT 361.035 177.155 361.205 178.205 ;
      RECT 359.605 177.155 359.775 178.205 ;
      RECT 361.035 178.435 361.205 178.765 ;
      RECT 359.605 178.435 359.775 178.765 ;
      RECT 356.085 179.885 356.255 182.595 ;
      RECT 356.085 179.385 356.255 179.715 ;
      RECT 357.845 179.885 358.015 182.595 ;
      RECT 357.845 179.385 358.015 179.715 ;
      RECT 361.035 179.885 361.205 182.595 ;
      RECT 359.605 179.885 359.775 182.595 ;
      RECT 361.035 179.385 361.205 179.715 ;
      RECT 359.605 179.385 359.775 179.715 ;
      RECT 361.915 179.85 362.085 182.9 ;
      RECT 361.915 177.155 362.085 179.32 ;
      RECT 361.915 179.32 362.34 179.85 ;
      RECT 362.735 179.035 363.9 179.205 ;
      RECT 362.85 176.985 363.12 179.035 ;
      RECT 362.17 176.655 363.12 176.985 ;
      RECT 363.29 177.785 365.1 177.955 ;
      RECT 363.29 177.955 363.46 178.455 ;
      RECT 364.93 177.955 365.1 178.455 ;
      RECT 362.51 177.155 362.68 178.595 ;
      RECT 365.765 179.3 366.005 180.975 ;
      RECT 365.765 178.795 365.935 179.3 ;
      RECT 365.435 178.625 365.935 178.795 ;
      RECT 365.435 177.955 365.62 178.625 ;
      RECT 365.435 177.785 366.615 177.955 ;
      RECT 366.445 177.675 366.615 177.785 ;
      RECT 366.445 177.955 366.615 178.685 ;
      RECT 364.07 178.965 365.595 179.455 ;
      RECT 364.07 178.125 364.24 178.965 ;
      RECT 364.07 179.455 364.24 180.975 ;
      RECT 366.105 178.455 366.275 178.855 ;
      RECT 366.105 178.855 366.415 179.13 ;
      RECT 366.175 179.13 366.415 179.965 ;
      RECT 365.79 178.125 366.275 178.455 ;
      RECT 366.175 179.965 366.525 180.975 ;
      RECT 367.015 179.395 367.525 179.725 ;
      RECT 367.265 178.685 367.525 179.395 ;
      RECT 367.225 177.675 367.525 178.685 ;
      RECT 366.65 179.185 366.845 179.795 ;
      RECT 366.585 178.855 367.095 179.185 ;
      RECT 366.65 179.795 366.86 179.815 ;
      RECT 366.65 179.815 366.87 179.835 ;
      RECT 366.65 179.835 366.885 179.845 ;
      RECT 366.665 179.845 366.89 179.865 ;
      RECT 366.675 179.865 366.89 179.885 ;
      RECT 366.695 179.885 366.89 179.895 ;
      RECT 366.695 179.895 367.885 180.36 ;
      RECT 155.895 188.86 158.85 192.62 ;
      RECT 106.33 188.775 121.065 189.945 ;
      RECT 140.25 188.01 158.85 188.86 ;
      RECT 47.2 187.62 48.05 189.19 ;
      RECT 80.13 187.62 101.37 189.19 ;
      RECT 47.2 187.45 101.37 187.62 ;
      RECT 106.335 186.22 121.065 188.775 ;
      RECT 80.13 186.22 101.37 187.45 ;
      RECT 80.13 185.67 121.065 186.22 ;
      RECT 47.2 185.67 48.05 187.45 ;
      RECT 155.895 184.375 158.85 188.01 ;
      RECT 47.2 183.71 121.065 185.67 ;
      RECT 140.25 183.525 158.85 184.375 ;
      RECT 96.485 180.515 121.065 183.71 ;
      RECT 96.485 180.175 122.34 180.515 ;
      RECT 96.485 179.155 158.85 180.175 ;
      RECT 155.895 180.175 158.85 183.525 ;
      RECT 122.91 181.545 137.86 181.715 ;
      RECT 138.08 182.155 138.59 182.185 ;
      RECT 133.88 181.885 138.59 182.155 ;
      RECT 138.08 181.855 138.59 181.885 ;
      RECT 124.41 181.885 133.71 182.325 ;
      RECT 122.91 182.325 137.86 182.495 ;
      RECT 124.41 180.935 133.71 181.375 ;
      RECT 122.91 180.765 137.86 180.935 ;
      RECT 139.46 181.885 144.17 182.155 ;
      RECT 139.46 182.155 139.97 182.185 ;
      RECT 139.46 181.855 139.97 181.885 ;
      RECT 139.46 181.105 142.02 181.375 ;
      RECT 139.46 181.375 139.97 181.405 ;
      RECT 139.46 181.075 139.97 181.105 ;
      RECT 136.03 181.105 138.59 181.375 ;
      RECT 138.08 181.375 138.59 181.405 ;
      RECT 138.08 181.075 138.59 181.105 ;
      RECT 138.76 181.56 139.29 182.73 ;
      RECT 121.235 182.73 139.29 185.07 ;
      RECT 121.235 185.07 122.525 187.295 ;
      RECT 138.76 185.07 139.29 187.295 ;
      RECT 121.235 187.295 139.29 189.635 ;
      RECT 121.235 189.635 121.92 190.805 ;
      RECT 138.76 189.635 139.29 190.805 ;
      RECT 139.12 181.235 139.29 181.56 ;
      RECT 138.76 181.235 138.93 181.56 ;
      RECT 144.34 181.885 153.64 182.325 ;
      RECT 140.19 182.325 155.14 182.495 ;
      RECT 144.34 180.935 153.64 181.375 ;
      RECT 140.19 180.765 155.14 180.935 ;
      RECT 140.19 181.545 155.14 181.715 ;
      RECT 168.555 175.785 169.225 175.955 ;
      RECT 168.555 176.325 169.225 176.495 ;
      RECT 168.555 177.995 169.225 178.165 ;
      RECT 168.555 178.535 169.225 178.705 ;
      RECT 168.555 180.205 169.225 180.375 ;
      RECT 168.555 180.745 169.225 180.915 ;
      RECT 168.555 182.415 169.225 188.785 ;
      RECT 172.405 181.435 174.095 184.885 ;
      RECT 215.91 181.435 217.6 184.885 ;
      RECT 220.78 175.785 221.45 175.955 ;
      RECT 220.78 176.325 221.45 176.495 ;
      RECT 220.78 177.995 221.45 178.165 ;
      RECT 220.78 178.535 221.45 178.705 ;
      RECT 220.78 180.205 221.45 180.375 ;
      RECT 220.78 180.745 221.45 180.915 ;
      RECT 220.78 182.415 221.45 188.785 ;
      RECT 234.865 181.545 249.815 181.715 ;
      RECT 250.035 182.155 250.545 182.185 ;
      RECT 245.835 181.885 250.545 182.155 ;
      RECT 250.035 181.855 250.545 181.885 ;
      RECT 236.365 181.885 245.665 182.325 ;
      RECT 234.865 182.325 249.815 182.495 ;
      RECT 236.365 180.935 245.665 181.375 ;
      RECT 234.865 180.765 249.815 180.935 ;
      RECT 247.985 181.105 250.545 181.375 ;
      RECT 250.035 181.375 250.545 181.405 ;
      RECT 250.035 181.075 250.545 181.105 ;
      RECT 251.415 181.885 256.125 182.155 ;
      RECT 251.415 182.155 251.925 182.185 ;
      RECT 251.415 181.855 251.925 181.885 ;
      RECT 251.415 181.105 253.975 181.375 ;
      RECT 251.415 181.375 251.925 181.405 ;
      RECT 251.415 181.075 251.925 181.105 ;
      RECT 250.715 181.56 251.245 182.73 ;
      RECT 250.715 182.73 268.77 185.07 ;
      RECT 250.715 185.07 251.245 187.295 ;
      RECT 267.48 185.07 268.77 187.295 ;
      RECT 250.715 187.295 268.77 189.635 ;
      RECT 250.715 189.635 251.245 190.805 ;
      RECT 268.085 189.635 268.77 190.805 ;
      RECT 250.715 181.235 250.885 181.56 ;
      RECT 251.075 181.235 251.245 181.56 ;
      RECT 256.295 180.935 265.595 181.375 ;
      RECT 252.145 180.765 267.095 180.935 ;
      RECT 252.145 181.545 267.095 181.715 ;
      RECT 256.295 181.885 265.595 182.325 ;
      RECT 252.145 182.325 267.095 182.495 ;
      RECT 275.845 195.44 342.805 195.445 ;
      RECT 231.155 194.595 342.805 195.44 ;
      RECT 288.635 194.5 342.805 194.595 ;
      RECT 305.32 193.91 308.105 194.08 ;
      RECT 305.32 194.08 308.03 194.5 ;
      RECT 231.155 193.515 283.67 194.595 ;
      RECT 309.875 192.985 310.045 194.5 ;
      RECT 322.385 192.985 342.805 194.5 ;
      RECT 231.155 192.95 234.11 193.515 ;
      RECT 309.875 192.815 342.805 192.985 ;
      RECT 231.155 192.62 235.245 192.95 ;
      RECT 288.635 191.955 303.89 194.5 ;
      RECT 246.5 191.905 283.67 193.515 ;
      RECT 341.955 191.1 342.805 192.815 ;
      RECT 288.635 191.1 309.875 191.955 ;
      RECT 288.635 190.93 342.805 191.1 ;
      RECT 268.94 189.945 283.67 191.905 ;
      RECT 288.635 189.36 309.875 190.93 ;
      RECT 341.955 189.36 342.805 190.93 ;
      RECT 288.635 189.19 342.805 189.36 ;
      RECT 231.155 188.86 234.11 192.62 ;
      RECT 268.94 188.775 283.675 189.945 ;
      RECT 231.155 188.01 249.755 188.86 ;
      RECT 341.955 187.62 342.805 189.19 ;
      RECT 288.635 187.62 309.875 189.19 ;
      RECT 288.635 187.45 342.805 187.62 ;
      RECT 288.635 186.22 309.875 187.45 ;
      RECT 268.94 186.22 283.67 188.775 ;
      RECT 268.94 185.67 309.875 186.22 ;
      RECT 341.955 185.67 342.805 187.45 ;
      RECT 231.155 184.375 234.11 188.01 ;
      RECT 268.94 183.71 342.805 185.67 ;
      RECT 23 182.465 23.425 182.795 ;
      RECT 23.255 182.795 23.425 183.275 ;
      RECT 23.14 183.275 23.425 183.945 ;
      RECT 23.255 183.945 23.425 184.645 ;
      RECT 23.255 184.645 23.61 185.655 ;
      RECT 31.11 177.155 31.28 182.9 ;
      RECT 31.38 176.655 32.77 176.985 ;
      RECT 31.38 183.065 32.77 183.395 ;
      RECT 31.45 176.985 31.82 183.065 ;
      RECT 32.33 176.985 32.7 183.065 ;
      RECT 30.5 176.655 31.01 176.985 ;
      RECT 30.5 183.065 31.01 183.395 ;
      RECT 30.57 176.985 30.94 183.065 ;
      RECT 27.92 179.85 28.09 182.9 ;
      RECT 27.92 177.155 28.09 179.32 ;
      RECT 27.665 179.32 28.09 179.85 ;
      RECT 29.68 177.155 29.85 182.9 ;
      RECT 28.26 176.985 28.63 183.065 ;
      RECT 28.19 183.065 28.7 183.395 ;
      RECT 28.19 176.69 28.72 176.86 ;
      RECT 28.19 176.86 28.7 176.985 ;
      RECT 28.19 176.655 28.7 176.69 ;
      RECT 29.14 176.985 29.51 183.065 ;
      RECT 29.07 176.655 29.58 176.985 ;
      RECT 29.07 183.065 29.58 183.395 ;
      RECT 26.105 179.035 27.27 179.205 ;
      RECT 26.885 176.985 27.155 179.035 ;
      RECT 26.885 176.655 27.835 176.985 ;
      RECT 28.8 177.155 28.97 178.205 ;
      RECT 27.325 177.155 27.495 178.595 ;
      RECT 28.8 178.435 28.97 178.765 ;
      RECT 30.23 177.155 30.4 178.205 ;
      RECT 30.23 178.435 30.4 178.765 ;
      RECT 26.28 182.795 26.45 183.275 ;
      RECT 26.28 183.945 26.45 184.675 ;
      RECT 26.09 182.465 26.45 182.795 ;
      RECT 25.92 183.275 26.45 183.945 ;
      RECT 26.28 184.675 26.66 185.685 ;
      RECT 26.12 181.885 27.54 182.265 ;
      RECT 26.705 182.265 27.54 182.795 ;
      RECT 27.295 179.575 27.465 179.625 ;
      RECT 27.295 179.625 27.495 180.825 ;
      RECT 27.325 180.825 27.495 180.975 ;
      RECT 28.8 179.885 28.97 182.595 ;
      RECT 28.8 179.385 28.97 179.715 ;
      RECT 30.23 179.885 30.4 182.595 ;
      RECT 30.23 179.385 30.4 179.715 ;
      RECT 35.605 176.6 42.115 176.77 ;
      RECT 37.075 176.77 42.115 176.8 ;
      RECT 33.14 176.655 33.65 176.985 ;
      RECT 33.14 183.065 33.65 183.395 ;
      RECT 33.21 176.985 33.58 183.065 ;
      RECT 33.75 177.155 33.92 178.205 ;
      RECT 33.75 179.885 33.92 182.595 ;
      RECT 32.87 177.155 33.04 182.9 ;
      RECT 31.99 179.885 32.16 182.595 ;
      RECT 31.99 179.385 32.16 179.715 ;
      RECT 33.75 179.385 33.92 179.715 ;
      RECT 31.99 178.435 32.16 178.765 ;
      RECT 33.75 178.435 33.92 178.765 ;
      RECT 31.99 177.155 32.16 178.205 ;
      RECT 35.38 177.27 35.55 179.98 ;
      RECT 35.38 180.74 35.55 183.45 ;
      RECT 36.16 177.27 36.33 183.45 ;
      RECT 36.94 177.27 37.11 179.98 ;
      RECT 36.94 180.74 37.11 183.45 ;
      RECT 37.49 180.74 37.66 183.45 ;
      RECT 42.17 180.74 42.34 183.45 ;
      RECT 37.49 177.27 37.66 179.98 ;
      RECT 42.17 177.27 42.34 179.98 ;
      RECT 39.05 180.74 39.22 183.45 ;
      RECT 40.61 180.74 40.78 183.45 ;
      RECT 38.27 180.15 41.56 180.57 ;
      RECT 38.27 180.57 38.44 183.45 ;
      RECT 39.83 180.57 40 183.45 ;
      RECT 41.39 180.57 41.56 183.45 ;
      RECT 38.27 177.27 38.44 180.15 ;
      RECT 39.83 177.27 40 180.15 ;
      RECT 41.39 177.27 41.56 180.15 ;
      RECT 39.05 177.27 39.22 179.98 ;
      RECT 40.61 177.27 40.78 179.98 ;
      RECT 43.485 251.735 164.155 251.76 ;
      RECT 43.485 247.105 165.29 251.735 ;
      RECT 153.06 244.355 165.29 247.105 ;
      RECT 164.44 242.435 165.29 244.355 ;
      RECT 164.44 241.585 172.95 242.435 ;
      RECT 43.485 220.085 47.855 247.105 ;
      RECT 140.05 220.085 140.9 247.105 ;
      RECT 172.1 220.065 172.95 241.585 ;
      RECT 43.485 220.065 140.9 220.085 ;
      RECT 43.485 219.215 172.95 220.065 ;
      RECT 158.33 218.74 172.95 219.215 ;
      RECT 43.485 216.295 51.3 219.215 ;
      RECT 158.33 214.785 164.21 218.74 ;
      RECT 170.18 207.37 172.95 218.74 ;
      RECT 158.33 209.275 159.93 214.785 ;
      RECT 46.28 199.885 51.3 216.295 ;
      RECT 158.33 197.275 159.18 209.275 ;
      RECT 80.19 197.275 81.04 219.215 ;
      RECT 172.1 197.275 172.95 207.37 ;
      RECT 45.3 197.275 51.3 199.885 ;
      RECT 45.3 196.425 172.95 197.275 ;
      RECT 45.3 182.95 46.44 196.425 ;
      RECT 159.95 178.905 160.8 196.425 ;
      RECT 45.3 178.905 95.64 182.95 ;
      RECT 45.3 178.21 160.8 178.905 ;
      RECT 91.155 176.905 160.8 178.21 ;
      RECT 47.2 195.44 114.16 195.445 ;
      RECT 47.2 194.595 158.85 195.44 ;
      RECT 47.2 194.5 101.37 194.595 ;
      RECT 81.9 193.91 84.685 194.08 ;
      RECT 81.975 194.08 84.685 194.5 ;
      RECT 106.335 193.515 158.85 194.595 ;
      RECT 47.2 192.985 67.62 194.5 ;
      RECT 79.96 192.985 80.13 194.5 ;
      RECT 155.895 192.95 158.85 193.515 ;
      RECT 154.76 192.62 158.85 192.95 ;
      RECT 47.2 192.815 80.13 192.985 ;
      RECT 106.335 191.905 143.505 193.515 ;
      RECT 86.115 191.955 101.37 194.5 ;
      RECT 47.2 191.1 48.05 192.815 ;
      RECT 80.13 191.1 101.37 191.955 ;
      RECT 47.2 190.93 101.37 191.1 ;
      RECT 106.335 189.945 121.065 191.905 ;
      RECT 47.2 189.36 48.05 190.93 ;
      RECT 80.13 189.36 101.37 190.93 ;
      RECT 47.2 189.19 101.37 189.36 ;
      RECT 364.53 169.58 366.14 169.75 ;
      RECT 367.26 169.58 369.97 169.75 ;
      RECT 366.56 169.58 367.09 169.75 ;
      RECT 364.03 169.34 364.36 169.41 ;
      RECT 364.03 168.9 364.36 168.97 ;
      RECT 364.03 168.97 370.77 169.34 ;
      RECT 370.44 169.34 370.77 169.41 ;
      RECT 370.44 168.9 370.77 168.97 ;
      RECT 364.655 170.46 370.275 170.63 ;
      RECT 361.955 170.46 363.02 170.63 ;
      RECT 364.03 171.17 364.36 171.24 ;
      RECT 364.03 170.73 364.36 170.8 ;
      RECT 364.03 170.8 370.77 171.17 ;
      RECT 370.44 170.73 370.77 170.8 ;
      RECT 370.44 171.17 370.77 171.26 ;
      RECT 364.655 172.77 370.275 172.94 ;
      RECT 364.03 172.6 364.36 172.67 ;
      RECT 364.03 172.16 364.36 172.23 ;
      RECT 364.03 172.23 370.77 172.6 ;
      RECT 370.44 172.16 370.77 172.23 ;
      RECT 370.44 172.6 370.77 172.69 ;
      RECT 364.53 173.65 366.14 173.82 ;
      RECT 367.26 173.65 369.97 173.82 ;
      RECT 366.56 173.65 367.09 173.82 ;
      RECT 370.955 173.02 371.125 173.04 ;
      RECT 363.765 173.48 364.36 173.555 ;
      RECT 363.765 173.025 364.36 173.11 ;
      RECT 370.44 173.48 371.125 173.55 ;
      RECT 363.765 173.11 371.125 173.48 ;
      RECT 370.44 173.04 371.125 173.11 ;
      RECT 361.97 173.65 363.02 173.82 ;
      RECT 387.7 168.645 388.03 169.295 ;
      RECT 388.96 168.645 389.29 169.295 ;
      RECT 388.33 168.645 388.66 169.295 ;
      RECT 389.59 168.645 389.92 169.295 ;
      RECT 390.22 168.645 390.55 169.295 ;
      RECT 387.7 167.615 388.03 168.265 ;
      RECT 390.22 167.615 390.55 168.265 ;
      RECT 389.59 167.615 389.92 168.265 ;
      RECT 388.33 167.615 388.66 168.265 ;
      RECT 388.96 167.615 389.29 168.265 ;
      RECT 396.2 168.535 399.77 168.865 ;
      RECT 396.2 174.495 399.77 174.825 ;
      RECT 395.76 169.315 395.93 174.165 ;
      RECT 390.85 168.645 391.18 169.295 ;
      RECT 390.85 167.615 391.18 168.265 ;
      RECT 400.48 168.535 404.05 168.865 ;
      RECT 400.48 174.495 404.05 174.825 ;
      RECT 400.04 169.315 400.21 174.165 ;
      RECT 404.32 169.315 404.49 174.165 ;
      RECT 413.66 168.535 417.23 168.865 ;
      RECT 409.38 168.535 412.95 168.865 ;
      RECT 413.66 174.495 417.23 174.825 ;
      RECT 409.38 174.495 412.95 174.825 ;
      RECT 413.22 169.315 413.39 174.165 ;
      RECT 408.94 169.315 409.11 174.165 ;
      RECT 417.5 169.315 417.67 174.165 ;
      RECT 450.32 171.825 456.455 172.355 ;
      RECT 450.32 167.395 456.455 167.925 ;
      RECT 450.32 171.115 454.735 171.645 ;
      RECT 450.32 170.21 455.595 170.74 ;
      RECT 450.32 174.64 454.305 175.17 ;
      RECT 448.865 171.71 449.875 171.88 ;
      RECT 448.865 170.83 449.875 171 ;
      RECT 448.865 169.03 458.585 169.295 ;
      RECT 448.865 169.95 449.875 170.12 ;
      RECT 448.865 172.535 458.585 172.8 ;
      RECT 448.865 173.46 458.585 173.725 ;
      RECT 448.865 174.38 449.875 174.55 ;
      RECT 448.865 167.28 449.875 167.45 ;
      RECT 448.865 168.105 458.585 168.37 ;
      RECT 457.565 169.895 459.345 170.175 ;
      RECT 459.095 168.88 459.345 169.895 ;
      RECT 459.095 171.935 459.345 172.95 ;
      RECT 457.565 171.655 459.345 171.935 ;
      RECT 459.095 170.175 459.345 171.655 ;
      RECT 456.695 170.775 458.575 171.055 ;
      RECT 457.565 174.325 459.345 174.605 ;
      RECT 459.095 173.31 459.345 174.325 ;
      RECT 459.095 176.365 459.345 177.38 ;
      RECT 457.565 176.085 459.345 176.365 ;
      RECT 459.095 174.605 459.345 176.085 ;
      RECT 456.675 169.51 457.345 169.68 ;
      RECT 456.675 173.94 457.345 174.11 ;
      RECT 22.48 178.685 22.74 179.395 ;
      RECT 22.48 179.395 22.99 179.725 ;
      RECT 22.48 177.675 22.78 178.685 ;
      RECT 23.73 178.455 23.9 178.855 ;
      RECT 23.59 178.855 23.9 179.13 ;
      RECT 23.59 179.13 23.83 179.965 ;
      RECT 23.73 178.125 24.215 178.455 ;
      RECT 23.48 179.965 23.83 180.975 ;
      RECT 24.905 177.785 26.715 177.955 ;
      RECT 24.905 177.955 25.075 178.455 ;
      RECT 26.545 177.955 26.715 178.455 ;
      RECT 24.385 177.955 24.57 178.625 ;
      RECT 24.07 178.625 24.57 178.795 ;
      RECT 24.07 178.795 24.24 179.3 ;
      RECT 24 179.3 24.24 180.975 ;
      RECT 23.39 177.785 24.57 177.955 ;
      RECT 23.39 177.675 23.56 177.785 ;
      RECT 23.39 177.955 23.56 178.685 ;
      RECT 23.115 179.885 23.31 179.895 ;
      RECT 23.115 179.865 23.33 179.885 ;
      RECT 23.115 179.845 23.34 179.865 ;
      RECT 23.12 179.835 23.355 179.845 ;
      RECT 23.135 179.815 23.355 179.835 ;
      RECT 23.145 179.795 23.355 179.815 ;
      RECT 23.16 179.185 23.355 179.795 ;
      RECT 22.91 178.855 23.42 179.185 ;
      RECT 22.12 179.455 22.29 179.895 ;
      RECT 22.12 179.895 23.31 180.36 ;
      RECT 22.12 180.36 22.87 180.975 ;
      RECT 25.54 184.585 26.11 184.915 ;
      RECT 25.54 181.885 25.71 183.385 ;
      RECT 23.665 183.385 25.71 183.555 ;
      RECT 25.09 183.555 25.71 183.725 ;
      RECT 25.54 183.725 25.71 184.585 ;
      RECT 25.94 184.915 26.11 184.975 ;
      RECT 23.07 181.885 24.83 182.265 ;
      RECT 23.78 182.265 24.83 182.895 ;
      RECT 24.41 178.965 25.935 179.455 ;
      RECT 25.765 178.125 25.935 178.965 ;
      RECT 25.765 179.455 25.935 180.975 ;
      RECT 24.985 181.145 26.715 181.315 ;
      RECT 24.985 179.625 25.155 181.145 ;
      RECT 26.545 179.625 26.715 181.145 ;
      RECT 352.245 170.74 352.415 171.115 ;
      RECT 348.6 171.555 349.005 171.885 ;
      RECT 348.6 172.935 349.005 173.265 ;
      RECT 348.6 171.885 348.77 172.935 ;
      RECT 348.305 167.295 351.015 167.465 ;
      RECT 347.425 168.075 351.015 168.245 ;
      RECT 348.305 168.855 351.015 169.025 ;
      RECT 348.305 169.635 351.325 169.97 ;
      RECT 347.395 169.175 347.565 169.355 ;
      RECT 347.395 168.825 347.565 169.005 ;
      RECT 344.475 169.005 347.565 169.175 ;
      RECT 348.305 170.31 351.015 170.355 ;
      RECT 348.305 170.14 355.775 170.31 ;
      RECT 348.305 171.065 351.015 171.235 ;
      RECT 349.505 171.235 349.675 171.655 ;
      RECT 347.395 170.735 347.565 170.915 ;
      RECT 347.395 170.385 347.565 170.565 ;
      RECT 344.475 170.565 347.565 170.735 ;
      RECT 348.94 172.575 351.3 172.745 ;
      RECT 348.94 172.415 349.61 172.575 ;
      RECT 347.395 172.295 347.565 172.475 ;
      RECT 347.395 171.945 347.565 172.125 ;
      RECT 344.475 172.125 347.565 172.295 ;
      RECT 348.305 173.585 351.015 173.755 ;
      RECT 349.99 173.165 350.16 173.585 ;
      RECT 347.395 173.505 347.565 173.685 ;
      RECT 347.395 174.465 351.015 174.635 ;
      RECT 344.475 173.685 347.565 173.855 ;
      RECT 347.395 173.855 347.565 174.465 ;
      RECT 352.535 168.02 352.865 168.575 ;
      RECT 353.065 167.8 356.025 167.97 ;
      RECT 352.725 167.56 352.895 167.665 ;
      RECT 352.725 167.39 356.97 167.56 ;
      RECT 350.74 167.665 352.895 167.835 ;
      RECT 356.64 167.56 356.97 168.225 ;
      RECT 351.485 168.515 352.155 168.685 ;
      RECT 351.965 168.155 352.135 168.515 ;
      RECT 352.245 169.33 352.415 169.595 ;
      RECT 351.485 169.16 352.415 169.33 ;
      RECT 352.245 168.93 352.415 169.16 ;
      RECT 353.065 169.36 356.025 169.53 ;
      RECT 351.565 169.635 351.945 169.97 ;
      RECT 357.11 169.19 357.44 169.2 ;
      RECT 354.28 168.92 357.44 169.19 ;
      RECT 357.11 168.69 357.44 168.92 ;
      RECT 353.065 168.58 355.775 168.75 ;
      RECT 350.65 171.555 351.815 171.885 ;
      RECT 351.485 171.455 351.815 171.555 ;
      RECT 351.485 170.915 351.815 171.285 ;
      RECT 351.485 171.285 354.59 171.455 ;
      RECT 350.39 172.075 351.06 172.405 ;
      RECT 353.065 171.7 355.775 171.87 ;
      RECT 353.065 170.92 356.025 171.09 ;
      RECT 353.335 173.63 356.045 173.8 ;
      RECT 350.38 173.06 351.815 173.265 ;
      RECT 350.38 172.935 354.87 173.06 ;
      RECT 351.485 172.89 354.87 172.935 ;
      RECT 351.485 173.265 351.815 173.85 ;
      RECT 353.065 172.48 356.025 172.65 ;
      RECT 352.245 173.46 352.415 173.79 ;
      RECT 363.19 173.48 363.52 173.55 ;
      RECT 363.19 173.04 363.52 173.11 ;
      RECT 356.78 173.48 357.11 173.55 ;
      RECT 356.78 173.46 363.52 173.48 ;
      RECT 352.245 173.26 363.52 173.46 ;
      RECT 356.78 173.11 363.52 173.26 ;
      RECT 356.78 173.04 357.11 173.11 ;
      RECT 351.855 174.02 370.25 174.22 ;
      RECT 359.83 167.555 360.16 167.81 ;
      RECT 359.83 167.385 363.02 167.555 ;
      RECT 360.64 167.555 361.31 167.67 ;
      RECT 362.01 167.2 363.02 167.385 ;
      RECT 359.25 167.98 362.34 168.15 ;
      RECT 359.25 168.15 360.59 168.32 ;
      RECT 360.42 168.32 360.59 168.54 ;
      RECT 362.01 167.75 362.34 167.98 ;
      RECT 359.25 169.03 360.26 169.2 ;
      RECT 359.25 168.67 360.25 169.03 ;
      RECT 362.82 167.78 362.99 168.32 ;
      RECT 361.12 168.32 362.99 168.49 ;
      RECT 361.21 170.46 361.785 170.63 ;
      RECT 357.58 170.46 360.29 170.63 ;
      RECT 360.46 170.46 360.79 170.63 ;
      RECT 356.78 170.29 357.11 170.36 ;
      RECT 356.78 169.85 357.11 169.92 ;
      RECT 356.78 169.92 363.52 170.29 ;
      RECT 363.19 170.29 363.52 170.37 ;
      RECT 363.19 169.84 363.52 169.92 ;
      RECT 357.275 169.5 363.86 169.67 ;
      RECT 363.69 169.67 363.86 169.85 ;
      RECT 357.275 169.67 363.02 169.75 ;
      RECT 370.44 170.29 370.77 170.36 ;
      RECT 370.44 169.85 370.77 169.92 ;
      RECT 363.69 170.29 364.36 170.36 ;
      RECT 363.69 169.85 364.36 169.92 ;
      RECT 363.69 169.92 370.77 170.29 ;
      RECT 357.275 171.34 362.895 171.51 ;
      RECT 356.78 172.05 357.11 172.12 ;
      RECT 356.78 171.61 357.11 171.68 ;
      RECT 356.78 171.82 366.71 171.99 ;
      RECT 356.78 171.99 363.52 172.05 ;
      RECT 363.19 172.05 363.52 172.12 ;
      RECT 356.78 171.68 363.52 171.82 ;
      RECT 363.19 171.61 363.52 171.68 ;
      RECT 364.53 171.99 366.71 172.06 ;
      RECT 363.69 171.24 363.86 171.41 ;
      RECT 363.69 171.41 366.71 171.58 ;
      RECT 356.78 171.17 357.11 171.24 ;
      RECT 356.78 170.73 357.11 170.8 ;
      RECT 363.19 171.17 363.86 171.24 ;
      RECT 356.78 170.8 363.86 171.17 ;
      RECT 363.19 170.73 363.86 170.8 ;
      RECT 364.53 171.34 366.71 171.41 ;
      RECT 357.58 172.22 360.29 172.39 ;
      RECT 361.2 172.22 363.02 172.39 ;
      RECT 357.275 172.745 357.58 172.77 ;
      RECT 357.275 172.77 363.02 172.94 ;
      RECT 356.325 172.415 357.41 172.56 ;
      RECT 356.325 172.56 357.58 172.745 ;
      RECT 357.58 173.65 360.29 173.82 ;
      RECT 361.21 173.65 361.74 173.82 ;
      RECT 360.46 173.65 360.79 173.82 ;
      RECT 364.53 167.68 366.14 167.85 ;
      RECT 367.26 167.68 370.275 167.85 ;
      RECT 364.53 168.63 369 168.8 ;
      RECT 366.56 167.68 367.09 167.85 ;
      RECT 362 169.03 362.89 169.2 ;
      RECT 26.485 173.46 33.225 173.48 ;
      RECT 32.895 173.48 33.225 173.55 ;
      RECT 26.485 173.11 33.225 173.26 ;
      RECT 32.895 173.04 33.225 173.11 ;
      RECT 26.985 173.65 28.035 173.82 ;
      RECT 29.715 173.65 32.425 173.82 ;
      RECT 28.265 173.65 28.795 173.82 ;
      RECT 29.215 173.65 29.545 173.82 ;
      RECT 37.14 168.02 37.47 168.575 ;
      RECT 33.035 167.39 37.28 167.56 ;
      RECT 37.11 167.56 37.28 167.665 ;
      RECT 37.11 167.665 39.265 167.835 ;
      RECT 33.035 167.56 33.365 168.225 ;
      RECT 33.98 167.8 36.94 167.97 ;
      RECT 34.23 168.58 36.94 168.75 ;
      RECT 32.565 169.19 32.895 169.2 ;
      RECT 32.565 168.69 32.895 168.92 ;
      RECT 32.565 168.92 35.725 169.19 ;
      RECT 33.98 169.36 36.94 169.53 ;
      RECT 34.23 170.14 41.7 170.31 ;
      RECT 38.99 170.31 41.7 170.355 ;
      RECT 33.98 172.48 36.94 172.65 ;
      RECT 38.19 171.455 38.52 171.555 ;
      RECT 38.19 171.555 39.355 171.885 ;
      RECT 35.415 171.285 38.52 171.455 ;
      RECT 38.19 170.915 38.52 171.285 ;
      RECT 34.23 171.7 36.94 171.87 ;
      RECT 33.98 170.92 36.94 171.09 ;
      RECT 33.96 173.63 36.67 173.8 ;
      RECT 38.19 173.06 39.625 173.265 ;
      RECT 35.135 172.935 39.625 173.06 ;
      RECT 35.135 172.89 38.52 172.935 ;
      RECT 38.19 173.265 38.52 173.85 ;
      RECT 37.59 170.54 42.27 170.74 ;
      RECT 42.1 170.74 42.27 171.29 ;
      RECT 42.1 168.58 42.27 170.54 ;
      RECT 37.59 170.74 37.76 171.115 ;
      RECT 41 171.555 41.405 171.885 ;
      RECT 41 172.935 41.405 173.265 ;
      RECT 41.235 171.885 41.405 172.935 ;
      RECT 38.99 167.295 41.7 167.465 ;
      RECT 38.99 168.075 42.58 168.245 ;
      RECT 38.99 168.855 41.7 169.025 ;
      RECT 37.85 168.515 38.52 168.685 ;
      RECT 37.87 168.155 38.04 168.515 ;
      RECT 42.44 169.175 42.61 169.355 ;
      RECT 42.44 168.825 42.61 169.005 ;
      RECT 42.44 169.005 45.53 169.175 ;
      RECT 37.59 169.16 38.52 169.33 ;
      RECT 37.59 169.33 37.76 169.595 ;
      RECT 37.59 168.93 37.76 169.16 ;
      RECT 38.68 169.635 41.7 169.97 ;
      RECT 38.06 169.635 38.44 169.97 ;
      RECT 42.44 170.735 42.61 170.915 ;
      RECT 42.44 170.385 42.61 170.565 ;
      RECT 42.44 170.565 45.53 170.735 ;
      RECT 38.99 171.065 41.7 171.235 ;
      RECT 40.33 171.235 40.5 171.655 ;
      RECT 42.44 172.295 42.61 172.475 ;
      RECT 42.44 171.945 42.61 172.125 ;
      RECT 42.44 172.125 45.53 172.295 ;
      RECT 38.705 172.575 41.065 172.745 ;
      RECT 40.395 172.415 41.065 172.575 ;
      RECT 38.945 172.075 39.615 172.405 ;
      RECT 38.99 173.585 41.7 173.755 ;
      RECT 39.845 173.165 40.015 173.585 ;
      RECT 38.99 174.465 42.61 174.635 ;
      RECT 42.44 173.505 42.61 173.685 ;
      RECT 42.44 173.685 45.53 173.855 ;
      RECT 42.44 173.855 42.61 174.465 ;
      RECT 49.625 169.345 50.325 175.24 ;
      RECT 49.625 175.24 61.085 175.94 ;
      RECT 49.625 168.645 61.085 169.345 ;
      RECT 60.385 169.345 61.085 175.24 ;
      RECT 51.085 170.805 51.785 173.78 ;
      RECT 51.085 173.78 59.625 174.48 ;
      RECT 51.085 170.105 59.625 170.805 ;
      RECT 58.915 170.805 59.625 173.78 ;
      RECT 52.655 171.28 58.05 171.82 ;
      RECT 52.655 172.755 58.05 173.295 ;
      RECT 58.22 171.625 58.63 172.95 ;
      RECT 75.615 167.825 76.145 168.355 ;
      RECT 75.615 168.88 76.145 169.41 ;
      RECT 63.355 161.46 88.445 162.31 ;
      RECT 63.355 162.31 64.205 174.99 ;
      RECT 87.595 162.31 88.445 174.99 ;
      RECT 63.355 174.99 88.445 175.84 ;
      RECT 168.555 174.115 169.225 174.285 ;
      RECT 168.555 173.755 169.225 173.925 ;
      RECT 168.625 173.705 169.155 173.755 ;
      RECT 169.76 173.655 171.78 174.405 ;
      RECT 172.405 174.15 174.095 174.32 ;
      RECT 172.405 173.755 174.095 173.925 ;
      RECT 172.405 174.32 174.09 174.355 ;
      RECT 172.405 173.925 174.09 174.15 ;
      RECT 215.91 174.15 217.6 174.32 ;
      RECT 215.91 173.755 217.6 173.925 ;
      RECT 215.915 174.32 217.6 174.355 ;
      RECT 215.915 173.925 217.6 174.15 ;
      RECT 220.78 174.115 221.45 174.285 ;
      RECT 220.78 173.755 221.45 173.925 ;
      RECT 220.85 173.705 221.38 173.755 ;
      RECT 218.225 173.655 220.245 174.405 ;
      RECT 301.56 161.46 326.65 162.31 ;
      RECT 325.8 162.31 326.65 174.99 ;
      RECT 301.56 162.31 302.41 174.99 ;
      RECT 301.56 174.99 326.65 175.84 ;
      RECT 313.86 167.825 314.39 168.355 ;
      RECT 313.86 168.88 314.39 169.41 ;
      RECT 331.375 171.625 331.785 172.95 ;
      RECT 328.92 169.345 329.62 175.24 ;
      RECT 328.92 175.24 340.38 175.94 ;
      RECT 328.92 168.645 340.38 169.345 ;
      RECT 339.68 169.345 340.38 175.24 ;
      RECT 330.38 170.805 331.09 173.78 ;
      RECT 330.38 173.78 338.92 174.48 ;
      RECT 330.38 170.105 338.92 170.805 ;
      RECT 338.22 170.805 338.92 173.78 ;
      RECT 331.955 171.28 337.35 171.82 ;
      RECT 331.955 172.755 337.35 173.295 ;
      RECT 351.485 174.28 351.685 174.405 ;
      RECT 351.485 174.405 368.96 174.605 ;
      RECT 347.735 174.08 351.685 174.28 ;
      RECT 347.735 171.57 347.905 174.08 ;
      RECT 347.735 170.54 352.415 170.74 ;
      RECT 347.735 170.74 347.905 171.29 ;
      RECT 347.735 168.58 347.905 170.54 ;
      RECT 438.24 160.345 438.57 160.995 ;
      RECT 440.67 160.345 441 160.995 ;
      RECT 437.43 160.345 437.76 160.995 ;
      RECT 439.86 160.345 440.19 160.995 ;
      RECT 439.05 160.345 439.38 160.995 ;
      RECT 450.32 162.965 455.165 163.495 ;
      RECT 450.32 162.255 456.025 162.785 ;
      RECT 450.32 166.685 454.735 167.215 ;
      RECT 450.32 161.35 455.595 161.88 ;
      RECT 450.32 165.78 454.305 166.31 ;
      RECT 448.865 162.85 449.875 163.02 ;
      RECT 448.865 161.97 449.875 162.14 ;
      RECT 448.865 160.17 458.585 160.435 ;
      RECT 448.865 161.09 449.875 161.26 ;
      RECT 448.865 163.675 458.585 163.94 ;
      RECT 448.865 166.4 449.875 166.57 ;
      RECT 448.865 164.6 458.585 164.865 ;
      RECT 448.865 165.52 449.875 165.69 ;
      RECT 456.695 166.345 458.575 166.625 ;
      RECT 457.565 165.465 459.345 165.745 ;
      RECT 459.095 164.45 459.345 165.465 ;
      RECT 459.095 167.505 459.345 168.52 ;
      RECT 457.565 167.225 459.345 167.505 ;
      RECT 459.095 165.745 459.345 167.225 ;
      RECT 457.565 161.035 459.345 161.315 ;
      RECT 459.095 160.02 459.345 161.035 ;
      RECT 459.095 163.075 459.345 164.09 ;
      RECT 457.565 162.795 459.345 163.075 ;
      RECT 459.095 161.315 459.345 162.795 ;
      RECT 456.695 161.915 458.575 162.195 ;
      RECT 456.675 160.65 457.345 160.82 ;
      RECT 456.675 165.08 457.345 165.25 ;
      RECT 19.73 170.46 25.35 170.63 ;
      RECT 19.73 172.77 25.35 172.94 ;
      RECT 26.145 169.67 26.315 169.85 ;
      RECT 26.145 169.5 32.73 169.67 ;
      RECT 19.235 170.29 19.565 170.36 ;
      RECT 19.235 169.85 19.565 169.92 ;
      RECT 26.985 169.67 32.73 169.75 ;
      RECT 25.645 170.29 26.315 170.36 ;
      RECT 19.235 169.92 26.315 170.29 ;
      RECT 25.645 169.85 26.315 169.92 ;
      RECT 18.88 173.02 19.05 173.04 ;
      RECT 18.88 173.48 19.565 173.55 ;
      RECT 18.88 173.04 19.565 173.11 ;
      RECT 18.88 173.11 26.24 173.48 ;
      RECT 25.645 173.48 26.24 173.555 ;
      RECT 25.645 173.025 26.24 173.11 ;
      RECT 19.235 170.73 19.565 170.8 ;
      RECT 19.235 170.8 25.975 171.17 ;
      RECT 25.645 171.17 25.975 171.24 ;
      RECT 25.645 170.73 25.975 170.8 ;
      RECT 19.235 171.17 19.565 171.26 ;
      RECT 19.235 172.16 19.565 172.23 ;
      RECT 19.235 172.23 25.975 172.6 ;
      RECT 25.645 172.6 25.975 172.67 ;
      RECT 25.645 172.16 25.975 172.23 ;
      RECT 19.235 172.6 19.565 172.69 ;
      RECT 19.235 169.34 19.565 169.41 ;
      RECT 19.235 168.9 19.565 168.97 ;
      RECT 19.235 168.97 25.975 169.34 ;
      RECT 25.645 169.34 25.975 169.41 ;
      RECT 25.645 168.9 25.975 168.97 ;
      RECT 19.73 167.68 22.745 167.85 ;
      RECT 19.755 174.02 38.15 174.22 ;
      RECT 23.865 167.68 25.475 167.85 ;
      RECT 22.915 167.68 23.445 167.85 ;
      RECT 21.005 168.63 25.475 168.8 ;
      RECT 20.035 169.58 22.745 169.75 ;
      RECT 23.865 169.58 25.475 169.75 ;
      RECT 22.915 169.58 23.445 169.75 ;
      RECT 23.295 171.41 26.315 171.58 ;
      RECT 26.145 171.24 26.315 171.41 ;
      RECT 32.895 171.17 33.225 171.24 ;
      RECT 32.895 170.73 33.225 170.8 ;
      RECT 23.295 171.34 25.475 171.41 ;
      RECT 26.145 171.17 26.815 171.24 ;
      RECT 26.145 170.73 26.815 170.8 ;
      RECT 26.145 170.8 33.225 171.17 ;
      RECT 26.485 172.05 26.815 172.12 ;
      RECT 26.485 171.61 26.815 171.68 ;
      RECT 32.895 172.05 33.225 172.12 ;
      RECT 32.895 171.61 33.225 171.68 ;
      RECT 23.295 171.99 25.475 172.06 ;
      RECT 26.485 171.99 33.225 172.05 ;
      RECT 26.485 171.68 33.225 171.82 ;
      RECT 23.295 171.82 33.225 171.99 ;
      RECT 20.035 173.65 22.745 173.82 ;
      RECT 23.865 173.65 25.475 173.82 ;
      RECT 22.915 173.65 23.445 173.82 ;
      RECT 21.045 174.405 38.52 174.605 ;
      RECT 38.32 174.28 38.52 174.405 ;
      RECT 42.1 171.57 42.27 174.08 ;
      RECT 38.32 174.08 42.27 174.28 ;
      RECT 27.11 171.34 32.73 171.51 ;
      RECT 26.985 172.77 32.73 172.94 ;
      RECT 32.425 172.745 32.73 172.77 ;
      RECT 32.425 172.56 33.68 172.745 ;
      RECT 32.595 172.415 33.68 172.56 ;
      RECT 27.665 167.98 30.755 168.15 ;
      RECT 29.415 168.15 30.755 168.32 ;
      RECT 29.415 168.32 29.585 168.54 ;
      RECT 27.665 167.75 27.995 167.98 ;
      RECT 26.985 167.385 30.175 167.555 ;
      RECT 28.695 167.555 29.365 167.67 ;
      RECT 29.845 167.555 30.175 167.81 ;
      RECT 26.985 167.2 27.995 167.385 ;
      RECT 27.015 168.32 28.885 168.49 ;
      RECT 27.015 167.78 27.185 168.32 ;
      RECT 27.115 169.03 28.005 169.2 ;
      RECT 29.745 169.03 30.755 169.2 ;
      RECT 29.755 168.67 30.755 169.03 ;
      RECT 26.985 170.46 28.05 170.63 ;
      RECT 26.485 169.92 33.225 170.29 ;
      RECT 32.895 170.29 33.225 170.36 ;
      RECT 32.895 169.85 33.225 169.92 ;
      RECT 26.485 170.29 26.815 170.37 ;
      RECT 26.485 169.84 26.815 169.92 ;
      RECT 29.715 170.46 32.425 170.63 ;
      RECT 28.22 170.46 28.795 170.63 ;
      RECT 29.215 170.46 29.545 170.63 ;
      RECT 26.985 172.22 28.805 172.39 ;
      RECT 29.715 172.22 32.425 172.39 ;
      RECT 26.485 173.48 26.815 173.55 ;
      RECT 26.485 173.04 26.815 173.11 ;
      RECT 37.59 173.46 37.76 173.79 ;
      RECT 26.485 173.26 37.76 173.46 ;
      RECT 352.245 167.16 352.415 167.495 ;
      RECT 352.245 166.965 352.415 166.99 ;
      RECT 351.485 163.965 352.155 164.135 ;
      RECT 351.955 162.645 352.155 163.965 ;
      RECT 351.955 162.445 369.46 162.645 ;
      RECT 368.87 162.645 369.46 162.86 ;
      RECT 359.25 167.03 359.63 167.74 ;
      RECT 359.25 166.58 360.26 167.03 ;
      RECT 357.11 166.41 360.26 166.58 ;
      RECT 359.25 165.98 360.26 166.07 ;
      RECT 352.565 166.24 360.26 166.41 ;
      RECT 357.11 166.07 360.26 166.24 ;
      RECT 353.065 164.68 356.025 164.85 ;
      RECT 353.065 163.12 356.025 163.29 ;
      RECT 357.11 163.45 357.44 163.46 ;
      RECT 354.28 163.46 357.44 163.73 ;
      RECT 357.11 163.73 357.44 163.96 ;
      RECT 352.725 165.09 356.97 165.26 ;
      RECT 352.725 164.985 352.895 165.09 ;
      RECT 350.44 164.815 352.895 164.985 ;
      RECT 356.64 164.425 356.97 165.09 ;
      RECT 353.065 167.02 355.775 167.19 ;
      RECT 353.065 165.46 355.775 165.63 ;
      RECT 353.065 163.9 355.775 164.07 ;
      RECT 353.265 163.885 353.795 163.9 ;
      RECT 357.97 164.015 358.14 165.025 ;
      RECT 359.25 163.27 360.16 164.105 ;
      RECT 359.25 164.105 359.63 164.69 ;
      RECT 363.52 163.875 363.69 164.89 ;
      RECT 363.52 164.89 370.275 165.06 ;
      RECT 364.53 164.82 370.275 164.89 ;
      RECT 364.03 166.08 364.36 166.15 ;
      RECT 364.03 165.71 370.77 166.08 ;
      RECT 370.44 166.08 370.77 166.15 ;
      RECT 370.44 165.64 370.77 165.71 ;
      RECT 360.51 163.705 363.69 163.875 ;
      RECT 360.51 163.875 361.09 164.06 ;
      RECT 360.51 163.53 361.09 163.705 ;
      RECT 364.03 165.06 364.36 165.71 ;
      RECT 359.83 164.36 363.05 164.53 ;
      RECT 359.83 164.53 360.16 164.72 ;
      RECT 360.64 164.53 361.31 164.89 ;
      RECT 362.04 164.15 363.05 164.36 ;
      RECT 359.25 165.1 362.28 165.27 ;
      RECT 360.75 165.27 361.09 165.72 ;
      RECT 361.95 164.7 362.34 164.87 ;
      RECT 361.95 164.87 362.28 165.1 ;
      RECT 360.75 165.72 360.92 167.145 ;
      RECT 361.49 165.78 361.74 166.44 ;
      RECT 361.49 165.47 362.99 165.78 ;
      RECT 362.82 164.73 362.99 165.47 ;
      RECT 363.52 166.99 363.69 168.02 ;
      RECT 361.15 166.305 361.32 166.82 ;
      RECT 361.15 166.82 363.69 166.99 ;
      RECT 370.44 168.46 370.77 168.53 ;
      RECT 363.52 168.02 364.36 168.09 ;
      RECT 364.03 168.46 364.36 168.53 ;
      RECT 370.44 168.02 370.77 168.09 ;
      RECT 363.52 168.09 370.77 168.19 ;
      RECT 364.03 168.19 370.77 168.46 ;
      RECT 364.53 167.13 370.275 167.3 ;
      RECT 364.53 165.37 370.275 165.54 ;
      RECT 364.53 163.06 370.275 163.23 ;
      RECT 364.53 163.84 365.58 163.94 ;
      RECT 364.03 163.77 365.58 163.84 ;
      RECT 370.44 163.77 370.77 163.84 ;
      RECT 370.44 163.33 370.77 163.4 ;
      RECT 364.53 163.94 366.14 164.11 ;
      RECT 364.03 163.4 370.77 163.77 ;
      RECT 364.03 163.33 364.36 163.4 ;
      RECT 362 163.27 363.05 163.44 ;
      RECT 367.26 163.94 369.97 164.11 ;
      RECT 366.76 163.94 367.09 164.11 ;
      RECT 364.19 164.19 364.36 164.21 ;
      RECT 364.03 164.65 364.36 164.72 ;
      RECT 364.03 164.21 364.36 164.28 ;
      RECT 364.03 164.28 370.77 164.65 ;
      RECT 370.44 164.65 370.77 164.72 ;
      RECT 370.44 164.21 370.77 164.28 ;
      RECT 362 166.15 363.02 166.32 ;
      RECT 362.01 166.32 363.02 166.51 ;
      RECT 362.01 165.98 363.02 166.15 ;
      RECT 364.03 166.96 364.36 167.03 ;
      RECT 364.03 166.52 364.36 166.59 ;
      RECT 364.03 166.59 370.77 166.96 ;
      RECT 370.44 166.96 370.77 167.03 ;
      RECT 370.44 166.52 370.77 166.59 ;
      RECT 364.53 166.25 366.14 166.42 ;
      RECT 367.26 166.25 369.97 166.42 ;
      RECT 366.56 166.25 367.09 166.42 ;
      RECT 371.425 165.335 371.935 165.425 ;
      RECT 367.26 171.34 369.97 171.43 ;
      RECT 367.26 171.99 369.97 172.06 ;
      RECT 370.94 171.99 371.935 172.1 ;
      RECT 367.26 171.43 371.935 171.99 ;
      RECT 370.94 165.425 371.935 171.43 ;
      RECT 396.2 162.575 399.77 162.905 ;
      RECT 395.76 163.355 395.93 168.205 ;
      RECT 400.48 162.575 404.05 162.905 ;
      RECT 400.04 163.355 400.21 168.205 ;
      RECT 404.625 162.575 406.33 162.905 ;
      RECT 406.16 162.315 406.33 162.575 ;
      RECT 404.32 163.355 404.49 168.205 ;
      RECT 409.38 162.575 412.95 162.905 ;
      RECT 413.66 162.575 417.23 162.905 ;
      RECT 408.94 163.355 409.11 168.205 ;
      RECT 413.22 163.355 413.39 168.205 ;
      RECT 417.5 163.355 417.67 168.205 ;
      RECT 423.66 160.345 423.99 160.995 ;
      RECT 425.28 160.345 425.61 160.995 ;
      RECT 422.85 160.345 423.18 160.995 ;
      RECT 422.04 160.345 422.37 160.995 ;
      RECT 424.47 160.345 424.8 160.995 ;
      RECT 430.14 160.345 430.47 160.995 ;
      RECT 430.95 160.345 431.28 160.995 ;
      RECT 426.9 160.345 427.23 160.995 ;
      RECT 426.09 160.345 426.42 160.995 ;
      RECT 429.33 160.345 429.66 160.995 ;
      RECT 428.52 160.345 428.85 160.995 ;
      RECT 427.71 160.345 428.04 160.995 ;
      RECT 431.76 160.345 432.09 160.995 ;
      RECT 432.57 160.345 432.9 160.995 ;
      RECT 434.19 160.345 434.52 160.995 ;
      RECT 435 160.345 435.33 160.995 ;
      RECT 433.38 160.345 433.71 160.995 ;
      RECT 435.81 160.345 436.14 160.995 ;
      RECT 436.62 160.345 436.95 160.995 ;
      RECT 26.315 166.82 28.855 166.99 ;
      RECT 28.685 166.305 28.855 166.82 ;
      RECT 19.235 168.46 19.565 168.53 ;
      RECT 25.645 168.02 26.485 168.09 ;
      RECT 25.645 168.46 25.975 168.53 ;
      RECT 19.235 168.02 19.565 168.09 ;
      RECT 19.235 168.09 26.485 168.19 ;
      RECT 19.235 168.19 25.975 168.46 ;
      RECT 27.015 164.73 27.185 165.47 ;
      RECT 27.015 165.47 28.515 165.78 ;
      RECT 28.265 165.78 28.515 166.44 ;
      RECT 30.375 167.03 30.755 167.74 ;
      RECT 29.745 166.41 32.895 166.58 ;
      RECT 29.745 166.58 30.755 167.03 ;
      RECT 29.745 165.98 30.755 166.07 ;
      RECT 29.745 166.24 37.44 166.41 ;
      RECT 29.745 166.07 32.895 166.24 ;
      RECT 31.315 166.82 33.76 167.09 ;
      RECT 33.43 166.795 33.76 166.82 ;
      RECT 33.43 166.785 39.27 166.795 ;
      RECT 38.99 166.515 41.7 166.58 ;
      RECT 33.43 166.58 41.7 166.785 ;
      RECT 31.315 167.09 31.645 169.2 ;
      RECT 31.865 164.015 32.035 165.025 ;
      RECT 32.565 163.45 32.895 163.46 ;
      RECT 32.565 163.73 32.895 163.96 ;
      RECT 32.565 163.46 35.725 163.73 ;
      RECT 37.11 163.175 37.44 163.73 ;
      RECT 33.035 165.09 37.28 165.26 ;
      RECT 37.11 164.985 37.28 165.09 ;
      RECT 37.11 164.815 39.565 164.985 ;
      RECT 33.035 164.425 33.365 165.09 ;
      RECT 33.98 164.68 36.94 164.85 ;
      RECT 33.98 163.12 36.94 163.29 ;
      RECT 34.23 167.02 36.94 167.19 ;
      RECT 34.23 165.46 36.94 165.63 ;
      RECT 34.23 163.9 36.94 164.07 ;
      RECT 36.21 163.885 36.74 163.9 ;
      RECT 38.99 162.845 41.7 163.015 ;
      RECT 42.02 163.57 42.19 164.1 ;
      RECT 41.92 162.9 42.19 163.57 ;
      RECT 42.46 163.625 43.04 164.015 ;
      RECT 42.46 163.295 46.915 163.625 ;
      RECT 42.46 164.015 46.915 164.345 ;
      RECT 37.46 164.305 41.7 164.575 ;
      RECT 38.99 163.625 41.7 163.795 ;
      RECT 39.94 164.815 46.915 164.985 ;
      RECT 42.46 164.985 46.915 165.065 ;
      RECT 42.46 164.735 46.915 164.815 ;
      RECT 38.99 165.185 41.7 165.355 ;
      RECT 41.92 165.41 42.19 166.08 ;
      RECT 42.46 165.785 43.04 166.175 ;
      RECT 42.46 165.455 46.915 165.785 ;
      RECT 42.46 166.175 46.915 166.505 ;
      RECT 37.59 166.99 38.52 167.16 ;
      RECT 37.59 167.16 37.76 167.495 ;
      RECT 37.59 166.965 37.76 166.99 ;
      RECT 39.66 166.955 46.915 167.125 ;
      RECT 42.46 167.125 46.915 167.225 ;
      RECT 42.46 166.895 46.915 166.955 ;
      RECT 47.165 166.175 55.535 166.505 ;
      RECT 47.165 164.015 55.535 164.345 ;
      RECT 47.165 166.895 55.535 167.225 ;
      RECT 47.165 164.735 55.535 165.065 ;
      RECT 47.165 165.455 55.535 165.785 ;
      RECT 47.165 163.295 55.535 163.625 ;
      RECT 43.185 162.755 59.495 163.075 ;
      RECT 56.685 163.075 58.295 163.125 ;
      RECT 59.66 166.505 60.24 166.895 ;
      RECT 55.785 166.895 60.24 167.225 ;
      RECT 55.785 166.175 60.24 166.505 ;
      RECT 59.66 164.345 60.24 164.735 ;
      RECT 55.785 164.735 60.24 165.065 ;
      RECT 55.785 164.015 60.24 164.345 ;
      RECT 64.445 166.45 64.615 170.85 ;
      RECT 75.615 160.565 76.145 160.895 ;
      RECT 86.325 160.565 86.855 160.895 ;
      RECT 87.185 166.45 87.355 170.85 ;
      RECT 303.15 160.565 303.68 160.895 ;
      RECT 302.65 166.45 302.82 170.85 ;
      RECT 313.86 160.565 314.39 160.895 ;
      RECT 325.39 166.45 325.56 170.85 ;
      RECT 330.51 162.755 346.82 163.075 ;
      RECT 331.71 163.075 333.32 163.125 ;
      RECT 329.765 166.505 330.345 166.895 ;
      RECT 329.765 166.895 334.22 167.225 ;
      RECT 329.765 166.175 334.22 166.505 ;
      RECT 329.765 164.345 330.345 164.735 ;
      RECT 329.765 164.735 334.22 165.065 ;
      RECT 329.765 164.015 334.22 164.345 ;
      RECT 334.47 166.895 342.84 167.225 ;
      RECT 334.47 166.175 342.84 166.505 ;
      RECT 334.47 165.455 342.84 165.785 ;
      RECT 334.47 164.735 342.84 165.065 ;
      RECT 334.47 164.015 342.84 164.345 ;
      RECT 334.47 163.295 342.84 163.625 ;
      RECT 346.965 165.785 347.545 166.175 ;
      RECT 343.09 166.175 347.545 166.505 ;
      RECT 343.09 165.455 347.545 165.785 ;
      RECT 346.965 163.625 347.545 164.015 ;
      RECT 343.09 164.015 347.545 164.345 ;
      RECT 343.09 163.295 347.545 163.625 ;
      RECT 343.09 167.125 347.545 167.225 ;
      RECT 343.09 166.895 347.545 166.955 ;
      RECT 343.09 166.955 350.345 167.125 ;
      RECT 343.09 164.985 347.545 165.065 ;
      RECT 343.09 164.735 347.545 164.815 ;
      RECT 343.09 164.815 350.065 164.985 ;
      RECT 348.305 163.625 351.015 163.795 ;
      RECT 348.305 162.845 351.015 163.015 ;
      RECT 348.305 166.515 351.015 166.58 ;
      RECT 348.305 166.58 356.575 166.785 ;
      RECT 350.735 166.785 356.575 166.795 ;
      RECT 356.245 166.795 356.575 166.82 ;
      RECT 356.245 166.82 358.69 167.09 ;
      RECT 358.36 167.09 358.69 169.2 ;
      RECT 348.305 166.07 351.015 166.135 ;
      RECT 348.305 165.83 356.575 166.07 ;
      RECT 356.245 165.56 358.69 165.83 ;
      RECT 358.36 163.45 358.69 165.56 ;
      RECT 348.305 165.185 351.015 165.355 ;
      RECT 348.305 164.305 352.545 164.575 ;
      RECT 347.815 165.41 348.085 166.08 ;
      RECT 347.815 163.57 347.985 164.1 ;
      RECT 347.815 162.9 348.085 163.57 ;
      RECT 352.565 163.175 352.895 163.73 ;
      RECT 351.485 166.99 352.415 167.16 ;
      RECT 407.57 180.955 419.04 181.135 ;
      RECT 407.57 162.575 408.805 162.905 ;
      RECT 407.57 157.045 408.33 162.575 ;
      RECT 407.57 174.495 408.805 174.825 ;
      RECT 417.805 162.575 419.04 162.905 ;
      RECT 417.805 174.495 419.04 174.825 ;
      RECT 418.28 168.865 419.04 174.495 ;
      RECT 417.805 168.535 419.04 168.865 ;
      RECT 418.28 162.905 419.04 168.535 ;
      RECT 418.28 180.785 419.04 180.955 ;
      RECT 418.28 174.825 419.04 180.455 ;
      RECT 407.57 174.825 408.33 180.455 ;
      RECT 407.57 180.785 408.33 180.955 ;
      RECT 407.57 168.865 408.33 174.495 ;
      RECT 407.57 168.535 408.805 168.865 ;
      RECT 407.57 162.905 408.33 168.535 ;
      RECT 418.28 157.045 419.04 162.575 ;
      RECT 417.805 180.455 419.04 180.785 ;
      RECT 407.57 180.455 408.805 180.785 ;
      RECT 412.75 155.16 413.08 155.67 ;
      RECT 412.83 155.09 413 155.16 ;
      RECT 411.97 155.16 412.3 155.67 ;
      RECT 412.05 155.09 412.22 155.16 ;
      RECT 413.53 155.16 413.86 155.67 ;
      RECT 413.61 155.09 413.78 155.16 ;
      RECT 410.88 155.16 411.52 155.67 ;
      RECT 410.88 153.4 411.05 155.16 ;
      RECT 413.22 157.395 413.39 162.245 ;
      RECT 408.94 157.395 409.11 162.245 ;
      RECT 414.78 153.4 414.95 154.75 ;
      RECT 414 153.4 414.17 154.75 ;
      RECT 414.31 155.16 414.64 155.67 ;
      RECT 414.39 155.09 414.56 155.16 ;
      RECT 415.09 155.16 415.73 155.67 ;
      RECT 415.56 153.4 415.73 155.16 ;
      RECT 417.5 157.395 417.67 162.245 ;
      RECT 450.32 154.105 455.165 154.635 ;
      RECT 450.32 158.535 455.165 159.065 ;
      RECT 450.32 153.395 454.735 153.925 ;
      RECT 450.32 157.825 456.025 158.355 ;
      RECT 450.32 152.49 455.595 153.02 ;
      RECT 450.32 156.92 454.305 157.45 ;
      RECT 448.865 153.99 449.875 154.16 ;
      RECT 448.865 153.11 449.875 153.28 ;
      RECT 448.865 152.23 449.875 152.4 ;
      RECT 448.865 154.815 458.585 155.08 ;
      RECT 448.865 158.42 449.875 158.59 ;
      RECT 448.865 157.54 449.875 157.71 ;
      RECT 448.865 155.74 458.585 156.005 ;
      RECT 448.865 156.66 449.875 156.83 ;
      RECT 448.865 159.245 458.585 159.51 ;
      RECT 456.695 153.055 458.575 153.335 ;
      RECT 457.565 156.605 459.345 156.885 ;
      RECT 459.095 155.59 459.345 156.605 ;
      RECT 459.095 158.645 459.345 159.66 ;
      RECT 457.565 158.365 459.345 158.645 ;
      RECT 459.095 156.885 459.345 158.365 ;
      RECT 456.695 157.485 458.575 157.765 ;
      RECT 456.675 151.79 457.345 151.96 ;
      RECT 456.675 156.22 457.345 156.39 ;
      RECT 24.425 163.84 25.475 163.94 ;
      RECT 19.235 163.77 19.565 163.84 ;
      RECT 19.235 163.33 19.565 163.4 ;
      RECT 24.425 163.77 25.975 163.84 ;
      RECT 23.865 163.94 25.475 164.11 ;
      RECT 25.645 163.33 25.975 163.4 ;
      RECT 19.235 163.4 25.975 163.77 ;
      RECT 19.235 166.96 19.565 167.03 ;
      RECT 19.235 166.52 19.565 166.59 ;
      RECT 19.235 166.59 25.975 166.96 ;
      RECT 25.645 166.96 25.975 167.03 ;
      RECT 25.645 166.52 25.975 166.59 ;
      RECT 19.73 164.89 26.485 165.06 ;
      RECT 26.315 163.875 26.485 164.89 ;
      RECT 19.235 166.08 19.565 166.15 ;
      RECT 19.235 165.64 19.565 165.71 ;
      RECT 19.235 165.71 25.975 166.08 ;
      RECT 25.645 166.08 25.975 166.15 ;
      RECT 19.73 164.82 25.475 164.89 ;
      RECT 28.915 163.875 29.495 164.06 ;
      RECT 28.915 163.53 29.495 163.705 ;
      RECT 26.315 163.705 29.495 163.875 ;
      RECT 25.645 165.06 25.975 165.71 ;
      RECT 19.235 164.65 19.565 164.72 ;
      RECT 19.235 164.21 19.565 164.28 ;
      RECT 25.645 164.19 25.815 164.21 ;
      RECT 19.235 164.28 25.975 164.65 ;
      RECT 25.645 164.65 25.975 164.72 ;
      RECT 25.645 164.21 25.975 164.28 ;
      RECT 18.07 165.335 18.58 165.425 ;
      RECT 20.035 171.34 22.745 171.43 ;
      RECT 20.035 171.99 22.745 172.06 ;
      RECT 18.07 171.99 19.065 172.1 ;
      RECT 18.07 171.43 22.745 171.99 ;
      RECT 18.07 165.425 19.065 171.43 ;
      RECT 19.73 167.13 25.475 167.3 ;
      RECT 19.73 165.37 25.475 165.54 ;
      RECT 19.73 163.06 25.475 163.23 ;
      RECT 20.545 162.645 21.135 162.86 ;
      RECT 20.545 162.445 38.05 162.645 ;
      RECT 37.85 162.645 38.05 163.965 ;
      RECT 37.85 163.965 38.52 164.135 ;
      RECT 20.035 163.94 22.745 164.11 ;
      RECT 22.915 163.94 23.245 164.11 ;
      RECT 23.865 166.25 25.475 166.42 ;
      RECT 20.035 166.25 22.745 166.42 ;
      RECT 22.915 166.25 23.445 166.42 ;
      RECT 26.955 164.36 30.175 164.53 ;
      RECT 26.955 164.15 27.965 164.36 ;
      RECT 28.695 164.53 29.365 164.89 ;
      RECT 29.845 164.53 30.175 164.72 ;
      RECT 26.955 163.27 28.005 163.44 ;
      RECT 29.845 163.27 30.755 164.105 ;
      RECT 30.375 164.105 30.755 164.69 ;
      RECT 31.315 165.56 33.76 165.83 ;
      RECT 38.99 166.07 41.7 166.135 ;
      RECT 33.43 165.83 41.7 166.07 ;
      RECT 31.315 163.45 31.645 165.56 ;
      RECT 27.725 164.87 28.055 165.1 ;
      RECT 27.665 164.7 28.055 164.87 ;
      RECT 27.725 165.1 30.755 165.27 ;
      RECT 28.915 165.27 29.255 165.72 ;
      RECT 29.085 165.72 29.255 167.145 ;
      RECT 26.985 166.15 28.005 166.32 ;
      RECT 26.985 166.32 27.995 166.51 ;
      RECT 26.985 165.98 27.995 166.15 ;
      RECT 26.315 166.99 26.485 168.02 ;
      RECT 342.28 155.295 344.99 155.465 ;
      RECT 342.28 156.855 344.99 157.025 ;
      RECT 345.75 157.25 346.28 157.42 ;
      RECT 345.75 157.42 345.92 157.65 ;
      RECT 345.75 156.3 345.92 157.25 ;
      RECT 345.21 154.87 345.92 155.54 ;
      RECT 345.21 155.54 345.38 157.58 ;
      RECT 346.47 157.635 349.18 157.805 ;
      RECT 346.185 156.075 349.18 156.245 ;
      RECT 346.14 153.215 349.14 153.385 ;
      RECT 346.47 156.855 349.18 157.025 ;
      RECT 346.14 155.525 349.15 155.695 ;
      RECT 346.14 153.765 348.92 153.935 ;
      RECT 344.865 153.765 345.395 153.935 ;
      RECT 345.21 153.24 345.38 153.765 ;
      RECT 344.79 152.32 345.38 152.49 ;
      RECT 345.21 152.49 345.38 152.63 ;
      RECT 345.21 151.96 345.38 152.32 ;
      RECT 355.16 159.1 356.85 159.27 ;
      RECT 355.715 151.67 360.565 151.84 ;
      RECT 355.715 151.84 355.885 154.735 ;
      RECT 357.275 151.84 357.445 154.735 ;
      RECT 358.835 151.84 359.005 154.735 ;
      RECT 360.395 151.84 360.565 154.735 ;
      RECT 354.935 152.01 355.105 154.72 ;
      RECT 354.935 156.345 355.465 156.875 ;
      RECT 354.935 156.875 355.105 158.88 ;
      RECT 354.935 155.975 355.105 156.345 ;
      RECT 354.355 147.88 354.525 159.775 ;
      RECT 354.355 147.71 369.515 147.88 ;
      RECT 354.355 159.775 369.515 159.945 ;
      RECT 369.345 147.88 369.515 159.775 ;
      RECT 354.415 147.69 369.515 147.71 ;
      RECT 358.055 152.01 358.225 154.72 ;
      RECT 361.175 152.01 361.345 154.735 ;
      RECT 359.615 152.01 359.785 154.72 ;
      RECT 356.495 152.01 356.665 154.72 ;
      RECT 356.215 155.83 358.145 156 ;
      RECT 356.215 156 356.385 158.88 ;
      RECT 357.975 156 358.145 158.88 ;
      RECT 357.095 159.045 357.625 159.575 ;
      RECT 357.095 156.17 357.265 159.045 ;
      RECT 358.2 159.1 361.59 159.27 ;
      RECT 358.315 158.675 358.845 159.1 ;
      RECT 359.805 156.17 359.975 158.88 ;
      RECT 358.895 156.455 359.425 156.985 ;
      RECT 359.255 156.985 359.425 158.88 ;
      RECT 359.255 156.17 359.425 156.455 ;
      RECT 361.565 156.17 361.735 158.88 ;
      RECT 360.685 155.945 360.855 158.88 ;
      RECT 364.55 155.44 364.72 158.88 ;
      RECT 363.71 155.105 364.72 155.44 ;
      RECT 361.725 152.01 361.895 154.72 ;
      RECT 364.365 152.01 364.535 154.865 ;
      RECT 366.125 155.015 368.055 155.06 ;
      RECT 366.125 154.89 368.06 155.015 ;
      RECT 366.125 152.01 366.295 154.89 ;
      RECT 367.885 152.01 368.055 152.89 ;
      RECT 367.885 152.89 368.06 154.89 ;
      RECT 367.005 152.01 367.175 154.72 ;
      RECT 365.245 152.01 365.415 154.72 ;
      RECT 363.485 152.01 363.655 154.72 ;
      RECT 361.88 155.27 362.55 155.44 ;
      RECT 361.76 159.1 362.29 159.27 ;
      RECT 361.905 159.27 362.115 159.44 ;
      RECT 361.905 155.44 362.115 159.1 ;
      RECT 363.295 155.7 363.925 155.87 ;
      RECT 363.295 155.44 363.465 155.7 ;
      RECT 362.795 155.27 363.465 155.44 ;
      RECT 363.755 155.87 363.925 156.845 ;
      RECT 365.47 155.27 368.86 155.44 ;
      RECT 366.35 158.74 366.88 159.27 ;
      RECT 366.71 155.44 366.88 158.74 ;
      RECT 364.705 159.1 365.375 159.27 ;
      RECT 367.265 159.1 367.935 159.27 ;
      RECT 367.365 159.27 367.895 159.285 ;
      RECT 365.43 156.17 365.6 158.88 ;
      RECT 363.325 156.17 363.495 158.88 ;
      RECT 362.605 152.01 362.775 154.72 ;
      RECT 362.445 155.945 362.615 158.88 ;
      RECT 368.765 152.01 368.935 154.72 ;
      RECT 367.99 156.17 368.16 158.88 ;
      RECT 387.7 158.57 388.03 159.22 ;
      RECT 390.22 158.57 390.55 159.22 ;
      RECT 389.59 158.57 389.92 159.22 ;
      RECT 388.33 158.57 388.66 159.22 ;
      RECT 388.96 158.57 389.29 159.22 ;
      RECT 387.7 157.54 388.03 158.19 ;
      RECT 388.96 157.54 389.29 158.19 ;
      RECT 389.59 157.54 389.92 158.19 ;
      RECT 390.22 157.54 390.55 158.19 ;
      RECT 388.33 157.54 388.66 158.19 ;
      RECT 394.39 156.865 405.86 157.045 ;
      RECT 394.39 180.955 405.86 181.135 ;
      RECT 394.39 162.575 395.625 162.905 ;
      RECT 405.1 157.045 405.86 162.32 ;
      RECT 405.68 163.075 405.86 163.17 ;
      RECT 394.39 174.495 395.625 174.825 ;
      RECT 404.625 174.495 405.86 174.825 ;
      RECT 405.1 168.865 405.86 174.495 ;
      RECT 404.625 168.535 405.86 168.865 ;
      RECT 405.1 163.17 405.86 168.535 ;
      RECT 405.1 180.785 405.86 180.955 ;
      RECT 405.1 174.825 405.86 180.455 ;
      RECT 394.39 180.785 395.15 180.955 ;
      RECT 394.39 174.825 395.15 180.455 ;
      RECT 394.39 168.865 395.15 174.495 ;
      RECT 394.39 168.535 395.625 168.865 ;
      RECT 394.39 162.905 395.15 168.535 ;
      RECT 394.39 157.045 395.15 162.575 ;
      RECT 404.625 180.455 405.86 180.785 ;
      RECT 394.39 180.455 395.625 180.785 ;
      RECT 392.91 155.42 395.015 155.75 ;
      RECT 392.91 155.16 393.08 155.42 ;
      RECT 395.94 155.42 397.47 155.75 ;
      RECT 395.76 157.395 395.93 162.245 ;
      RECT 390.85 158.57 391.18 159.22 ;
      RECT 390.85 157.54 391.18 158.19 ;
      RECT 400.5 155.42 402.03 155.75 ;
      RECT 398.22 155.42 399.75 155.75 ;
      RECT 400.04 157.395 400.21 162.245 ;
      RECT 402.78 155.42 404.31 155.75 ;
      RECT 404.32 157.395 404.49 162.245 ;
      RECT 413.22 153.375 413.39 154.75 ;
      RECT 412.44 153.4 412.61 154.75 ;
      RECT 411.66 153.4 411.83 154.75 ;
      RECT 407.57 156.865 419.04 157.045 ;
      RECT 21.145 155.27 24.535 155.44 ;
      RECT 23.125 158.74 23.655 159.27 ;
      RECT 23.125 155.44 23.295 158.74 ;
      RECT 20.49 147.71 35.65 147.88 ;
      RECT 35.48 147.88 35.65 159.775 ;
      RECT 20.49 159.775 35.65 159.945 ;
      RECT 20.49 147.88 20.66 159.775 ;
      RECT 20.49 147.69 35.59 147.71 ;
      RECT 24.63 159.1 25.3 159.27 ;
      RECT 22.07 159.1 22.74 159.27 ;
      RECT 22.11 159.27 22.64 159.285 ;
      RECT 21.845 156.17 22.015 158.88 ;
      RECT 24.405 156.17 24.575 158.88 ;
      RECT 28.11 152.01 28.28 154.72 ;
      RECT 26.35 152.01 26.52 154.72 ;
      RECT 28.66 152.01 28.83 154.735 ;
      RECT 30.22 152.01 30.39 154.72 ;
      RECT 29.44 151.67 34.29 151.84 ;
      RECT 31 151.84 31.17 154.735 ;
      RECT 29.44 151.84 29.61 154.735 ;
      RECT 32.56 151.84 32.73 154.735 ;
      RECT 34.12 151.84 34.29 154.735 ;
      RECT 27.455 155.27 28.125 155.44 ;
      RECT 27.715 159.1 28.245 159.27 ;
      RECT 27.89 159.27 28.1 159.44 ;
      RECT 27.89 155.44 28.1 159.1 ;
      RECT 26.08 155.7 26.71 155.87 ;
      RECT 26.54 155.44 26.71 155.7 ;
      RECT 26.54 155.27 27.21 155.44 ;
      RECT 26.08 155.87 26.25 156.845 ;
      RECT 28.415 159.1 31.805 159.27 ;
      RECT 31.16 158.675 31.69 159.1 ;
      RECT 30.58 156.455 31.11 156.985 ;
      RECT 30.58 156.985 30.75 158.88 ;
      RECT 30.58 156.17 30.75 156.455 ;
      RECT 30.03 156.17 30.2 158.88 ;
      RECT 26.51 156.17 26.68 158.88 ;
      RECT 27.23 152.01 27.4 154.72 ;
      RECT 29.15 155.945 29.32 158.88 ;
      RECT 27.39 155.945 27.56 158.88 ;
      RECT 28.27 156.17 28.44 158.88 ;
      RECT 33.155 159.1 34.845 159.27 ;
      RECT 31.78 152.01 31.95 154.72 ;
      RECT 34.9 152.01 35.07 154.72 ;
      RECT 33.34 152.01 33.51 154.72 ;
      RECT 31.86 155.83 33.79 156 ;
      RECT 31.86 156 32.03 158.88 ;
      RECT 33.62 156 33.79 158.88 ;
      RECT 34.54 156.345 35.07 156.875 ;
      RECT 34.9 156.875 35.07 158.88 ;
      RECT 34.9 155.975 35.07 156.345 ;
      RECT 32.38 159.045 32.91 159.575 ;
      RECT 32.74 156.17 32.91 159.045 ;
      RECT 40.825 157.635 43.535 157.805 ;
      RECT 40.825 156.075 43.82 156.245 ;
      RECT 40.865 153.215 43.865 153.385 ;
      RECT 40.825 156.855 43.535 157.025 ;
      RECT 40.855 155.525 43.865 155.695 ;
      RECT 41.085 153.765 43.865 153.935 ;
      RECT 43.725 157.25 44.255 157.42 ;
      RECT 44.085 157.42 44.255 157.65 ;
      RECT 44.085 156.3 44.255 157.25 ;
      RECT 44.085 154.87 44.795 155.54 ;
      RECT 44.625 155.54 44.795 157.58 ;
      RECT 45.345 151.805 48.055 151.975 ;
      RECT 47.895 154.685 48.065 156.075 ;
      RECT 47.895 156.245 48.065 157.635 ;
      RECT 45.015 154.515 48.065 154.685 ;
      RECT 45.015 156.075 48.065 156.245 ;
      RECT 45.015 157.635 48.065 157.805 ;
      RECT 45.345 153.965 48.055 154.135 ;
      RECT 45.015 155.295 47.725 155.465 ;
      RECT 45.015 156.855 47.725 157.025 ;
      RECT 44.61 153.765 45.14 153.935 ;
      RECT 44.625 153.24 44.795 153.765 ;
      RECT 44.625 152.32 45.215 152.49 ;
      RECT 44.625 152.49 44.795 152.63 ;
      RECT 44.625 151.96 44.795 152.32 ;
      RECT 57.655 151.465 57.985 152.865 ;
      RECT 57.025 151.465 57.355 152.865 ;
      RECT 55.765 151.465 56.095 152.865 ;
      RECT 56.395 151.465 56.725 152.865 ;
      RECT 58.285 151.465 58.615 152.865 ;
      RECT 60.175 151.465 60.505 152.865 ;
      RECT 59.545 151.465 59.875 152.865 ;
      RECT 58.915 151.465 59.245 152.865 ;
      RECT 57.025 157.265 57.985 157.775 ;
      RECT 55.765 157.265 56.725 157.775 ;
      RECT 59.545 157.265 60.505 157.775 ;
      RECT 58.285 157.265 59.245 157.775 ;
      RECT 64.6 157.01 72.88 157.18 ;
      RECT 60.805 151.465 61.135 152.865 ;
      RECT 62.065 151.465 62.395 152.865 ;
      RECT 62.695 151.465 63.025 152.865 ;
      RECT 60.805 157.265 61.765 157.775 ;
      RECT 61.435 151.465 61.765 152.865 ;
      RECT 62.065 157.265 63.025 157.775 ;
      RECT 73.16 157.01 77.16 157.18 ;
      RECT 77.57 157.01 85.72 157.18 ;
      RECT 304.285 157.01 312.435 157.18 ;
      RECT 312.845 157.01 316.845 157.18 ;
      RECT 317.125 157.01 325.405 157.18 ;
      RECT 327.61 151.465 327.94 152.865 ;
      RECT 326.98 151.465 327.31 152.865 ;
      RECT 328.87 151.465 329.2 152.865 ;
      RECT 329.5 151.465 329.83 152.865 ;
      RECT 330.13 151.465 330.46 152.865 ;
      RECT 328.24 151.465 328.57 152.865 ;
      RECT 332.02 151.465 332.35 152.865 ;
      RECT 332.65 151.465 332.98 152.865 ;
      RECT 330.76 151.465 331.09 152.865 ;
      RECT 331.39 151.465 331.72 152.865 ;
      RECT 326.98 157.265 327.94 157.775 ;
      RECT 328.24 157.265 329.2 157.775 ;
      RECT 329.5 157.265 330.46 157.775 ;
      RECT 330.76 157.265 331.72 157.775 ;
      RECT 332.02 157.265 332.98 157.775 ;
      RECT 333.91 151.465 334.24 152.865 ;
      RECT 333.28 151.465 333.61 152.865 ;
      RECT 333.28 157.265 334.24 157.775 ;
      RECT 341.95 151.805 344.66 151.975 ;
      RECT 341.94 154.685 342.11 156.075 ;
      RECT 341.94 156.245 342.11 157.635 ;
      RECT 341.94 154.515 344.99 154.685 ;
      RECT 341.94 156.075 344.99 156.245 ;
      RECT 341.94 157.635 344.99 157.805 ;
      RECT 341.95 153.965 344.66 154.135 ;
      RECT 346.14 151.455 348.85 151.625 ;
      RECT 345.75 150.575 348.85 150.745 ;
      RECT 345.75 149.85 345.92 150.575 ;
      RECT 345.44 151.455 345.97 151.625 ;
      RECT 345.75 151.625 345.92 154.59 ;
      RECT 345.75 151.2 345.92 151.455 ;
      RECT 354.935 148.79 355.105 151.5 ;
      RECT 355.715 148.63 355.885 151.5 ;
      RECT 359.615 148.79 359.785 151.5 ;
      RECT 361.175 148.79 361.345 151.5 ;
      RECT 356.495 148.79 356.665 151.5 ;
      RECT 357.275 148.63 357.445 151.5 ;
      RECT 358.835 148.63 359.005 151.5 ;
      RECT 360.395 148.63 360.565 151.5 ;
      RECT 358.055 148.79 358.225 151.5 ;
      RECT 363.515 148.63 363.685 151.5 ;
      RECT 365.075 148.63 365.245 151.5 ;
      RECT 366.635 148.63 366.805 151.5 ;
      RECT 364.295 148.79 364.465 151.5 ;
      RECT 365.855 148.79 366.025 151.5 ;
      RECT 367.415 148.63 367.585 151.5 ;
      RECT 362.735 148.79 362.905 151.5 ;
      RECT 361.955 148.63 362.125 151.5 ;
      RECT 365.705 144.1 368.455 144.27 ;
      RECT 365.705 143.67 368.415 143.84 ;
      RECT 386.27 144.955 386.6 145.605 ;
      RECT 386.9 144.955 387.23 145.605 ;
      RECT 388.79 144.955 389.12 145.605 ;
      RECT 388.16 144.955 388.49 145.605 ;
      RECT 387.53 144.955 387.86 145.605 ;
      RECT 389.42 144.955 389.75 145.605 ;
      RECT 390.05 144.955 390.38 145.605 ;
      RECT 387.7 148.495 388.03 149.145 ;
      RECT 388.96 148.495 389.29 149.145 ;
      RECT 389.59 148.495 389.92 149.145 ;
      RECT 390.22 148.495 390.55 149.145 ;
      RECT 388.33 148.495 388.66 149.145 ;
      RECT 391.55 148.085 391.73 198.9 ;
      RECT 387.15 147.725 391.73 148.085 ;
      RECT 387.15 148.085 387.33 198.9 ;
      RECT 387.15 198.9 391.73 199.2 ;
      RECT 395.48 148.22 395.65 155.23 ;
      RECT 394.2 148.24 394.37 155.23 ;
      RECT 390.68 144.955 391.01 145.605 ;
      RECT 391.31 144.955 391.64 145.605 ;
      RECT 391.94 144.955 392.27 145.605 ;
      RECT 392.57 144.955 392.9 145.605 ;
      RECT 393.2 144.955 393.53 145.605 ;
      RECT 393.83 144.955 394.16 145.605 ;
      RECT 394.46 144.955 394.79 145.605 ;
      RECT 390.85 148.495 391.18 149.145 ;
      RECT 400.04 148.22 400.21 155.23 ;
      RECT 397.76 148.24 397.93 155.23 ;
      RECT 396.46 147.345 399.87 147.515 ;
      RECT 400.135 144.89 401.825 145.285 ;
      RECT 397.855 144.89 399.545 145.285 ;
      RECT 396.515 146.115 397.045 147.145 ;
      RECT 399.635 146.115 400.165 147.145 ;
      RECT 398.595 145.7 398.765 146.115 ;
      RECT 397.475 145.53 398.765 145.7 ;
      RECT 398.595 146.115 399.205 147.125 ;
      RECT 397.475 144.815 397.645 145.53 ;
      RECT 397.475 145.7 397.645 147.125 ;
      RECT 397.895 146.115 398.425 147.145 ;
      RECT 402.32 148.24 402.49 155.23 ;
      RECT 404.6 148.22 404.77 155.23 ;
      RECT 404.695 144.89 406.385 145.285 ;
      RECT 402.415 144.89 404.105 145.285 ;
      RECT 407.57 145.91 413 146.08 ;
      RECT 407.175 146.3 407.345 155.175 ;
      RECT 405.235 155.42 406.05 155.75 ;
      RECT 405.88 148.22 406.05 155.42 ;
      RECT 407.665 146.3 408.415 155.305 ;
      RECT 409.515 146.3 410.27 152.785 ;
      RECT 409.515 152.785 409.685 155.175 ;
      RECT 411.985 144.89 413.675 145.285 ;
      RECT 409.705 144.89 411.395 145.285 ;
      RECT 413.61 145.91 419.04 146.08 ;
      RECT 408.735 146.3 408.905 155.175 ;
      RECT 410.88 146.33 411.05 152.35 ;
      RECT 412.44 146.33 412.61 152.35 ;
      RECT 411.37 146.3 412.12 152.785 ;
      RECT 412.93 146.3 413.68 152.785 ;
      RECT 419.265 146.3 419.435 155.175 ;
      RECT 416.34 146.3 417.095 152.785 ;
      RECT 416.925 152.785 417.095 155.175 ;
      RECT 416.545 144.89 418.235 145.285 ;
      RECT 414.265 144.89 415.955 145.285 ;
      RECT 418.195 146.3 418.945 155.305 ;
      RECT 417.705 146.3 417.875 155.175 ;
      RECT 414 146.33 414.17 152.35 ;
      RECT 414.49 146.3 415.24 152.785 ;
      RECT 415.56 146.33 415.73 152.35 ;
      RECT 447.765 144.475 460.045 145.045 ;
      RECT 447.765 143.695 460.045 144.265 ;
      RECT 450.32 149.675 455.165 150.205 ;
      RECT 450.32 148.965 454.735 149.495 ;
      RECT 450.32 148.06 454.305 148.59 ;
      RECT 448.865 151.31 458.585 151.575 ;
      RECT 448.865 149.56 449.875 149.73 ;
      RECT 448.865 148.68 449.875 148.85 ;
      RECT 448.865 146.88 458.585 147.145 ;
      RECT 448.865 147.8 449.875 147.97 ;
      RECT 448.865 150.385 458.585 150.65 ;
      RECT 457.565 147.745 459.345 148.025 ;
      RECT 459.095 146.73 459.345 147.745 ;
      RECT 459.095 149.785 459.345 150.8 ;
      RECT 457.565 149.505 459.345 149.785 ;
      RECT 459.095 148.025 459.345 149.505 ;
      RECT 456.695 148.625 458.575 148.905 ;
      RECT 456.675 147.36 457.345 147.53 ;
      RECT 457.565 153.935 459.345 154.215 ;
      RECT 459.095 154.215 459.345 155.23 ;
      RECT 459.095 152.455 459.345 153.935 ;
      RECT 457.565 152.175 459.345 152.455 ;
      RECT 459.095 151.16 459.345 152.175 ;
      RECT 25.285 155.44 25.455 158.88 ;
      RECT 25.285 155.105 26.295 155.44 ;
      RECT 21.95 155.015 23.88 155.06 ;
      RECT 21.945 154.89 23.88 155.015 ;
      RECT 21.95 152.01 22.12 152.89 ;
      RECT 23.71 152.01 23.88 154.89 ;
      RECT 21.945 152.89 22.12 154.89 ;
      RECT 25.47 152.01 25.64 154.865 ;
      RECT 21.07 152.01 21.24 154.72 ;
      RECT 22.83 152.01 23 154.72 ;
      RECT 24.59 152.01 24.76 154.72 ;
      RECT 457.335 138.375 460.045 138.545 ;
      RECT 460.595 141 460.765 144.62 ;
      RECT 24.76 148.63 24.93 151.5 ;
      RECT 23.2 148.63 23.37 151.5 ;
      RECT 25.54 148.79 25.71 151.5 ;
      RECT 23.98 148.79 24.15 151.5 ;
      RECT 22.42 148.63 22.59 151.5 ;
      RECT 21.55 144.1 24.3 144.27 ;
      RECT 21.59 143.67 24.3 143.84 ;
      RECT 30.22 148.79 30.39 151.5 ;
      RECT 28.66 148.79 28.83 151.5 ;
      RECT 27.1 148.79 27.27 151.5 ;
      RECT 31 148.63 31.17 151.5 ;
      RECT 29.44 148.63 29.61 151.5 ;
      RECT 27.88 148.63 28.05 151.5 ;
      RECT 26.32 148.63 26.49 151.5 ;
      RECT 33.34 148.79 33.51 151.5 ;
      RECT 34.9 148.79 35.07 151.5 ;
      RECT 34.12 148.63 34.29 151.5 ;
      RECT 32.56 148.63 32.73 151.5 ;
      RECT 31.78 148.79 31.95 151.5 ;
      RECT 41.115 144.405 46.255 144.575 ;
      RECT 46.085 144.01 46.255 144.405 ;
      RECT 44.455 144.575 46.255 145.44 ;
      RECT 41.03 145.725 43.865 145.895 ;
      RECT 41.155 146.605 43.865 146.775 ;
      RECT 41.155 147.485 43.865 147.655 ;
      RECT 41.155 149.795 43.865 149.965 ;
      RECT 41.155 149.245 43.865 149.415 ;
      RECT 41.155 151.455 43.865 151.625 ;
      RECT 41.155 150.575 44.255 150.745 ;
      RECT 44.085 149.85 44.255 150.575 ;
      RECT 44.625 148.35 45.155 148.52 ;
      RECT 44.625 148.52 44.795 149.025 ;
      RECT 44.625 147.675 44.795 148.35 ;
      RECT 44.085 149.335 44.795 149.505 ;
      RECT 44.625 149.505 44.795 149.78 ;
      RECT 44.625 150.31 44.795 150.87 ;
      RECT 44.085 147.84 44.255 149.335 ;
      RECT 44.6 149.78 44.795 150.31 ;
      RECT 43.665 145.285 44.255 145.455 ;
      RECT 44.035 145.455 44.255 146.96 ;
      RECT 45.22 146.455 48.055 146.625 ;
      RECT 44.265 147.335 44.795 147.505 ;
      RECT 44.625 146.61 44.795 147.335 ;
      RECT 47.045 145.905 48.055 146.075 ;
      RECT 45.22 149.645 48.055 149.815 ;
      RECT 45.22 149.095 48.055 149.265 ;
      RECT 44.035 151.455 44.565 151.625 ;
      RECT 44.085 151.625 44.255 154.59 ;
      RECT 44.085 151.2 44.255 151.455 ;
      RECT 45.345 148.215 48.055 148.385 ;
      RECT 51.89 146.815 54.26 146.985 ;
      RECT 50.955 158.215 86.525 158.385 ;
      RECT 50.955 145.325 51.125 158.215 ;
      RECT 86.355 145.325 86.525 158.215 ;
      RECT 55.165 145.325 55.335 158.215 ;
      RECT 50.955 145.155 86.525 145.325 ;
      RECT 63.395 145.325 63.985 158.215 ;
      RECT 58.215 146.39 58.745 146.555 ;
      RECT 57.655 146.555 58.745 146.56 ;
      RECT 57.655 146.56 58.615 147.065 ;
      RECT 56.395 146.555 57.355 147.065 ;
      RECT 55.565 146.39 56.095 146.56 ;
      RECT 55.765 146.56 56.095 147.065 ;
      RECT 60.735 146.39 61.265 146.555 ;
      RECT 60.175 146.555 61.265 146.56 ;
      RECT 60.175 146.56 61.135 147.065 ;
      RECT 58.915 146.555 59.875 147.065 ;
      RECT 64.715 146.36 68.485 146.53 ;
      RECT 61.435 146.555 62.395 147.065 ;
      RECT 62.695 146.39 63.225 146.56 ;
      RECT 62.695 146.56 63.025 147.065 ;
      RECT 68.995 146.36 72.765 146.53 ;
      RECT 73.315 146.36 77.045 146.53 ;
      RECT 77.555 146.36 81.32 146.53 ;
      RECT 81.835 146.36 85.605 146.53 ;
      RECT 338.88 145.325 339.05 158.215 ;
      RECT 303.48 145.325 303.65 158.215 ;
      RECT 303.48 158.215 339.05 158.385 ;
      RECT 303.48 145.155 339.05 145.325 ;
      RECT 334.67 145.325 334.84 158.215 ;
      RECT 326.02 145.325 326.61 158.215 ;
      RECT 304.4 146.36 308.17 146.53 ;
      RECT 308.685 146.36 312.45 146.53 ;
      RECT 312.96 146.36 316.69 146.53 ;
      RECT 317.24 146.36 321.01 146.53 ;
      RECT 321.52 146.36 325.29 146.53 ;
      RECT 326.78 146.39 327.31 146.56 ;
      RECT 326.98 146.56 327.31 147.065 ;
      RECT 331.26 146.39 331.79 146.555 ;
      RECT 331.26 146.555 332.35 146.56 ;
      RECT 331.39 146.56 332.35 147.065 ;
      RECT 332.65 146.555 333.61 147.065 ;
      RECT 328.74 146.39 329.27 146.555 ;
      RECT 328.74 146.555 329.83 146.56 ;
      RECT 328.87 146.56 329.83 147.065 ;
      RECT 330.13 146.555 331.09 147.065 ;
      RECT 327.61 146.555 328.57 147.065 ;
      RECT 335.745 146.815 338.115 146.985 ;
      RECT 333.91 146.39 334.44 146.56 ;
      RECT 333.91 146.56 334.24 147.065 ;
      RECT 343.75 144.405 348.89 144.575 ;
      RECT 343.75 144.01 343.92 144.405 ;
      RECT 343.75 144.575 345.55 145.44 ;
      RECT 341.95 146.455 344.785 146.625 ;
      RECT 341.95 145.905 342.96 146.075 ;
      RECT 341.95 149.645 344.785 149.815 ;
      RECT 341.95 149.095 344.785 149.265 ;
      RECT 341.95 148.215 344.66 148.385 ;
      RECT 344.85 148.35 345.38 148.52 ;
      RECT 345.21 148.52 345.38 149.025 ;
      RECT 345.21 147.675 345.38 148.35 ;
      RECT 345.21 149.335 345.92 149.505 ;
      RECT 345.21 149.505 345.38 149.78 ;
      RECT 345.21 150.31 345.38 150.87 ;
      RECT 345.75 147.84 345.92 149.335 ;
      RECT 345.21 149.78 345.405 150.31 ;
      RECT 345.75 145.285 346.34 145.455 ;
      RECT 345.75 145.455 345.97 146.96 ;
      RECT 346.14 145.725 348.975 145.895 ;
      RECT 346.14 146.605 348.85 146.775 ;
      RECT 346.14 147.485 348.85 147.655 ;
      RECT 345.21 147.335 345.74 147.505 ;
      RECT 345.21 146.61 345.38 147.335 ;
      RECT 346.14 149.795 348.85 149.965 ;
      RECT 346.14 149.245 348.85 149.415 ;
      RECT 316.685 141.94 317.645 142.45 ;
      RECT 317.945 141.94 318.905 142.45 ;
      RECT 319.205 141.94 320.165 142.45 ;
      RECT 320.595 141.94 321.555 142.45 ;
      RECT 315.425 141.94 316.385 142.45 ;
      RECT 325.005 136.43 325.965 136.94 ;
      RECT 326.265 136.43 327.225 136.94 ;
      RECT 323.745 136.43 324.705 136.94 ;
      RECT 322.485 136.43 323.445 136.94 ;
      RECT 321.225 136.43 322.185 136.94 ;
      RECT 324.375 141.94 325.335 142.45 ;
      RECT 323.115 141.94 324.075 142.45 ;
      RECT 321.855 141.94 322.815 142.45 ;
      RECT 325.635 141.94 326.595 142.45 ;
      RECT 326.895 141.94 327.855 142.45 ;
      RECT 327.525 136.43 328.485 136.94 ;
      RECT 328.785 136.43 329.745 136.94 ;
      RECT 329.195 136.94 329.365 137 ;
      RECT 332.565 136.43 333.525 136.94 ;
      RECT 331.305 136.43 332.265 136.94 ;
      RECT 330.045 136.43 331.005 136.94 ;
      RECT 331.935 141.94 332.895 142.45 ;
      RECT 330.675 141.94 331.635 142.45 ;
      RECT 329.415 141.94 330.375 142.45 ;
      RECT 328.155 141.94 329.115 142.45 ;
      RECT 337.605 136.43 337.935 136.94 ;
      RECT 337.685 136.94 337.855 137 ;
      RECT 333.195 141.94 334.155 142.45 ;
      RECT 333.825 136.43 334.785 136.94 ;
      RECT 335.085 136.43 336.045 136.94 ;
      RECT 336.345 136.43 337.305 136.94 ;
      RECT 334.455 141.94 335.415 142.45 ;
      RECT 335.715 141.94 336.675 142.45 ;
      RECT 336.975 141.94 337.935 142.45 ;
      RECT 341.95 143.3 342.96 143.795 ;
      RECT 342.85 142.93 343.38 143.1 ;
      RECT 343.21 143.1 343.38 145.85 ;
      RECT 344.14 143.3 348.89 143.795 ;
      RECT 364.565 142.93 364.735 144.58 ;
      RECT 364.565 142.76 368.865 142.93 ;
      RECT 368.695 142.93 368.865 144.58 ;
      RECT 364.565 144.58 368.865 144.75 ;
      RECT 364.985 143.27 365.515 143.44 ;
      RECT 364.985 143.44 365.155 144.135 ;
      RECT 365.705 143.24 368.455 143.41 ;
      RECT 379.515 136.14 379.845 136.73 ;
      RECT 397.475 137.855 397.645 144.645 ;
      RECT 402.035 137.855 402.205 144.645 ;
      RECT 399.755 137.855 399.925 144.645 ;
      RECT 406.595 137.855 406.765 144.645 ;
      RECT 404.315 137.855 404.485 144.645 ;
      RECT 409.325 137.855 409.495 144.645 ;
      RECT 411.605 137.855 411.775 144.645 ;
      RECT 418.445 137.855 418.615 144.645 ;
      RECT 413.885 137.855 414.055 144.645 ;
      RECT 416.165 137.855 416.335 144.645 ;
      RECT 421.645 139.65 422.995 139.83 ;
      RECT 424.75 138.345 424.92 139.355 ;
      RECT 423.66 141.155 423.99 141.805 ;
      RECT 425.28 141.155 425.61 141.805 ;
      RECT 422.85 141.155 423.18 141.805 ;
      RECT 422.04 141.155 422.37 141.805 ;
      RECT 424.47 141.155 424.8 141.805 ;
      RECT 423.115 136.72 423.285 139.43 ;
      RECT 421.31 180.755 430.39 180.925 ;
      RECT 421.31 140.415 441.73 140.585 ;
      RECT 421.31 140.585 421.48 180.755 ;
      RECT 441.56 140.585 441.73 199.94 ;
      RECT 430.22 180.925 430.39 199.94 ;
      RECT 430.22 199.94 441.73 200.115 ;
      RECT 421.355 136.72 421.525 139.43 ;
      RECT 422.235 136.72 422.405 139.43 ;
      RECT 424.805 137.925 425.475 138.095 ;
      RECT 428.005 139.415 433.185 139.585 ;
      RECT 433.005 137.945 433.185 138.355 ;
      RECT 428.005 138.355 433.185 138.525 ;
      RECT 426.955 139.995 433.185 140.175 ;
      RECT 426.955 137.765 433.185 137.945 ;
      RECT 433.005 139.585 433.185 139.995 ;
      RECT 433.005 138.525 433.185 139.415 ;
      RECT 426.955 137.945 427.135 139.995 ;
      RECT 428.005 138.885 432.755 139.055 ;
      RECT 425.53 138.345 425.7 139.355 ;
      RECT 426.9 141.155 427.23 141.805 ;
      RECT 426.09 141.155 426.42 141.805 ;
      RECT 430.14 141.155 430.47 141.805 ;
      RECT 430.95 141.155 431.28 141.805 ;
      RECT 429.33 141.155 429.66 141.805 ;
      RECT 428.52 141.155 428.85 141.805 ;
      RECT 427.71 141.155 428.04 141.805 ;
      RECT 427.325 138.635 427.83 139.305 ;
      RECT 431.76 141.155 432.09 141.805 ;
      RECT 432.57 141.155 432.9 141.805 ;
      RECT 434.19 141.155 434.52 141.805 ;
      RECT 433.38 141.155 433.71 141.805 ;
      RECT 435 141.155 435.33 141.805 ;
      RECT 435.81 141.155 436.14 141.805 ;
      RECT 436.62 141.155 436.95 141.805 ;
      RECT 440.67 141.155 441 141.805 ;
      RECT 439.86 141.155 440.19 141.805 ;
      RECT 439.05 141.155 439.38 141.805 ;
      RECT 438.24 141.155 438.57 141.805 ;
      RECT 437.43 141.155 437.76 141.805 ;
      RECT 447.215 139.155 447.385 139.175 ;
      RECT 447.165 139.085 447.495 139.155 ;
      RECT 447.165 138.645 447.495 138.715 ;
      RECT 447.165 138.715 460.845 139.085 ;
      RECT 460.515 139.085 460.845 139.155 ;
      RECT 460.515 138.645 460.845 138.715 ;
      RECT 447.215 137.745 447.385 137.765 ;
      RECT 447.165 138.205 447.495 138.275 ;
      RECT 447.165 137.765 447.495 137.835 ;
      RECT 447.165 137.835 460.845 138.205 ;
      RECT 460.515 138.205 460.845 138.275 ;
      RECT 460.515 137.765 460.845 137.835 ;
      RECT 447.665 139.255 460.35 139.425 ;
      RECT 447.665 138.375 448.715 138.545 ;
      RECT 447.665 137.495 460.35 137.665 ;
      RECT 447.755 139.99 449.145 140.16 ;
      RECT 447.755 136.76 449.145 136.93 ;
      RECT 447.215 141 447.385 144.62 ;
      RECT 447.765 140.575 460.045 141.145 ;
      RECT 447.765 135.775 460.045 136.345 ;
      RECT 447.765 141.355 460.045 141.925 ;
      RECT 447.765 142.135 460.045 142.705 ;
      RECT 447.765 142.915 460.045 143.485 ;
      RECT 448.945 138.375 449.275 138.545 ;
      RECT 431.25 135.19 432.35 135.36 ;
      RECT 437.08 128.035 437.41 128.725 ;
      RECT 440.16 128.035 440.49 128.725 ;
      RECT 439.39 128.035 439.72 128.725 ;
      RECT 440.93 128.035 441.26 128.725 ;
      RECT 441.7 128.035 442.03 128.725 ;
      RECT 437.85 128.035 438.18 128.725 ;
      RECT 439.39 135.19 440.49 135.36 ;
      RECT 440.93 135.19 442.03 135.36 ;
      RECT 437.08 134.945 438.18 135.4 ;
      RECT 447.215 132.3 447.385 135.92 ;
      RECT 447.765 131.875 460.045 132.445 ;
      RECT 447.765 130.965 460.045 131.535 ;
      RECT 447.765 134.995 460.045 135.565 ;
      RECT 447.765 134.215 460.045 134.785 ;
      RECT 447.765 133.435 460.045 134.005 ;
      RECT 447.765 132.655 460.045 133.225 ;
      RECT 447.765 128.625 460.045 129.195 ;
      RECT 447.765 129.405 460.045 129.975 ;
      RECT 447.765 130.185 460.045 130.755 ;
      RECT 460.595 132.3 460.765 135.92 ;
      RECT 10.16 136.14 10.49 136.73 ;
      RECT 21.14 142.93 21.31 144.58 ;
      RECT 21.14 142.76 25.44 142.93 ;
      RECT 21.14 144.58 25.44 144.75 ;
      RECT 25.27 142.93 25.44 144.58 ;
      RECT 24.49 143.27 25.02 143.44 ;
      RECT 24.85 143.44 25.02 144.135 ;
      RECT 21.55 143.24 24.3 143.41 ;
      RECT 41.115 143.3 45.865 143.795 ;
      RECT 47.045 143.3 48.055 143.795 ;
      RECT 46.625 142.93 47.155 143.1 ;
      RECT 46.625 143.1 46.795 145.85 ;
      RECT 54.59 141.94 55.55 142.45 ;
      RECT 53.33 141.94 54.29 142.45 ;
      RECT 52.07 141.94 53.03 142.45 ;
      RECT 52.07 136.43 52.4 136.94 ;
      RECT 52.15 136.94 52.32 137 ;
      RECT 53.96 136.43 54.92 136.94 ;
      RECT 52.7 136.43 53.66 136.94 ;
      RECT 55.22 136.43 56.18 136.94 ;
      RECT 56.48 136.43 57.44 136.94 ;
      RECT 57.74 136.43 58.7 136.94 ;
      RECT 59 136.43 59.96 136.94 ;
      RECT 60.26 136.43 61.22 136.94 ;
      RECT 60.64 136.94 60.81 137 ;
      RECT 55.85 141.94 56.81 142.45 ;
      RECT 57.11 141.94 58.07 142.45 ;
      RECT 58.37 141.94 59.33 142.45 ;
      RECT 59.63 141.94 60.59 142.45 ;
      RECT 64.04 136.43 65 136.94 ;
      RECT 62.78 136.43 63.74 136.94 ;
      RECT 61.52 136.43 62.48 136.94 ;
      RECT 65.3 136.43 66.26 136.94 ;
      RECT 64.67 141.94 65.63 142.45 ;
      RECT 65.93 141.94 66.89 142.45 ;
      RECT 63.41 141.94 64.37 142.45 ;
      RECT 62.15 141.94 63.11 142.45 ;
      RECT 60.89 141.94 61.85 142.45 ;
      RECT 66.56 136.43 67.52 136.94 ;
      RECT 67.82 136.43 68.78 136.94 ;
      RECT 69.08 136.43 69.41 136.94 ;
      RECT 69.16 136.94 69.33 137 ;
      RECT 69.84 136.43 70.17 136.94 ;
      RECT 69.92 136.94 70.09 137 ;
      RECT 71.73 136.43 72.69 136.94 ;
      RECT 70.47 136.43 71.43 136.94 ;
      RECT 71.1 141.94 72.06 142.45 ;
      RECT 69.84 141.94 70.8 142.45 ;
      RECT 67.19 141.94 68.15 142.45 ;
      RECT 68.45 141.94 69.41 142.45 ;
      RECT 74.25 136.43 75.21 136.94 ;
      RECT 75.51 136.43 76.47 136.94 ;
      RECT 76.77 136.43 77.73 136.94 ;
      RECT 72.99 136.43 73.95 136.94 ;
      RECT 73.62 141.94 74.58 142.45 ;
      RECT 72.36 141.94 73.32 142.45 ;
      RECT 74.88 141.94 75.84 142.45 ;
      RECT 76.14 141.94 77.1 142.45 ;
      RECT 77.4 141.94 78.36 142.45 ;
      RECT 78.03 136.43 78.99 136.94 ;
      RECT 78.41 136.94 78.58 137 ;
      RECT 81.81 136.43 82.77 136.94 ;
      RECT 80.55 136.43 81.51 136.94 ;
      RECT 79.29 136.43 80.25 136.94 ;
      RECT 83.07 136.43 84.03 136.94 ;
      RECT 82.44 141.94 83.4 142.45 ;
      RECT 81.18 141.94 82.14 142.45 ;
      RECT 79.92 141.94 80.88 142.45 ;
      RECT 78.66 141.94 79.62 142.45 ;
      RECT 85.59 136.43 86.55 136.94 ;
      RECT 86.85 136.43 87.18 136.94 ;
      RECT 86.93 136.94 87.1 137 ;
      RECT 83.7 141.94 84.66 142.45 ;
      RECT 84.96 141.94 85.92 142.45 ;
      RECT 86.22 141.94 87.18 142.45 ;
      RECT 84.33 136.43 85.29 136.94 ;
      RECT 302.825 141.94 303.785 142.45 ;
      RECT 303.455 136.43 304.415 136.94 ;
      RECT 302.825 136.43 303.155 136.94 ;
      RECT 302.905 136.94 303.075 137 ;
      RECT 307.235 136.43 308.195 136.94 ;
      RECT 308.495 136.43 309.455 136.94 ;
      RECT 305.975 136.43 306.935 136.94 ;
      RECT 304.715 136.43 305.675 136.94 ;
      RECT 306.605 141.94 307.565 142.45 ;
      RECT 305.345 141.94 306.305 142.45 ;
      RECT 304.085 141.94 305.045 142.45 ;
      RECT 307.865 141.94 308.825 142.45 ;
      RECT 309.125 141.94 310.085 142.45 ;
      RECT 309.755 136.43 310.715 136.94 ;
      RECT 311.015 136.43 311.975 136.94 ;
      RECT 311.425 136.94 311.595 137 ;
      RECT 314.795 136.43 315.755 136.94 ;
      RECT 313.535 136.43 314.495 136.94 ;
      RECT 312.275 136.43 313.235 136.94 ;
      RECT 314.165 141.94 315.125 142.45 ;
      RECT 312.905 141.94 313.865 142.45 ;
      RECT 311.645 141.94 312.605 142.45 ;
      RECT 310.385 141.94 311.345 142.45 ;
      RECT 320.595 136.43 320.925 136.94 ;
      RECT 320.675 136.94 320.845 137 ;
      RECT 319.835 136.43 320.165 136.94 ;
      RECT 319.915 136.94 320.085 137 ;
      RECT 316.055 136.43 317.015 136.94 ;
      RECT 317.315 136.43 318.275 136.94 ;
      RECT 318.575 136.43 319.535 136.94 ;
      RECT 304.085 135.54 305.045 136.05 ;
      RECT 314.795 130.03 315.755 130.54 ;
      RECT 313.535 130.03 314.495 130.54 ;
      RECT 312.275 130.03 313.235 130.54 ;
      RECT 311.015 130.03 311.975 130.54 ;
      RECT 311.425 130.54 311.595 130.6 ;
      RECT 309.755 130.03 310.715 130.54 ;
      RECT 310.385 135.54 311.345 136.05 ;
      RECT 314.165 135.54 315.125 136.05 ;
      RECT 312.905 135.54 313.865 136.05 ;
      RECT 311.645 135.54 312.605 136.05 ;
      RECT 320.595 130.03 320.925 130.54 ;
      RECT 320.675 130.54 320.845 130.6 ;
      RECT 319.835 130.03 320.165 130.54 ;
      RECT 319.915 130.54 320.085 130.6 ;
      RECT 316.055 130.03 317.015 130.54 ;
      RECT 317.315 130.03 318.275 130.54 ;
      RECT 318.575 130.03 319.535 130.54 ;
      RECT 315.425 135.54 316.385 136.05 ;
      RECT 316.685 135.54 317.645 136.05 ;
      RECT 317.945 135.54 318.905 136.05 ;
      RECT 319.205 135.54 320.165 136.05 ;
      RECT 320.595 135.54 321.555 136.05 ;
      RECT 326.265 130.03 327.225 130.54 ;
      RECT 323.745 130.03 324.705 130.54 ;
      RECT 322.485 130.03 323.445 130.54 ;
      RECT 321.225 130.03 322.185 130.54 ;
      RECT 325.005 130.03 325.965 130.54 ;
      RECT 324.375 135.54 325.335 136.05 ;
      RECT 325.635 135.54 326.595 136.05 ;
      RECT 326.895 135.54 327.855 136.05 ;
      RECT 323.115 135.54 324.075 136.05 ;
      RECT 321.855 135.54 322.815 136.05 ;
      RECT 327.525 130.03 328.485 130.54 ;
      RECT 328.785 130.03 329.745 130.54 ;
      RECT 329.195 130.54 329.365 130.6 ;
      RECT 332.565 130.03 333.525 130.54 ;
      RECT 331.305 130.03 332.265 130.54 ;
      RECT 330.045 130.03 331.005 130.54 ;
      RECT 331.935 135.54 332.895 136.05 ;
      RECT 330.675 135.54 331.635 136.05 ;
      RECT 329.415 135.54 330.375 136.05 ;
      RECT 328.155 135.54 329.115 136.05 ;
      RECT 333.195 135.54 334.155 136.05 ;
      RECT 333.825 130.03 334.785 130.54 ;
      RECT 335.085 130.03 336.045 130.54 ;
      RECT 336.345 130.03 337.305 130.54 ;
      RECT 334.455 135.54 335.415 136.05 ;
      RECT 335.715 135.54 336.675 136.05 ;
      RECT 336.975 135.54 337.935 136.05 ;
      RECT 337.605 130.03 337.935 130.54 ;
      RECT 337.685 130.54 337.855 130.6 ;
      RECT 341.43 129.45 356.68 129.62 ;
      RECT 356.51 129.62 356.68 131.49 ;
      RECT 356.51 131.66 356.68 142.95 ;
      RECT 341.43 129.62 341.6 131.49 ;
      RECT 341.43 131.49 356.68 131.66 ;
      RECT 341.43 147.335 344.935 147.505 ;
      RECT 341.43 131.66 341.6 147.335 ;
      RECT 349.62 142.95 356.68 143.12 ;
      RECT 341.43 150.925 344.66 151.095 ;
      RECT 341.43 147.505 341.6 150.925 ;
      RECT 346.14 148.365 349.79 148.535 ;
      RECT 349.62 143.12 349.79 148.365 ;
      RECT 341.43 152.855 341.6 158.215 ;
      RECT 341.43 152.685 344.66 152.855 ;
      RECT 341.43 151.095 341.6 152.685 ;
      RECT 346.14 152.335 349.79 152.505 ;
      RECT 349.62 148.535 349.79 152.335 ;
      RECT 349.62 154.815 349.79 158.215 ;
      RECT 346.14 154.645 349.79 154.815 ;
      RECT 349.62 152.505 349.79 154.645 ;
      RECT 341.43 158.215 349.79 158.59 ;
      RECT 352.87 130.03 355.585 130.2 ;
      RECT 352.87 130.91 355.585 131.08 ;
      RECT 356.085 130.57 356.255 130.91 ;
      RECT 355.625 130.4 356.255 130.57 ;
      RECT 356.085 130.24 356.255 130.4 ;
      RECT 363.105 128.155 363.275 132.905 ;
      RECT 362.225 128.155 362.395 132.905 ;
      RECT 362.45 133.415 363.12 133.585 ;
      RECT 362.49 133.405 363.06 133.415 ;
      RECT 365.745 128.135 365.915 132.905 ;
      RECT 363.985 128.135 364.155 132.905 ;
      RECT 364.865 128.155 365.035 132.905 ;
      RECT 366.625 128.155 366.795 132.905 ;
      RECT 370.145 128.155 370.315 132.905 ;
      RECT 369.265 128.135 369.435 132.905 ;
      RECT 367.505 128.135 367.675 132.905 ;
      RECT 368.385 128.155 368.555 132.905 ;
      RECT 400.135 129.815 401.825 129.985 ;
      RECT 397.855 129.815 399.545 129.985 ;
      RECT 402.035 130.205 402.205 137.215 ;
      RECT 397.475 130.205 397.645 137.215 ;
      RECT 399.755 130.205 399.925 137.215 ;
      RECT 404.695 129.815 406.385 129.985 ;
      RECT 402.415 129.815 404.105 129.985 ;
      RECT 406.595 130.205 406.765 137.215 ;
      RECT 404.315 130.205 404.485 137.215 ;
      RECT 411.985 129.815 413.675 129.985 ;
      RECT 409.705 129.815 411.395 129.985 ;
      RECT 409.325 130.205 409.495 137.215 ;
      RECT 411.605 130.205 411.775 137.215 ;
      RECT 414.265 129.815 415.955 129.985 ;
      RECT 416.545 129.815 418.235 129.985 ;
      RECT 413.885 130.205 414.055 137.215 ;
      RECT 418.445 130.205 418.615 137.215 ;
      RECT 416.165 130.205 416.335 137.215 ;
      RECT 422.735 129.99 423.065 130.58 ;
      RECT 422.035 129.99 422.365 130.58 ;
      RECT 424.835 133.915 425.165 134.875 ;
      RECT 424.135 133.915 424.465 134.875 ;
      RECT 423.435 133.915 423.765 134.875 ;
      RECT 421.415 134.355 421.585 134.365 ;
      RECT 421.415 134.875 421.585 134.885 ;
      RECT 421.335 134.365 421.665 134.875 ;
      RECT 430.48 128.035 430.81 128.725 ;
      RECT 429.71 128.035 430.04 128.725 ;
      RECT 429.71 135.19 430.81 135.36 ;
      RECT 426.235 133.91 426.565 134.875 ;
      RECT 425.555 133.915 425.865 134.365 ;
      RECT 425.535 134.365 425.865 134.875 ;
      RECT 431.25 128.035 431.58 128.725 ;
      RECT 432.02 128.035 432.35 128.725 ;
      RECT 433.56 128.035 433.89 128.725 ;
      RECT 434.33 128.035 434.66 128.725 ;
      RECT 433.56 134.945 434.66 135.4 ;
      RECT 447.765 120.705 460.045 121.275 ;
      RECT 448.945 124.865 449.275 125.035 ;
      RECT 457.335 124.865 460.045 125.035 ;
      RECT 447.765 127.845 460.045 128.415 ;
      RECT 460.595 127.49 460.765 131.11 ;
      RECT 19.69 128.155 19.86 132.905 ;
      RECT 20.57 128.135 20.74 132.905 ;
      RECT 22.33 128.135 22.5 132.905 ;
      RECT 24.09 128.135 24.26 132.905 ;
      RECT 24.97 128.155 25.14 132.905 ;
      RECT 23.21 128.155 23.38 132.905 ;
      RECT 21.45 128.155 21.62 132.905 ;
      RECT 26.73 128.155 26.9 132.905 ;
      RECT 27.61 128.155 27.78 132.905 ;
      RECT 26.885 133.415 27.555 133.585 ;
      RECT 26.945 133.405 27.515 133.415 ;
      RECT 25.85 128.135 26.02 132.905 ;
      RECT 33.325 129.62 33.495 131.49 ;
      RECT 33.325 129.45 48.575 129.62 ;
      RECT 33.325 131.66 33.495 142.95 ;
      RECT 48.405 129.62 48.575 131.49 ;
      RECT 33.325 131.49 48.575 131.66 ;
      RECT 45.07 147.335 48.575 147.505 ;
      RECT 48.405 131.66 48.575 147.335 ;
      RECT 33.325 142.95 40.385 143.12 ;
      RECT 45.345 150.925 48.575 151.095 ;
      RECT 48.405 147.505 48.575 150.925 ;
      RECT 40.215 148.365 43.865 148.535 ;
      RECT 40.215 143.12 40.385 148.365 ;
      RECT 48.405 152.855 48.575 158.215 ;
      RECT 45.345 152.685 48.575 152.855 ;
      RECT 48.405 151.095 48.575 152.685 ;
      RECT 40.215 152.335 43.865 152.505 ;
      RECT 40.215 148.535 40.385 152.335 ;
      RECT 40.215 154.815 40.385 158.215 ;
      RECT 40.215 154.645 43.865 154.815 ;
      RECT 40.215 152.505 40.385 154.645 ;
      RECT 40.215 158.215 48.575 158.59 ;
      RECT 34.42 130.03 37.135 130.2 ;
      RECT 34.42 130.91 37.135 131.08 ;
      RECT 33.75 130.57 33.92 130.91 ;
      RECT 33.75 130.4 34.38 130.57 ;
      RECT 33.75 130.24 33.92 130.4 ;
      RECT 52.07 130.03 52.4 130.54 ;
      RECT 52.15 130.54 52.32 130.6 ;
      RECT 53.96 130.03 54.92 130.54 ;
      RECT 52.7 130.03 53.66 130.54 ;
      RECT 54.59 135.54 55.55 136.05 ;
      RECT 53.33 135.54 54.29 136.05 ;
      RECT 52.07 135.54 53.03 136.05 ;
      RECT 55.22 130.03 56.18 130.54 ;
      RECT 56.48 130.03 57.44 130.54 ;
      RECT 57.74 130.03 58.7 130.54 ;
      RECT 59 130.03 59.96 130.54 ;
      RECT 60.26 130.03 61.22 130.54 ;
      RECT 60.64 130.54 60.81 130.6 ;
      RECT 55.85 135.54 56.81 136.05 ;
      RECT 57.11 135.54 58.07 136.05 ;
      RECT 58.37 135.54 59.33 136.05 ;
      RECT 59.63 135.54 60.59 136.05 ;
      RECT 64.04 130.03 65 130.54 ;
      RECT 62.78 130.03 63.74 130.54 ;
      RECT 61.52 130.03 62.48 130.54 ;
      RECT 65.3 130.03 66.26 130.54 ;
      RECT 64.67 135.54 65.63 136.05 ;
      RECT 65.93 135.54 66.89 136.05 ;
      RECT 63.41 135.54 64.37 136.05 ;
      RECT 62.15 135.54 63.11 136.05 ;
      RECT 60.89 135.54 61.85 136.05 ;
      RECT 71.73 130.03 72.69 130.54 ;
      RECT 70.47 130.03 71.43 130.54 ;
      RECT 66.56 130.03 67.52 130.54 ;
      RECT 67.82 130.03 68.78 130.54 ;
      RECT 69.08 130.03 69.41 130.54 ;
      RECT 69.16 130.54 69.33 130.6 ;
      RECT 69.84 130.03 70.17 130.54 ;
      RECT 69.92 130.54 70.09 130.6 ;
      RECT 71.1 135.54 72.06 136.05 ;
      RECT 69.84 135.54 70.8 136.05 ;
      RECT 67.19 135.54 68.15 136.05 ;
      RECT 68.45 135.54 69.41 136.05 ;
      RECT 72.99 130.03 73.95 130.54 ;
      RECT 74.25 130.03 75.21 130.54 ;
      RECT 75.51 130.03 76.47 130.54 ;
      RECT 76.77 130.03 77.73 130.54 ;
      RECT 73.62 135.54 74.58 136.05 ;
      RECT 74.88 135.54 75.84 136.05 ;
      RECT 76.14 135.54 77.1 136.05 ;
      RECT 77.4 135.54 78.36 136.05 ;
      RECT 72.36 135.54 73.32 136.05 ;
      RECT 80.55 130.03 81.51 130.54 ;
      RECT 79.29 130.03 80.25 130.54 ;
      RECT 78.03 130.03 78.99 130.54 ;
      RECT 78.41 130.54 78.58 130.6 ;
      RECT 83.07 130.03 84.03 130.54 ;
      RECT 81.81 130.03 82.77 130.54 ;
      RECT 82.44 135.54 83.4 136.05 ;
      RECT 81.18 135.54 82.14 136.05 ;
      RECT 79.92 135.54 80.88 136.05 ;
      RECT 78.66 135.54 79.62 136.05 ;
      RECT 84.33 130.03 85.29 130.54 ;
      RECT 85.59 130.03 86.55 130.54 ;
      RECT 86.85 130.03 87.18 130.54 ;
      RECT 86.93 130.54 87.1 130.6 ;
      RECT 83.7 135.54 84.66 136.05 ;
      RECT 84.96 135.54 85.92 136.05 ;
      RECT 86.22 135.54 87.18 136.05 ;
      RECT 51.495 129.45 87.79 129.62 ;
      RECT 51.495 129.62 51.665 142.385 ;
      RECT 87.62 129.62 87.79 142.385 ;
      RECT 51.525 129.415 87.73 129.45 ;
      RECT 303.455 130.03 304.415 130.54 ;
      RECT 302.825 130.03 303.155 130.54 ;
      RECT 302.905 130.54 303.075 130.6 ;
      RECT 302.825 135.54 303.785 136.05 ;
      RECT 302.215 129.45 338.51 129.62 ;
      RECT 338.34 129.62 338.51 142.385 ;
      RECT 302.215 129.62 302.385 142.385 ;
      RECT 302.275 129.415 338.48 129.45 ;
      RECT 305.975 130.03 306.935 130.54 ;
      RECT 304.715 130.03 305.675 130.54 ;
      RECT 307.235 130.03 308.195 130.54 ;
      RECT 308.495 130.03 309.455 130.54 ;
      RECT 306.605 135.54 307.565 136.05 ;
      RECT 307.865 135.54 308.825 136.05 ;
      RECT 309.125 135.54 310.085 136.05 ;
      RECT 305.345 135.54 306.305 136.05 ;
      RECT 364.45 125.695 369.2 125.865 ;
      RECT 364.45 127.255 369.2 127.425 ;
      RECT 364.45 126.475 369.2 126.645 ;
      RECT 364.53 126.645 369.12 126.65 ;
      RECT 369.42 125.92 369.59 127.2 ;
      RECT 386.27 125.48 386.6 126.13 ;
      RECT 387.53 125.48 387.86 126.13 ;
      RECT 386.9 125.48 387.23 126.13 ;
      RECT 388.79 125.48 389.12 126.13 ;
      RECT 388.16 125.48 388.49 126.13 ;
      RECT 389.42 125.48 389.75 126.13 ;
      RECT 390.05 125.48 390.38 126.13 ;
      RECT 386.27 126.51 386.6 127.16 ;
      RECT 387.53 126.51 387.86 127.16 ;
      RECT 386.9 126.51 387.23 127.16 ;
      RECT 388.79 126.51 389.12 127.16 ;
      RECT 388.16 126.51 388.49 127.16 ;
      RECT 389.42 126.51 389.75 127.16 ;
      RECT 390.05 126.51 390.38 127.16 ;
      RECT 390.68 125.48 391.01 126.13 ;
      RECT 391.94 125.48 392.27 126.13 ;
      RECT 390.68 126.51 391.01 127.16 ;
      RECT 391.31 126.51 391.64 127.16 ;
      RECT 391.94 126.51 392.27 127.16 ;
      RECT 392.57 126.51 392.9 127.16 ;
      RECT 391.31 125.48 391.64 126.13 ;
      RECT 392.65 125.54 392.82 125.62 ;
      RECT 392.57 125.62 392.9 126.13 ;
      RECT 393.2 125.48 393.53 126.13 ;
      RECT 393.2 126.51 393.53 127.16 ;
      RECT 394.46 125.48 394.79 126.13 ;
      RECT 393.83 126.51 394.16 127.16 ;
      RECT 394.46 126.51 394.79 127.16 ;
      RECT 393.83 125.48 394.16 126.13 ;
      RECT 397.855 122.165 399.545 122.335 ;
      RECT 400.135 122.165 401.825 122.335 ;
      RECT 402.05 121.025 402.72 121.195 ;
      RECT 400.87 121.025 401.54 121.195 ;
      RECT 399.69 121.025 400.36 121.195 ;
      RECT 396.635 145.115 397.305 145.285 ;
      RECT 396.695 122.165 397.42 122.335 ;
      RECT 396.695 129.815 397.42 129.985 ;
      RECT 396.695 137.465 397.42 137.635 ;
      RECT 396.695 122.335 396.865 129.815 ;
      RECT 396.695 129.985 396.865 137.465 ;
      RECT 396.695 137.635 396.865 145.115 ;
      RECT 402.035 122.555 402.205 129.565 ;
      RECT 397.475 122.555 397.645 129.565 ;
      RECT 399.755 122.555 399.925 129.565 ;
      RECT 402.415 122.165 404.105 122.335 ;
      RECT 404.695 122.165 406.385 122.335 ;
      RECT 405.59 121.025 406.26 121.195 ;
      RECT 404.41 121.025 405.08 121.195 ;
      RECT 403.23 121.025 403.9 121.195 ;
      RECT 406.82 122.165 407.545 122.335 ;
      RECT 406.82 129.815 407.545 129.985 ;
      RECT 406.82 137.465 407.545 137.635 ;
      RECT 406.82 145.115 407.545 145.285 ;
      RECT 407.375 122.335 407.545 129.815 ;
      RECT 407.375 129.985 407.545 137.465 ;
      RECT 407.375 137.635 407.545 145.115 ;
      RECT 406.595 122.555 406.765 129.565 ;
      RECT 404.315 122.555 404.485 129.565 ;
      RECT 409.705 122.165 411.395 122.335 ;
      RECT 411.985 122.165 413.675 122.335 ;
      RECT 408.545 122.165 409.27 122.335 ;
      RECT 408.545 129.815 409.27 129.985 ;
      RECT 408.545 137.465 409.27 137.635 ;
      RECT 408.545 145.115 409.27 145.285 ;
      RECT 408.545 122.335 408.715 129.815 ;
      RECT 408.545 129.985 408.715 137.465 ;
      RECT 408.545 137.635 408.715 145.115 ;
      RECT 409.83 121.025 410.5 121.195 ;
      RECT 411.01 121.025 411.68 121.195 ;
      RECT 412.19 121.025 412.86 121.195 ;
      RECT 413.37 121.025 414.04 121.195 ;
      RECT 409.325 122.555 409.495 129.565 ;
      RECT 411.605 122.555 411.775 129.465 ;
      RECT 414.265 122.165 415.955 122.335 ;
      RECT 416.545 122.165 418.235 122.335 ;
      RECT 418.67 122.165 419.395 122.335 ;
      RECT 418.67 129.815 419.395 129.985 ;
      RECT 418.67 137.465 419.395 137.635 ;
      RECT 418.67 145.115 419.395 145.285 ;
      RECT 419.225 122.335 419.395 129.815 ;
      RECT 419.225 129.985 419.395 137.465 ;
      RECT 419.225 137.635 419.395 145.115 ;
      RECT 414.55 121.025 415.22 121.195 ;
      RECT 415.73 121.025 416.4 121.195 ;
      RECT 413.885 122.555 414.055 129.565 ;
      RECT 418.445 122.555 418.615 129.565 ;
      RECT 416.165 122.555 416.335 129.565 ;
      RECT 430.48 120.88 430.81 121.57 ;
      RECT 429.71 120.88 430.04 121.57 ;
      RECT 431.25 120.88 431.58 121.57 ;
      RECT 432.02 120.88 432.35 121.57 ;
      RECT 433.56 120.88 433.89 121.57 ;
      RECT 434.225 120.88 434.755 121.05 ;
      RECT 434.33 121.05 434.66 121.57 ;
      RECT 436.985 120.88 437.515 121.05 ;
      RECT 437.08 121.05 437.41 121.57 ;
      RECT 440.16 120.88 440.49 121.57 ;
      RECT 439.39 120.88 439.72 121.57 ;
      RECT 440.93 120.88 441.26 121.57 ;
      RECT 441.7 120.88 442.03 121.57 ;
      RECT 437.85 120.88 438.18 121.57 ;
      RECT 447.215 125.645 447.385 125.665 ;
      RECT 447.165 125.575 447.495 125.645 ;
      RECT 447.165 125.135 447.495 125.205 ;
      RECT 447.165 125.205 460.845 125.575 ;
      RECT 460.515 125.575 460.845 125.645 ;
      RECT 460.515 125.135 460.845 125.205 ;
      RECT 447.215 124.235 447.385 124.255 ;
      RECT 447.165 124.695 447.495 124.765 ;
      RECT 447.165 124.255 447.495 124.325 ;
      RECT 447.165 124.325 460.845 124.695 ;
      RECT 460.515 124.695 460.845 124.765 ;
      RECT 460.515 124.255 460.845 124.325 ;
      RECT 447.665 125.745 460.35 125.915 ;
      RECT 447.665 124.865 448.715 125.035 ;
      RECT 447.665 123.985 460.35 124.155 ;
      RECT 447.755 123.25 449.145 123.42 ;
      RECT 447.755 126.48 449.145 126.65 ;
      RECT 447.215 127.49 447.385 131.11 ;
      RECT 447.765 122.265 460.045 122.835 ;
      RECT 447.765 127.065 460.045 127.635 ;
      RECT 447.765 121.485 460.045 122.055 ;
      RECT 303.815 124.61 303.985 124.67 ;
      RECT 303.815 124 303.985 124.44 ;
      RECT 302.215 115.305 309.585 116.07 ;
      RECT 302.215 124.44 303.985 124.61 ;
      RECT 302.215 122.38 303.525 122.55 ;
      RECT 302.215 122.55 302.385 124.44 ;
      RECT 302.215 116.07 302.385 122.38 ;
      RECT 305.535 113.55 315.165 113.72 ;
      RECT 304.555 116.77 304.725 126.62 ;
      RECT 308.835 116.77 309.005 126.62 ;
      RECT 302.855 123.66 303.985 123.83 ;
      RECT 303.815 117.65 303.985 123.66 ;
      RECT 304.78 116.43 308.78 116.6 ;
      RECT 304.78 126.98 308.78 127.15 ;
      RECT 304.895 116.6 308.665 126.98 ;
      RECT 313.245 116.43 317.245 116.6 ;
      RECT 313.245 126.98 317.245 127.15 ;
      RECT 313.36 116.6 317.13 126.98 ;
      RECT 312.34 124.02 313.19 126.81 ;
      RECT 312.3 119.145 313.19 124.02 ;
      RECT 312.34 116.9 313.19 119.145 ;
      RECT 312.34 116.79 312.51 116.9 ;
      RECT 318.675 116.43 322.675 116.6 ;
      RECT 318.675 126.98 322.675 127.15 ;
      RECT 318.79 116.6 322.56 126.98 ;
      RECT 317.3 116.9 318.62 126.81 ;
      RECT 322.955 116.43 326.955 116.6 ;
      RECT 322.955 126.98 326.955 127.15 ;
      RECT 323.07 116.6 326.84 126.98 ;
      RECT 322.73 116.96 322.9 126.81 ;
      RECT 328.255 116.43 332.385 116.6 ;
      RECT 328.255 126.98 332.385 127.15 ;
      RECT 328.5 116.6 332.27 126.98 ;
      RECT 327.01 116.9 328.33 126.81 ;
      RECT 332.44 119.145 333.33 124.02 ;
      RECT 332.44 124.02 333.29 126.81 ;
      RECT 332.44 116.9 333.29 119.145 ;
      RECT 333.12 116.79 333.29 116.9 ;
      RECT 337.045 116.43 341.045 116.6 ;
      RECT 337.045 126.98 341.045 127.15 ;
      RECT 337.16 116.6 340.93 126.98 ;
      RECT 336.1 118.025 336.99 122.9 ;
      RECT 336.14 122.9 336.99 126.81 ;
      RECT 336.14 116.9 336.99 118.025 ;
      RECT 336.14 116.79 336.31 116.9 ;
      RECT 342.475 116.43 346.475 116.6 ;
      RECT 342.475 126.98 346.475 127.15 ;
      RECT 342.72 116.6 346.36 126.98 ;
      RECT 341.1 116.9 342.42 126.81 ;
      RECT 346.755 116.43 350.755 116.6 ;
      RECT 346.755 126.98 350.755 127.15 ;
      RECT 347 116.6 350.64 126.98 ;
      RECT 346.53 116.96 346.7 126.81 ;
      RECT 352.185 116.43 356.185 116.6 ;
      RECT 352.185 126.98 356.185 127.15 ;
      RECT 352.3 116.6 356.07 126.98 ;
      RECT 350.81 116.9 352.13 126.81 ;
      RECT 356.24 118.025 357.13 122.9 ;
      RECT 356.24 122.9 357.09 126.81 ;
      RECT 356.24 116.9 357.09 118.025 ;
      RECT 356.92 116.79 357.09 116.9 ;
      RECT 362.225 117.835 362.395 124.625 ;
      RECT 365.095 113.725 365.265 116.765 ;
      RECT 363.035 113.005 363.985 113.175 ;
      RECT 363.035 116.655 363.985 116.825 ;
      RECT 363.815 113.175 363.985 116.655 ;
      RECT 363.035 113.175 363.205 116.655 ;
      RECT 366.375 113.725 366.545 116.435 ;
      RECT 364.455 113.205 364.625 116.655 ;
      RECT 364.155 116.655 364.925 116.825 ;
      RECT 365.735 113.205 365.905 116.655 ;
      RECT 367.02 113.205 367.19 116.655 ;
      RECT 365.435 116.655 366.205 116.825 ;
      RECT 366.715 116.655 367.485 116.825 ;
      RECT 368.295 113.205 368.465 116.655 ;
      RECT 367.995 116.655 368.765 116.825 ;
      RECT 364.235 113.175 364.845 113.205 ;
      RECT 365.515 113.175 366.125 113.205 ;
      RECT 366.8 113.175 367.41 113.205 ;
      RECT 368.075 113.175 368.685 113.205 ;
      RECT 364.155 113.005 368.765 113.175 ;
      RECT 363.345 112.465 364.115 112.635 ;
      RECT 370.475 118.465 370.675 123.88 ;
      RECT 370.505 123.88 370.675 124.625 ;
      RECT 370.505 117.835 370.675 118.465 ;
      RECT 367.655 113.725 367.825 116.765 ;
      RECT 368.935 113.725 369.105 116.435 ;
      RECT 369.715 113.725 369.885 116.435 ;
      RECT 393.83 119.155 394.16 119.805 ;
      RECT 391.31 119.155 391.64 119.805 ;
      RECT 392.57 119.155 392.9 119.805 ;
      RECT 430.48 113.725 430.81 114.415 ;
      RECT 429.71 113.725 430.04 114.415 ;
      RECT 431.25 113.725 431.58 114.415 ;
      RECT 431.935 114.065 432.435 114.415 ;
      RECT 431.935 113.61 433.205 114.065 ;
      RECT 433.56 113.725 433.89 114.415 ;
      RECT 434.33 113.725 434.66 114.415 ;
      RECT 437.08 113.725 437.41 114.415 ;
      RECT 440.16 113.725 440.49 114.415 ;
      RECT 439.305 114.065 439.805 114.415 ;
      RECT 438.535 113.61 439.805 114.065 ;
      RECT 440.93 113.725 441.26 114.415 ;
      RECT 441.7 113.725 442.03 114.415 ;
      RECT 437.85 113.725 438.18 114.415 ;
      RECT 447.665 112.235 460.35 112.405 ;
      RECT 447.755 112.97 449.145 113.14 ;
      RECT 447.215 113.98 447.385 117.6 ;
      RECT 447.215 118.79 447.385 122.41 ;
      RECT 447.765 117.455 460.045 118.025 ;
      RECT 447.765 118.365 460.045 118.935 ;
      RECT 447.765 113.555 460.045 114.125 ;
      RECT 447.765 119.145 460.045 119.715 ;
      RECT 447.765 114.335 460.045 114.905 ;
      RECT 447.765 115.115 460.045 115.685 ;
      RECT 447.765 115.895 460.045 116.465 ;
      RECT 447.765 116.675 460.045 117.245 ;
      RECT 447.765 119.925 460.045 120.495 ;
      RECT 460.595 113.98 460.765 117.6 ;
      RECT 460.595 118.79 460.765 122.41 ;
      RECT 20.805 125.695 25.555 125.865 ;
      RECT 20.805 127.255 25.555 127.425 ;
      RECT 20.805 126.475 25.555 126.645 ;
      RECT 20.885 126.645 25.475 126.65 ;
      RECT 20.415 125.92 20.585 127.2 ;
      RECT 86.37 121.1 87.26 121.27 ;
      RECT 302.745 121.1 303.635 121.27 ;
      RECT 32.915 122.9 33.765 126.81 ;
      RECT 32.915 116.9 33.765 118.025 ;
      RECT 32.915 116.79 33.085 116.9 ;
      RECT 39.25 116.43 43.25 116.6 ;
      RECT 39.25 126.98 43.25 127.15 ;
      RECT 39.365 116.6 43.005 126.98 ;
      RECT 37.875 116.9 39.195 126.81 ;
      RECT 43.53 116.43 47.53 116.6 ;
      RECT 43.53 126.98 47.53 127.15 ;
      RECT 43.645 116.6 47.285 126.98 ;
      RECT 47.585 116.9 48.905 126.81 ;
      RECT 43.305 116.96 43.475 126.81 ;
      RECT 48.96 116.43 52.96 116.6 ;
      RECT 48.96 126.98 52.96 127.15 ;
      RECT 49.075 116.6 52.845 126.98 ;
      RECT 53.015 118.025 53.905 122.9 ;
      RECT 53.015 122.9 53.865 126.81 ;
      RECT 53.015 116.9 53.865 118.025 ;
      RECT 53.695 116.79 53.865 116.9 ;
      RECT 57.62 116.43 61.75 116.6 ;
      RECT 57.62 126.98 61.75 127.15 ;
      RECT 57.735 116.6 61.505 126.98 ;
      RECT 56.675 119.145 57.565 124.02 ;
      RECT 56.715 124.02 57.565 126.81 ;
      RECT 56.715 116.9 57.565 119.145 ;
      RECT 56.715 116.79 56.885 116.9 ;
      RECT 63.05 116.43 67.05 116.6 ;
      RECT 63.05 126.98 67.05 127.15 ;
      RECT 63.165 116.6 66.935 126.98 ;
      RECT 61.675 116.9 62.995 126.81 ;
      RECT 67.33 116.43 71.33 116.6 ;
      RECT 67.33 126.98 71.33 127.15 ;
      RECT 67.445 116.6 71.215 126.98 ;
      RECT 71.385 116.9 72.705 126.81 ;
      RECT 67.105 116.96 67.275 126.81 ;
      RECT 74.84 113.55 84.47 113.72 ;
      RECT 72.76 116.43 76.76 116.6 ;
      RECT 72.76 126.98 76.76 127.15 ;
      RECT 72.875 116.6 76.645 126.98 ;
      RECT 76.815 124.02 77.665 126.81 ;
      RECT 76.815 119.145 77.705 124.02 ;
      RECT 76.815 116.9 77.665 119.145 ;
      RECT 77.495 116.79 77.665 116.9 ;
      RECT 80.42 116.07 80.59 126.79 ;
      RECT 73.13 113.96 87.79 114.13 ;
      RECT 79.72 114.715 87.79 115.305 ;
      RECT 80.42 114.13 87.79 114.715 ;
      RECT 86.02 124.61 86.19 124.67 ;
      RECT 86.02 124 86.19 124.44 ;
      RECT 80.42 115.305 87.79 116.07 ;
      RECT 86.02 124.44 87.79 124.61 ;
      RECT 86.48 122.38 87.79 122.55 ;
      RECT 87.62 122.55 87.79 124.44 ;
      RECT 87.62 116.07 87.79 122.38 ;
      RECT 87.62 124.61 87.79 126.48 ;
      RECT 81 116.77 81.17 126.62 ;
      RECT 81.225 116.43 85.225 116.6 ;
      RECT 81.225 126.98 85.225 127.15 ;
      RECT 81.34 116.6 85.11 126.98 ;
      RECT 87.13 117.43 87.3 117.79 ;
      RECT 86.48 117.26 87.3 117.43 ;
      RECT 86.48 119.82 87.37 119.99 ;
      RECT 86.48 116.48 87.15 116.65 ;
      RECT 86.38 113.55 87.455 113.72 ;
      RECT 86.37 118.54 87.26 118.71 ;
      RECT 85.72 116.325 86.25 116.495 ;
      RECT 86.02 116.495 86.19 117.09 ;
      RECT 85.28 116.77 85.45 126.62 ;
      RECT 86.02 123.66 87.15 123.83 ;
      RECT 86.02 117.65 86.19 123.66 ;
      RECT 95.705 113.195 96.375 113.525 ;
      RECT 95.775 113.165 96.305 113.195 ;
      RECT 102.165 113.195 102.835 113.525 ;
      RECT 104.725 113.195 105.395 113.525 ;
      RECT 111.185 113.195 111.855 113.525 ;
      RECT 113.745 113.195 114.415 113.525 ;
      RECT 122.765 113.195 123.435 113.525 ;
      RECT 120.205 113.195 120.875 113.525 ;
      RECT 129.225 113.195 129.895 113.525 ;
      RECT 131.785 113.195 132.455 113.525 ;
      RECT 138.245 113.195 138.915 113.525 ;
      RECT 140.805 113.195 141.475 113.525 ;
      RECT 147.265 113.195 147.935 113.525 ;
      RECT 149.825 113.195 150.495 113.525 ;
      RECT 156.285 113.195 156.955 113.525 ;
      RECT 158.845 113.195 159.515 113.525 ;
      RECT 167.865 113.195 168.535 113.525 ;
      RECT 165.305 113.195 165.975 113.525 ;
      RECT 174.325 113.195 174.995 113.525 ;
      RECT 176.885 113.195 177.555 113.525 ;
      RECT 183.345 113.195 184.015 113.525 ;
      RECT 183.415 113.165 183.945 113.195 ;
      RECT 205.99 113.195 206.66 113.525 ;
      RECT 206.06 113.165 206.59 113.195 ;
      RECT 215.01 113.195 215.68 113.525 ;
      RECT 212.45 113.195 213.12 113.525 ;
      RECT 221.47 113.195 222.14 113.525 ;
      RECT 224.03 113.195 224.7 113.525 ;
      RECT 233.05 113.195 233.72 113.525 ;
      RECT 230.49 113.195 231.16 113.525 ;
      RECT 239.51 113.195 240.18 113.525 ;
      RECT 242.07 113.195 242.74 113.525 ;
      RECT 251.09 113.195 251.76 113.525 ;
      RECT 248.53 113.195 249.2 113.525 ;
      RECT 260.11 113.195 260.78 113.525 ;
      RECT 257.55 113.195 258.22 113.525 ;
      RECT 266.57 113.195 267.24 113.525 ;
      RECT 269.13 113.195 269.8 113.525 ;
      RECT 278.15 113.195 278.82 113.525 ;
      RECT 275.59 113.195 276.26 113.525 ;
      RECT 284.61 113.195 285.28 113.525 ;
      RECT 287.17 113.195 287.84 113.525 ;
      RECT 293.63 113.195 294.3 113.525 ;
      RECT 293.7 113.165 294.23 113.195 ;
      RECT 302.635 119.82 303.525 119.99 ;
      RECT 302.705 117.43 302.875 117.79 ;
      RECT 302.705 117.26 303.525 117.43 ;
      RECT 302.855 116.48 303.525 116.65 ;
      RECT 302.55 113.55 303.625 113.72 ;
      RECT 302.745 118.54 303.635 118.71 ;
      RECT 303.755 116.325 304.285 116.495 ;
      RECT 303.815 116.495 303.985 117.09 ;
      RECT 309.415 116.07 309.585 126.79 ;
      RECT 302.215 113.96 316.875 114.13 ;
      RECT 302.215 124.61 302.385 126.48 ;
      RECT 302.215 114.715 310.285 115.305 ;
      RECT 302.215 114.13 309.585 114.715 ;
      RECT 388.79 107.035 389.12 107.685 ;
      RECT 388.16 107.035 388.49 107.685 ;
      RECT 389.42 107.035 389.75 107.685 ;
      RECT 390.05 107.035 390.38 107.685 ;
      RECT 390.68 106.005 391.01 106.655 ;
      RECT 391.31 106.005 391.64 106.655 ;
      RECT 391.94 106.005 392.27 106.655 ;
      RECT 393.2 106.005 393.53 106.655 ;
      RECT 392.57 106.005 392.9 106.655 ;
      RECT 393.83 106.005 394.16 106.655 ;
      RECT 394.46 106.005 394.79 106.655 ;
      RECT 390.68 107.035 391.01 107.685 ;
      RECT 391.94 107.035 392.27 107.685 ;
      RECT 393.2 107.035 393.53 107.685 ;
      RECT 394.46 107.035 394.79 107.685 ;
      RECT 399.1 108.295 402.83 108.465 ;
      RECT 399.69 110.375 406.26 110.545 ;
      RECT 400.53 110.545 400.7 120.655 ;
      RECT 405.25 110.545 405.42 120.655 ;
      RECT 402.89 110.545 403.06 120.655 ;
      RECT 398.165 109.115 398.755 109.435 ;
      RECT 398.165 109.435 398.59 110.595 ;
      RECT 407.66 108.295 411.39 108.465 ;
      RECT 403.38 108.295 407.11 108.465 ;
      RECT 407.195 109.115 408.895 109.435 ;
      RECT 408.305 109.435 408.73 111.295 ;
      RECT 407.36 109.435 407.785 111.295 ;
      RECT 413.26 108.295 416.99 108.465 ;
      RECT 409.83 110.375 416.4 110.545 ;
      RECT 410.67 110.545 410.84 120.655 ;
      RECT 413.03 110.545 413.2 120.655 ;
      RECT 415.39 110.545 415.56 120.655 ;
      RECT 417.56 108.295 419.25 108.465 ;
      RECT 417.5 109.435 417.925 111.38 ;
      RECT 417.335 109.115 417.925 109.435 ;
      RECT 419.84 108.295 421.53 108.465 ;
      RECT 422.12 108.295 423.81 108.465 ;
      RECT 421.415 112.135 421.585 112.145 ;
      RECT 421.415 112.655 421.585 112.665 ;
      RECT 421.335 112.145 421.665 112.655 ;
      RECT 420.75 111.555 427.15 111.735 ;
      RECT 420.75 111.735 420.93 135.285 ;
      RECT 420.75 135.285 427.15 135.465 ;
      RECT 423.695 136.04 423.875 140.06 ;
      RECT 420.75 140.06 423.875 140.24 ;
      RECT 426.97 111.735 427.15 135.285 ;
      RECT 420.75 135.465 423.875 136.04 ;
      RECT 420.75 136.04 420.93 140.06 ;
      RECT 424.835 112.145 425.165 113.105 ;
      RECT 424.135 112.145 424.465 113.105 ;
      RECT 423.435 112.145 423.765 113.105 ;
      RECT 422.735 112.145 423.065 113.105 ;
      RECT 422.035 112.145 422.365 113.105 ;
      RECT 430.48 106.57 430.81 107.26 ;
      RECT 429.71 106.57 430.04 107.26 ;
      RECT 426.235 112.145 426.565 113.105 ;
      RECT 425.535 112.145 425.865 113.105 ;
      RECT 431.25 107.09 431.58 107.26 ;
      RECT 431.25 106.57 431.58 106.74 ;
      RECT 431.335 106.74 431.505 107.09 ;
      RECT 431.935 106.57 433.205 107.26 ;
      RECT 433.56 106.57 433.89 107.26 ;
      RECT 434.33 106.57 434.66 107.26 ;
      RECT 437.08 106.57 437.41 107.26 ;
      RECT 440.16 107.09 440.49 107.26 ;
      RECT 440.16 106.57 440.49 106.74 ;
      RECT 440.235 106.74 440.405 107.09 ;
      RECT 438.535 106.57 439.805 107.26 ;
      RECT 440.93 106.57 441.26 107.26 ;
      RECT 441.7 106.57 442.03 107.26 ;
      RECT 437.85 106.57 438.18 107.26 ;
      RECT 447.215 112.135 447.385 112.155 ;
      RECT 447.165 112.065 447.495 112.135 ;
      RECT 447.165 111.625 447.495 111.695 ;
      RECT 447.165 111.695 460.845 112.065 ;
      RECT 460.515 112.065 460.845 112.135 ;
      RECT 460.515 111.625 460.845 111.695 ;
      RECT 447.215 110.725 447.385 110.745 ;
      RECT 447.165 111.185 447.495 111.255 ;
      RECT 447.165 110.745 447.495 110.815 ;
      RECT 447.165 110.815 460.845 111.185 ;
      RECT 460.515 111.185 460.845 111.255 ;
      RECT 460.515 110.745 460.845 110.815 ;
      RECT 447.665 111.355 448.715 111.525 ;
      RECT 447.665 110.475 460.35 110.645 ;
      RECT 447.755 109.74 449.145 109.91 ;
      RECT 447.215 105.28 447.385 108.9 ;
      RECT 447.765 108.755 460.045 109.325 ;
      RECT 447.765 104.855 460.045 105.425 ;
      RECT 447.765 107.975 460.045 108.545 ;
      RECT 447.765 107.195 460.045 107.765 ;
      RECT 447.765 106.415 460.045 106.985 ;
      RECT 447.765 105.635 460.045 106.205 ;
      RECT 448.945 111.355 449.275 111.525 ;
      RECT 457.335 111.355 460.045 111.525 ;
      RECT 460.595 105.28 460.765 108.9 ;
      RECT 19.33 118.465 19.53 123.88 ;
      RECT 19.33 123.88 19.5 124.625 ;
      RECT 19.33 117.835 19.5 118.465 ;
      RECT 22.18 113.725 22.35 116.765 ;
      RECT 23.46 113.725 23.63 116.435 ;
      RECT 20.9 113.725 21.07 116.435 ;
      RECT 24.74 113.725 24.91 116.765 ;
      RECT 20.12 113.725 20.29 116.435 ;
      RECT 25.38 113.205 25.55 116.655 ;
      RECT 25.08 116.655 25.85 116.825 ;
      RECT 24.1 113.205 24.27 116.655 ;
      RECT 22.815 113.205 22.985 116.655 ;
      RECT 21.54 113.205 21.71 116.655 ;
      RECT 23.8 116.655 24.57 116.825 ;
      RECT 22.52 116.655 23.29 116.825 ;
      RECT 21.24 116.655 22.01 116.825 ;
      RECT 25.16 113.175 25.77 113.205 ;
      RECT 21.32 113.175 21.93 113.205 ;
      RECT 21.24 113.005 25.85 113.175 ;
      RECT 23.88 113.175 24.49 113.205 ;
      RECT 22.595 113.175 23.205 113.205 ;
      RECT 27.61 117.835 27.78 124.625 ;
      RECT 26.02 113.005 26.97 113.175 ;
      RECT 26.02 116.655 26.97 116.825 ;
      RECT 26.02 113.175 26.19 116.655 ;
      RECT 26.8 113.175 26.97 116.655 ;
      RECT 25.89 112.465 26.66 112.635 ;
      RECT 33.82 116.43 37.82 116.6 ;
      RECT 33.82 126.98 37.82 127.15 ;
      RECT 33.935 116.6 37.705 126.98 ;
      RECT 32.875 118.025 33.765 122.9 ;
      RECT 312.825 108.34 312.995 113.205 ;
      RECT 314.635 106.95 315.305 107.12 ;
      RECT 313.12 105.455 313.29 105.76 ;
      RECT 313.115 105.76 313.29 106.425 ;
      RECT 313.115 106.425 313.285 106.77 ;
      RECT 311.545 108.34 311.715 113.09 ;
      RECT 314.105 108.34 314.275 113.09 ;
      RECT 314.295 105.76 314.465 107.065 ;
      RECT 320.645 108.17 320.815 113.55 ;
      RECT 320.235 110.28 320.415 111.17 ;
      RECT 320.245 108 320.895 108.17 ;
      RECT 320.245 113.55 320.895 113.72 ;
      RECT 320.245 108.17 320.415 110.28 ;
      RECT 320.245 111.17 320.415 113.55 ;
      RECT 321.025 108.34 321.195 113.09 ;
      RECT 315.385 108.34 315.555 113.205 ;
      RECT 316.665 108.34 316.835 113.55 ;
      RECT 315.61 113.55 316.835 113.72 ;
      RECT 315.475 105.455 315.645 106.77 ;
      RECT 302.225 104.77 316.875 104.94 ;
      RECT 302.225 107.58 316.875 107.75 ;
      RECT 316.055 104.94 316.225 107.58 ;
      RECT 302.225 104.94 312.705 107.58 ;
      RECT 319.665 107.76 319.835 113.96 ;
      RECT 319.665 113.96 356.795 114.13 ;
      RECT 319.665 107.59 356.795 107.76 ;
      RECT 356.625 107.76 356.795 113.96 ;
      RECT 325.305 108.34 325.475 113.09 ;
      RECT 325.53 108 329.53 108.17 ;
      RECT 325.53 113.55 329.53 113.72 ;
      RECT 326.885 108.17 328.18 113.55 ;
      RECT 321.25 108 325.25 108.17 ;
      RECT 321.25 113.55 325.25 113.72 ;
      RECT 322.605 108.17 323.9 113.55 ;
      RECT 329.585 108.34 329.755 113.09 ;
      RECT 329.81 108 333.81 108.17 ;
      RECT 329.81 113.55 333.81 113.72 ;
      RECT 331.165 108.17 332.46 113.55 ;
      RECT 333.865 108.34 334.035 113.09 ;
      RECT 338.145 108.34 338.315 113.09 ;
      RECT 334.09 108 338.09 108.17 ;
      RECT 334.09 113.55 338.09 113.72 ;
      RECT 335.445 108.17 336.74 113.55 ;
      RECT 338.37 108 342.37 108.17 ;
      RECT 338.37 113.55 342.37 113.72 ;
      RECT 339.725 108.17 341.02 113.55 ;
      RECT 342.425 108.34 342.595 113.09 ;
      RECT 342.65 108 346.65 108.17 ;
      RECT 342.65 113.55 346.65 113.72 ;
      RECT 344.005 108.17 345.3 113.55 ;
      RECT 346.705 108.34 346.875 113.09 ;
      RECT 346.93 108 350.93 108.17 ;
      RECT 346.93 113.55 350.93 113.72 ;
      RECT 348.285 108.17 349.58 113.55 ;
      RECT 355.265 108.34 355.435 113.09 ;
      RECT 350.985 108.34 351.155 113.09 ;
      RECT 355.665 108.17 355.835 113.55 ;
      RECT 355.585 108 356.215 108.17 ;
      RECT 355.585 113.55 356.215 113.72 ;
      RECT 356.045 110.28 356.225 111.17 ;
      RECT 356.045 111.17 356.215 113.55 ;
      RECT 356.045 108.17 356.215 110.28 ;
      RECT 351.21 108 355.21 108.17 ;
      RECT 351.21 113.55 355.21 113.72 ;
      RECT 352.565 108.17 353.86 113.55 ;
      RECT 364.16 104.51 369.13 104.68 ;
      RECT 362.615 106.46 363.285 106.63 ;
      RECT 362.105 105.82 362.275 106.49 ;
      RECT 362.615 105.675 363.285 105.85 ;
      RECT 364.16 106.07 369.13 106.24 ;
      RECT 364.16 105.29 369.12 105.46 ;
      RECT 363.77 107.46 363.94 107.575 ;
      RECT 363.77 106.68 363.94 107.19 ;
      RECT 363.77 106.41 369.59 106.68 ;
      RECT 363.77 104.85 369.59 105.12 ;
      RECT 363.77 104.675 363.94 104.85 ;
      RECT 363.77 107.19 369.59 107.46 ;
      RECT 369.42 105.9 369.59 106.41 ;
      RECT 369.42 105.12 369.59 105.63 ;
      RECT 363.77 105.9 363.94 106.41 ;
      RECT 363.77 105.63 369.59 105.9 ;
      RECT 363.77 105.12 363.94 105.63 ;
      RECT 369.42 104.73 369.59 104.85 ;
      RECT 369.42 107.46 369.59 107.57 ;
      RECT 369.42 106.68 369.59 107.19 ;
      RECT 364.16 107.63 369.13 107.8 ;
      RECT 365.56 111.685 365.735 111.915 ;
      RECT 365.565 108.815 366.675 108.985 ;
      RECT 365.56 112.465 366.675 112.635 ;
      RECT 365.56 111.915 365.73 112.465 ;
      RECT 365.565 108.985 365.735 111.685 ;
      RECT 366.845 108.815 367.955 108.985 ;
      RECT 366.845 112.465 367.955 112.635 ;
      RECT 366.845 108.985 367.015 112.465 ;
      RECT 362.565 109.995 363.175 110.165 ;
      RECT 363.005 110.165 363.175 111.915 ;
      RECT 363.005 109.205 363.175 109.995 ;
      RECT 364.285 108.815 365.395 108.985 ;
      RECT 364.285 112.465 365.39 112.635 ;
      RECT 364.285 108.985 364.455 112.465 ;
      RECT 362.225 112.465 362.95 112.635 ;
      RECT 362.225 108.815 362.395 112.465 ;
      RECT 364.16 106.85 369.12 107.02 ;
      RECT 363.345 108.815 364.115 108.985 ;
      RECT 363.425 108.985 364.035 109.015 ;
      RECT 369.63 108.815 370.3 108.985 ;
      RECT 369.815 108.985 369.985 113.005 ;
      RECT 369.375 113.175 369.545 116.655 ;
      RECT 369.16 116.655 369.83 116.825 ;
      RECT 369.815 108.535 369.985 108.815 ;
      RECT 369.16 113.005 369.985 113.175 ;
      RECT 368.125 108.815 369.235 108.985 ;
      RECT 368.125 112.465 369.235 112.635 ;
      RECT 368.545 108.985 369.155 109.015 ;
      RECT 368.125 108.985 368.295 112.465 ;
      RECT 369.405 109.205 369.575 111.915 ;
      RECT 370.185 109.205 370.355 111.915 ;
      RECT 386.27 106.005 386.6 106.655 ;
      RECT 387.53 106.005 387.86 106.655 ;
      RECT 386.9 106.005 387.23 106.655 ;
      RECT 388.79 106.005 389.12 106.655 ;
      RECT 388.16 106.005 388.49 106.655 ;
      RECT 389.42 106.005 389.75 106.655 ;
      RECT 390.05 106.005 390.38 106.655 ;
      RECT 386.27 107.035 386.6 107.685 ;
      RECT 387.53 107.035 387.86 107.685 ;
      RECT 386.9 107.035 387.23 107.685 ;
      RECT 91.795 111.435 92.645 166.535 ;
      RECT 122.32 106.36 122.85 106.53 ;
      RECT 122.32 106.53 122.49 106.75 ;
      RECT 122.32 105.4 122.49 106.36 ;
      RECT 122.42 105.04 138.91 105.21 ;
      RECT 122.95 105.21 127.7 105.28 ;
      RECT 128.555 105.21 133.305 105.28 ;
      RECT 134.16 105.21 138.91 105.28 ;
      RECT 122.95 106.87 127.77 106.92 ;
      RECT 128.19 106.87 133.375 106.92 ;
      RECT 133.795 106.87 138.91 106.92 ;
      RECT 121.91 104.53 139.43 104.7 ;
      RECT 122.95 106.92 138.91 107.065 ;
      RECT 122.95 107.065 139.43 107.09 ;
      RECT 139.26 104.7 139.43 107.065 ;
      RECT 121.91 104.7 122.08 107.09 ;
      RECT 121.91 107.09 139.43 107.62 ;
      RECT 122.95 105.99 127.7 106.16 ;
      RECT 127.815 106.36 128.345 106.53 ;
      RECT 127.895 106.53 128.065 106.75 ;
      RECT 127.895 105.4 128.065 106.36 ;
      RECT 128.555 105.99 133.305 106.16 ;
      RECT 133.42 106.36 133.95 106.53 ;
      RECT 133.5 106.53 133.67 106.75 ;
      RECT 133.5 105.4 133.67 106.36 ;
      RECT 134.16 105.99 138.91 106.16 ;
      RECT 141.13 107.45 153.065 107.62 ;
      RECT 141.13 104.53 153.065 104.7 ;
      RECT 152.895 104.7 153.065 107.45 ;
      RECT 141.13 104.7 141.3 107.45 ;
      RECT 146.61 106.36 147.14 106.53 ;
      RECT 146.88 106.53 147.05 106.75 ;
      RECT 146.88 105.4 147.05 106.36 ;
      RECT 141.65 105.035 152.555 105.205 ;
      RECT 147.255 105.205 152.005 105.28 ;
      RECT 141.65 105.205 146.4 105.28 ;
      RECT 141.65 106.94 152.555 107.11 ;
      RECT 147.255 106.87 152.005 106.94 ;
      RECT 141.65 106.87 146.4 106.94 ;
      RECT 147.255 105.99 152.005 106.16 ;
      RECT 141.65 105.99 146.4 106.16 ;
      RECT 152.125 106.36 152.655 106.53 ;
      RECT 152.485 106.53 152.655 106.725 ;
      RECT 152.485 105.375 152.655 106.36 ;
      RECT 148.625 112.085 149.155 112.255 ;
      RECT 148.635 112.255 149.145 112.33 ;
      RECT 148.635 112 149.145 112.085 ;
      RECT 159.335 112.085 159.865 112.255 ;
      RECT 159.345 112.255 159.855 112.33 ;
      RECT 159.345 112 159.855 112.085 ;
      RECT 168.6 106.195 171.465 106.365 ;
      RECT 168.6 104.635 171.465 104.805 ;
      RECT 168.6 105.415 171.465 105.585 ;
      RECT 175.995 105.9 176.545 106.07 ;
      RECT 175.995 106.07 176.465 106.545 ;
      RECT 175.995 105.87 176.465 105.9 ;
      RECT 202.1 110.585 298.21 111.435 ;
      RECT 202.1 166.535 298.21 167.385 ;
      RECT 202.1 111.435 202.95 166.535 ;
      RECT 297.36 111.435 298.21 166.535 ;
      RECT 213.46 105.9 214.01 106.07 ;
      RECT 213.54 106.07 214.01 106.545 ;
      RECT 213.54 105.87 214.01 105.9 ;
      RECT 218.54 106.195 221.405 106.365 ;
      RECT 218.54 104.635 221.405 104.805 ;
      RECT 218.54 105.415 221.405 105.585 ;
      RECT 230.14 112.085 230.67 112.255 ;
      RECT 230.15 112.255 230.66 112.33 ;
      RECT 230.15 112 230.66 112.085 ;
      RECT 237.35 106.36 237.88 106.53 ;
      RECT 237.35 106.53 237.52 106.725 ;
      RECT 237.35 105.375 237.52 106.36 ;
      RECT 237.45 105.035 248.355 105.205 ;
      RECT 238 105.205 242.75 105.28 ;
      RECT 243.605 105.205 248.355 105.28 ;
      RECT 237.45 106.94 248.355 107.11 ;
      RECT 238 106.87 242.75 106.94 ;
      RECT 243.605 106.87 248.355 106.94 ;
      RECT 238 105.99 242.75 106.16 ;
      RECT 236.94 104.7 237.11 107.45 ;
      RECT 236.94 107.45 248.875 107.62 ;
      RECT 236.94 104.53 248.875 104.7 ;
      RECT 248.705 104.7 248.875 107.45 ;
      RECT 242.865 106.36 243.395 106.53 ;
      RECT 242.955 106.53 243.125 106.75 ;
      RECT 242.955 105.4 243.125 106.36 ;
      RECT 240.85 112.085 241.38 112.255 ;
      RECT 240.86 112.255 241.37 112.33 ;
      RECT 240.86 112 241.37 112.085 ;
      RECT 243.605 105.99 248.355 106.16 ;
      RECT 251.095 105.04 267.585 105.21 ;
      RECT 251.095 105.21 255.845 105.28 ;
      RECT 256.7 105.21 261.45 105.28 ;
      RECT 262.305 105.21 267.055 105.28 ;
      RECT 251.095 106.87 256.21 106.92 ;
      RECT 256.63 106.87 261.815 106.92 ;
      RECT 262.235 106.87 267.055 106.92 ;
      RECT 250.575 104.53 268.095 104.7 ;
      RECT 251.095 106.92 267.055 107.065 ;
      RECT 250.575 107.065 267.055 107.09 ;
      RECT 250.575 104.7 250.745 107.065 ;
      RECT 267.925 104.7 268.095 107.09 ;
      RECT 250.575 107.09 268.095 107.62 ;
      RECT 251.095 105.99 255.845 106.16 ;
      RECT 256.055 106.36 256.585 106.53 ;
      RECT 256.335 106.53 256.505 106.75 ;
      RECT 256.335 105.4 256.505 106.36 ;
      RECT 256.7 105.99 261.45 106.16 ;
      RECT 261.66 106.36 262.19 106.53 ;
      RECT 261.94 106.53 262.11 106.75 ;
      RECT 261.94 105.4 262.11 106.36 ;
      RECT 262.305 105.99 267.055 106.16 ;
      RECT 267.155 106.36 267.685 106.53 ;
      RECT 267.515 106.53 267.685 106.75 ;
      RECT 267.515 105.4 267.685 106.36 ;
      RECT 302.615 104.35 303.625 104.52 ;
      RECT 302.255 108.34 302.425 113.205 ;
      RECT 303.035 108.34 303.205 113.09 ;
      RECT 305.145 108.34 305.315 113.205 ;
      RECT 304.365 113.55 305.09 113.72 ;
      RECT 304.365 108.34 304.535 113.55 ;
      RECT 307.705 108.34 307.875 113.205 ;
      RECT 303.815 108.34 303.985 113.205 ;
      RECT 305.535 104.36 315.165 104.53 ;
      RECT 306.425 108.34 306.595 113.09 ;
      RECT 308.985 108.34 309.155 113.09 ;
      RECT 310.265 108.34 310.435 113.205 ;
      RECT 20.02 113.005 20.845 113.175 ;
      RECT 19.65 109.205 19.82 111.915 ;
      RECT 20.875 104.51 25.845 104.68 ;
      RECT 20.875 106.07 25.845 106.24 ;
      RECT 20.885 105.29 25.845 105.46 ;
      RECT 26.065 104.675 26.235 104.85 ;
      RECT 20.415 105.9 20.585 106.41 ;
      RECT 20.415 107.46 20.585 107.57 ;
      RECT 20.415 106.68 20.585 107.19 ;
      RECT 20.415 106.41 26.235 106.68 ;
      RECT 20.415 105.12 20.585 105.63 ;
      RECT 20.415 104.85 26.235 105.12 ;
      RECT 20.415 104.73 20.585 104.85 ;
      RECT 26.065 105.9 26.235 106.41 ;
      RECT 20.415 105.63 26.235 105.9 ;
      RECT 26.065 105.12 26.235 105.63 ;
      RECT 26.065 107.46 26.235 107.575 ;
      RECT 20.415 107.19 26.235 107.46 ;
      RECT 26.065 106.68 26.235 107.19 ;
      RECT 20.875 107.63 25.845 107.8 ;
      RECT 24.27 111.685 24.445 111.915 ;
      RECT 23.33 108.815 24.44 108.985 ;
      RECT 23.33 112.465 24.445 112.635 ;
      RECT 24.275 111.915 24.445 112.465 ;
      RECT 24.27 108.985 24.44 111.685 ;
      RECT 22.05 108.815 23.16 108.985 ;
      RECT 22.05 112.465 23.16 112.635 ;
      RECT 22.99 108.985 23.16 112.465 ;
      RECT 24.61 108.815 25.72 108.985 ;
      RECT 24.615 112.465 25.72 112.635 ;
      RECT 25.55 108.985 25.72 112.465 ;
      RECT 20.77 108.815 21.88 108.985 ;
      RECT 20.77 112.465 21.88 112.635 ;
      RECT 20.85 108.985 21.46 109.015 ;
      RECT 21.71 108.985 21.88 112.465 ;
      RECT 20.43 109.205 20.6 111.915 ;
      RECT 20.885 106.85 25.845 107.02 ;
      RECT 26.72 106.46 27.39 106.63 ;
      RECT 27.73 105.82 27.9 106.49 ;
      RECT 26.72 105.675 27.39 105.85 ;
      RECT 26.83 109.995 27.44 110.165 ;
      RECT 26.83 110.165 27 111.915 ;
      RECT 26.83 109.205 27 109.995 ;
      RECT 27.055 112.465 27.78 112.635 ;
      RECT 27.61 108.815 27.78 112.465 ;
      RECT 25.89 108.815 26.66 108.985 ;
      RECT 25.97 108.985 26.58 109.015 ;
      RECT 34.57 108.34 34.74 113.09 ;
      RECT 34.17 108.17 34.34 113.55 ;
      RECT 33.78 110.28 33.96 111.17 ;
      RECT 33.79 108 34.42 108.17 ;
      RECT 33.79 113.55 34.42 113.72 ;
      RECT 33.79 108.17 33.96 110.28 ;
      RECT 33.79 111.17 33.96 113.55 ;
      RECT 34.795 108 38.795 108.17 ;
      RECT 34.795 113.55 38.795 113.72 ;
      RECT 36.145 108.17 37.44 113.55 ;
      RECT 33.21 107.76 33.38 113.96 ;
      RECT 33.21 107.59 70.34 107.76 ;
      RECT 33.21 113.96 70.34 114.13 ;
      RECT 70.17 107.76 70.34 113.96 ;
      RECT 38.85 108.34 39.02 113.09 ;
      RECT 39.075 108 43.075 108.17 ;
      RECT 39.075 113.55 43.075 113.72 ;
      RECT 40.425 108.17 41.72 113.55 ;
      RECT 47.41 108.34 47.58 113.09 ;
      RECT 43.13 108.34 43.3 113.09 ;
      RECT 43.355 108 47.355 108.17 ;
      RECT 43.355 113.55 47.355 113.72 ;
      RECT 44.705 108.17 46 113.55 ;
      RECT 47.635 108 51.635 108.17 ;
      RECT 47.635 113.55 51.635 113.72 ;
      RECT 48.985 108.17 50.28 113.55 ;
      RECT 51.69 108.34 51.86 113.09 ;
      RECT 51.915 108 55.915 108.17 ;
      RECT 51.915 113.55 55.915 113.72 ;
      RECT 53.265 108.17 54.56 113.55 ;
      RECT 55.97 108.34 56.14 113.09 ;
      RECT 60.25 108.34 60.42 113.09 ;
      RECT 56.195 108 60.195 108.17 ;
      RECT 56.195 113.55 60.195 113.72 ;
      RECT 57.545 108.17 58.84 113.55 ;
      RECT 60.475 108 64.475 108.17 ;
      RECT 60.475 113.55 64.475 113.72 ;
      RECT 61.825 108.17 63.12 113.55 ;
      RECT 64.53 108.34 64.7 113.09 ;
      RECT 64.755 108 68.755 108.17 ;
      RECT 64.755 113.55 68.755 113.72 ;
      RECT 66.105 108.17 67.4 113.55 ;
      RECT 69.19 108.17 69.36 113.55 ;
      RECT 69.59 110.28 69.77 111.17 ;
      RECT 69.11 108 69.76 108.17 ;
      RECT 69.11 113.55 69.76 113.72 ;
      RECT 69.59 108.17 69.76 110.28 ;
      RECT 69.59 111.17 69.76 113.55 ;
      RECT 68.81 108.34 68.98 113.09 ;
      RECT 77.01 108.34 77.18 113.205 ;
      RECT 74.7 106.95 75.37 107.12 ;
      RECT 74.84 104.36 84.47 104.53 ;
      RECT 74.45 108.34 74.62 113.205 ;
      RECT 73.17 108.34 73.34 113.55 ;
      RECT 73.17 113.55 74.395 113.72 ;
      RECT 74.36 105.455 74.53 106.77 ;
      RECT 76.715 105.455 76.885 105.76 ;
      RECT 76.715 105.76 76.89 106.425 ;
      RECT 76.72 106.425 76.89 106.77 ;
      RECT 75.73 108.34 75.9 113.09 ;
      RECT 75.54 105.76 75.71 107.065 ;
      RECT 73.13 104.77 87.78 104.94 ;
      RECT 73.13 107.58 87.78 107.75 ;
      RECT 73.78 104.94 73.95 107.58 ;
      RECT 77.3 104.94 87.78 107.58 ;
      RECT 79.57 108.34 79.74 113.205 ;
      RECT 82.13 108.34 82.3 113.205 ;
      RECT 83.41 108.34 83.58 113.09 ;
      RECT 80.85 108.34 81.02 113.09 ;
      RECT 78.29 108.34 78.46 113.09 ;
      RECT 84.915 113.55 85.64 113.72 ;
      RECT 85.47 108.34 85.64 113.55 ;
      RECT 84.69 108.34 84.86 113.205 ;
      RECT 86.38 104.35 87.39 104.52 ;
      RECT 87.58 108.34 87.75 113.205 ;
      RECT 86.02 108.34 86.19 113.205 ;
      RECT 86.8 108.34 86.97 113.09 ;
      RECT 91.795 110.585 187.905 111.435 ;
      RECT 91.795 166.535 187.905 167.385 ;
      RECT 187.055 111.435 187.905 166.535 ;
      RECT 319.665 98.56 319.835 104.76 ;
      RECT 319.665 98.39 356.795 98.56 ;
      RECT 319.665 104.76 356.795 104.93 ;
      RECT 356.625 98.56 356.795 104.76 ;
      RECT 325.305 99.14 325.475 103.89 ;
      RECT 321.25 98.8 325.25 98.97 ;
      RECT 321.25 104.35 325.25 104.52 ;
      RECT 322.605 98.97 323.9 104.35 ;
      RECT 325.53 98.8 329.53 98.97 ;
      RECT 325.53 104.35 329.53 104.52 ;
      RECT 326.885 98.97 328.18 104.35 ;
      RECT 329.585 99.14 329.755 103.89 ;
      RECT 329.81 98.8 333.81 98.97 ;
      RECT 329.81 104.35 333.81 104.52 ;
      RECT 331.165 98.97 332.46 104.35 ;
      RECT 338.145 99.14 338.315 103.89 ;
      RECT 333.865 99.14 334.035 103.89 ;
      RECT 334.09 98.8 338.09 98.97 ;
      RECT 334.09 104.35 338.09 104.52 ;
      RECT 335.445 98.97 336.74 104.35 ;
      RECT 338.37 98.8 342.37 98.97 ;
      RECT 338.37 104.35 342.37 104.52 ;
      RECT 339.725 98.97 341.02 104.35 ;
      RECT 342.425 99.14 342.595 103.89 ;
      RECT 342.65 98.8 346.65 98.97 ;
      RECT 342.65 104.35 346.65 104.52 ;
      RECT 344.005 98.97 345.3 104.35 ;
      RECT 346.705 99.14 346.875 103.89 ;
      RECT 346.93 98.8 350.93 98.97 ;
      RECT 346.93 104.35 350.93 104.52 ;
      RECT 348.285 98.97 349.58 104.35 ;
      RECT 355.265 99.14 355.435 103.89 ;
      RECT 350.985 99.14 351.155 103.89 ;
      RECT 351.21 98.8 355.21 98.97 ;
      RECT 351.21 104.35 355.21 104.52 ;
      RECT 352.565 98.97 353.86 104.35 ;
      RECT 355.665 98.97 355.835 104.35 ;
      RECT 355.585 98.8 356.215 98.97 ;
      RECT 355.585 104.35 356.215 104.52 ;
      RECT 356.045 101.08 356.225 101.97 ;
      RECT 356.045 101.97 356.215 104.35 ;
      RECT 356.045 98.97 356.215 101.08 ;
      RECT 362.225 103.265 362.95 103.435 ;
      RECT 362.225 99.615 362.95 99.785 ;
      RECT 362.225 99.785 362.395 103.265 ;
      RECT 362.565 100.795 363.175 100.965 ;
      RECT 363.005 100.965 363.175 102.715 ;
      RECT 363.005 100.005 363.175 100.795 ;
      RECT 364.285 103.265 365.39 103.435 ;
      RECT 364.285 99.615 365.395 99.785 ;
      RECT 364.285 99.785 364.455 103.265 ;
      RECT 365.56 102.715 365.73 103.375 ;
      RECT 365.56 102.485 365.735 102.715 ;
      RECT 365.565 99.615 366.675 99.785 ;
      RECT 365.565 99.785 365.735 102.485 ;
      RECT 366.845 103.265 367.955 103.435 ;
      RECT 366.845 99.615 367.955 99.785 ;
      RECT 366.845 99.785 367.015 103.265 ;
      RECT 363.345 99.615 364.115 99.785 ;
      RECT 363.425 99.785 364.035 99.815 ;
      RECT 365.905 103.265 366.675 103.435 ;
      RECT 363.345 103.265 364.115 103.435 ;
      RECT 369.405 99.615 370.355 99.785 ;
      RECT 369.405 103.265 370.355 103.435 ;
      RECT 369.405 99.785 369.575 103.265 ;
      RECT 370.185 99.785 370.355 103.265 ;
      RECT 368.125 99.615 369.235 99.785 ;
      RECT 368.125 103.265 369.235 103.435 ;
      RECT 368.545 99.785 369.155 99.815 ;
      RECT 368.125 99.785 368.295 103.265 ;
      RECT 400.46 97.43 401.47 97.6 ;
      RECT 401.64 97.43 404.57 97.61 ;
      RECT 404.74 97.43 405.75 97.6 ;
      RECT 405.92 97.43 408.85 97.61 ;
      RECT 409.02 97.43 410.03 97.6 ;
      RECT 414.62 97.43 415.63 97.6 ;
      RECT 417.9 97.43 418.91 97.6 ;
      RECT 415.8 97.43 417.73 97.61 ;
      RECT 419.08 97.43 420.01 97.61 ;
      RECT 420.18 97.43 421.19 97.6 ;
      RECT 422.46 97.43 423.47 97.6 ;
      RECT 421.36 97.43 422.29 97.61 ;
      RECT 430.48 99.415 430.81 100.105 ;
      RECT 429.71 99.415 430.04 100.105 ;
      RECT 431.25 99.415 431.58 100.105 ;
      RECT 431.935 99.895 433.205 100.145 ;
      RECT 431.935 99.415 432.435 99.895 ;
      RECT 433.56 99.415 433.89 100.105 ;
      RECT 434.33 99.415 434.66 100.105 ;
      RECT 437.08 99.415 437.41 100.105 ;
      RECT 440.16 99.415 440.49 100.105 ;
      RECT 438.535 99.895 439.805 100.145 ;
      RECT 439.305 99.415 439.805 99.895 ;
      RECT 440.93 99.415 441.26 100.105 ;
      RECT 441.7 99.415 442.03 100.105 ;
      RECT 437.85 99.415 438.18 100.105 ;
      RECT 447.215 98.625 447.385 98.645 ;
      RECT 447.165 98.555 447.495 98.625 ;
      RECT 447.165 98.115 447.495 98.185 ;
      RECT 447.165 98.185 460.845 98.555 ;
      RECT 460.515 98.555 460.845 98.625 ;
      RECT 460.515 98.115 460.845 98.185 ;
      RECT 447.215 97.215 447.385 97.235 ;
      RECT 447.165 97.675 447.495 97.745 ;
      RECT 447.165 97.235 447.495 97.305 ;
      RECT 447.165 97.305 460.845 97.675 ;
      RECT 460.515 97.675 460.845 97.745 ;
      RECT 460.515 97.235 460.845 97.305 ;
      RECT 447.665 98.725 460.35 98.895 ;
      RECT 447.665 97.845 448.715 98.015 ;
      RECT 447.665 96.965 460.35 97.135 ;
      RECT 447.755 99.46 449.145 99.63 ;
      RECT 447.215 100.47 447.385 104.09 ;
      RECT 447.765 100.045 460.045 100.615 ;
      RECT 447.765 103.945 460.045 104.515 ;
      RECT 447.765 100.825 460.045 101.395 ;
      RECT 447.765 101.605 460.045 102.175 ;
      RECT 447.765 102.385 460.045 102.955 ;
      RECT 447.765 103.165 460.045 103.735 ;
      RECT 448.945 97.845 449.275 98.015 ;
      RECT 457.335 97.845 460.045 98.015 ;
      RECT 460.595 100.47 460.765 104.09 ;
      RECT 19.705 108.815 20.375 108.985 ;
      RECT 20.02 108.985 20.19 113.005 ;
      RECT 20.46 113.175 20.63 116.655 ;
      RECT 20.175 116.655 20.845 116.825 ;
      RECT 20.02 108.535 20.19 108.815 ;
      RECT 25.89 103.265 26.66 103.435 ;
      RECT 34.57 99.14 34.74 103.89 ;
      RECT 34.17 98.97 34.34 104.35 ;
      RECT 33.78 101.08 33.96 101.97 ;
      RECT 33.79 104.35 34.42 104.52 ;
      RECT 33.79 98.8 34.42 98.97 ;
      RECT 33.79 101.97 33.96 104.35 ;
      RECT 33.79 98.97 33.96 101.08 ;
      RECT 34.795 98.8 38.795 98.97 ;
      RECT 34.795 104.35 38.795 104.52 ;
      RECT 36.145 98.97 37.44 104.35 ;
      RECT 33.21 98.56 33.38 104.76 ;
      RECT 33.21 98.39 70.34 98.56 ;
      RECT 33.21 104.76 70.34 104.93 ;
      RECT 70.17 98.56 70.34 104.76 ;
      RECT 38.85 99.14 39.02 103.89 ;
      RECT 39.075 98.8 43.075 98.97 ;
      RECT 39.075 104.35 43.075 104.52 ;
      RECT 40.425 98.97 41.72 104.35 ;
      RECT 47.41 99.14 47.58 103.89 ;
      RECT 43.13 99.14 43.3 103.89 ;
      RECT 43.355 98.8 47.355 98.97 ;
      RECT 43.355 104.35 47.355 104.52 ;
      RECT 44.705 98.97 46 104.35 ;
      RECT 47.635 98.8 51.635 98.97 ;
      RECT 47.635 104.35 51.635 104.52 ;
      RECT 48.985 98.97 50.28 104.35 ;
      RECT 51.69 99.14 51.86 103.89 ;
      RECT 51.915 98.8 55.915 98.97 ;
      RECT 51.915 104.35 55.915 104.52 ;
      RECT 53.265 98.97 54.56 104.35 ;
      RECT 60.25 99.14 60.42 103.89 ;
      RECT 55.97 99.14 56.14 103.89 ;
      RECT 56.195 98.8 60.195 98.97 ;
      RECT 56.195 104.35 60.195 104.52 ;
      RECT 57.545 98.97 58.84 104.35 ;
      RECT 60.475 98.8 64.475 98.97 ;
      RECT 60.475 104.35 64.475 104.52 ;
      RECT 61.825 98.97 63.12 104.35 ;
      RECT 64.53 99.14 64.7 103.89 ;
      RECT 64.755 98.8 68.755 98.97 ;
      RECT 64.755 104.35 68.755 104.52 ;
      RECT 66.105 98.97 67.4 104.35 ;
      RECT 69.19 98.97 69.36 104.35 ;
      RECT 69.59 101.08 69.77 101.97 ;
      RECT 69.11 104.35 69.76 104.52 ;
      RECT 69.11 98.8 69.76 98.97 ;
      RECT 69.59 101.97 69.76 104.35 ;
      RECT 69.59 98.97 69.76 101.08 ;
      RECT 68.81 99.14 68.98 103.89 ;
      RECT 74.445 103.89 74.615 104.005 ;
      RECT 74.445 100.235 74.62 103.89 ;
      RECT 74.45 99.14 74.62 100.235 ;
      RECT 77.01 99.14 77.18 104.005 ;
      RECT 73.17 99.14 73.34 104.36 ;
      RECT 73.17 104.36 74.395 104.53 ;
      RECT 75.73 99.14 75.9 103.89 ;
      RECT 82.13 99.14 82.3 104.005 ;
      RECT 79.57 99.14 79.74 104.005 ;
      RECT 78.29 99.14 78.46 103.89 ;
      RECT 80.85 99.14 81.02 103.89 ;
      RECT 83.41 99.14 83.58 103.89 ;
      RECT 84.69 99.14 84.86 104.005 ;
      RECT 84.915 104.36 85.64 104.53 ;
      RECT 85.47 99.14 85.64 104.36 ;
      RECT 87.58 99.14 87.75 103.89 ;
      RECT 86.02 99.14 86.19 103.89 ;
      RECT 86.8 99.14 86.97 103.89 ;
      RECT 168.6 99.085 171.49 99.255 ;
      RECT 168.6 99.865 171.49 100.035 ;
      RECT 168.6 101.975 171.49 102.145 ;
      RECT 168.6 100.415 171.52 100.585 ;
      RECT 168.6 102.525 171.465 102.695 ;
      RECT 168.6 104.085 171.465 104.255 ;
      RECT 168.6 101.195 171.525 101.365 ;
      RECT 166.82 97.825 173.07 98.675 ;
      RECT 166.82 106.775 173.07 107.625 ;
      RECT 166.82 98.675 167.67 106.775 ;
      RECT 172.22 98.675 173.07 106.775 ;
      RECT 168.6 103.305 171.465 103.475 ;
      RECT 176.05 102.785 176.38 102.955 ;
      RECT 176.05 102.445 176.38 102.615 ;
      RECT 176.13 102.615 176.3 102.785 ;
      RECT 176.13 102.425 176.3 102.445 ;
      RECT 171.735 99.215 172.04 106.14 ;
      RECT 213.625 102.785 213.955 102.955 ;
      RECT 213.625 102.445 213.955 102.615 ;
      RECT 213.705 102.615 213.875 102.785 ;
      RECT 213.705 102.425 213.875 102.445 ;
      RECT 217.965 99.215 218.27 106.14 ;
      RECT 218.515 99.085 221.405 99.255 ;
      RECT 218.515 99.865 221.405 100.035 ;
      RECT 218.515 101.975 221.405 102.145 ;
      RECT 218.485 100.415 221.405 100.585 ;
      RECT 218.54 102.525 221.405 102.695 ;
      RECT 218.54 104.085 221.405 104.255 ;
      RECT 218.48 101.195 221.405 101.365 ;
      RECT 216.935 97.825 223.185 98.675 ;
      RECT 216.935 106.775 223.185 107.625 ;
      RECT 216.935 98.675 217.785 106.775 ;
      RECT 222.335 98.675 223.185 106.775 ;
      RECT 218.54 103.305 221.405 103.475 ;
      RECT 302.255 99.14 302.425 103.89 ;
      RECT 303.035 99.14 303.205 103.89 ;
      RECT 304.365 104.36 305.09 104.53 ;
      RECT 304.365 99.14 304.535 104.36 ;
      RECT 305.145 99.14 305.315 104.005 ;
      RECT 303.815 99.14 303.985 103.89 ;
      RECT 307.705 99.14 307.875 104.005 ;
      RECT 308.985 99.14 309.155 103.89 ;
      RECT 306.425 99.14 306.595 103.89 ;
      RECT 312.825 99.14 312.995 104.005 ;
      RECT 310.265 99.14 310.435 104.005 ;
      RECT 311.545 99.14 311.715 103.89 ;
      RECT 314.105 99.14 314.275 103.89 ;
      RECT 320.645 98.97 320.815 104.35 ;
      RECT 320.235 101.08 320.415 101.97 ;
      RECT 320.245 104.35 320.895 104.52 ;
      RECT 320.245 98.8 320.895 98.97 ;
      RECT 320.245 101.97 320.415 104.35 ;
      RECT 320.245 98.97 320.415 101.08 ;
      RECT 321.025 99.14 321.195 103.89 ;
      RECT 315.39 103.89 315.56 104.005 ;
      RECT 315.385 100.235 315.56 103.89 ;
      RECT 315.385 99.14 315.555 100.235 ;
      RECT 316.665 99.14 316.835 104.36 ;
      RECT 315.61 104.36 316.835 104.53 ;
      RECT 53.015 94.495 53.865 95.62 ;
      RECT 53.015 85.71 53.865 89.62 ;
      RECT 86.02 88.69 87.15 88.86 ;
      RECT 86.02 88.86 86.19 94.87 ;
      RECT 86.48 95.87 87.15 96.04 ;
      RECT 86.495 96.04 87.025 96.09 ;
      RECT 86.48 95.09 87.425 95.26 ;
      RECT 87.255 94.73 87.425 95.09 ;
      RECT 86.48 92.53 87.37 92.7 ;
      RECT 86.37 91.25 87.26 91.42 ;
      RECT 86.37 93.81 87.26 93.98 ;
      RECT 85.705 95.92 86.235 96.09 ;
      RECT 86.02 96.09 86.19 96.1 ;
      RECT 86.02 95.43 86.19 95.92 ;
      RECT 102.56 89.715 103.115 89.885 ;
      RECT 102.56 89.885 102.73 89.98 ;
      RECT 102.56 89.65 102.73 89.715 ;
      RECT 286.89 89.715 287.445 89.885 ;
      RECT 287.275 89.885 287.445 89.98 ;
      RECT 287.275 89.65 287.445 89.715 ;
      RECT 302.58 95.09 303.525 95.26 ;
      RECT 302.58 94.73 302.75 95.09 ;
      RECT 302.635 92.53 303.525 92.7 ;
      RECT 302.855 88.69 303.985 88.86 ;
      RECT 303.815 88.86 303.985 94.87 ;
      RECT 302.855 95.87 303.525 96.04 ;
      RECT 302.98 96.04 303.51 96.09 ;
      RECT 302.745 93.81 303.635 93.98 ;
      RECT 302.745 91.25 303.635 91.42 ;
      RECT 303.77 95.92 304.3 96.09 ;
      RECT 303.815 96.09 303.985 96.1 ;
      RECT 303.815 95.43 303.985 95.92 ;
      RECT 336.14 95.62 336.31 95.73 ;
      RECT 336.1 89.62 336.99 94.495 ;
      RECT 336.14 94.495 336.99 95.62 ;
      RECT 336.14 85.71 336.99 89.62 ;
      RECT 341.1 85.71 342.42 95.62 ;
      RECT 346.53 85.71 346.7 95.56 ;
      RECT 350.81 85.71 352.13 95.62 ;
      RECT 356.92 95.62 357.09 95.73 ;
      RECT 356.24 94.495 357.09 95.62 ;
      RECT 356.24 89.62 357.13 94.495 ;
      RECT 356.24 85.71 357.09 89.62 ;
      RECT 365.095 95.485 365.265 98.855 ;
      RECT 363.035 95.425 363.985 95.595 ;
      RECT 363.035 99.075 363.985 99.245 ;
      RECT 363.815 95.595 363.985 99.075 ;
      RECT 363.035 95.595 363.205 99.075 ;
      RECT 366.375 96.145 366.545 98.855 ;
      RECT 366.715 95.425 367.485 95.595 ;
      RECT 364.455 95.595 364.625 99.045 ;
      RECT 364.155 95.425 364.925 95.595 ;
      RECT 365.435 95.425 366.205 95.595 ;
      RECT 368.295 95.595 368.465 99.045 ;
      RECT 367.995 95.425 368.765 95.595 ;
      RECT 367.02 95.595 367.19 99.045 ;
      RECT 366.8 99.045 367.41 99.075 ;
      RECT 364.235 99.045 364.845 99.075 ;
      RECT 365.515 99.045 366.125 99.075 ;
      RECT 368.075 99.045 368.685 99.075 ;
      RECT 365.735 95.595 365.905 99.045 ;
      RECT 364.155 99.075 368.765 99.245 ;
      RECT 368.935 95.425 369.885 95.595 ;
      RECT 368.935 99.075 369.885 99.245 ;
      RECT 368.935 95.595 369.105 99.075 ;
      RECT 369.715 95.595 369.885 99.075 ;
      RECT 367.655 95.485 367.825 98.855 ;
      RECT 430.385 92.78 430.915 92.95 ;
      RECT 430.48 92.26 430.81 92.78 ;
      RECT 429.71 92.26 430.04 92.95 ;
      RECT 431.145 92.47 431.665 93.08 ;
      RECT 431.145 92.085 432.435 92.47 ;
      RECT 434.33 92.26 434.66 92.95 ;
      RECT 431.935 92.74 432.435 97.165 ;
      RECT 431.935 97.165 433.205 97.61 ;
      RECT 432.705 97.61 433.205 99.625 ;
      RECT 432.79 92.26 433.12 92.95 ;
      RECT 433.56 92.26 433.89 92.95 ;
      RECT 436.225 92.26 436.755 92.43 ;
      RECT 434.985 92.26 435.515 92.43 ;
      RECT 437.85 92.26 438.18 92.95 ;
      RECT 437.08 92.26 437.41 92.95 ;
      RECT 440.075 92.47 440.595 93.08 ;
      RECT 439.305 92.085 440.595 92.47 ;
      RECT 439.305 92.74 439.805 97.165 ;
      RECT 438.535 97.165 439.805 97.61 ;
      RECT 438.535 97.61 439.035 99.625 ;
      RECT 440.825 92.78 441.355 92.95 ;
      RECT 440.93 92.26 441.26 92.78 ;
      RECT 441.7 92.26 442.03 92.95 ;
      RECT 438.62 92.26 438.95 92.95 ;
      RECT 447.755 96.23 449.145 96.4 ;
      RECT 447.215 91.77 447.385 95.39 ;
      RECT 447.765 95.245 460.045 95.815 ;
      RECT 447.765 91.345 460.045 91.915 ;
      RECT 447.765 94.465 460.045 95.035 ;
      RECT 447.765 93.685 460.045 94.255 ;
      RECT 447.765 92.905 460.045 93.475 ;
      RECT 447.765 92.125 460.045 92.695 ;
      RECT 460.595 91.77 460.765 95.39 ;
      RECT 19.65 103.265 20.6 103.435 ;
      RECT 19.65 99.615 20.6 99.785 ;
      RECT 20.43 99.785 20.6 103.265 ;
      RECT 19.65 99.785 19.82 103.265 ;
      RECT 20.77 99.615 21.88 99.785 ;
      RECT 20.77 103.265 21.88 103.435 ;
      RECT 20.85 99.785 21.46 99.815 ;
      RECT 21.71 99.785 21.88 103.265 ;
      RECT 24.615 103.265 25.72 103.435 ;
      RECT 24.61 99.615 25.72 99.785 ;
      RECT 25.55 99.785 25.72 103.265 ;
      RECT 24.275 102.715 24.445 103.375 ;
      RECT 24.27 102.485 24.445 102.715 ;
      RECT 23.33 99.615 24.44 99.785 ;
      RECT 24.27 99.785 24.44 102.485 ;
      RECT 22.05 103.265 23.16 103.435 ;
      RECT 22.05 99.615 23.16 99.785 ;
      RECT 22.99 99.785 23.16 103.265 ;
      RECT 23.33 103.265 24.1 103.435 ;
      RECT 27.055 103.265 27.78 103.435 ;
      RECT 27.055 99.615 27.78 99.785 ;
      RECT 27.61 99.785 27.78 103.265 ;
      RECT 26.83 100.795 27.44 100.965 ;
      RECT 26.83 100.965 27 102.715 ;
      RECT 26.83 100.005 27 100.795 ;
      RECT 25.89 99.615 26.66 99.785 ;
      RECT 25.97 99.785 26.58 99.815 ;
      RECT 363.71 127.905 370.075 127.935 ;
      RECT 363.71 125.185 370.075 125.215 ;
      RECT 361.715 127.04 363.94 127.705 ;
      RECT 361.715 125.415 363.94 126.035 ;
      RECT 361.72 104.365 363.445 105.115 ;
      RECT 361.72 103.825 361.915 104.365 ;
      RECT 369.845 125.415 371.155 127.705 ;
      RECT 361.72 107.84 361.915 108.45 ;
      RECT 361.72 107.09 363.445 107.84 ;
      RECT 361.72 105.115 361.915 107.09 ;
      RECT 361.715 117.4 361.915 125.365 ;
      RECT 361.745 108.45 361.915 117.4 ;
      RECT 370.985 86.19 371.155 104.255 ;
      RECT 361.715 126.035 363.91 127.04 ;
      RECT 361.715 127.705 371.155 127.755 ;
      RECT 361.715 125.365 371.155 125.415 ;
      RECT 370.985 127.905 371.155 133.775 ;
      RECT 363.71 127.755 371.155 127.905 ;
      RECT 370.985 107.995 371.155 125.215 ;
      RECT 363.71 125.215 371.155 125.365 ;
      RECT 361.745 133.775 371.155 133.945 ;
      RECT 361.715 127.755 361.915 133.1 ;
      RECT 362.105 85.42 362.275 86.4 ;
      RECT 370.475 88.31 370.675 93.725 ;
      RECT 370.505 93.725 370.675 94.355 ;
      RECT 370.505 87.565 370.675 88.31 ;
      RECT 386.27 86.53 386.6 87.18 ;
      RECT 387.53 86.53 387.86 87.18 ;
      RECT 386.9 86.53 387.23 87.18 ;
      RECT 388.79 86.53 389.12 87.18 ;
      RECT 388.16 86.53 388.49 87.18 ;
      RECT 389.42 86.53 389.75 87.18 ;
      RECT 390.05 86.53 390.38 87.18 ;
      RECT 386.27 87.56 386.6 88.21 ;
      RECT 386.9 87.56 387.23 88.21 ;
      RECT 387.53 87.56 387.86 88.21 ;
      RECT 388.79 87.56 389.12 88.21 ;
      RECT 388.16 87.56 388.49 88.21 ;
      RECT 389.42 87.56 389.75 88.21 ;
      RECT 390.05 87.56 390.38 88.21 ;
      RECT 390.68 86.53 391.01 87.18 ;
      RECT 391.31 86.53 391.64 87.18 ;
      RECT 391.94 86.53 392.27 87.18 ;
      RECT 393.2 86.53 393.53 87.18 ;
      RECT 392.57 86.53 392.9 87.18 ;
      RECT 393.83 86.53 394.16 87.18 ;
      RECT 394.46 86.53 394.79 87.18 ;
      RECT 390.68 87.56 391.01 88.21 ;
      RECT 391.31 87.56 391.64 88.21 ;
      RECT 391.94 87.56 392.27 88.21 ;
      RECT 393.2 87.56 393.53 88.21 ;
      RECT 392.57 87.56 392.9 88.21 ;
      RECT 393.83 87.56 394.16 88.21 ;
      RECT 394.46 87.56 394.79 88.21 ;
      RECT 400.46 86.33 401.47 86.5 ;
      RECT 401.64 86.33 404.57 86.51 ;
      RECT 404.74 86.33 405.75 86.5 ;
      RECT 405.92 86.33 408.85 86.51 ;
      RECT 409.02 86.33 410.03 86.5 ;
      RECT 417.9 86.33 418.91 86.5 ;
      RECT 414.62 86.33 415.63 86.5 ;
      RECT 415.8 86.33 417.73 86.51 ;
      RECT 419.08 86.33 420.01 86.51 ;
      RECT 422.46 86.33 423.47 86.5 ;
      RECT 420.18 86.33 421.19 86.5 ;
      RECT 421.36 86.33 422.29 86.51 ;
      RECT 430.48 85.105 430.81 85.795 ;
      RECT 429.71 85.105 430.04 85.795 ;
      RECT 436.31 85.105 436.64 85.795 ;
      RECT 434.33 85.105 434.66 85.795 ;
      RECT 431.25 85.395 432.35 85.795 ;
      RECT 431.25 84.8 433.89 85.395 ;
      RECT 432.79 85.585 433.89 85.925 ;
      RECT 435.1 85.105 435.43 85.795 ;
      RECT 437.85 85.585 438.95 85.925 ;
      RECT 437.08 85.105 437.41 85.795 ;
      RECT 439.39 85.395 440.49 85.795 ;
      RECT 437.85 84.8 440.49 85.395 ;
      RECT 440.93 85.105 441.26 85.795 ;
      RECT 441.7 85.105 442.03 85.795 ;
      RECT 453.22 85.635 456.36 85.805 ;
      RECT 457.755 82.24 458.265 82.57 ;
      RECT 457.825 82.57 458.195 84.045 ;
      RECT 457.825 84.045 458.355 84.215 ;
      RECT 457.755 86.185 458.265 86.515 ;
      RECT 457.825 84.61 458.195 86.185 ;
      RECT 457.825 84.44 458.355 84.61 ;
      RECT 459.245 82.74 459.415 84.045 ;
      RECT 458.885 84.045 459.415 84.215 ;
      RECT 458.365 82.74 458.535 83.75 ;
      RECT 457.485 82.74 457.655 83.79 ;
      RECT 459.245 84.61 459.415 86.015 ;
      RECT 458.885 84.44 459.415 84.61 ;
      RECT 458.365 84.965 458.535 86.015 ;
      RECT 20.12 95.425 21.07 95.595 ;
      RECT 20.12 99.075 21.07 99.245 ;
      RECT 20.9 95.595 21.07 99.075 ;
      RECT 20.12 95.595 20.29 99.075 ;
      RECT 24.74 95.485 24.91 98.855 ;
      RECT 23.46 96.145 23.63 98.855 ;
      RECT 22.18 95.485 22.35 98.855 ;
      RECT 21.54 95.595 21.71 99.045 ;
      RECT 21.24 95.425 22.01 95.595 ;
      RECT 25.38 95.595 25.55 99.045 ;
      RECT 22.52 95.425 23.29 95.595 ;
      RECT 25.08 95.425 25.85 95.595 ;
      RECT 23.8 95.425 24.57 95.595 ;
      RECT 21.32 99.045 21.93 99.075 ;
      RECT 22.595 99.045 23.205 99.075 ;
      RECT 25.16 99.045 25.77 99.075 ;
      RECT 21.24 99.075 25.85 99.245 ;
      RECT 23.88 99.045 24.49 99.075 ;
      RECT 22.815 95.595 22.985 99.045 ;
      RECT 24.1 95.595 24.27 99.045 ;
      RECT 26.02 95.425 26.97 95.595 ;
      RECT 26.02 99.075 26.97 99.245 ;
      RECT 26.02 95.595 26.19 99.075 ;
      RECT 26.8 95.595 26.97 99.075 ;
      RECT 32.915 95.62 33.085 95.73 ;
      RECT 32.915 94.495 33.765 95.62 ;
      RECT 32.875 89.62 33.765 94.495 ;
      RECT 32.915 85.71 33.765 89.62 ;
      RECT 37.875 85.71 39.195 95.62 ;
      RECT 43.305 85.71 43.475 95.56 ;
      RECT 47.585 85.71 48.905 95.62 ;
      RECT 53.695 95.62 53.865 95.73 ;
      RECT 53.015 89.62 53.905 94.495 ;
      RECT 287.945 83 288.115 84.335 ;
      RECT 286.89 88.725 287.445 88.895 ;
      RECT 287.275 88.895 287.445 88.94 ;
      RECT 287.275 88.61 287.445 88.725 ;
      RECT 287.215 83.765 287.385 86.475 ;
      RECT 287.345 88.205 289.565 88.425 ;
      RECT 287.565 82.81 287.765 86.995 ;
      RECT 287.58 86.995 287.75 87.34 ;
      RECT 287.565 82.14 288.53 82.81 ;
      RECT 286.435 83.765 286.605 86.475 ;
      RECT 288.825 83 288.995 84.01 ;
      RECT 288.56 84.535 289.23 84.705 ;
      RECT 288.56 84.705 289.09 84.735 ;
      RECT 302.215 98.39 316.875 98.56 ;
      RECT 309.415 85.73 309.585 96.45 ;
      RECT 303.815 88.08 303.985 88.52 ;
      RECT 303.815 87.85 303.985 87.91 ;
      RECT 302.215 86.04 302.385 87.36 ;
      RECT 302.215 97.225 310.285 97.815 ;
      RECT 302.215 97.815 309.585 98.39 ;
      RECT 302.215 87.91 303.985 88.08 ;
      RECT 302.215 87.53 302.385 87.91 ;
      RECT 302.215 87.36 303.745 87.53 ;
      RECT 302.215 89.97 303.525 90.14 ;
      RECT 302.215 88.08 302.385 89.97 ;
      RECT 302.215 90.14 302.385 96.45 ;
      RECT 302.215 96.45 309.585 97.225 ;
      RECT 302.725 86.08 303.745 86.25 ;
      RECT 299.795 82.265 301.815 83.015 ;
      RECT 305.11 81.61 305.92 81.78 ;
      RECT 306.39 81.61 307.2 81.78 ;
      RECT 306.51 81.18 307.04 81.61 ;
      RECT 307.67 81.61 308.48 81.78 ;
      RECT 307.79 81.18 308.32 81.61 ;
      RECT 308.95 81.61 309.76 81.78 ;
      RECT 309.07 81.18 309.6 81.61 ;
      RECT 304.555 85.71 304.725 95.56 ;
      RECT 305.25 82.615 305.78 82.785 ;
      RECT 308.835 85.71 309.005 95.56 ;
      RECT 303.945 86.305 304.115 87.305 ;
      RECT 304.78 85.37 308.78 85.54 ;
      RECT 304.78 95.92 308.78 96.09 ;
      RECT 304.895 85.54 308.665 95.92 ;
      RECT 310.23 81.61 311.04 81.78 ;
      RECT 310.35 81.18 310.88 81.61 ;
      RECT 311.51 81.61 312.32 81.78 ;
      RECT 311.63 81.18 312.16 81.61 ;
      RECT 312.79 81.61 313.6 81.78 ;
      RECT 312.91 81.18 313.44 81.61 ;
      RECT 314.07 81.61 314.88 81.78 ;
      RECT 314.19 81.18 314.72 81.61 ;
      RECT 313.245 85.37 317.245 85.54 ;
      RECT 313.245 95.92 317.245 96.09 ;
      RECT 313.36 85.54 317.13 95.92 ;
      RECT 312.34 95.62 312.51 95.73 ;
      RECT 312.3 88.5 313.19 93.375 ;
      RECT 312.34 93.375 313.19 95.62 ;
      RECT 312.34 85.71 313.19 88.5 ;
      RECT 320.47 81.61 321.28 81.78 ;
      RECT 320.59 81.18 321.12 81.61 ;
      RECT 315.35 81.61 316.16 81.78 ;
      RECT 315.47 81.18 316 81.61 ;
      RECT 316.63 81.61 317.44 81.78 ;
      RECT 316.75 81.18 317.28 81.61 ;
      RECT 317.91 81.61 318.72 81.78 ;
      RECT 318.03 81.18 318.56 81.61 ;
      RECT 319.19 81.61 320 81.78 ;
      RECT 319.31 81.18 319.84 81.61 ;
      RECT 318.675 85.37 322.675 85.54 ;
      RECT 318.675 95.92 322.675 96.09 ;
      RECT 318.79 85.54 322.56 95.92 ;
      RECT 317.3 85.71 318.62 95.62 ;
      RECT 326.87 81.61 327.68 81.78 ;
      RECT 326.99 81.18 327.52 81.61 ;
      RECT 321.75 81.61 322.56 81.78 ;
      RECT 321.87 81.18 322.4 81.61 ;
      RECT 323.03 81.61 323.84 81.78 ;
      RECT 323.15 81.18 323.68 81.61 ;
      RECT 324.31 81.61 325.12 81.78 ;
      RECT 324.43 81.18 324.96 81.61 ;
      RECT 325.59 81.61 326.4 81.78 ;
      RECT 325.71 81.18 326.24 81.61 ;
      RECT 322.955 85.37 326.955 85.54 ;
      RECT 322.955 95.92 326.955 96.09 ;
      RECT 323.07 85.54 326.84 95.92 ;
      RECT 322.73 85.71 322.9 95.56 ;
      RECT 328.15 81.61 328.96 81.78 ;
      RECT 328.27 81.18 328.8 81.61 ;
      RECT 329.43 81.61 330.24 81.78 ;
      RECT 329.55 81.18 330.08 81.61 ;
      RECT 330.71 81.61 331.52 81.78 ;
      RECT 330.83 81.18 331.36 81.61 ;
      RECT 331.99 81.61 332.8 81.78 ;
      RECT 332.11 81.18 332.64 81.61 ;
      RECT 328.385 85.37 332.385 85.54 ;
      RECT 328.385 95.92 332.385 96.09 ;
      RECT 328.5 85.54 332.27 95.92 ;
      RECT 332.44 88.5 333.33 93.375 ;
      RECT 332.44 93.375 333.29 95.62 ;
      RECT 332.44 85.71 333.29 88.5 ;
      RECT 333.12 95.62 333.29 95.73 ;
      RECT 327.01 85.71 328.33 95.62 ;
      RECT 333.27 81.61 334.08 81.78 ;
      RECT 333.39 81.18 333.92 81.61 ;
      RECT 337.045 85.37 341.245 85.54 ;
      RECT 337.045 95.92 341.245 96.09 ;
      RECT 337.16 85.54 340.93 95.92 ;
      RECT 338.57 82.39 339.1 82.56 ;
      RECT 342.475 85.37 346.475 85.54 ;
      RECT 342.475 95.92 346.475 96.09 ;
      RECT 342.59 85.54 346.36 95.92 ;
      RECT 345.83 81.61 346.54 81.78 ;
      RECT 345.985 80.88 346.155 81.61 ;
      RECT 346.755 85.37 350.755 85.54 ;
      RECT 346.755 95.92 350.755 96.09 ;
      RECT 346.87 85.54 350.64 95.92 ;
      RECT 352.185 85.37 356.185 85.54 ;
      RECT 352.185 95.92 356.185 96.09 ;
      RECT 352.3 85.54 356.07 95.92 ;
      RECT 362.225 87.565 362.395 94.355 ;
      RECT 362.495 85.175 365.205 85.345 ;
      RECT 362.495 86.455 365.205 86.625 ;
      RECT 361.745 84.375 371.155 84.545 ;
      RECT 365.825 84.545 371.155 86.19 ;
      RECT 361.745 84.545 361.915 103.825 ;
      RECT 361.745 133.1 361.915 133.775 ;
      RECT 369.815 104.255 371.155 107.995 ;
      RECT 259.13 85.15 260.14 85.32 ;
      RECT 262.165 87.005 265.935 87.175 ;
      RECT 262.165 87 265.895 87.005 ;
      RECT 257.945 87.005 261.715 87.175 ;
      RECT 257.97 87 261.7 87.005 ;
      RECT 262.045 85.15 263.735 85.32 ;
      RECT 261.14 81.95 261.31 84.85 ;
      RECT 259.95 81.335 260.62 81.57 ;
      RECT 261.63 84.07 262.16 84.24 ;
      RECT 261.63 84.24 261.8 84.93 ;
      RECT 261.63 82.22 261.8 84.07 ;
      RECT 258.65 83.29 259.18 83.46 ;
      RECT 258.83 83.46 259 84.93 ;
      RECT 258.83 82.22 259 83.29 ;
      RECT 259.95 83.29 260.56 83.46 ;
      RECT 260.39 83.46 260.56 84.93 ;
      RECT 260.39 82.22 260.56 83.29 ;
      RECT 262.41 82.2 262.58 84.93 ;
      RECT 258.05 82.14 258.22 84.93 ;
      RECT 261.83 85.77 262 86.78 ;
      RECT 266.875 87 267.885 87.17 ;
      RECT 267.05 85.34 267.7 87 ;
      RECT 268.165 87 269.175 87.17 ;
      RECT 268.335 86.58 268.985 87 ;
      RECT 268.335 84.74 268.69 86.58 ;
      RECT 268.335 84.57 268.865 84.74 ;
      RECT 268.235 83.09 268.905 83.49 ;
      RECT 264.275 81.49 265.165 81.51 ;
      RECT 264.215 81.32 264.885 81.34 ;
      RECT 264.215 81.34 265.165 81.49 ;
      RECT 265.28 81.95 265.45 84.85 ;
      RECT 265.96 86.58 266.49 86.75 ;
      RECT 266.11 86.75 266.28 86.78 ;
      RECT 266.11 85.77 266.28 86.58 ;
      RECT 266.12 90.46 288.2 90.7 ;
      RECT 256.7 89.69 267.165 89.87 ;
      RECT 266.12 90.11 267.165 90.46 ;
      RECT 266.37 88.61 267.165 89.69 ;
      RECT 246.24 89.87 267.165 90.11 ;
      RECT 267.94 84.07 268.11 86.78 ;
      RECT 266.66 84.97 267.19 85.14 ;
      RECT 266.66 85.14 266.83 86.78 ;
      RECT 266.66 84.07 266.83 84.97 ;
      RECT 263.97 82.2 264.14 84.93 ;
      RECT 264.39 84.07 264.92 84.24 ;
      RECT 264.75 84.24 264.92 84.93 ;
      RECT 264.75 82.22 264.92 84.07 ;
      RECT 265.205 88.075 268.6 88.36 ;
      RECT 246.315 89.285 266.11 89.455 ;
      RECT 267.405 89.285 287.22 89.455 ;
      RECT 265.205 88.36 265.87 89.285 ;
      RECT 267.895 88.36 268.6 89.285 ;
      RECT 268.86 85.34 269.39 85.51 ;
      RECT 269.22 85.51 269.39 86.78 ;
      RECT 269.22 84.07 269.39 85.34 ;
      RECT 274.235 87.275 276.805 87.475 ;
      RECT 270.075 87.17 272.765 87.175 ;
      RECT 270.05 87 272.76 87.005 ;
      RECT 270.05 87.005 272.765 87.17 ;
      RECT 273.37 83.61 273.54 86.76 ;
      RECT 269.38 83.09 272.77 83.51 ;
      RECT 269.77 83.73 273.06 83.9 ;
      RECT 270.01 83.69 273.06 83.73 ;
      RECT 269.77 83.9 269.94 86.78 ;
      RECT 272.89 83.9 273.06 86.78 ;
      RECT 271.33 83.9 271.5 86.78 ;
      RECT 273.2 82.61 277.95 82.78 ;
      RECT 273.85 84.275 274.02 87.055 ;
      RECT 271.92 84.97 272.45 85.14 ;
      RECT 272.11 85.14 272.28 86.78 ;
      RECT 272.11 84.07 272.28 84.97 ;
      RECT 270.36 85.34 270.89 85.51 ;
      RECT 270.55 85.51 270.72 86.78 ;
      RECT 270.55 84.07 270.72 85.34 ;
      RECT 274.455 81.725 278.09 81.73 ;
      RECT 273.2 81.73 278.09 81.895 ;
      RECT 273.2 81.895 277.95 81.9 ;
      RECT 274.45 85.23 274.98 85.4 ;
      RECT 274.63 85.4 274.8 87.055 ;
      RECT 274.63 84.345 274.8 85.23 ;
      RECT 273.2 80.85 277.95 81.02 ;
      RECT 280.445 87.275 282.475 87.445 ;
      RECT 280.505 87.445 282.415 87.455 ;
      RECT 277.885 87.275 279.915 87.445 ;
      RECT 277.945 87.445 279.855 87.455 ;
      RECT 279.245 81.805 281.955 81.975 ;
      RECT 279.36 81.775 280.62 81.805 ;
      RECT 280.08 84.215 280.25 86.925 ;
      RECT 277.52 84.215 277.69 86.925 ;
      RECT 276.97 84.275 277.14 87.055 ;
      RECT 275.41 84.275 275.58 87.055 ;
      RECT 280.935 81.095 282.145 81.1 ;
      RECT 279.245 80.925 281.955 80.93 ;
      RECT 279.245 80.93 282.145 81.095 ;
      RECT 278.275 83.8 278.865 83.97 ;
      RECT 278.275 81.955 278.6 83.8 ;
      RECT 275.99 86.68 276.52 86.85 ;
      RECT 276.19 86.85 276.36 87.055 ;
      RECT 276.19 84.345 276.36 86.68 ;
      RECT 278.6 85.23 279.13 85.4 ;
      RECT 278.8 85.4 278.97 86.925 ;
      RECT 278.8 84.215 278.97 85.23 ;
      RECT 279.475 82.625 282.125 83.565 ;
      RECT 284.985 83.755 285.155 85.105 ;
      RECT 283.645 83.815 284.045 86.825 ;
      RECT 283.705 83.755 283.875 83.815 ;
      RECT 285.055 85.74 285.225 86.825 ;
      RECT 282.64 84.215 282.81 86.925 ;
      RECT 285.655 83.765 285.825 86.475 ;
      RECT 283.93 83.365 284.93 83.535 ;
      RECT 283.99 83.535 284.87 83.625 ;
      RECT 283.08 87.015 285 87.21 ;
      RECT 284 87.21 285 87.215 ;
      RECT 282.825 83.8 283.415 83.97 ;
      RECT 283.08 83.97 283.415 87.015 ;
      RECT 281.185 86.68 281.715 86.85 ;
      RECT 281.36 86.85 281.53 86.925 ;
      RECT 281.36 84.215 281.53 86.68 ;
      RECT 285.88 83.375 287.16 83.545 ;
      RECT 287.945 81.435 288.115 81.965 ;
      RECT 289.19 85.03 289.775 85.2 ;
      RECT 289.19 85.2 289.36 85.935 ;
      RECT 289.19 84.925 289.36 85.03 ;
      RECT 288.41 84.925 288.58 85.935 ;
      RECT 289.7 83.09 289.875 83.945 ;
      RECT 289.705 83.945 289.875 84.01 ;
      RECT 289.705 83 289.875 83.09 ;
      RECT 221.875 81.48 222.545 81.65 ;
      RECT 221.955 81.395 222.485 81.48 ;
      RECT 219.695 83.66 220.225 83.83 ;
      RECT 219.695 83.83 219.865 84.415 ;
      RECT 219.695 83.405 219.865 83.66 ;
      RECT 220.08 84.555 220.25 85.565 ;
      RECT 220.3 85.85 220.83 86.02 ;
      RECT 220.42 84.615 221.08 85.575 ;
      RECT 220.86 83.06 221.08 84.615 ;
      RECT 220.86 82.05 221.135 83.06 ;
      RECT 220.42 85.575 220.83 85.85 ;
      RECT 221 85.87 221.67 86.04 ;
      RECT 221.25 84.485 221.42 85.87 ;
      RECT 221.555 84.07 222.445 84.24 ;
      RECT 221.555 83.735 222.085 84.07 ;
      RECT 221.33 83.31 222.68 83.48 ;
      RECT 221.64 84.595 222.25 84.765 ;
      RECT 221.64 84.765 221.81 85.565 ;
      RECT 221.64 84.555 221.81 84.595 ;
      RECT 226.195 81.77 226.725 81.94 ;
      RECT 226.365 81.94 226.535 83.06 ;
      RECT 224.205 81.395 224.795 81.94 ;
      RECT 224.205 81.94 224.375 83.06 ;
      RECT 226.98 83.29 229.31 83.46 ;
      RECT 222.9 84.745 229.69 84.915 ;
      RECT 226.98 83.46 229.25 84.745 ;
      RECT 223.065 83.895 226.54 84.405 ;
      RECT 223.065 82.05 223.435 83.895 ;
      RECT 225.125 82.05 225.91 83.895 ;
      RECT 223.605 83.31 224.955 83.48 ;
      RECT 225.165 81.43 227.875 81.6 ;
      RECT 222.755 81.395 223.425 81.565 ;
      RECT 226.11 83.31 226.78 83.48 ;
      RECT 228.165 81.77 228.695 81.94 ;
      RECT 228.525 81.94 228.695 83.06 ;
      RECT 227.445 82.05 227.615 83.06 ;
      RECT 231.765 84.56 234.475 84.715 ;
      RECT 230.935 84.545 234.475 84.56 ;
      RECT 230.935 81.285 231.105 84.38 ;
      RECT 230.935 84.38 234.46 84.545 ;
      RECT 232.09 80.77 232.62 80.94 ;
      RECT 232.265 80.94 232.435 83.995 ;
      RECT 233.465 80.77 233.995 80.94 ;
      RECT 233.825 80.94 233.995 83.995 ;
      RECT 230.935 84.95 231.105 85.465 ;
      RECT 230.935 84.78 231.525 84.95 ;
      RECT 229.795 84.01 230.325 84.18 ;
      RECT 230.155 84.465 230.765 84.795 ;
      RECT 230.155 84.18 230.325 84.465 ;
      RECT 230.155 81.285 230.325 84.01 ;
      RECT 233.045 81.285 233.215 83.995 ;
      RECT 238.26 87.15 240.29 87.32 ;
      RECT 237.97 83.29 238.5 83.46 ;
      RECT 237.97 83.46 238.14 86.64 ;
      RECT 237.97 81.89 238.14 83.29 ;
      RECT 236.4 81.285 236.57 86.27 ;
      RECT 234.84 81.285 235.01 86.27 ;
      RECT 235.96 80.895 236.63 81.065 ;
      RECT 236.04 80.8 236.57 80.895 ;
      RECT 234.78 80.895 235.45 81.065 ;
      RECT 234.84 80.8 235.37 80.895 ;
      RECT 238.85 81.89 239.02 86.64 ;
      RECT 239.56 83.29 240.09 83.46 ;
      RECT 239.73 83.46 239.9 86.64 ;
      RECT 239.73 81.89 239.9 83.29 ;
      RECT 243.78 86.43 244.94 86.94 ;
      RECT 242.18 86.43 243.34 86.94 ;
      RECT 245.46 83.29 246.01 83.46 ;
      RECT 245.46 83.46 245.63 86.64 ;
      RECT 245.46 81.89 245.63 83.29 ;
      RECT 240.61 81.89 240.78 86.64 ;
      RECT 241.11 83.29 241.66 83.46 ;
      RECT 241.49 83.46 241.66 86.64 ;
      RECT 241.49 81.89 241.66 83.29 ;
      RECT 245.595 87.15 246.265 87.32 ;
      RECT 240.855 87.15 241.525 87.32 ;
      RECT 249.9 81.45 250.57 81.94 ;
      RECT 250.25 87.15 251.6 87.32 ;
      RECT 247.205 81.3 248.215 81.47 ;
      RECT 247.455 80.875 247.985 81.3 ;
      RECT 245.925 81.3 246.935 81.47 ;
      RECT 246.175 80.875 246.705 81.3 ;
      RECT 246.83 87.15 248.86 87.32 ;
      RECT 249.47 85.82 249.65 86.35 ;
      RECT 249.47 86.35 249.64 86.765 ;
      RECT 249.47 81.95 249.64 85.82 ;
      RECT 249.96 82.18 250.13 86.93 ;
      RECT 248.62 83.29 249.15 83.46 ;
      RECT 248.98 83.46 249.15 86.64 ;
      RECT 248.98 81.89 249.15 83.29 ;
      RECT 246.34 81.89 246.51 86.64 ;
      RECT 246.09 88.895 246.62 89.065 ;
      RECT 246.09 88.61 246.26 88.895 ;
      RECT 248.1 81.89 248.27 86.64 ;
      RECT 247.03 83.29 247.56 83.46 ;
      RECT 247.22 83.46 247.39 86.64 ;
      RECT 247.22 81.89 247.39 83.29 ;
      RECT 251.98 81.43 252.65 81.6 ;
      RECT 251.98 81.4 252.51 81.43 ;
      RECT 254.82 85.15 256.17 85.32 ;
      RECT 255.205 81.03 256.215 81.545 ;
      RECT 257.07 85.76 257.24 85.77 ;
      RECT 257.07 85.77 257.72 86.78 ;
      RECT 251.72 82.18 251.89 86.93 ;
      RECT 252.24 83.69 252.77 83.86 ;
      RECT 252.6 83.86 252.77 86.93 ;
      RECT 252.6 82.18 252.77 83.69 ;
      RECT 253.16 81.95 253.33 84.85 ;
      RECT 256.78 81.95 256.95 84.85 ;
      RECT 253.715 81.325 254.385 81.57 ;
      RECT 256.465 81.33 257.135 81.5 ;
      RECT 257.27 83.29 257.88 83.46 ;
      RECT 257.27 83.46 257.44 84.93 ;
      RECT 257.27 82.22 257.44 83.29 ;
      RECT 254.53 83.3 255.23 83.47 ;
      RECT 254.53 83.47 254.7 84.93 ;
      RECT 254.53 82.22 254.7 83.3 ;
      RECT 255.76 83.3 256.46 83.47 ;
      RECT 256.29 83.47 256.46 84.93 ;
      RECT 256.29 82.22 256.46 83.3 ;
      RECT 255.41 82.14 255.58 84.93 ;
      RECT 261.49 81.805 262.81 81.94 ;
      RECT 261.46 81.335 262.81 81.805 ;
      RECT 257.53 81.335 258.54 81.505 ;
      RECT 257.53 81.19 258.115 81.335 ;
      RECT 257.585 81.02 258.115 81.19 ;
      RECT 257.665 85.15 258.675 85.32 ;
      RECT 133.545 83.3 134.245 83.47 ;
      RECT 133.545 83.47 133.715 84.93 ;
      RECT 133.545 82.22 133.715 83.3 ;
      RECT 131.785 82.14 131.955 84.93 ;
      RECT 134.425 82.14 134.595 84.93 ;
      RECT 137.355 81.43 138.025 81.6 ;
      RECT 137.495 81.4 138.025 81.43 ;
      RECT 139.435 81.45 140.105 81.94 ;
      RECT 138.405 87.15 139.755 87.32 ;
      RECT 141.145 87.15 143.175 87.32 ;
      RECT 140.355 85.82 140.535 86.35 ;
      RECT 140.365 86.35 140.535 86.765 ;
      RECT 140.365 81.95 140.535 85.82 ;
      RECT 138.115 82.18 138.285 86.93 ;
      RECT 139.875 82.18 140.045 86.93 ;
      RECT 137.235 83.69 137.765 83.86 ;
      RECT 137.235 83.86 137.405 86.93 ;
      RECT 137.235 82.18 137.405 83.69 ;
      RECT 140.855 83.29 141.385 83.46 ;
      RECT 140.855 83.46 141.025 86.64 ;
      RECT 140.855 81.89 141.025 83.29 ;
      RECT 136.675 81.95 136.845 84.85 ;
      RECT 145.065 86.43 146.225 86.94 ;
      RECT 141.79 81.3 142.8 81.47 ;
      RECT 142.02 80.875 142.55 81.3 ;
      RECT 143.07 81.3 144.08 81.47 ;
      RECT 143.3 80.875 143.83 81.3 ;
      RECT 146.665 86.43 147.825 86.94 ;
      RECT 143.495 81.89 143.665 86.64 ;
      RECT 143.995 83.29 144.545 83.46 ;
      RECT 144.375 83.46 144.545 86.64 ;
      RECT 144.375 81.89 144.545 83.29 ;
      RECT 143.74 87.15 144.41 87.32 ;
      RECT 143.385 88.895 143.915 89.065 ;
      RECT 143.745 88.61 143.915 88.895 ;
      RECT 141.735 81.89 141.905 86.64 ;
      RECT 142.445 83.29 142.975 83.46 ;
      RECT 142.615 83.46 142.785 86.64 ;
      RECT 142.615 81.89 142.785 83.29 ;
      RECT 149.715 87.15 151.745 87.32 ;
      RECT 151.505 83.29 152.035 83.46 ;
      RECT 151.865 83.46 152.035 86.64 ;
      RECT 151.865 81.89 152.035 83.29 ;
      RECT 149.225 81.89 149.395 86.64 ;
      RECT 148.345 83.29 148.895 83.46 ;
      RECT 148.345 83.46 148.515 86.64 ;
      RECT 148.345 81.89 148.515 83.29 ;
      RECT 148.48 87.15 149.15 87.32 ;
      RECT 150.985 81.89 151.155 86.64 ;
      RECT 149.915 83.29 150.445 83.46 ;
      RECT 150.105 83.46 150.275 86.64 ;
      RECT 150.105 81.89 150.275 83.29 ;
      RECT 155.53 84.56 158.24 84.715 ;
      RECT 155.53 84.545 159.07 84.56 ;
      RECT 158.9 81.285 159.07 84.38 ;
      RECT 155.545 84.38 159.07 84.545 ;
      RECT 157.385 80.77 157.915 80.94 ;
      RECT 157.57 80.94 157.74 83.995 ;
      RECT 156.01 80.77 156.54 80.94 ;
      RECT 156.01 80.94 156.18 83.995 ;
      RECT 158.9 84.95 159.07 85.465 ;
      RECT 158.48 84.78 159.07 84.95 ;
      RECT 153.435 81.285 153.605 86.27 ;
      RECT 154.995 81.285 155.165 86.27 ;
      RECT 153.375 80.895 154.045 81.065 ;
      RECT 153.435 80.8 153.965 80.895 ;
      RECT 154.555 80.895 155.225 81.065 ;
      RECT 154.635 80.8 155.165 80.895 ;
      RECT 156.79 81.285 156.96 83.995 ;
      RECT 160.695 83.29 163.025 83.46 ;
      RECT 160.315 84.745 167.105 84.915 ;
      RECT 160.755 83.46 163.025 84.745 ;
      RECT 161.31 81.77 161.84 81.94 ;
      RECT 161.31 81.94 161.48 83.06 ;
      RECT 159.68 84.01 160.21 84.18 ;
      RECT 159.24 84.465 159.85 84.795 ;
      RECT 159.68 84.18 159.85 84.465 ;
      RECT 159.68 81.285 159.85 84.01 ;
      RECT 164.095 82.05 164.88 83.895 ;
      RECT 166.57 82.05 166.94 83.895 ;
      RECT 163.465 83.895 166.94 84.405 ;
      RECT 163.28 81.77 163.81 81.94 ;
      RECT 163.47 81.94 163.64 83.06 ;
      RECT 162.13 81.43 164.84 81.6 ;
      RECT 163.225 83.31 163.895 83.48 ;
      RECT 162.39 82.05 162.56 83.06 ;
      RECT 169.175 85.85 169.705 86.02 ;
      RECT 168.87 82.05 169.145 83.06 ;
      RECT 169.175 85.575 169.585 85.85 ;
      RECT 168.925 83.06 169.145 84.615 ;
      RECT 168.925 84.615 169.585 85.575 ;
      RECT 165.21 81.395 165.8 81.94 ;
      RECT 165.63 81.94 165.8 83.06 ;
      RECT 167.43 81.82 167.96 81.99 ;
      RECT 167.79 81.99 167.96 83.06 ;
      RECT 167.46 81.48 168.13 81.65 ;
      RECT 167.52 81.395 168.05 81.48 ;
      RECT 166.58 81.395 167.25 81.565 ;
      RECT 168.34 81.395 169.53 81.565 ;
      RECT 169.36 84.03 169.95 84.2 ;
      RECT 169.36 84.2 169.53 84.415 ;
      RECT 169.36 81.565 169.53 84.03 ;
      RECT 165.05 83.31 166.4 83.48 ;
      RECT 167.325 83.31 168.675 83.48 ;
      RECT 167.92 83.735 168.45 84.07 ;
      RECT 167.56 84.07 168.45 84.24 ;
      RECT 167.755 84.595 168.365 84.765 ;
      RECT 168.195 84.555 168.365 84.595 ;
      RECT 168.195 84.765 168.365 85.565 ;
      RECT 168.335 85.87 169.005 86.04 ;
      RECT 168.585 84.485 168.755 85.87 ;
      RECT 169.78 83.66 170.31 83.83 ;
      RECT 170.14 83.83 170.31 84.415 ;
      RECT 170.14 83.405 170.31 83.66 ;
      RECT 169.755 84.555 169.925 85.565 ;
      RECT 173.185 81.37 173.715 81.94 ;
      RECT 172.165 81.285 172.675 81.615 ;
      RECT 172.305 81.615 172.675 84.93 ;
      RECT 216.29 81.37 216.82 81.94 ;
      RECT 217.33 81.285 217.84 81.615 ;
      RECT 217.33 81.615 217.7 84.93 ;
      RECT 220.475 81.395 221.665 81.565 ;
      RECT 220.475 81.565 220.645 84.03 ;
      RECT 220.475 84.2 220.645 84.415 ;
      RECT 220.055 84.03 220.645 84.2 ;
      RECT 222.045 81.82 222.575 81.99 ;
      RECT 222.045 81.99 222.215 83.06 ;
      RECT 103.4 83.765 103.57 86.475 ;
      RECT 102.845 83.375 104.125 83.545 ;
      RECT 107.53 87.275 109.56 87.445 ;
      RECT 107.59 87.445 109.5 87.455 ;
      RECT 110.09 87.275 112.12 87.445 ;
      RECT 110.15 87.445 112.06 87.455 ;
      RECT 112.055 82.61 116.805 82.78 ;
      RECT 108.05 81.805 110.76 81.975 ;
      RECT 109.385 81.775 110.645 81.805 ;
      RECT 107.195 84.215 107.365 86.925 ;
      RECT 109.755 84.215 109.925 86.925 ;
      RECT 112.315 84.215 112.485 86.925 ;
      RECT 107.86 81.095 109.07 81.1 ;
      RECT 108.05 80.925 110.76 80.93 ;
      RECT 107.86 80.93 110.76 81.095 ;
      RECT 111.915 81.725 115.55 81.73 ;
      RECT 111.915 81.73 116.805 81.895 ;
      RECT 112.055 81.895 116.805 81.9 ;
      RECT 108.29 86.68 108.82 86.85 ;
      RECT 108.475 86.85 108.645 86.925 ;
      RECT 108.475 84.215 108.645 86.68 ;
      RECT 111.14 83.8 111.73 83.97 ;
      RECT 111.405 81.955 111.73 83.8 ;
      RECT 110.875 85.23 111.405 85.4 ;
      RECT 111.035 85.4 111.205 86.925 ;
      RECT 111.035 84.215 111.205 85.23 ;
      RECT 112.055 80.85 116.805 81.02 ;
      RECT 107.88 82.625 110.53 83.565 ;
      RECT 113.2 87.275 115.77 87.475 ;
      RECT 117.24 87.17 119.93 87.175 ;
      RECT 117.245 87 119.955 87.005 ;
      RECT 117.24 87.005 119.955 87.17 ;
      RECT 116.465 83.61 116.635 86.76 ;
      RECT 117.235 83.09 120.625 83.51 ;
      RECT 116.945 83.73 120.235 83.9 ;
      RECT 116.945 83.69 119.995 83.73 ;
      RECT 116.945 83.9 117.115 86.78 ;
      RECT 120.065 83.9 120.235 86.78 ;
      RECT 118.505 83.9 118.675 86.78 ;
      RECT 112.865 84.275 113.035 87.055 ;
      RECT 114.425 84.275 114.595 87.055 ;
      RECT 115.985 84.275 116.155 87.055 ;
      RECT 117.555 84.97 118.085 85.14 ;
      RECT 117.725 85.14 117.895 86.78 ;
      RECT 117.725 84.07 117.895 84.97 ;
      RECT 115.025 85.23 115.555 85.4 ;
      RECT 115.205 85.4 115.375 87.055 ;
      RECT 115.205 84.345 115.375 85.23 ;
      RECT 113.485 86.68 114.015 86.85 ;
      RECT 113.645 86.85 113.815 87.055 ;
      RECT 113.645 84.345 113.815 86.68 ;
      RECT 122.12 87 123.13 87.17 ;
      RECT 122.305 85.34 122.955 87 ;
      RECT 120.83 87 121.84 87.17 ;
      RECT 121.02 86.58 121.67 87 ;
      RECT 121.315 84.74 121.67 86.58 ;
      RECT 121.14 84.57 121.67 84.74 ;
      RECT 124.07 87.005 127.84 87.175 ;
      RECT 124.11 87 127.84 87.005 ;
      RECT 121.1 83.09 121.77 83.49 ;
      RECT 123.515 86.58 124.045 86.75 ;
      RECT 123.725 86.75 123.895 86.78 ;
      RECT 123.725 85.77 123.895 86.58 ;
      RECT 101.805 90.46 123.885 90.7 ;
      RECT 122.84 89.69 133.305 89.87 ;
      RECT 122.84 90.11 123.885 90.46 ;
      RECT 122.84 88.61 123.635 89.69 ;
      RECT 122.84 89.87 143.765 90.11 ;
      RECT 120.615 85.34 121.145 85.51 ;
      RECT 120.615 85.51 120.785 86.78 ;
      RECT 120.615 84.07 120.785 85.34 ;
      RECT 121.895 84.07 122.065 86.78 ;
      RECT 122.815 84.97 123.345 85.14 ;
      RECT 123.175 85.14 123.345 86.78 ;
      RECT 123.175 84.07 123.345 84.97 ;
      RECT 121.405 88.075 124.8 88.36 ;
      RECT 102.785 89.285 122.6 89.455 ;
      RECT 123.895 89.285 143.69 89.455 ;
      RECT 121.405 88.36 122.11 89.285 ;
      RECT 124.135 88.36 124.8 89.285 ;
      RECT 119.115 85.34 119.645 85.51 ;
      RECT 119.285 85.51 119.455 86.78 ;
      RECT 119.285 84.07 119.455 85.34 ;
      RECT 127.195 81.805 128.515 81.94 ;
      RECT 127.195 81.335 128.545 81.805 ;
      RECT 129.865 85.15 130.875 85.32 ;
      RECT 128.29 87.005 132.06 87.175 ;
      RECT 128.305 87 132.035 87.005 ;
      RECT 126.27 85.15 127.96 85.32 ;
      RECT 124.84 81.49 125.73 81.51 ;
      RECT 125.12 81.32 125.79 81.34 ;
      RECT 124.84 81.34 125.79 81.49 ;
      RECT 128.695 81.95 128.865 84.85 ;
      RECT 124.555 81.95 124.725 84.85 ;
      RECT 129.385 81.335 130.055 81.57 ;
      RECT 127.845 84.07 128.375 84.24 ;
      RECT 128.205 84.24 128.375 84.93 ;
      RECT 128.205 82.22 128.375 84.07 ;
      RECT 125.865 82.2 126.035 84.93 ;
      RECT 125.085 84.07 125.615 84.24 ;
      RECT 125.085 84.24 125.255 84.93 ;
      RECT 125.085 82.22 125.255 84.07 ;
      RECT 129.445 83.29 130.055 83.46 ;
      RECT 129.445 83.46 129.615 84.93 ;
      RECT 129.445 82.22 129.615 83.29 ;
      RECT 127.425 82.2 127.595 84.93 ;
      RECT 128.005 85.77 128.175 86.78 ;
      RECT 133.835 85.15 135.185 85.32 ;
      RECT 131.465 81.335 132.475 81.505 ;
      RECT 131.89 81.19 132.475 81.335 ;
      RECT 131.89 81.02 132.42 81.19 ;
      RECT 131.33 85.15 132.34 85.32 ;
      RECT 133.79 81.03 134.8 81.545 ;
      RECT 132.765 85.76 132.935 85.77 ;
      RECT 132.285 85.77 132.935 86.78 ;
      RECT 133.055 81.95 133.225 84.85 ;
      RECT 135.62 81.325 136.29 81.57 ;
      RECT 132.87 81.33 133.54 81.5 ;
      RECT 132.125 83.29 132.735 83.46 ;
      RECT 132.565 83.46 132.735 84.93 ;
      RECT 132.565 82.22 132.735 83.29 ;
      RECT 130.825 83.29 131.355 83.46 ;
      RECT 131.005 83.46 131.175 84.93 ;
      RECT 131.005 82.22 131.175 83.29 ;
      RECT 134.775 83.3 135.475 83.47 ;
      RECT 135.305 83.47 135.475 84.93 ;
      RECT 135.305 82.22 135.475 83.3 ;
      RECT 49.075 85.54 52.845 95.92 ;
      RECT 43.53 85.37 47.53 85.54 ;
      RECT 43.53 95.92 47.53 96.09 ;
      RECT 43.645 85.54 47.415 95.92 ;
      RECT 50.905 82.39 51.435 82.56 ;
      RECT 59.765 81.61 60.575 81.78 ;
      RECT 59.925 81.18 60.455 81.61 ;
      RECT 58.485 81.61 59.295 81.78 ;
      RECT 58.645 81.18 59.175 81.61 ;
      RECT 57.205 81.61 58.015 81.78 ;
      RECT 57.365 81.18 57.895 81.61 ;
      RECT 55.925 81.61 56.735 81.78 ;
      RECT 56.085 81.18 56.615 81.61 ;
      RECT 57.62 85.37 61.62 85.54 ;
      RECT 57.62 95.92 61.62 96.09 ;
      RECT 57.735 85.54 61.505 95.92 ;
      RECT 56.715 95.62 56.885 95.73 ;
      RECT 56.675 88.5 57.565 93.375 ;
      RECT 56.715 93.375 57.565 95.62 ;
      RECT 56.715 85.71 57.565 88.5 ;
      RECT 62.325 81.61 63.135 81.78 ;
      RECT 62.485 81.18 63.015 81.61 ;
      RECT 61.045 81.61 61.855 81.78 ;
      RECT 61.205 81.18 61.735 81.61 ;
      RECT 64.885 81.61 65.695 81.78 ;
      RECT 65.045 81.18 65.575 81.61 ;
      RECT 63.605 81.61 64.415 81.78 ;
      RECT 63.765 81.18 64.295 81.61 ;
      RECT 66.165 81.61 66.975 81.78 ;
      RECT 66.325 81.18 66.855 81.61 ;
      RECT 63.05 85.37 67.05 85.54 ;
      RECT 63.05 95.92 67.05 96.09 ;
      RECT 63.165 85.54 66.935 95.92 ;
      RECT 61.675 85.71 62.995 95.62 ;
      RECT 68.725 81.61 69.535 81.78 ;
      RECT 68.885 81.18 69.415 81.61 ;
      RECT 67.445 81.61 68.255 81.78 ;
      RECT 67.605 81.18 68.135 81.61 ;
      RECT 71.285 81.61 72.095 81.78 ;
      RECT 71.445 81.18 71.975 81.61 ;
      RECT 70.005 81.61 70.815 81.78 ;
      RECT 70.165 81.18 70.695 81.61 ;
      RECT 67.33 85.37 71.33 85.54 ;
      RECT 67.33 95.92 71.33 96.09 ;
      RECT 67.445 85.54 71.215 95.92 ;
      RECT 67.105 85.71 67.275 95.56 ;
      RECT 71.385 85.71 72.705 95.62 ;
      RECT 73.845 81.61 74.655 81.78 ;
      RECT 74.005 81.18 74.535 81.61 ;
      RECT 72.565 81.61 73.375 81.78 ;
      RECT 72.725 81.18 73.255 81.61 ;
      RECT 77.685 81.61 78.495 81.78 ;
      RECT 77.845 81.18 78.375 81.61 ;
      RECT 76.405 81.61 77.215 81.78 ;
      RECT 76.565 81.18 77.095 81.61 ;
      RECT 75.125 81.61 75.935 81.78 ;
      RECT 75.285 81.18 75.815 81.61 ;
      RECT 72.76 85.37 76.76 85.54 ;
      RECT 72.76 95.92 76.76 96.09 ;
      RECT 72.875 85.54 76.645 95.92 ;
      RECT 77.495 95.62 77.665 95.73 ;
      RECT 76.815 88.5 77.705 93.375 ;
      RECT 76.815 93.375 77.665 95.62 ;
      RECT 76.815 85.71 77.665 88.5 ;
      RECT 78.965 81.61 79.775 81.78 ;
      RECT 79.125 81.18 79.655 81.61 ;
      RECT 82.805 81.61 83.615 81.78 ;
      RECT 82.965 81.18 83.495 81.61 ;
      RECT 81.525 81.61 82.335 81.78 ;
      RECT 81.685 81.18 82.215 81.61 ;
      RECT 80.245 81.61 81.055 81.78 ;
      RECT 80.405 81.18 80.935 81.61 ;
      RECT 81 85.71 81.17 95.56 ;
      RECT 80.42 85.73 80.59 96.45 ;
      RECT 73.13 98.39 87.79 98.56 ;
      RECT 79.72 97.225 87.79 97.815 ;
      RECT 80.42 97.815 87.79 98.39 ;
      RECT 86.02 88.08 86.19 88.52 ;
      RECT 86.02 87.85 86.19 87.91 ;
      RECT 80.42 96.45 87.79 97.225 ;
      RECT 86.02 87.91 87.79 88.08 ;
      RECT 86.48 89.97 87.79 90.14 ;
      RECT 87.62 90.14 87.79 96.45 ;
      RECT 87.62 88.08 87.79 89.97 ;
      RECT 86.26 87.36 87.79 87.53 ;
      RECT 87.62 87.53 87.79 87.91 ;
      RECT 87.62 86.04 87.79 87.36 ;
      RECT 81.225 85.37 85.225 85.54 ;
      RECT 81.225 95.92 85.225 96.09 ;
      RECT 81.34 85.54 85.11 95.92 ;
      RECT 84.085 81.61 84.895 81.78 ;
      RECT 86.26 86.08 87.28 86.25 ;
      RECT 88.19 82.265 90.21 83.015 ;
      RECT 85.28 85.71 85.45 95.56 ;
      RECT 84.225 82.615 84.755 82.785 ;
      RECT 85.89 86.305 86.06 87.305 ;
      RECT 100.23 85.03 100.815 85.2 ;
      RECT 100.645 85.2 100.815 85.935 ;
      RECT 100.645 84.925 100.815 85.03 ;
      RECT 100.13 83.09 100.305 83.945 ;
      RECT 100.13 83.945 100.3 84.01 ;
      RECT 100.13 83 100.3 83.09 ;
      RECT 100.44 88.205 102.66 88.425 ;
      RECT 101.01 83 101.18 84.01 ;
      RECT 100.775 84.535 101.445 84.705 ;
      RECT 100.915 84.705 101.445 84.735 ;
      RECT 104.85 83.755 105.02 85.105 ;
      RECT 105.96 83.815 106.36 86.825 ;
      RECT 106.13 83.755 106.3 83.815 ;
      RECT 101.89 81.435 102.06 81.965 ;
      RECT 104.78 85.74 104.95 86.825 ;
      RECT 101.425 84.925 101.595 85.935 ;
      RECT 101.89 83 102.06 84.335 ;
      RECT 102.56 88.725 103.115 88.895 ;
      RECT 102.56 88.895 102.73 88.94 ;
      RECT 102.56 88.61 102.73 88.725 ;
      RECT 102.62 83.765 102.79 86.475 ;
      RECT 104.18 83.765 104.35 86.475 ;
      RECT 102.24 82.81 102.44 86.995 ;
      RECT 102.255 86.995 102.425 87.34 ;
      RECT 101.475 82.14 102.44 82.81 ;
      RECT 105.075 83.365 106.075 83.535 ;
      RECT 105.135 83.535 106.015 83.625 ;
      RECT 105.005 87.015 106.925 87.21 ;
      RECT 105.005 87.21 106.005 87.215 ;
      RECT 106.59 83.8 107.18 83.97 ;
      RECT 106.59 83.97 106.925 87.015 ;
      RECT 458.635 74.8 459.145 75.13 ;
      RECT 458.725 75.13 459.095 77.85 ;
      RECT 453.395 77.85 459.095 78.22 ;
      RECT 457.755 74.8 458.265 75.13 ;
      RECT 457.825 73.325 458.195 74.8 ;
      RECT 457.825 73.155 458.355 73.325 ;
      RECT 457.485 73.58 457.655 74.63 ;
      RECT 458.365 73.62 458.535 74.63 ;
      RECT 459.245 73.325 459.415 74.63 ;
      RECT 458.885 73.155 459.415 73.325 ;
      RECT 455.145 80.565 455.705 80.885 ;
      RECT 455.35 80.885 455.52 85.285 ;
      RECT 455.35 80.535 455.52 80.565 ;
      RECT 455.94 81.145 456.475 81.465 ;
      RECT 456.13 81.465 456.3 85.285 ;
      RECT 456.13 80.535 456.3 81.145 ;
      RECT 454.415 81.725 454.98 82.045 ;
      RECT 454.57 82.045 454.74 85.285 ;
      RECT 454.57 80.535 454.74 81.725 ;
      RECT 457.03 79.855 457.655 80.025 ;
      RECT 457.03 79.825 457.2 79.855 ;
      RECT 457.03 85.005 457.655 86.015 ;
      RECT 457.03 80.025 457.2 85.005 ;
      RECT 459.645 79.325 460.175 79.495 ;
      RECT 459.805 79.495 460.175 86.185 ;
      RECT 459.805 79.32 460.175 79.325 ;
      RECT 458.635 86.185 460.175 86.515 ;
      RECT 455.575 79.855 456.245 80.025 ;
      RECT 455.575 77.345 456.245 77.515 ;
      RECT 454.625 79.855 455.295 80.025 ;
      RECT 454.625 77.345 455.295 77.515 ;
      RECT 462.425 79.855 462.955 80.025 ;
      RECT 462.425 80.025 462.935 80.105 ;
      RECT 462.425 79.775 462.935 79.855 ;
      RECT 461.545 79.775 462.055 80.105 ;
      RECT 461.615 84.44 462.145 84.61 ;
      RECT 461.615 80.105 461.985 84.44 ;
      RECT 462.425 77.345 462.955 77.515 ;
      RECT 462.425 77.515 462.935 77.595 ;
      RECT 462.425 77.265 462.935 77.345 ;
      RECT 463.035 84.44 463.565 84.61 ;
      RECT 463.035 80.27 463.205 84.44 ;
      RECT 462.155 80.575 462.325 83.285 ;
      RECT 461.18 80.27 461.445 83.285 ;
      RECT 461.18 79.755 461.35 80.27 ;
      RECT 462.155 74.085 462.325 76.795 ;
      RECT 461.18 74.085 461.445 77.1 ;
      RECT 461.18 77.1 461.35 77.615 ;
      RECT 467.555 79.775 468.065 80.105 ;
      RECT 467.625 80.105 467.995 84.1 ;
      RECT 468.435 79.855 468.945 80.105 ;
      RECT 468.415 78.815 468.945 79.855 ;
      RECT 467.555 77.265 468.065 77.595 ;
      RECT 467.625 73.27 467.995 77.265 ;
      RECT 468.435 77.265 468.945 77.515 ;
      RECT 468.415 77.515 468.945 78.555 ;
      RECT 469.485 81.145 470.045 81.465 ;
      RECT 469.65 81.465 469.82 85.285 ;
      RECT 469.65 80.535 469.82 81.145 ;
      RECT 471.21 80.535 471.38 85.285 ;
      RECT 466.925 83.65 467.455 83.82 ;
      RECT 466.845 79.855 467.375 80.025 ;
      RECT 467.205 80.27 467.455 83.65 ;
      RECT 467.205 80.025 467.375 80.27 ;
      RECT 468.165 80.385 468.615 84.375 ;
      RECT 467.245 84.375 469.1 84.625 ;
      RECT 468.85 84.625 469.1 85.635 ;
      RECT 468.85 85.635 471.42 85.885 ;
      RECT 469.045 80.27 469.215 84.1 ;
      RECT 466.925 73.55 467.455 73.72 ;
      RECT 466.845 77.345 467.375 77.515 ;
      RECT 467.205 73.72 467.455 77.1 ;
      RECT 467.205 77.1 467.375 77.345 ;
      RECT 469.045 73.27 469.215 77.1 ;
      RECT 470.2 80.565 470.76 80.885 ;
      RECT 470.43 80.885 470.6 85.285 ;
      RECT 470.43 80.535 470.6 80.565 ;
      RECT 470.655 79.855 471.325 80.025 ;
      RECT 470.735 78.815 471.265 79.855 ;
      RECT 470.655 77.345 471.325 77.515 ;
      RECT 470.735 77.515 471.265 78.555 ;
      RECT 469.705 79.855 470.375 80.025 ;
      RECT 469.705 77.345 470.375 77.515 ;
      RECT 19.33 88.31 19.53 93.725 ;
      RECT 19.33 93.725 19.5 94.355 ;
      RECT 19.33 87.565 19.5 88.31 ;
      RECT 18.85 84.375 28.26 84.545 ;
      RECT 18.85 84.545 24.18 86.19 ;
      RECT 28.09 84.545 28.26 103.825 ;
      RECT 28.09 133.1 28.26 133.775 ;
      RECT 18.85 104.255 20.19 107.995 ;
      RECT 19.93 127.905 26.295 127.935 ;
      RECT 19.93 125.185 26.295 125.215 ;
      RECT 26.065 127.04 28.29 127.705 ;
      RECT 26.065 125.415 28.29 126.035 ;
      RECT 26.56 107.09 28.285 107.84 ;
      RECT 28.09 107.84 28.285 108.45 ;
      RECT 18.85 125.415 20.16 127.705 ;
      RECT 28.09 105.115 28.285 107.09 ;
      RECT 26.56 104.365 28.285 105.115 ;
      RECT 28.09 103.825 28.285 104.365 ;
      RECT 28.09 117.4 28.29 125.365 ;
      RECT 28.09 108.45 28.26 117.4 ;
      RECT 18.85 86.19 19.02 104.255 ;
      RECT 26.095 126.035 28.29 127.04 ;
      RECT 18.85 127.705 28.29 127.755 ;
      RECT 18.85 125.365 28.29 125.415 ;
      RECT 18.85 127.905 19.02 133.775 ;
      RECT 18.85 127.755 26.295 127.905 ;
      RECT 18.85 107.995 19.02 125.215 ;
      RECT 18.85 125.215 26.295 125.365 ;
      RECT 18.85 133.775 28.26 133.945 ;
      RECT 28.09 127.755 28.29 133.1 ;
      RECT 24.8 85.175 27.51 85.345 ;
      RECT 24.8 86.455 27.51 86.625 ;
      RECT 27.61 87.565 27.78 94.355 ;
      RECT 27.73 85.42 27.9 86.4 ;
      RECT 33.82 85.37 37.82 85.54 ;
      RECT 33.82 95.92 37.82 96.09 ;
      RECT 33.935 85.54 37.705 95.92 ;
      RECT 39.25 85.37 43.25 85.54 ;
      RECT 39.25 95.92 43.25 96.09 ;
      RECT 39.365 85.54 43.135 95.92 ;
      RECT 43.465 81.61 44.175 81.78 ;
      RECT 43.85 80.88 44.02 81.61 ;
      RECT 48.76 85.37 52.96 85.54 ;
      RECT 48.76 95.92 52.96 96.09 ;
      RECT 336.025 77.05 336.205 80.46 ;
      RECT 336.035 80.46 336.205 81.15 ;
      RECT 336.035 76.4 336.205 77.05 ;
      RECT 336.375 80.75 336.645 81.32 ;
      RECT 337.155 80.75 337.425 81.32 ;
      RECT 337.935 80.75 338.205 81.32 ;
      RECT 338.715 81.315 339.1 81.32 ;
      RECT 338.715 80.75 338.985 81.315 ;
      RECT 336.26 81.32 339.1 81.78 ;
      RECT 338.375 76.4 338.545 81.15 ;
      RECT 336.815 76.4 336.985 81.15 ;
      RECT 337.595 76.4 337.765 81.15 ;
      RECT 332.925 76.4 333.095 81.15 ;
      RECT 343.03 77.05 343.23 80.86 ;
      RECT 343.045 80.86 343.215 81.15 ;
      RECT 343.045 76.4 343.215 77.05 ;
      RECT 340.47 77.05 340.67 80.86 ;
      RECT 340.485 80.86 340.655 81.15 ;
      RECT 340.485 76.4 340.655 77.05 ;
      RECT 339.69 77.05 339.89 80.86 ;
      RECT 339.705 76.4 339.875 77.05 ;
      RECT 339.705 81.61 340.43 81.78 ;
      RECT 339.705 80.86 339.875 81.61 ;
      RECT 341.75 77.11 341.95 80.92 ;
      RECT 340.71 81.555 345.55 81.835 ;
      RECT 344.31 77.11 344.51 80.92 ;
      RECT 341.765 76.4 341.935 77.11 ;
      RECT 344.325 76.4 344.495 77.11 ;
      RECT 341.765 80.92 341.935 81.555 ;
      RECT 344.325 80.92 344.495 81.555 ;
      RECT 339.155 76.4 339.325 81.15 ;
      RECT 345.57 77.05 345.775 80.25 ;
      RECT 345.605 76.4 345.775 77.05 ;
      RECT 345.605 80.25 345.775 81.15 ;
      RECT 346.37 77.11 346.57 80.65 ;
      RECT 346.385 80.65 346.555 81.15 ;
      RECT 346.385 76.4 346.555 77.11 ;
      RECT 352.18 74.405 352.35 79.155 ;
      RECT 353.46 74.405 353.63 79.155 ;
      RECT 353.94 74.155 354.11 80.16 ;
      RECT 351.7 74.155 351.87 80.16 ;
      RECT 351.7 73.985 354.11 74.155 ;
      RECT 351.7 80.16 354.11 80.36 ;
      RECT 352.475 79.665 353.285 79.835 ;
      RECT 354.675 76.64 356.795 78.76 ;
      RECT 354.675 73.725 355.955 76.64 ;
      RECT 355.105 79.595 366.875 82.42 ;
      RECT 354.675 79.19 366.875 79.595 ;
      RECT 354.675 78.93 366.815 79.19 ;
      RECT 366.705 76.64 366.875 78.76 ;
      RECT 354.675 78.76 366.875 78.93 ;
      RECT 359.455 78.35 361.485 78.52 ;
      RECT 361.015 77.07 361.185 78.35 ;
      RECT 358.825 75.82 360.875 75.99 ;
      RECT 360.705 75.12 360.875 75.82 ;
      RECT 359.105 76.62 359.275 77.97 ;
      RECT 358.485 74.59 358.655 77.66 ;
      RECT 357.205 76.65 357.375 77.66 ;
      RECT 357.205 74.59 357.375 75.6 ;
      RECT 359.765 74.59 359.935 75.6 ;
      RECT 360.265 74.59 361.215 74.76 ;
      RECT 361.045 75.99 361.215 76.62 ;
      RECT 361.045 75.82 362.115 75.99 ;
      RECT 361.045 74.76 361.215 75.82 ;
      RECT 360.385 76.79 360.555 77.97 ;
      RECT 360.385 76.62 361.215 76.79 ;
      RECT 356.625 74.08 356.795 75.58 ;
      RECT 366.705 74.08 366.875 75.58 ;
      RECT 356.625 73.91 366.875 74.08 ;
      RECT 361.645 74.08 361.815 75.58 ;
      RECT 361.665 76.62 361.835 77.97 ;
      RECT 362.015 78.35 364.045 78.52 ;
      RECT 362.315 77.07 362.485 78.35 ;
      RECT 362.645 75.82 364.675 75.99 ;
      RECT 364.225 76.62 364.395 77.97 ;
      RECT 364.845 74.59 365.015 77.66 ;
      RECT 366.125 76.65 366.295 77.66 ;
      RECT 363.565 74.59 363.735 75.6 ;
      RECT 366.125 74.59 366.295 75.6 ;
      RECT 362.285 74.59 363.235 74.76 ;
      RECT 362.285 74.56 362.455 74.59 ;
      RECT 362.285 74.76 362.455 75.12 ;
      RECT 362.285 75.65 362.455 76.62 ;
      RECT 362.945 76.79 363.115 77.97 ;
      RECT 362.285 76.62 363.115 76.79 ;
      RECT 361.985 75.12 362.455 75.65 ;
      RECT 367.485 80.16 369.875 80.33 ;
      RECT 367.485 73.91 369.875 74.08 ;
      RECT 369.705 74.08 369.875 80.16 ;
      RECT 367.485 74.08 367.655 80.16 ;
      RECT 367.825 79.69 369.05 79.86 ;
      RECT 368.065 74.51 368.235 79.47 ;
      RECT 369.125 74.51 369.295 79.47 ;
      RECT 368.595 74.72 368.765 79.47 ;
      RECT 400.46 75.235 401.47 75.405 ;
      RECT 401.64 75.235 404.57 75.415 ;
      RECT 404.74 75.235 405.75 75.405 ;
      RECT 405.92 75.235 408.85 75.415 ;
      RECT 409.02 75.235 410.03 75.405 ;
      RECT 417.9 75.235 418.91 75.405 ;
      RECT 414.62 75.235 415.63 75.405 ;
      RECT 419.08 75.235 420.01 75.415 ;
      RECT 415.8 75.235 417.73 75.415 ;
      RECT 422.46 75.235 423.47 75.405 ;
      RECT 420.18 75.235 421.19 75.405 ;
      RECT 421.36 75.235 422.29 75.415 ;
      RECT 430.48 77.95 430.81 78.64 ;
      RECT 429.71 77.95 430.04 78.64 ;
      RECT 436.31 77.95 436.64 78.64 ;
      RECT 434.33 77.95 434.66 78.64 ;
      RECT 431.25 77.95 433.89 78.64 ;
      RECT 435.1 77.95 435.43 78.64 ;
      RECT 437.85 77.95 440.49 78.64 ;
      RECT 437.08 77.95 437.41 78.64 ;
      RECT 440.93 77.95 441.26 78.64 ;
      RECT 441.7 77.95 442.03 78.64 ;
      RECT 453.17 80.535 453.34 85.285 ;
      RECT 453.755 80.565 454.315 80.885 ;
      RECT 453.95 80.885 454.12 85.285 ;
      RECT 453.95 80.535 454.12 80.565 ;
      RECT 453.395 79.52 453.765 79.855 ;
      RECT 453.24 79.855 453.91 80.025 ;
      RECT 458.635 82.24 459.145 82.57 ;
      RECT 458.725 79.52 459.095 82.24 ;
      RECT 453.395 79.15 459.095 79.52 ;
      RECT 453.395 77.515 453.765 77.85 ;
      RECT 453.24 77.345 453.91 77.515 ;
      RECT 288.17 80.16 290.32 80.405 ;
      RECT 289.905 80.405 290.32 82.14 ;
      RECT 290.055 82.81 290.32 86.93 ;
      RECT 288.355 86.93 290.32 87.285 ;
      RECT 289.29 82.14 290.32 82.81 ;
      RECT 214.085 252.535 348.425 253.385 ;
      RECT 347.575 249.375 348.425 252.535 ;
      RECT 347.575 248.525 364.855 249.375 ;
      RECT 223.105 244.045 223.955 252.535 ;
      RECT 214.085 244.045 215.845 252.535 ;
      RECT 214.085 243.195 223.955 244.045 ;
      RECT 364.005 226.45 364.855 248.525 ;
      RECT 347.575 226.44 348.425 248.525 ;
      RECT 364.005 226.44 371.14 226.45 ;
      RECT 347.575 225.59 371.14 226.44 ;
      RECT 347.575 215.97 348.425 225.59 ;
      RECT 344.63 215.53 348.425 215.97 ;
      RECT 370.28 204.335 371.14 225.59 ;
      RECT 344.485 204.335 348.425 215.53 ;
      RECT 344.485 203.475 371.14 204.335 ;
      RECT 344.485 200.645 348.425 203.475 ;
      RECT 214.085 195.155 216.005 243.195 ;
      RECT 214.085 194.305 227.965 195.155 ;
      RECT 345.47 184.19 348.425 200.645 ;
      RECT 345.47 177.45 346.32 184.19 ;
      RECT 299.78 176.6 346.32 177.45 ;
      RECT 227.115 176.145 227.965 194.305 ;
      RECT 299.78 176.145 300.63 176.6 ;
      RECT 214.085 174.305 214.985 194.305 ;
      RECT 199.68 173.235 214.985 174.305 ;
      RECT 227.115 173.235 300.63 176.145 ;
      RECT 199.68 168.145 300.63 173.235 ;
      RECT 327.41 160.22 328.26 176.6 ;
      RECT 299.78 160 300.63 168.145 ;
      RECT 301.865 160 351.405 160.22 ;
      RECT 299.78 159.15 351.405 160 ;
      RECT 339.815 157.925 340.665 159.15 ;
      RECT 350.555 154.015 351.405 159.15 ;
      RECT 339.81 152.475 340.7 157.925 ;
      RECT 350.535 152.35 351.425 154.015 ;
      RECT 350.555 151.61 351.405 152.35 ;
      RECT 339.815 151.055 340.665 152.475 ;
      RECT 350.535 150.57 351.425 151.61 ;
      RECT 350.555 149.94 351.405 150.57 ;
      RECT 339.81 148.365 340.7 151.055 ;
      RECT 350.535 148.365 351.425 149.94 ;
      RECT 350.555 147.6 351.405 148.365 ;
      RECT 339.815 147.135 340.665 148.365 ;
      RECT 350.535 147.07 351.425 147.6 ;
      RECT 339.81 146.79 340.7 147.135 ;
      RECT 350.555 145.1 351.405 147.07 ;
      RECT 299.78 143.905 302.715 159.15 ;
      RECT 339.815 143.905 340.665 146.79 ;
      RECT 350.555 143.885 358.295 145.1 ;
      RECT 299.78 143.735 340.665 143.905 ;
      RECT 357.445 128.205 358.295 143.885 ;
      RECT 299.78 128.205 300.97 143.735 ;
      RECT 340.015 128.205 340.665 143.735 ;
      RECT 299.78 127.885 358.6 128.205 ;
      RECT 310.83 115.675 311 127.885 ;
      RECT 334.63 115.675 334.8 127.885 ;
      RECT 358.43 115.675 358.6 127.885 ;
      RECT 310.83 115.375 358.6 115.675 ;
      RECT 199.68 109.585 200.53 168.145 ;
      RECT 299.78 109.585 300.97 127.885 ;
      RECT 199.68 108.735 300.97 109.585 ;
      RECT 223.95 108.38 271.97 108.735 ;
      RECT 358.43 106.36 358.6 115.375 ;
      RECT 318.25 106.36 318.42 115.375 ;
      RECT 318.25 106.16 358.6 106.36 ;
      RECT 268.86 103.77 271.97 108.38 ;
      RECT 223.95 103.77 236.175 108.38 ;
      RECT 249.64 103.77 249.81 108.38 ;
      RECT 223.95 102.92 271.97 103.77 ;
      RECT 199.73 101.9 212.41 108.735 ;
      RECT 215.275 101.9 216.125 108.735 ;
      RECT 318.25 97.145 318.42 106.16 ;
      RECT 358.43 97.145 358.6 106.16 ;
      RECT 199.73 97.095 216.125 101.9 ;
      RECT 199.735 97.045 216.125 97.095 ;
      RECT 223.95 97.045 235.725 102.92 ;
      RECT 199.735 96.88 235.725 97.045 ;
      RECT 310.83 96.855 358.6 97.145 ;
      RECT 199.735 95.985 215.7 95.995 ;
      RECT 199.735 95.995 215.825 96.03 ;
      RECT 216.125 95.995 222.875 96.03 ;
      RECT 199.73 96.03 235.725 96.88 ;
      RECT 300.8 84.825 300.97 108.735 ;
      RECT 310.83 84.825 311 96.855 ;
      RECT 334.63 84.825 334.8 96.855 ;
      RECT 358.43 84.825 358.6 96.855 ;
      RECT 300.8 83.975 358.6 84.825 ;
      RECT 302.285 82.955 348.75 83.975 ;
      RECT 302.285 75.12 303.575 82.955 ;
      RECT 347.895 75.12 348.75 82.955 ;
      RECT 302.285 74.465 348.75 75.12 ;
      RECT 308.605 76.4 308.775 81.15 ;
      RECT 306.045 76.4 306.215 81.15 ;
      RECT 304.765 76.4 304.935 81.15 ;
      RECT 304.185 76.05 304.355 82.02 ;
      RECT 346.95 77.11 347.15 80.65 ;
      RECT 304.185 75.88 347.135 76.05 ;
      RECT 346.965 80.65 347.135 82.02 ;
      RECT 346.965 76.05 347.135 77.11 ;
      RECT 304.185 82.02 347.135 82.19 ;
      RECT 307.325 76.4 307.495 81.15 ;
      RECT 313.725 76.4 313.895 81.15 ;
      RECT 311.165 76.4 311.335 81.15 ;
      RECT 315.005 76.4 315.175 81.15 ;
      RECT 312.445 76.4 312.615 81.15 ;
      RECT 309.885 76.4 310.055 81.15 ;
      RECT 316.285 76.4 316.455 81.15 ;
      RECT 318.845 76.4 319.015 81.15 ;
      RECT 320.125 76.4 320.295 81.15 ;
      RECT 317.565 76.4 317.735 81.15 ;
      RECT 326.525 76.4 326.695 81.15 ;
      RECT 323.965 76.4 324.135 81.15 ;
      RECT 321.405 76.4 321.575 81.15 ;
      RECT 325.245 76.4 325.415 81.15 ;
      RECT 322.685 76.4 322.855 81.15 ;
      RECT 331.645 76.4 331.815 81.15 ;
      RECT 329.085 76.4 329.255 81.15 ;
      RECT 327.805 76.4 327.975 81.15 ;
      RECT 330.365 76.4 330.535 81.15 ;
      RECT 334.205 76.4 334.375 81.15 ;
      RECT 334.55 81.61 335.655 81.78 ;
      RECT 335.485 76.4 335.655 81.61 ;
      RECT 254.945 77.7 255.615 77.87 ;
      RECT 261.46 77.68 262.81 77.85 ;
      RECT 257.61 76.42 261.01 76.59 ;
      RECT 260.84 76.59 261.01 77.155 ;
      RECT 257.91 76.37 260.24 76.42 ;
      RECT 261.97 75.16 262.5 75.33 ;
      RECT 262.06 75.33 262.39 75.69 ;
      RECT 262.835 75.16 263.365 75.33 ;
      RECT 262.94 75.33 263.27 75.69 ;
      RECT 258.615 80.95 259.78 81.12 ;
      RECT 259.44 84.28 259.97 84.45 ;
      RECT 259.61 84.45 259.78 84.93 ;
      RECT 258.615 78.07 258.785 80.95 ;
      RECT 259.61 81.12 259.78 84.28 ;
      RECT 257.735 78.07 257.905 80.78 ;
      RECT 257.61 77.2 260.32 77.37 ;
      RECT 257.91 77.08 260.24 77.2 ;
      RECT 261.17 79.055 261.87 79.225 ;
      RECT 261.17 79.225 261.34 80.78 ;
      RECT 261.17 78.07 261.34 79.055 ;
      RECT 262.76 79.055 263.29 79.225 ;
      RECT 262.93 79.225 263.1 80.78 ;
      RECT 262.93 78.07 263.1 79.055 ;
      RECT 259.495 78.07 259.665 80.78 ;
      RECT 259.66 74.79 260.25 74.96 ;
      RECT 260.08 74.96 260.25 75.77 ;
      RECT 260.08 74.76 260.25 74.79 ;
      RECT 261.63 76.22 261.8 77.36 ;
      RECT 257.86 77.68 258.53 77.85 ;
      RECT 258.86 77.68 259.53 77.85 ;
      RECT 260.145 78.09 260.695 81.09 ;
      RECT 258.8 75.18 259.34 75.35 ;
      RECT 258.8 74.76 258.97 75.18 ;
      RECT 258.8 75.35 258.97 75.77 ;
      RECT 262.05 80.95 263.36 81.165 ;
      RECT 262.96 84.07 263.49 84.24 ;
      RECT 263.19 84.24 263.36 84.93 ;
      RECT 262.05 78.07 262.22 80.95 ;
      RECT 263.19 81.165 263.36 84.07 ;
      RECT 263.22 77.68 264.57 77.85 ;
      RECT 268.08 81.77 268.61 81.94 ;
      RECT 268.08 81.94 268.25 82.87 ;
      RECT 268.08 78.12 268.25 81.77 ;
      RECT 268.96 78.12 269.13 82.87 ;
      RECT 265.28 78.13 265.45 81.05 ;
      RECT 264.16 79.055 264.86 79.225 ;
      RECT 264.69 79.225 264.86 80.78 ;
      RECT 264.69 78.07 264.86 79.055 ;
      RECT 263.53 76.22 263.7 77.36 ;
      RECT 263.81 78.07 263.98 80.78 ;
      RECT 273.2 79.09 277.95 79.26 ;
      RECT 271.24 81.77 271.77 81.94 ;
      RECT 271.6 81.94 271.77 82.87 ;
      RECT 271.6 78.12 271.77 81.77 ;
      RECT 273.29 77.08 273.82 77.25 ;
      RECT 273.29 77.25 273.46 77.475 ;
      RECT 273.29 74.765 273.46 77.08 ;
      RECT 274.32 79.965 278.09 79.97 ;
      RECT 273.2 79.97 278.09 80.135 ;
      RECT 273.2 80.135 277.95 80.14 ;
      RECT 270.72 78.12 270.89 82.87 ;
      RECT 269.67 81.77 270.2 81.94 ;
      RECT 269.84 81.94 270.01 82.87 ;
      RECT 269.84 78.12 270.01 81.77 ;
      RECT 279.545 74.405 280.555 74.575 ;
      RECT 279.66 74.575 279.83 75.69 ;
      RECT 280.34 74.575 280.51 75.69 ;
      RECT 277.82 74.405 278.95 74.575 ;
      RECT 277.9 74.575 278.07 75.69 ;
      RECT 278.78 74.575 278.95 75.69 ;
      RECT 275.18 73.865 276.19 74.035 ;
      RECT 275.24 73.6 276.13 73.865 ;
      RECT 279.245 79.265 282.145 79.435 ;
      RECT 279.245 80.045 281.955 80.215 ;
      RECT 276.45 77.08 276.98 77.25 ;
      RECT 276.81 77.25 276.98 77.475 ;
      RECT 276.81 74.765 276.98 77.08 ;
      RECT 279.82 77.08 280.35 77.25 ;
      RECT 280 77.25 280.17 77.475 ;
      RECT 280 74.765 280.17 77.08 ;
      RECT 278.06 77.08 278.59 77.25 ;
      RECT 278.24 77.25 278.41 77.475 ;
      RECT 278.24 74.765 278.41 77.08 ;
      RECT 274.87 77.08 275.4 77.25 ;
      RECT 275.05 77.25 275.22 77.475 ;
      RECT 275.05 74.765 275.22 77.08 ;
      RECT 278.77 83.31 279.3 83.48 ;
      RECT 278.77 81.675 278.995 83.31 ;
      RECT 278.43 79.315 278.995 81.675 ;
      RECT 281.405 74.405 282.415 74.575 ;
      RECT 281.465 74 282.355 74.405 ;
      RECT 281.7 77.08 282.23 77.25 ;
      RECT 281.76 77.25 281.93 77.475 ;
      RECT 281.76 74.765 281.93 77.08 ;
      RECT 284.155 73.865 285.505 74.035 ;
      RECT 284.205 73.6 285.455 73.865 ;
      RECT 285.305 74.405 286.655 74.575 ;
      RECT 285.49 74.575 285.66 75.69 ;
      RECT 286.17 74.575 286.34 75.69 ;
      RECT 283.19 74.765 283.36 77.645 ;
      RECT 283.19 77.645 286.88 77.815 ;
      RECT 284.95 74.765 285.12 77.645 ;
      RECT 286.71 74.765 286.88 77.645 ;
      RECT 285.47 77.08 286 77.25 ;
      RECT 285.83 77.25 286 77.475 ;
      RECT 285.83 74.765 286 77.08 ;
      RECT 282.525 79.26 282.695 79.99 ;
      RECT 282.51 80.27 282.71 82.645 ;
      RECT 282.51 82.645 286.87 82.845 ;
      RECT 283.63 82.845 286.87 82.855 ;
      RECT 283.405 79.755 283.575 82.465 ;
      RECT 284.29 79.525 284.46 79.755 ;
      RECT 284.285 80.54 284.455 82.465 ;
      RECT 284.285 79.755 284.46 80.54 ;
      RECT 285.165 79.755 285.335 82.465 ;
      RECT 286.05 79.525 286.22 79.755 ;
      RECT 286.045 80.54 286.215 82.465 ;
      RECT 286.045 79.755 286.22 80.54 ;
      RECT 288.75 80.615 289.07 81.925 ;
      RECT 288.825 80.595 288.995 80.615 ;
      RECT 287.945 80.595 288.115 81.18 ;
      RECT 287.625 78.89 288.485 79.42 ;
      RECT 287.625 79.42 288.155 79.96 ;
      RECT 289.095 78.83 289.265 79.42 ;
      RECT 286.925 79.755 287.095 82.465 ;
      RECT 290.07 78.225 290.4 79.61 ;
      RECT 288.405 79.61 290.4 79.945 ;
      RECT 237.72 78.41 238.14 78.75 ;
      RECT 237.72 77.4 238.14 78.24 ;
      RECT 238.215 76.37 241.945 76.54 ;
      RECT 239.96 77.4 240.13 78.75 ;
      RECT 239.96 79.54 240.13 81.08 ;
      RECT 238.66 75.1 242.05 75.27 ;
      RECT 241.475 75.27 242.005 75.33 ;
      RECT 238.105 79.12 238.67 79.29 ;
      RECT 238.105 79.29 238.615 79.405 ;
      RECT 238.105 79.075 238.615 79.12 ;
      RECT 234.305 78.35 234.835 78.52 ;
      RECT 234.48 78.52 234.65 78.875 ;
      RECT 234.48 76.165 234.65 78.35 ;
      RECT 243.8 78.95 244.39 79.12 ;
      RECT 243.8 83.29 245.03 83.46 ;
      RECT 243.8 83.46 244.13 83.83 ;
      RECT 243.8 79.12 244.13 83.29 ;
      RECT 244.61 81.92 244.94 83.29 ;
      RECT 242.73 78.95 243.32 79.12 ;
      RECT 242.09 83.29 243.32 83.46 ;
      RECT 242.99 83.46 243.32 83.83 ;
      RECT 242.99 79.12 243.32 83.29 ;
      RECT 242.18 81.92 242.51 83.29 ;
      RECT 243.8 78.24 244.39 78.41 ;
      RECT 243.8 78.41 244.13 78.44 ;
      RECT 243.8 74.92 244.13 78.24 ;
      RECT 242.73 78.24 243.32 78.41 ;
      RECT 242.99 78.41 243.32 78.44 ;
      RECT 242.99 74.92 243.32 78.24 ;
      RECT 244.685 79.73 245.16 81.08 ;
      RECT 244.685 78.75 244.855 79.73 ;
      RECT 244.685 78.24 245.59 78.41 ;
      RECT 244.685 78.41 245.16 78.75 ;
      RECT 244.685 77.4 245.16 78.24 ;
      RECT 241.96 79.73 242.435 81.08 ;
      RECT 242.265 78.75 242.435 79.73 ;
      RECT 241.53 78.24 242.435 78.41 ;
      RECT 241.96 78.41 242.435 78.75 ;
      RECT 241.96 77.4 242.435 78.24 ;
      RECT 245.175 76.37 248.905 76.54 ;
      RECT 244.7 74.4 244.87 74.93 ;
      RECT 244.7 75.43 244.87 76.02 ;
      RECT 242.25 74.4 242.42 74.93 ;
      RECT 242.25 75.43 242.42 76.02 ;
      RECT 245.07 75.1 248.46 75.27 ;
      RECT 245.115 75.27 245.645 75.33 ;
      RECT 245.115 79.11 245.645 79.28 ;
      RECT 245.125 79.28 245.635 79.405 ;
      RECT 245.125 79.075 245.635 79.11 ;
      RECT 241.475 79.11 242.005 79.28 ;
      RECT 241.485 79.28 241.995 79.405 ;
      RECT 241.485 79.075 241.995 79.11 ;
      RECT 249.57 74.4 249.74 81.02 ;
      RECT 250.87 73.83 252.19 74.37 ;
      RECT 250.785 74.37 254.905 74.54 ;
      RECT 248.98 74.42 249.15 76.02 ;
      RECT 251.25 74.79 251.78 74.96 ;
      RECT 251.44 74.96 251.61 75.77 ;
      RECT 251.44 74.76 251.61 74.79 ;
      RECT 245.925 77.01 246.935 77.18 ;
      RECT 246.005 76.895 246.535 77.01 ;
      RECT 247.205 77.01 248.215 77.18 ;
      RECT 247.285 76.895 247.815 77.01 ;
      RECT 246.99 77.4 247.16 78.75 ;
      RECT 246.99 79.54 247.16 81.08 ;
      RECT 248.45 79.12 249.015 79.29 ;
      RECT 248.505 79.29 249.015 79.405 ;
      RECT 248.505 79.075 249.015 79.12 ;
      RECT 249.23 78.75 249.4 79.73 ;
      RECT 248.98 79.73 249.4 81.08 ;
      RECT 248.98 78.41 249.4 78.75 ;
      RECT 248.56 78.24 249.4 78.41 ;
      RECT 248.98 77.4 249.4 78.24 ;
      RECT 251.17 76.42 256.07 76.59 ;
      RECT 252.32 74.76 253.03 75.77 ;
      RECT 252.49 75.77 253.03 76.42 ;
      RECT 255.78 74.54 256.07 76.42 ;
      RECT 255.78 74 259.98 74.54 ;
      RECT 251.17 77.3 256.45 77.48 ;
      RECT 255.92 77.48 256.45 78.01 ;
      RECT 252.835 77.48 253.725 77.62 ;
      RECT 256.24 76.07 256.41 77.3 ;
      RECT 256.24 78.01 256.41 80.82 ;
      RECT 250.74 81.43 251.01 81.6 ;
      RECT 250.67 83.69 251.2 83.86 ;
      RECT 250.74 78.075 250.91 81.43 ;
      RECT 250.84 83.86 251.01 86.93 ;
      RECT 250.84 81.6 251.01 83.69 ;
      RECT 251.62 78.075 251.79 80.785 ;
      RECT 250.865 77.7 251.535 77.87 ;
      RECT 250.47 77.08 251 77.25 ;
      RECT 250.49 76.575 250.66 77.08 ;
      RECT 251.65 76.02 252.32 76.065 ;
      RECT 251.27 76.19 252.16 76.235 ;
      RECT 251.27 76.065 252.32 76.19 ;
      RECT 254.56 73.405 255.09 73.575 ;
      RECT 254.08 74.76 254.78 75.77 ;
      RECT 254.25 75.77 254.78 76.25 ;
      RECT 252.96 73.405 253.51 73.575 ;
      RECT 252.98 73.12 253.51 73.405 ;
      RECT 253.2 74.79 253.73 74.96 ;
      RECT 253.2 74.96 253.37 75.77 ;
      RECT 253.2 74.76 253.37 74.79 ;
      RECT 255.28 73.405 255.65 73.575 ;
      RECT 254.96 74.93 255.13 75.77 ;
      RECT 255.28 73.575 255.61 74.76 ;
      RECT 254.96 74.76 255.61 74.93 ;
      RECT 257.33 74.79 257.86 74.96 ;
      RECT 257.52 74.96 257.69 75.77 ;
      RECT 257.52 74.76 257.69 74.79 ;
      RECT 256.24 75.16 256.77 75.33 ;
      RECT 256.24 75.33 256.41 75.77 ;
      RECT 256.24 74.76 256.41 75.16 ;
      RECT 253.82 78.07 253.99 80.78 ;
      RECT 252.5 78.075 252.67 80.785 ;
      RECT 253.16 78.13 253.33 81.05 ;
      RECT 251.865 77.7 252.535 77.87 ;
      RECT 253.945 77.7 254.615 77.87 ;
      RECT 253.41 76.02 254.08 76.19 ;
      RECT 257.12 75.99 257.65 76.16 ;
      RECT 257.12 76.16 257.29 80.82 ;
      RECT 253.65 81.81 254.87 81.98 ;
      RECT 253.65 84.28 254.18 84.45 ;
      RECT 253.65 84.45 253.82 84.93 ;
      RECT 254.7 78.07 254.87 81.81 ;
      RECT 253.65 81.98 253.82 84.28 ;
      RECT 255.58 78.07 255.75 80.78 ;
      RECT 165.365 79.14 166.17 79.31 ;
      RECT 166 79.31 166.17 80.475 ;
      RECT 169.99 73.855 171.34 74.17 ;
      RECT 168.87 79.54 169.04 80.985 ;
      RECT 169.355 78.34 169.885 78.51 ;
      RECT 169.715 78.51 169.885 78.875 ;
      RECT 169.715 76.165 169.885 78.34 ;
      RECT 166.595 78.34 167.125 78.51 ;
      RECT 166.595 78.51 166.765 78.875 ;
      RECT 166.595 76.165 166.765 78.34 ;
      RECT 166.045 76.165 166.215 78.875 ;
      RECT 167.965 78.34 168.495 78.51 ;
      RECT 168.155 78.51 168.325 78.875 ;
      RECT 168.155 76.165 168.325 78.34 ;
      RECT 170.935 80.165 171.155 81.175 ;
      RECT 170.935 81.175 171.105 82.38 ;
      RECT 170.935 82.38 171.255 85.09 ;
      RECT 171.865 79.54 172.035 81.175 ;
      RECT 172.845 80.66 173.795 81.175 ;
      RECT 173.625 80.165 173.795 80.66 ;
      RECT 172.845 81.175 173.015 85.09 ;
      RECT 170.665 77.48 173.715 78.01 ;
      RECT 170.785 78.01 173.675 79.185 ;
      RECT 170.785 75.265 173.675 77.48 ;
      RECT 171.275 81.37 171.785 81.7 ;
      RECT 171.325 80.66 171.695 81.37 ;
      RECT 216.21 80.66 217.16 81.175 ;
      RECT 216.21 80.165 216.38 80.66 ;
      RECT 216.99 81.175 217.16 85.09 ;
      RECT 216.29 77.48 219.34 78.01 ;
      RECT 216.33 78.01 219.22 79.185 ;
      RECT 216.33 75.265 219.22 77.48 ;
      RECT 219.87 79.14 220.76 79.24 ;
      RECT 219.85 79.31 220.25 83.06 ;
      RECT 219.85 79.24 220.76 79.31 ;
      RECT 220.415 75.775 223.415 75.945 ;
      RECT 222.46 75.945 222.63 78.875 ;
      RECT 220.9 75.945 221.07 78.875 ;
      RECT 219.53 75.275 236.8 75.525 ;
      RECT 219.53 75.525 219.7 79.145 ;
      RECT 236.63 75.525 236.8 79.145 ;
      RECT 218.665 73.855 220.015 74.17 ;
      RECT 220.965 79.54 221.135 80.985 ;
      RECT 220.12 78.34 220.65 78.51 ;
      RECT 220.12 78.51 220.29 78.875 ;
      RECT 220.12 76.165 220.29 78.34 ;
      RECT 218.85 80.165 219.07 81.175 ;
      RECT 218.9 81.175 219.07 82.38 ;
      RECT 218.75 82.38 219.07 85.09 ;
      RECT 217.97 79.54 218.14 81.175 ;
      RECT 218.22 81.37 218.73 81.7 ;
      RECT 218.31 80.66 218.68 81.37 ;
      RECT 221.51 78.34 222.04 78.51 ;
      RECT 221.68 78.51 221.85 78.875 ;
      RECT 221.68 76.165 221.85 78.34 ;
      RECT 227.21 79.14 229.9 79.25 ;
      RECT 227.205 79.25 229.915 79.595 ;
      RECT 224.085 75.775 226.795 75.945 ;
      RECT 224.395 78.34 224.925 78.51 ;
      RECT 225.96 78.34 226.49 78.51 ;
      RECT 224.57 78.51 224.74 78.875 ;
      RECT 226.13 78.51 226.3 78.875 ;
      RECT 224.57 75.945 224.74 78.34 ;
      RECT 226.13 75.945 226.3 78.34 ;
      RECT 223.835 79.14 224.64 79.31 ;
      RECT 223.835 79.31 224.005 80.475 ;
      RECT 228.115 79.9 228.285 80.475 ;
      RECT 223.285 80.79 227.875 80.96 ;
      RECT 224.485 80.96 227.875 81.205 ;
      RECT 224.485 80.695 227.875 80.79 ;
      RECT 223.285 80.96 223.455 80.985 ;
      RECT 223.285 79.635 223.455 80.79 ;
      RECT 222.88 78.34 223.41 78.51 ;
      RECT 223.24 78.51 223.41 78.875 ;
      RECT 223.24 76.165 223.41 78.34 ;
      RECT 226.91 76.165 227.08 78.875 ;
      RECT 223.79 76.165 223.96 78.875 ;
      RECT 225.35 76.165 225.52 78.875 ;
      RECT 227.33 78.34 227.86 78.51 ;
      RECT 227.69 78.51 227.86 78.875 ;
      RECT 227.69 76.165 227.86 78.34 ;
      RECT 230.37 75.87 230.9 75.955 ;
      RECT 230.17 75.7 230.84 75.785 ;
      RECT 230.17 75.785 230.9 75.87 ;
      RECT 231.15 75.775 232.16 75.945 ;
      RECT 232.37 79.14 232.945 79.31 ;
      RECT 232.37 76.165 232.54 79.14 ;
      RECT 233.7 79.62 235.79 79.79 ;
      RECT 233.245 75.775 234.255 75.945 ;
      RECT 235.62 79.79 235.79 86.035 ;
      RECT 233.7 75.945 233.87 79.62 ;
      RECT 228.605 80.695 231.655 80.865 ;
      RECT 229.245 80.865 229.775 83.07 ;
      RECT 231.485 80.865 231.655 83.995 ;
      RECT 231.59 76.165 231.76 78.875 ;
      RECT 230.81 78.265 231.42 78.435 ;
      RECT 230.81 78.435 230.98 78.875 ;
      RECT 230.81 76.165 230.98 78.265 ;
      RECT 230.03 76.165 230.2 78.875 ;
      RECT 232.92 78.35 233.45 78.52 ;
      RECT 232.92 78.52 233.09 78.875 ;
      RECT 232.92 76.165 233.09 78.35 ;
      RECT 228.47 76.165 228.64 78.875 ;
      RECT 229.08 78.34 229.61 78.51 ;
      RECT 229.25 78.51 229.42 78.875 ;
      RECT 229.25 76.165 229.42 78.34 ;
      RECT 235.68 78.35 236.21 78.52 ;
      RECT 234.805 75.775 236.21 75.945 ;
      RECT 236.04 78.52 236.21 78.875 ;
      RECT 236.04 75.945 236.21 78.35 ;
      RECT 235.26 79.14 236.46 79.37 ;
      RECT 236.26 80.145 236.565 80.475 ;
      RECT 236.26 79.37 236.46 80.145 ;
      RECT 235.26 76.165 235.43 79.14 ;
      RECT 238.965 77.18 239.79 79.15 ;
      RECT 238.905 77.01 241.195 77.18 ;
      RECT 238.965 79.15 241.195 79.32 ;
      RECT 240.3 77.18 241.195 79.15 ;
      RECT 238.965 79.32 239.79 81.25 ;
      RECT 238.965 81.25 241.195 81.3 ;
      RECT 240.3 79.32 241.195 81.25 ;
      RECT 238.905 81.3 241.195 81.47 ;
      RECT 237.97 74.42 238.14 76.02 ;
      RECT 237.38 74.4 237.55 81.02 ;
      RECT 237.72 79.73 238.14 81.08 ;
      RECT 237.72 78.75 237.89 79.73 ;
      RECT 237.72 78.24 238.56 78.41 ;
      RECT 142.19 76.895 142.72 77.01 ;
      RECT 145.615 78.95 146.205 79.12 ;
      RECT 144.975 83.29 146.205 83.46 ;
      RECT 145.875 83.46 146.205 83.83 ;
      RECT 145.875 79.12 146.205 83.29 ;
      RECT 145.065 81.92 145.395 83.29 ;
      RECT 146.685 78.95 147.275 79.12 ;
      RECT 146.685 83.29 147.915 83.46 ;
      RECT 146.685 83.46 147.015 83.83 ;
      RECT 146.685 79.12 147.015 83.29 ;
      RECT 147.495 81.92 147.825 83.29 ;
      RECT 145.615 78.24 146.205 78.41 ;
      RECT 145.875 78.41 146.205 78.44 ;
      RECT 145.875 74.92 146.205 78.24 ;
      RECT 146.685 78.24 147.275 78.41 ;
      RECT 146.685 78.41 147.015 78.44 ;
      RECT 146.685 74.92 147.015 78.24 ;
      RECT 144.845 79.73 145.32 81.08 ;
      RECT 145.15 78.75 145.32 79.73 ;
      RECT 144.415 78.24 145.32 78.41 ;
      RECT 144.845 78.41 145.32 78.75 ;
      RECT 144.845 77.4 145.32 78.24 ;
      RECT 145.135 74.4 145.305 74.93 ;
      RECT 145.135 75.43 145.305 76.02 ;
      RECT 142.845 77.4 143.015 78.75 ;
      RECT 142.845 79.54 143.015 81.08 ;
      RECT 144.36 79.11 144.89 79.28 ;
      RECT 144.37 79.28 144.88 79.405 ;
      RECT 144.37 79.075 144.88 79.11 ;
      RECT 148.81 77.18 149.705 79.15 ;
      RECT 148.81 77.01 151.1 77.18 ;
      RECT 148.81 79.15 151.04 79.32 ;
      RECT 150.215 77.18 151.04 79.15 ;
      RECT 148.81 79.32 149.705 81.25 ;
      RECT 148.81 81.25 151.04 81.3 ;
      RECT 150.215 79.32 151.04 81.25 ;
      RECT 148.81 81.3 151.1 81.47 ;
      RECT 152.455 74.4 152.625 81.02 ;
      RECT 151.865 79.73 152.285 81.08 ;
      RECT 152.115 78.75 152.285 79.73 ;
      RECT 151.445 78.24 152.285 78.41 ;
      RECT 151.865 78.41 152.285 78.75 ;
      RECT 151.865 77.4 152.285 78.24 ;
      RECT 147.57 79.73 148.045 81.08 ;
      RECT 147.57 78.75 147.74 79.73 ;
      RECT 147.57 78.24 148.475 78.41 ;
      RECT 147.57 78.41 148.045 78.75 ;
      RECT 147.57 77.4 148.045 78.24 ;
      RECT 151.865 74.42 152.035 76.02 ;
      RECT 148.06 76.37 151.79 76.54 ;
      RECT 147.585 74.4 147.755 74.93 ;
      RECT 147.585 75.43 147.755 76.02 ;
      RECT 149.875 77.4 150.045 78.75 ;
      RECT 149.875 79.54 150.045 81.08 ;
      RECT 147.955 75.1 151.345 75.27 ;
      RECT 148 75.27 148.53 75.33 ;
      RECT 148 79.11 148.53 79.28 ;
      RECT 148.01 79.28 148.52 79.405 ;
      RECT 148.01 79.075 148.52 79.11 ;
      RECT 151.335 79.12 151.9 79.29 ;
      RECT 151.39 79.29 151.9 79.405 ;
      RECT 151.39 79.075 151.9 79.12 ;
      RECT 157.845 75.775 158.855 75.945 ;
      RECT 157.06 79.14 157.635 79.31 ;
      RECT 157.465 76.165 157.635 79.14 ;
      RECT 154.215 79.62 156.305 79.79 ;
      RECT 155.75 75.775 156.76 75.945 ;
      RECT 154.215 79.79 154.385 86.035 ;
      RECT 156.135 75.945 156.305 79.62 ;
      RECT 153.795 78.35 154.325 78.52 ;
      RECT 153.795 75.775 155.2 75.945 ;
      RECT 153.795 78.52 153.965 78.875 ;
      RECT 153.795 75.945 153.965 78.35 ;
      RECT 153.545 79.14 154.745 79.37 ;
      RECT 153.44 80.145 153.745 80.475 ;
      RECT 153.545 79.37 153.745 80.145 ;
      RECT 154.575 76.165 154.745 79.14 ;
      RECT 153.205 75.275 170.475 75.525 ;
      RECT 153.205 75.525 153.375 79.145 ;
      RECT 170.305 75.525 170.475 79.145 ;
      RECT 158.35 80.695 161.4 80.865 ;
      RECT 160.23 80.865 160.76 83.07 ;
      RECT 158.35 80.865 158.52 83.995 ;
      RECT 158.245 76.165 158.415 78.875 ;
      RECT 155.17 78.35 155.7 78.52 ;
      RECT 155.355 78.52 155.525 78.875 ;
      RECT 155.355 76.165 155.525 78.35 ;
      RECT 156.555 78.35 157.085 78.52 ;
      RECT 156.915 78.52 157.085 78.875 ;
      RECT 156.915 76.165 157.085 78.35 ;
      RECT 158.585 78.265 159.195 78.435 ;
      RECT 159.025 76.165 159.195 78.265 ;
      RECT 159.025 78.435 159.195 78.875 ;
      RECT 159.105 75.87 159.635 75.955 ;
      RECT 159.165 75.7 159.835 75.785 ;
      RECT 159.105 75.785 159.835 75.87 ;
      RECT 160.105 79.14 162.795 79.25 ;
      RECT 160.09 79.25 162.8 79.595 ;
      RECT 163.21 75.775 165.92 75.945 ;
      RECT 163.515 78.34 164.045 78.51 ;
      RECT 165.08 78.34 165.61 78.51 ;
      RECT 163.705 78.51 163.875 78.875 ;
      RECT 165.265 78.51 165.435 78.875 ;
      RECT 163.705 75.945 163.875 78.34 ;
      RECT 165.265 75.945 165.435 78.34 ;
      RECT 161.72 79.9 161.89 80.475 ;
      RECT 162.13 80.79 166.72 80.96 ;
      RECT 162.13 80.96 165.52 81.205 ;
      RECT 162.13 80.695 165.52 80.79 ;
      RECT 166.55 80.96 166.72 80.985 ;
      RECT 166.55 79.635 166.72 80.79 ;
      RECT 159.805 76.165 159.975 78.875 ;
      RECT 162.925 76.165 163.095 78.875 ;
      RECT 160.395 78.34 160.925 78.51 ;
      RECT 160.585 78.51 160.755 78.875 ;
      RECT 160.585 76.165 160.755 78.34 ;
      RECT 161.365 76.165 161.535 78.875 ;
      RECT 164.485 76.165 164.655 78.875 ;
      RECT 162.145 78.34 162.675 78.51 ;
      RECT 162.145 78.51 162.315 78.875 ;
      RECT 162.145 76.165 162.315 78.34 ;
      RECT 169.245 79.14 170.135 79.24 ;
      RECT 169.755 79.31 170.155 83.06 ;
      RECT 169.245 79.24 170.155 79.31 ;
      RECT 166.59 75.775 169.59 75.945 ;
      RECT 167.375 75.945 167.545 78.875 ;
      RECT 168.935 75.945 169.105 78.875 ;
      RECT 121.755 78.12 121.925 81.77 ;
      RECT 120.875 78.12 121.045 82.87 ;
      RECT 119.115 78.12 119.285 82.87 ;
      RECT 119.805 81.77 120.335 81.94 ;
      RECT 119.995 81.94 120.165 82.87 ;
      RECT 119.995 78.12 120.165 81.77 ;
      RECT 127.195 77.68 128.545 77.85 ;
      RECT 125.435 77.68 126.785 77.85 ;
      RECT 124.555 78.13 124.725 81.05 ;
      RECT 128.995 76.42 132.395 76.59 ;
      RECT 128.995 76.59 129.165 77.155 ;
      RECT 129.765 76.37 132.095 76.42 ;
      RECT 127.505 75.16 128.035 75.33 ;
      RECT 127.615 75.33 127.945 75.69 ;
      RECT 126.64 75.16 127.17 75.33 ;
      RECT 126.735 75.33 127.065 75.69 ;
      RECT 129.685 77.2 132.395 77.37 ;
      RECT 129.765 77.08 132.095 77.2 ;
      RECT 128.135 79.055 128.835 79.225 ;
      RECT 128.665 79.225 128.835 80.78 ;
      RECT 128.665 78.07 128.835 79.055 ;
      RECT 126.715 79.055 127.245 79.225 ;
      RECT 126.905 79.225 127.075 80.78 ;
      RECT 126.905 78.07 127.075 79.055 ;
      RECT 125.145 79.055 125.845 79.225 ;
      RECT 125.145 79.225 125.315 80.78 ;
      RECT 125.145 78.07 125.315 79.055 ;
      RECT 129.755 74.79 130.345 74.96 ;
      RECT 129.755 74.96 129.925 75.77 ;
      RECT 129.755 74.76 129.925 74.79 ;
      RECT 126.305 76.22 126.475 77.36 ;
      RECT 128.205 76.22 128.375 77.36 ;
      RECT 129.31 78.09 129.86 81.09 ;
      RECT 126.645 80.95 127.955 81.165 ;
      RECT 126.515 84.07 127.045 84.24 ;
      RECT 126.645 84.24 126.815 84.93 ;
      RECT 127.785 78.07 127.955 80.95 ;
      RECT 126.645 81.165 126.815 84.07 ;
      RECT 126.025 78.07 126.195 80.78 ;
      RECT 133.935 74.54 134.225 76.42 ;
      RECT 133.935 76.42 138.835 76.59 ;
      RECT 136.975 74.76 137.685 75.77 ;
      RECT 136.975 75.77 137.515 76.42 ;
      RECT 130.025 74 134.225 74.54 ;
      RECT 132.145 74.79 132.675 74.96 ;
      RECT 132.315 74.96 132.485 75.77 ;
      RECT 132.315 74.76 132.485 74.79 ;
      RECT 130.665 75.18 131.205 75.35 ;
      RECT 131.035 74.76 131.205 75.18 ;
      RECT 131.035 75.35 131.205 75.77 ;
      RECT 133.235 75.16 133.765 75.33 ;
      RECT 133.595 75.33 133.765 75.77 ;
      RECT 133.595 74.76 133.765 75.16 ;
      RECT 134.915 73.405 135.445 73.575 ;
      RECT 135.1 74.37 139.22 74.54 ;
      RECT 137.815 73.83 139.135 74.37 ;
      RECT 134.355 73.405 134.725 73.575 ;
      RECT 134.875 74.93 135.045 75.77 ;
      RECT 134.395 73.575 134.725 74.76 ;
      RECT 134.395 74.76 135.045 74.93 ;
      RECT 135.225 74.76 135.925 75.77 ;
      RECT 135.225 75.77 135.755 76.25 ;
      RECT 132.355 75.99 132.885 76.16 ;
      RECT 132.715 76.16 132.885 80.82 ;
      RECT 133.555 77.3 138.835 77.48 ;
      RECT 133.555 77.48 134.085 78.01 ;
      RECT 133.595 76.07 133.765 77.3 ;
      RECT 136.28 77.48 137.17 77.62 ;
      RECT 133.595 78.01 133.765 80.82 ;
      RECT 130.225 80.95 131.39 81.12 ;
      RECT 130.035 84.28 130.565 84.45 ;
      RECT 130.225 84.45 130.395 84.93 ;
      RECT 131.22 78.07 131.39 80.95 ;
      RECT 130.225 81.12 130.395 84.28 ;
      RECT 130.34 78.07 130.51 80.78 ;
      RECT 132.1 78.07 132.27 80.78 ;
      RECT 131.475 77.68 132.145 77.85 ;
      RECT 130.475 77.68 131.145 77.85 ;
      RECT 135.135 81.81 136.355 81.98 ;
      RECT 135.825 84.28 136.355 84.45 ;
      RECT 136.185 84.45 136.355 84.93 ;
      RECT 135.135 78.07 135.305 81.81 ;
      RECT 136.185 81.98 136.355 84.28 ;
      RECT 134.255 78.07 134.425 80.78 ;
      RECT 134.39 77.7 135.06 77.87 ;
      RECT 135.39 77.7 136.06 77.87 ;
      RECT 140.265 74.4 140.435 81.02 ;
      RECT 136.495 73.405 137.045 73.575 ;
      RECT 136.495 73.12 137.025 73.405 ;
      RECT 136.275 74.79 136.805 74.96 ;
      RECT 136.635 74.96 136.805 75.77 ;
      RECT 136.635 74.76 136.805 74.79 ;
      RECT 135.925 76.02 136.595 76.19 ;
      RECT 140.855 74.42 141.025 76.02 ;
      RECT 138.225 74.79 138.755 74.96 ;
      RECT 138.395 74.96 138.565 75.77 ;
      RECT 138.395 74.76 138.565 74.79 ;
      RECT 139.005 77.08 139.535 77.25 ;
      RECT 139.345 76.575 139.515 77.08 ;
      RECT 137.845 76.19 138.735 76.235 ;
      RECT 137.685 76.02 138.355 76.065 ;
      RECT 137.685 76.065 138.735 76.19 ;
      RECT 141.1 76.37 144.83 76.54 ;
      RECT 141.545 75.1 144.935 75.27 ;
      RECT 144.36 75.27 144.89 75.33 ;
      RECT 136.015 78.07 136.185 80.78 ;
      RECT 136.675 78.13 136.845 81.05 ;
      RECT 140.605 79.73 141.025 81.08 ;
      RECT 140.605 78.75 140.775 79.73 ;
      RECT 140.605 78.24 141.445 78.41 ;
      RECT 140.605 78.41 141.025 78.75 ;
      RECT 140.605 77.4 141.025 78.24 ;
      RECT 140.99 79.12 141.555 79.29 ;
      RECT 140.99 79.29 141.5 79.405 ;
      RECT 140.99 79.075 141.5 79.12 ;
      RECT 138.995 81.43 139.265 81.6 ;
      RECT 138.805 83.69 139.335 83.86 ;
      RECT 139.095 78.075 139.265 81.43 ;
      RECT 138.995 83.86 139.165 86.93 ;
      RECT 138.995 81.6 139.165 83.69 ;
      RECT 138.215 78.075 138.385 80.785 ;
      RECT 137.335 78.075 137.505 80.785 ;
      RECT 138.47 77.7 139.14 77.87 ;
      RECT 137.47 77.7 138.14 77.87 ;
      RECT 143.07 77.01 144.08 77.18 ;
      RECT 143.47 76.895 144 77.01 ;
      RECT 141.79 77.01 142.8 77.18 ;
      RECT 43.45 76.4 43.62 77.11 ;
      RECT 49.335 77.05 49.535 80.86 ;
      RECT 49.35 80.86 49.52 81.15 ;
      RECT 49.35 76.4 49.52 77.05 ;
      RECT 50.115 77.05 50.315 80.86 ;
      RECT 50.13 76.4 50.3 77.05 ;
      RECT 49.575 81.61 50.3 81.78 ;
      RECT 50.13 80.86 50.3 81.61 ;
      RECT 50.68 76.4 50.85 81.15 ;
      RECT 53.8 77.05 53.98 80.46 ;
      RECT 53.8 80.46 53.97 81.15 ;
      RECT 53.8 76.4 53.97 77.05 ;
      RECT 54.35 81.61 55.455 81.78 ;
      RECT 54.35 76.4 54.52 81.61 ;
      RECT 51.02 80.75 51.29 81.315 ;
      RECT 50.905 81.315 51.29 81.32 ;
      RECT 51.8 80.75 52.07 81.32 ;
      RECT 52.58 80.75 52.85 81.32 ;
      RECT 53.36 80.75 53.63 81.32 ;
      RECT 50.905 81.32 53.745 81.78 ;
      RECT 51.46 76.4 51.63 81.15 ;
      RECT 53.02 76.4 53.19 81.15 ;
      RECT 52.24 76.4 52.41 81.15 ;
      RECT 58.19 76.4 58.36 81.15 ;
      RECT 55.63 76.4 55.8 81.15 ;
      RECT 56.91 76.4 57.08 81.15 ;
      RECT 59.47 76.4 59.64 81.15 ;
      RECT 60.75 76.4 60.92 81.15 ;
      RECT 63.31 76.4 63.48 81.15 ;
      RECT 65.87 76.4 66.04 81.15 ;
      RECT 64.59 76.4 64.76 81.15 ;
      RECT 62.03 76.4 62.2 81.15 ;
      RECT 70.99 76.4 71.16 81.15 ;
      RECT 68.43 76.4 68.6 81.15 ;
      RECT 69.71 76.4 69.88 81.15 ;
      RECT 67.15 76.4 67.32 81.15 ;
      RECT 73.55 76.4 73.72 81.15 ;
      RECT 76.11 76.4 76.28 81.15 ;
      RECT 72.27 76.4 72.44 81.15 ;
      RECT 74.83 76.4 75 81.15 ;
      RECT 77.39 76.4 77.56 81.15 ;
      RECT 81.23 76.4 81.4 81.15 ;
      RECT 78.67 76.4 78.84 81.15 ;
      RECT 82.51 76.4 82.68 81.15 ;
      RECT 79.95 76.4 80.12 81.15 ;
      RECT 85.07 76.4 85.24 81.15 ;
      RECT 83.79 76.4 83.96 81.15 ;
      RECT 100.935 80.615 101.255 81.925 ;
      RECT 101.01 80.595 101.18 80.615 ;
      RECT 100.74 78.83 100.91 79.42 ;
      RECT 99.605 79.61 101.6 79.945 ;
      RECT 99.605 78.225 99.935 79.61 ;
      RECT 99.685 80.405 100.1 82.14 ;
      RECT 99.685 80.16 101.835 80.405 ;
      RECT 99.685 82.81 99.95 86.93 ;
      RECT 99.685 86.93 101.65 87.285 ;
      RECT 99.685 82.14 100.715 82.81 ;
      RECT 103.35 74.405 104.7 74.575 ;
      RECT 104.345 74.575 104.515 75.69 ;
      RECT 103.665 74.575 103.835 75.69 ;
      RECT 104.5 73.865 105.85 74.035 ;
      RECT 104.55 73.6 105.8 73.865 ;
      RECT 101.89 80.595 102.06 81.18 ;
      RECT 101.52 78.89 102.38 79.42 ;
      RECT 101.85 79.42 102.38 79.96 ;
      RECT 106.645 74.765 106.815 77.645 ;
      RECT 103.125 77.645 106.815 77.815 ;
      RECT 104.885 74.765 105.055 77.645 ;
      RECT 103.125 74.765 103.295 77.645 ;
      RECT 106.43 79.755 106.6 82.465 ;
      RECT 102.91 79.755 103.08 82.465 ;
      RECT 104.005 77.08 104.535 77.25 ;
      RECT 104.005 77.25 104.175 77.475 ;
      RECT 104.005 74.765 104.175 77.08 ;
      RECT 105.545 79.525 105.715 79.755 ;
      RECT 105.55 80.54 105.72 82.465 ;
      RECT 105.545 79.755 105.72 80.54 ;
      RECT 104.67 79.755 104.84 82.465 ;
      RECT 103.785 79.525 103.955 79.755 ;
      RECT 103.79 80.54 103.96 82.465 ;
      RECT 103.785 79.755 103.96 80.54 ;
      RECT 107.59 74.405 108.6 74.575 ;
      RECT 107.65 74 108.54 74.405 ;
      RECT 109.45 74.405 110.46 74.575 ;
      RECT 110.175 74.575 110.345 75.69 ;
      RECT 109.495 74.575 109.665 75.69 ;
      RECT 111.055 74.405 112.185 74.575 ;
      RECT 111.055 74.575 111.225 75.69 ;
      RECT 111.935 74.575 112.105 75.69 ;
      RECT 107.775 77.08 108.305 77.25 ;
      RECT 108.075 77.25 108.245 77.475 ;
      RECT 108.075 74.765 108.245 77.08 ;
      RECT 109.655 77.08 110.185 77.25 ;
      RECT 109.835 77.25 110.005 77.475 ;
      RECT 109.835 74.765 110.005 77.08 ;
      RECT 111.415 77.08 111.945 77.25 ;
      RECT 111.595 77.25 111.765 77.475 ;
      RECT 111.595 74.765 111.765 77.08 ;
      RECT 107.86 79.265 110.76 79.435 ;
      RECT 108.05 80.045 110.76 80.215 ;
      RECT 110.705 83.31 111.235 83.48 ;
      RECT 111.01 81.675 111.235 83.31 ;
      RECT 111.01 79.315 111.575 81.675 ;
      RECT 107.31 79.26 107.48 79.99 ;
      RECT 107.295 80.27 107.495 82.645 ;
      RECT 103.135 82.645 107.495 82.845 ;
      RECT 103.135 82.845 106.375 82.855 ;
      RECT 112.055 79.09 116.805 79.26 ;
      RECT 111.915 79.965 115.685 79.97 ;
      RECT 111.915 79.97 116.805 80.135 ;
      RECT 112.055 80.135 116.805 80.14 ;
      RECT 113.815 73.865 114.825 74.035 ;
      RECT 113.875 73.6 114.765 73.865 ;
      RECT 118.235 81.77 118.765 81.94 ;
      RECT 118.235 81.94 118.405 82.87 ;
      RECT 118.235 78.12 118.405 81.77 ;
      RECT 113.025 77.08 113.555 77.25 ;
      RECT 113.025 77.25 113.195 77.475 ;
      RECT 113.025 74.765 113.195 77.08 ;
      RECT 116.185 77.08 116.715 77.25 ;
      RECT 116.545 77.25 116.715 77.475 ;
      RECT 116.545 74.765 116.715 77.08 ;
      RECT 114.605 77.08 115.135 77.25 ;
      RECT 114.785 77.25 114.955 77.475 ;
      RECT 114.785 74.765 114.955 77.08 ;
      RECT 121.395 81.77 121.925 81.94 ;
      RECT 121.755 81.94 121.925 82.87 ;
      RECT 28.79 75.99 28.96 76.62 ;
      RECT 27.89 75.82 28.96 75.99 ;
      RECT 28.79 74.76 28.96 75.82 ;
      RECT 29.45 76.79 29.62 77.97 ;
      RECT 28.79 76.62 29.62 76.79 ;
      RECT 28.17 76.62 28.34 77.97 ;
      RECT 36.375 74.405 36.545 79.155 ;
      RECT 32.63 76.65 32.8 77.66 ;
      RECT 32.63 74.59 32.8 75.6 ;
      RECT 35.895 74.155 36.065 80.16 ;
      RECT 38.135 74.155 38.305 80.16 ;
      RECT 35.895 73.985 38.305 74.155 ;
      RECT 35.895 80.16 38.305 80.36 ;
      RECT 36.72 79.665 37.53 79.835 ;
      RECT 42.855 77.11 43.055 80.65 ;
      RECT 85.65 76.05 85.82 82.02 ;
      RECT 42.87 80.65 43.04 82.02 ;
      RECT 42.87 76.05 43.04 77.11 ;
      RECT 42.87 75.88 85.82 76.05 ;
      RECT 42.87 82.02 85.82 82.19 ;
      RECT 41.58 252.535 175.92 253.385 ;
      RECT 41.58 249.375 42.43 252.535 ;
      RECT 25.15 248.525 42.43 249.375 ;
      RECT 166.05 244.045 166.9 252.535 ;
      RECT 174.16 244.045 175.92 252.535 ;
      RECT 166.05 243.195 175.92 244.045 ;
      RECT 25.15 226.45 26 248.525 ;
      RECT 41.58 226.44 42.43 248.525 ;
      RECT 18.865 226.44 26 226.45 ;
      RECT 18.865 225.59 42.43 226.44 ;
      RECT 41.58 215.97 42.43 225.59 ;
      RECT 41.58 215.53 45.375 215.97 ;
      RECT 18.865 204.335 19.725 225.59 ;
      RECT 41.58 204.335 45.52 215.53 ;
      RECT 18.865 203.475 45.52 204.335 ;
      RECT 41.58 200.645 45.52 203.475 ;
      RECT 174 195.155 175.92 243.195 ;
      RECT 162.04 194.305 175.92 195.155 ;
      RECT 41.58 184.19 44.535 200.645 ;
      RECT 43.685 177.45 44.535 184.19 ;
      RECT 43.685 176.6 90.225 177.45 ;
      RECT 162.04 176.145 162.89 194.305 ;
      RECT 89.375 176.145 90.225 176.6 ;
      RECT 175.02 174.305 175.92 194.305 ;
      RECT 175.02 173.235 190.325 174.305 ;
      RECT 89.375 173.235 162.89 176.145 ;
      RECT 89.375 168.145 190.325 173.235 ;
      RECT 61.745 160.22 62.595 176.6 ;
      RECT 89.375 160 90.225 168.145 ;
      RECT 38.6 160 88.14 160.22 ;
      RECT 38.6 159.15 90.225 160 ;
      RECT 49.34 157.925 50.19 159.15 ;
      RECT 38.6 154.015 39.45 159.15 ;
      RECT 49.305 152.475 50.195 157.925 ;
      RECT 38.58 152.35 39.47 154.015 ;
      RECT 38.6 151.61 39.45 152.35 ;
      RECT 49.34 151.055 50.19 152.475 ;
      RECT 38.58 150.57 39.47 151.61 ;
      RECT 38.6 149.94 39.45 150.57 ;
      RECT 49.305 148.365 50.195 151.055 ;
      RECT 38.58 148.365 39.47 149.94 ;
      RECT 38.6 147.6 39.45 148.365 ;
      RECT 49.34 147.135 50.19 148.365 ;
      RECT 38.58 147.07 39.47 147.6 ;
      RECT 49.305 146.79 50.195 147.135 ;
      RECT 38.6 145.1 39.45 147.07 ;
      RECT 87.29 143.905 90.225 159.15 ;
      RECT 49.34 143.905 50.19 146.79 ;
      RECT 31.71 143.885 39.45 145.1 ;
      RECT 49.34 143.735 90.225 143.905 ;
      RECT 31.71 128.205 32.56 143.885 ;
      RECT 89.035 128.205 90.225 143.735 ;
      RECT 49.34 128.205 49.99 143.735 ;
      RECT 31.405 127.885 90.225 128.205 ;
      RECT 55.205 115.675 55.375 127.885 ;
      RECT 79.005 115.675 79.175 127.885 ;
      RECT 31.405 115.675 31.575 127.885 ;
      RECT 31.405 115.375 79.175 115.675 ;
      RECT 189.475 109.585 190.325 168.145 ;
      RECT 89.035 109.585 90.225 127.885 ;
      RECT 89.035 108.735 190.325 109.585 ;
      RECT 118.035 108.38 166.055 108.735 ;
      RECT 31.405 106.36 31.575 115.375 ;
      RECT 71.585 106.36 71.755 115.375 ;
      RECT 31.405 106.16 71.755 106.36 ;
      RECT 118.035 103.77 121.145 108.38 ;
      RECT 153.83 103.77 166.055 108.38 ;
      RECT 140.195 103.77 140.365 108.38 ;
      RECT 118.035 102.92 166.055 103.77 ;
      RECT 177.595 101.9 190.275 108.735 ;
      RECT 173.88 101.9 174.73 108.735 ;
      RECT 71.585 97.145 71.755 106.16 ;
      RECT 31.405 97.145 31.575 106.16 ;
      RECT 173.88 97.095 190.275 101.9 ;
      RECT 173.88 97.045 190.27 97.095 ;
      RECT 154.28 97.045 166.055 102.92 ;
      RECT 154.28 96.88 190.27 97.045 ;
      RECT 31.405 96.855 79.175 97.145 ;
      RECT 174.305 95.985 190.27 95.995 ;
      RECT 174.18 95.995 190.27 96.03 ;
      RECT 167.13 95.995 173.88 96.03 ;
      RECT 154.28 96.03 190.275 96.88 ;
      RECT 89.035 84.825 89.205 108.735 ;
      RECT 55.205 84.825 55.375 96.855 ;
      RECT 79.005 84.825 79.175 96.855 ;
      RECT 31.405 84.825 31.575 96.855 ;
      RECT 31.405 83.975 89.205 84.825 ;
      RECT 41.255 82.955 87.72 83.975 ;
      RECT 41.255 75.12 42.11 82.955 ;
      RECT 86.43 75.12 87.72 82.955 ;
      RECT 41.255 74.465 87.72 75.12 ;
      RECT 37.655 74.405 37.825 79.155 ;
      RECT 46.775 77.05 46.975 80.86 ;
      RECT 46.79 80.86 46.96 81.15 ;
      RECT 46.79 76.4 46.96 77.05 ;
      RECT 44.23 77.05 44.435 80.25 ;
      RECT 44.23 76.4 44.4 77.05 ;
      RECT 44.23 80.25 44.4 81.15 ;
      RECT 48.055 77.11 48.255 80.92 ;
      RECT 44.455 81.555 49.295 81.835 ;
      RECT 45.495 77.11 45.695 80.92 ;
      RECT 48.07 76.4 48.24 77.11 ;
      RECT 45.51 76.4 45.68 77.11 ;
      RECT 48.07 80.92 48.24 81.555 ;
      RECT 45.51 80.92 45.68 81.555 ;
      RECT 43.435 77.11 43.635 80.65 ;
      RECT 43.45 80.65 43.62 81.15 ;
      RECT 393.2 67.055 393.53 67.705 ;
      RECT 392.57 67.055 392.9 67.705 ;
      RECT 393.83 67.055 394.16 67.705 ;
      RECT 394.46 67.055 394.79 67.705 ;
      RECT 390.68 68.085 391.01 68.735 ;
      RECT 391.31 68.085 391.64 68.735 ;
      RECT 391.94 68.085 392.27 68.735 ;
      RECT 393.2 68.085 393.53 68.735 ;
      RECT 392.57 68.085 392.9 68.735 ;
      RECT 393.83 68.085 394.16 68.735 ;
      RECT 394.46 68.085 394.79 68.735 ;
      RECT 430.48 70.795 430.81 71.485 ;
      RECT 429.71 70.795 430.04 71.485 ;
      RECT 431.165 71.185 433.89 71.81 ;
      RECT 431.165 70.745 431.665 71.185 ;
      RECT 436.31 70.795 436.64 71.485 ;
      RECT 434.21 71.315 434.74 71.485 ;
      RECT 435.1 70.795 435.43 71.485 ;
      RECT 432.02 70.495 433.12 71.005 ;
      RECT 433.56 70.495 434.66 71.005 ;
      RECT 437 71.315 437.53 71.485 ;
      RECT 437.85 71.185 440.575 71.81 ;
      RECT 440.075 70.745 440.575 71.185 ;
      RECT 440.93 70.795 441.26 71.485 ;
      RECT 441.7 70.795 442.03 71.485 ;
      RECT 438.62 70.495 439.72 71.005 ;
      RECT 437.08 70.495 438.18 71.005 ;
      RECT 453.17 72.085 453.34 76.835 ;
      RECT 453.755 76.485 454.315 76.805 ;
      RECT 453.95 76.805 454.12 76.835 ;
      RECT 453.95 72.085 454.12 76.485 ;
      RECT 453.22 71.565 456.36 71.735 ;
      RECT 453.22 69.675 456.36 69.845 ;
      RECT 455.145 76.485 455.705 76.805 ;
      RECT 455.35 76.805 455.52 76.835 ;
      RECT 455.35 72.085 455.52 76.485 ;
      RECT 455.94 75.905 456.475 76.225 ;
      RECT 456.13 76.225 456.3 76.835 ;
      RECT 456.13 72.085 456.3 75.905 ;
      RECT 454.415 75.325 454.98 75.645 ;
      RECT 454.57 75.645 454.74 76.835 ;
      RECT 454.57 72.085 454.74 75.325 ;
      RECT 457.03 71.355 457.655 72.365 ;
      RECT 457.03 77.515 457.2 77.545 ;
      RECT 457.03 77.345 457.655 77.515 ;
      RECT 457.03 72.365 457.2 77.345 ;
      RECT 459.645 77.875 460.175 78.045 ;
      RECT 458.635 70.855 460.175 71.185 ;
      RECT 459.805 78.045 460.175 78.05 ;
      RECT 459.805 71.185 460.175 77.875 ;
      RECT 457.755 70.855 458.265 71.185 ;
      RECT 457.825 71.185 458.195 72.76 ;
      RECT 457.825 72.76 458.355 72.93 ;
      RECT 457.755 66.28 458.265 66.61 ;
      RECT 457.825 66.61 458.195 68.085 ;
      RECT 457.825 68.085 458.355 68.255 ;
      RECT 457.755 70.225 458.265 70.555 ;
      RECT 457.825 68.65 458.195 70.225 ;
      RECT 457.825 68.48 458.355 68.65 ;
      RECT 459.245 71.355 459.415 72.76 ;
      RECT 458.885 72.76 459.415 72.93 ;
      RECT 458.365 71.355 458.535 72.405 ;
      RECT 457.485 66.78 457.655 67.83 ;
      RECT 458.365 66.78 458.535 67.79 ;
      RECT 459.245 68.65 459.415 70.055 ;
      RECT 458.885 68.48 459.415 68.65 ;
      RECT 458.365 69.005 458.535 70.055 ;
      RECT 459.245 66.78 459.415 68.085 ;
      RECT 458.885 68.085 459.415 68.255 ;
      RECT 461.615 72.76 462.145 72.93 ;
      RECT 461.545 77.265 462.055 77.595 ;
      RECT 461.615 72.93 461.985 77.265 ;
      RECT 463.035 72.76 463.565 72.93 ;
      RECT 463.035 72.93 463.205 77.1 ;
      RECT 469.485 75.905 470.045 76.225 ;
      RECT 469.65 76.225 469.82 76.835 ;
      RECT 469.65 72.085 469.82 75.905 ;
      RECT 471.21 72.085 471.38 76.835 ;
      RECT 467.245 72.745 469.1 72.995 ;
      RECT 468.85 71.735 469.1 72.745 ;
      RECT 468.165 72.995 468.615 76.985 ;
      RECT 468.85 71.485 471.42 71.735 ;
      RECT 470.2 76.485 470.76 76.805 ;
      RECT 470.43 76.805 470.6 76.835 ;
      RECT 470.43 72.085 470.6 76.485 ;
      RECT 20.13 80.16 22.52 80.33 ;
      RECT 20.13 73.91 22.52 74.08 ;
      RECT 20.13 74.08 20.3 80.16 ;
      RECT 22.35 74.08 22.52 80.16 ;
      RECT 20.955 79.69 22.18 79.86 ;
      RECT 21.77 74.51 21.94 79.47 ;
      RECT 20.71 74.51 20.88 79.47 ;
      RECT 21.24 74.72 21.41 79.47 ;
      RECT 25.33 75.82 27.36 75.99 ;
      RECT 25.61 76.62 25.78 77.97 ;
      RECT 24.99 74.59 25.16 77.66 ;
      RECT 23.71 76.65 23.88 77.66 ;
      RECT 23.71 74.59 23.88 75.6 ;
      RECT 23.13 74.08 23.3 75.58 ;
      RECT 33.21 74.08 33.38 75.58 ;
      RECT 23.13 73.91 33.38 74.08 ;
      RECT 28.19 74.08 28.36 75.58 ;
      RECT 33.21 76.64 35.33 78.76 ;
      RECT 34.05 73.725 35.33 76.64 ;
      RECT 23.13 76.64 23.3 78.76 ;
      RECT 23.13 78.76 35.33 78.93 ;
      RECT 23.19 78.93 35.33 79.19 ;
      RECT 23.13 79.595 34.9 82.42 ;
      RECT 23.13 79.19 35.33 79.595 ;
      RECT 28.52 78.35 30.55 78.52 ;
      RECT 28.82 77.07 28.99 78.35 ;
      RECT 25.96 78.35 27.99 78.52 ;
      RECT 27.52 77.07 27.69 78.35 ;
      RECT 29.13 75.82 31.18 75.99 ;
      RECT 29.13 75.12 29.3 75.82 ;
      RECT 30.73 76.62 30.9 77.97 ;
      RECT 31.35 74.59 31.52 77.66 ;
      RECT 30.07 74.59 30.24 75.6 ;
      RECT 26.27 74.59 26.44 75.6 ;
      RECT 26.77 74.59 27.72 74.76 ;
      RECT 27.55 74.56 27.72 74.59 ;
      RECT 27.55 74.76 27.72 75.12 ;
      RECT 27.55 75.65 27.72 76.62 ;
      RECT 26.89 76.79 27.06 77.97 ;
      RECT 26.89 76.62 27.72 76.79 ;
      RECT 27.55 75.12 28.02 75.65 ;
      RECT 28.79 74.59 29.74 74.76 ;
      RECT 264.385 70.12 264.555 71.945 ;
      RECT 264.405 75.57 264.935 75.74 ;
      RECT 264.48 75.74 264.65 77.23 ;
      RECT 264.48 72.25 264.65 75.57 ;
      RECT 263.53 71.775 263.7 74.96 ;
      RECT 268.08 73.325 268.61 73.495 ;
      RECT 268.08 73.495 268.25 77.57 ;
      RECT 268.08 72.82 268.25 73.325 ;
      RECT 268.96 72.82 269.13 77.57 ;
      RECT 267.31 72.55 267.875 75.51 ;
      RECT 267.21 75.51 267.875 82.88 ;
      RECT 268.42 72.31 268.79 73.155 ;
      RECT 268.235 72.14 268.905 72.31 ;
      RECT 269.195 72.14 270.885 72.31 ;
      RECT 270.18 72.31 270.55 73.155 ;
      RECT 269.3 72.31 269.67 73.155 ;
      RECT 271.24 73.325 271.77 73.495 ;
      RECT 271.085 71.96 271.69 72.25 ;
      RECT 271.48 72.25 271.69 72.82 ;
      RECT 271.48 73.495 271.77 77.57 ;
      RECT 271.48 72.82 271.77 73.325 ;
      RECT 270.805 69.905 271.375 70.075 ;
      RECT 271.085 70.075 271.375 71.96 ;
      RECT 271.085 68.95 271.375 69.905 ;
      RECT 274.14 68.255 274.31 73.625 ;
      RECT 280.58 68.255 280.75 73.625 ;
      RECT 287.02 68.255 287.19 73.625 ;
      RECT 275.6 68.255 275.77 73.355 ;
      RECT 277.36 68.255 277.53 73.355 ;
      RECT 279.12 68.255 279.29 73.355 ;
      RECT 274.14 68.085 287.19 68.255 ;
      RECT 281.16 68.255 281.33 73.355 ;
      RECT 282.92 68.255 283.09 73.355 ;
      RECT 286.44 68.255 286.61 73.355 ;
      RECT 284.68 68.255 284.85 73.355 ;
      RECT 274.72 69.905 275.25 70.075 ;
      RECT 274.17 74.34 276.65 74.595 ;
      RECT 276.3 69.905 276.83 70.075 ;
      RECT 278.06 69.905 278.59 70.075 ;
      RECT 279.64 69.905 280.17 70.075 ;
      RECT 274.72 68.605 274.89 69.905 ;
      RECT 274.72 70.075 274.89 74.34 ;
      RECT 276.48 68.605 276.65 69.905 ;
      RECT 276.48 73.985 276.65 74.34 ;
      RECT 276.48 73.815 280.17 73.985 ;
      RECT 276.48 70.075 276.65 73.815 ;
      RECT 278.24 68.605 278.41 69.905 ;
      RECT 280 68.605 280.17 69.905 ;
      RECT 278.24 70.075 278.41 73.815 ;
      RECT 280 70.075 280.17 73.815 ;
      RECT 274.17 74.595 274.34 77.475 ;
      RECT 275.93 74.595 276.1 77.475 ;
      RECT 271.86 68.49 272.03 72.305 ;
      RECT 272.17 72.545 272.885 78.155 ;
      RECT 272.17 78.57 272.885 82.85 ;
      RECT 287.29 74.4 287.46 78.155 ;
      RECT 279.12 74.4 279.29 78.155 ;
      RECT 277.36 74.4 277.53 78.155 ;
      RECT 280.88 74.4 281.05 78.155 ;
      RECT 272.17 78.155 287.46 78.57 ;
      RECT 282.64 74.4 282.81 78.155 ;
      RECT 269.42 69.905 269.95 70.075 ;
      RECT 269.605 70.075 269.775 71.66 ;
      RECT 269.605 68.95 269.775 69.905 ;
      RECT 270.195 70.305 270.725 70.475 ;
      RECT 270.385 70.475 270.555 71.66 ;
      RECT 270.385 68.95 270.555 70.305 ;
      RECT 270.72 72.82 270.89 77.57 ;
      RECT 269.67 73.325 270.2 73.495 ;
      RECT 269.84 73.495 270.01 77.57 ;
      RECT 269.84 72.82 270.01 73.325 ;
      RECT 282.04 69.905 282.57 70.075 ;
      RECT 282.04 70.075 282.21 73.355 ;
      RECT 282.04 68.605 282.21 69.905 ;
      RECT 285.195 69.905 285.73 70.075 ;
      RECT 285.56 68.605 285.73 69.905 ;
      RECT 285.56 70.075 285.73 73.355 ;
      RECT 283.62 69.905 284.15 70.075 ;
      RECT 283.8 68.605 283.97 69.905 ;
      RECT 283.8 70.075 283.97 74.765 ;
      RECT 283.8 74.765 284.24 74.935 ;
      RECT 284.07 74.935 284.24 77.475 ;
      RECT 297.645 65.155 297.815 67.865 ;
      RECT 299.795 71.685 301.815 72.435 ;
      RECT 302.765 65.155 302.935 67.865 ;
      RECT 301.485 65.155 301.655 67.865 ;
      RECT 300.205 65.155 300.375 67.865 ;
      RECT 298.925 65.155 299.095 67.865 ;
      RECT 307.885 65.155 308.055 67.865 ;
      RECT 306.605 65.155 306.775 67.865 ;
      RECT 305.325 65.155 305.495 67.865 ;
      RECT 304.045 65.155 304.215 67.865 ;
      RECT 316.52 69.085 317.19 69.255 ;
      RECT 315.34 69.085 316.01 69.255 ;
      RECT 318.88 69.085 319.55 69.255 ;
      RECT 317.7 69.085 318.37 69.255 ;
      RECT 327.61 65.805 328.32 66.055 ;
      RECT 328.065 66.055 328.24 66.095 ;
      RECT 328.065 65.765 328.24 65.805 ;
      RECT 342.375 67.005 343.085 67.255 ;
      RECT 342.455 67.255 342.625 67.295 ;
      RECT 342.455 66.965 342.625 67.005 ;
      RECT 364.79 70.255 372.355 70.425 ;
      RECT 364.79 56.835 364.96 70.255 ;
      RECT 372.185 56.835 372.355 70.255 ;
      RECT 364.79 56.665 372.355 56.835 ;
      RECT 367.92 69.34 368.59 69.51 ;
      RECT 369.2 69.34 369.87 69.51 ;
      RECT 380.325 65.275 380.655 65.865 ;
      RECT 381.135 65.275 381.55 65.865 ;
      RECT 386.27 67.055 386.6 67.705 ;
      RECT 387.53 67.055 387.86 67.705 ;
      RECT 386.9 67.055 387.23 67.705 ;
      RECT 388.79 67.055 389.12 67.705 ;
      RECT 388.16 67.055 388.49 67.705 ;
      RECT 389.42 67.055 389.75 67.705 ;
      RECT 390.05 67.055 390.38 67.705 ;
      RECT 386.27 68.085 386.6 68.735 ;
      RECT 386.9 68.085 387.23 68.735 ;
      RECT 387.53 68.085 387.86 68.735 ;
      RECT 388.79 68.085 389.12 68.735 ;
      RECT 388.16 68.085 388.49 68.735 ;
      RECT 389.42 68.085 389.75 68.735 ;
      RECT 390.05 68.085 390.38 68.735 ;
      RECT 390.68 67.055 391.01 67.705 ;
      RECT 391.31 67.055 391.64 67.705 ;
      RECT 391.94 67.055 392.27 67.705 ;
      RECT 233.015 71.015 233.545 71.185 ;
      RECT 233.21 71.185 233.38 73.635 ;
      RECT 233.21 68.885 233.38 71.015 ;
      RECT 231.46 71.015 231.99 71.185 ;
      RECT 231.65 71.185 231.82 73.635 ;
      RECT 231.65 68.885 231.82 71.015 ;
      RECT 238.68 72.535 239.21 72.705 ;
      RECT 237.12 72.535 237.65 72.705 ;
      RECT 235.56 72.535 236.09 72.705 ;
      RECT 240.24 72.535 240.77 72.705 ;
      RECT 238.87 72.705 239.04 73.635 ;
      RECT 237.31 72.705 237.48 73.635 ;
      RECT 235.75 72.705 235.92 73.635 ;
      RECT 240.43 72.705 240.6 73.635 ;
      RECT 235.295 68.205 241.065 68.555 ;
      RECT 238.87 68.555 239.04 72.535 ;
      RECT 237.31 68.555 237.48 72.535 ;
      RECT 235.75 68.555 235.92 72.535 ;
      RECT 240.43 68.555 240.6 72.535 ;
      RECT 234.965 71.015 235.495 71.185 ;
      RECT 234.97 71.185 235.14 73.635 ;
      RECT 234.97 68.885 235.14 71.015 ;
      RECT 237.895 71.015 238.425 71.185 ;
      RECT 238.09 71.185 238.26 73.635 ;
      RECT 238.09 68.885 238.26 71.015 ;
      RECT 236.335 71.015 236.865 71.185 ;
      RECT 236.53 71.185 236.7 73.635 ;
      RECT 236.53 68.885 236.7 71.015 ;
      RECT 239.455 71.015 239.985 71.185 ;
      RECT 239.65 71.185 239.82 73.635 ;
      RECT 239.65 68.885 239.82 71.015 ;
      RECT 241.235 68.205 248.29 68.385 ;
      RECT 242.52 68.385 248.29 68.555 ;
      RECT 241.235 68.385 241.405 68.885 ;
      RECT 241.21 73.345 241.38 73.635 ;
      RECT 240.845 71.015 241.405 71.185 ;
      RECT 241.21 71.185 241.405 73.345 ;
      RECT 241.21 68.885 241.405 71.015 ;
      RECT 244.53 68.555 244.7 73.635 ;
      RECT 242.97 68.555 243.14 73.635 ;
      RECT 247.65 68.555 247.82 73.635 ;
      RECT 246.09 68.555 246.26 73.635 ;
      RECT 241.7 72.305 242.36 73.635 ;
      RECT 241.7 71.24 242.62 72.305 ;
      RECT 241.7 68.635 242.36 71.04 ;
      RECT 241.7 71.04 242.69 71.24 ;
      RECT 243.75 68.885 243.92 73.635 ;
      RECT 245.31 68.885 245.48 73.635 ;
      RECT 249.55 71.415 250.44 72.305 ;
      RECT 249.55 72.305 250.36 72.365 ;
      RECT 249.55 70.86 250.36 71.415 ;
      RECT 249.7 72.365 250.36 73.61 ;
      RECT 249.7 68.925 250.36 70.86 ;
      RECT 249.7 68.635 249.87 68.925 ;
      RECT 248.655 68.205 249.325 68.555 ;
      RECT 251.12 70.655 251.995 71.185 ;
      RECT 251.12 71.185 251.63 72.25 ;
      RECT 250.16 68.375 250.91 68.545 ;
      RECT 250.16 68.205 250.83 68.375 ;
      RECT 248.43 68.885 248.6 73.635 ;
      RECT 249.21 68.885 249.38 73.635 ;
      RECT 246.87 68.885 247.04 73.635 ;
      RECT 250.53 73.49 251.14 73.66 ;
      RECT 250.97 72.935 251.5 73.105 ;
      RECT 250.53 73.66 250.7 73.93 ;
      RECT 250.97 73.105 251.14 73.49 ;
      RECT 250.97 72.6 251.14 72.935 ;
      RECT 250.025 74 250.7 74.17 ;
      RECT 250.445 74.17 250.7 74.2 ;
      RECT 250.445 73.93 250.7 74 ;
      RECT 250.445 74.76 250.73 75.77 ;
      RECT 250.445 74.2 250.615 74.76 ;
      RECT 252.39 74 252.98 74.17 ;
      RECT 252.39 68.925 252.74 74 ;
      RECT 255.905 70.2 256.435 70.37 ;
      RECT 256 70.37 256.17 73.215 ;
      RECT 256 69.485 256.17 70.2 ;
      RECT 254.6 69.125 255.65 69.295 ;
      RECT 252.96 71.415 253.85 72.305 ;
      RECT 252.96 72.305 253.49 72.365 ;
      RECT 252.96 69.125 253.49 71.415 ;
      RECT 253.68 72.305 253.85 73.575 ;
      RECT 253.68 68.635 253.85 71.415 ;
      RECT 251.92 68.205 252.59 68.545 ;
      RECT 251.75 72.6 251.97 73.61 ;
      RECT 251.8 71.38 251.97 72.6 ;
      RECT 256.605 68.81 257.855 69.7 ;
      RECT 256.605 69.7 257.795 73.365 ;
      RECT 260.44 71.35 264.17 71.52 ;
      RECT 260.445 70.985 264.17 71.35 ;
      RECT 260.485 68.23 264.255 68.385 ;
      RECT 260.445 68.4 264.215 68.555 ;
      RECT 260.445 68.385 264.255 68.4 ;
      RECT 260.105 68.62 260.275 71.13 ;
      RECT 261.63 74 262.16 74.17 ;
      RECT 261.63 75.88 264.155 76.05 ;
      RECT 261.63 72.25 261.8 74 ;
      RECT 261.63 74.17 261.8 75.88 ;
      RECT 262.58 76.05 262.75 77.23 ;
      RECT 263.825 75.18 264.155 75.88 ;
      RECT 258.515 71.44 259.405 72.33 ;
      RECT 258.555 68.46 259.405 71.44 ;
      RECT 258.555 72.33 259.405 72.45 ;
      RECT 258.555 72.45 260.395 73.365 ;
      RECT 261.05 71.775 261.22 74.94 ;
      RECT 265.455 70.675 266.045 70.845 ;
      RECT 265.635 68.4 266.045 70.675 ;
      RECT 265.15 68.23 267.45 68.4 ;
      RECT 263.625 68.725 264.555 69.905 ;
      RECT 263.625 69.905 264.155 70.075 ;
      RECT 264.385 68.62 264.555 68.725 ;
      RECT 265.21 72.49 267.105 74.94 ;
      RECT 265.265 71.415 267.105 72.49 ;
      RECT 266.215 68.62 266.385 71.415 ;
      RECT 264.935 70.305 265.465 70.475 ;
      RECT 264.935 70.475 265.105 71.33 ;
      RECT 264.935 68.62 265.105 70.305 ;
      RECT 268.325 68.23 271.04 68.555 ;
      RECT 267.345 70.675 267.875 70.845 ;
      RECT 267.495 70.845 267.665 71.33 ;
      RECT 267.495 68.62 267.665 70.675 ;
      RECT 268.035 69.905 268.565 70.075 ;
      RECT 268.045 70.075 268.215 71.66 ;
      RECT 268.045 68.95 268.215 69.905 ;
      RECT 268.635 70.675 269.165 70.845 ;
      RECT 268.825 70.845 268.995 71.66 ;
      RECT 268.825 68.95 268.995 70.675 ;
      RECT 156.46 71.015 156.99 71.185 ;
      RECT 156.625 71.185 156.795 73.635 ;
      RECT 156.625 68.885 156.795 71.015 ;
      RECT 158.015 71.015 158.545 71.185 ;
      RECT 158.185 71.185 158.355 73.635 ;
      RECT 158.185 68.885 158.355 71.015 ;
      RECT 162.025 67.885 162.555 68.055 ;
      RECT 162.08 66.015 162.45 67.885 ;
      RECT 163.36 68.205 166.07 68.375 ;
      RECT 163.675 70.335 164.205 70.505 ;
      RECT 165.23 70.335 165.76 70.505 ;
      RECT 163.845 70.505 164.015 73.635 ;
      RECT 165.405 70.505 165.575 73.635 ;
      RECT 163.845 68.375 164.015 70.335 ;
      RECT 165.405 68.375 165.575 70.335 ;
      RECT 160.245 71.415 160.805 72.305 ;
      RECT 160.245 72.305 160.695 74.515 ;
      RECT 160.245 68.885 160.695 71.415 ;
      RECT 160.245 74.515 160.415 74.525 ;
      RECT 161.855 71.415 162.745 72.305 ;
      RECT 162.575 72.305 162.745 73.575 ;
      RECT 162.575 68.635 162.745 71.415 ;
      RECT 162.085 72.305 162.255 73.635 ;
      RECT 162.085 68.885 162.255 71.415 ;
      RECT 163.065 71.015 163.595 71.185 ;
      RECT 163.065 71.185 163.235 73.635 ;
      RECT 163.065 68.885 163.235 71.015 ;
      RECT 159.545 71.015 160.075 71.185 ;
      RECT 159.745 71.185 159.915 73.635 ;
      RECT 159.745 68.885 159.915 71.015 ;
      RECT 161.135 71.015 161.665 71.185 ;
      RECT 161.305 71.185 161.475 73.635 ;
      RECT 161.305 68.885 161.475 71.015 ;
      RECT 164.455 71.015 164.985 71.185 ;
      RECT 164.625 71.185 164.795 73.635 ;
      RECT 164.625 68.885 164.795 71.015 ;
      RECT 166.015 71.015 166.545 71.185 ;
      RECT 167.575 71.015 168.105 71.185 ;
      RECT 168.945 71.015 169.475 71.185 ;
      RECT 166.24 68.205 169.475 68.375 ;
      RECT 166.24 68.375 166.41 68.885 ;
      RECT 167.745 71.185 167.915 73.635 ;
      RECT 166.185 71.185 166.41 73.345 ;
      RECT 166.185 68.885 166.41 71.015 ;
      RECT 169.305 71.185 169.475 73.635 ;
      RECT 166.185 73.345 166.355 73.635 ;
      RECT 167.745 68.375 167.915 71.015 ;
      RECT 169.305 68.375 169.475 71.015 ;
      RECT 169.855 69.905 170.385 70.075 ;
      RECT 169.855 70.075 170.025 73.635 ;
      RECT 169.855 68.885 170.025 69.905 ;
      RECT 168.35 69.905 168.88 70.075 ;
      RECT 168.525 68.885 168.695 69.905 ;
      RECT 168.525 70.075 168.695 74.525 ;
      RECT 166.795 69.905 167.325 70.075 ;
      RECT 166.965 70.075 167.135 73.635 ;
      RECT 166.965 68.885 167.135 69.905 ;
      RECT 170.635 70.685 170.86 71.225 ;
      RECT 170.635 71.225 170.805 73.635 ;
      RECT 170.635 68.885 170.805 70.685 ;
      RECT 171.055 72.535 171.585 72.705 ;
      RECT 171.415 72.705 171.585 73.635 ;
      RECT 171.415 68.885 171.585 72.535 ;
      RECT 221.9 71.015 222.43 71.185 ;
      RECT 223.46 71.015 223.99 71.185 ;
      RECT 220.53 71.015 221.06 71.185 ;
      RECT 220.53 68.205 223.765 68.375 ;
      RECT 222.09 71.185 222.26 73.635 ;
      RECT 223.595 68.375 223.765 68.885 ;
      RECT 220.53 71.185 220.7 73.635 ;
      RECT 223.595 71.185 223.82 73.345 ;
      RECT 223.595 68.885 223.82 71.015 ;
      RECT 223.65 73.345 223.82 73.635 ;
      RECT 222.09 68.375 222.26 71.015 ;
      RECT 220.53 68.375 220.7 71.015 ;
      RECT 219.62 69.905 220.15 70.075 ;
      RECT 219.98 70.075 220.15 73.635 ;
      RECT 219.98 68.885 220.15 69.905 ;
      RECT 219.145 70.685 219.37 71.225 ;
      RECT 219.2 71.225 219.37 73.635 ;
      RECT 219.2 68.885 219.37 70.685 ;
      RECT 218.42 72.535 218.95 72.705 ;
      RECT 218.42 72.705 218.59 73.635 ;
      RECT 218.42 68.885 218.59 72.535 ;
      RECT 221.125 69.905 221.655 70.075 ;
      RECT 221.31 68.885 221.48 69.905 ;
      RECT 221.31 70.075 221.48 74.525 ;
      RECT 227.45 67.885 227.98 68.055 ;
      RECT 227.555 66.015 227.925 67.885 ;
      RECT 223.935 68.205 226.645 68.375 ;
      RECT 225.8 70.335 226.33 70.505 ;
      RECT 224.245 70.335 224.775 70.505 ;
      RECT 225.99 70.505 226.16 73.635 ;
      RECT 224.43 70.505 224.6 73.635 ;
      RECT 225.99 68.375 226.16 70.335 ;
      RECT 224.43 68.375 224.6 70.335 ;
      RECT 228.075 68.205 233.845 68.525 ;
      RECT 227.26 71.415 228.15 72.305 ;
      RECT 227.26 72.305 227.43 73.575 ;
      RECT 227.26 68.635 227.43 71.415 ;
      RECT 227.75 72.305 227.92 73.635 ;
      RECT 227.75 68.885 227.92 71.415 ;
      RECT 226.41 71.015 226.94 71.185 ;
      RECT 226.77 71.185 226.94 73.635 ;
      RECT 226.77 68.885 226.94 71.015 ;
      RECT 222.68 69.905 223.21 70.075 ;
      RECT 222.87 70.075 223.04 73.635 ;
      RECT 222.87 68.885 223.04 69.905 ;
      RECT 225.02 71.015 225.55 71.185 ;
      RECT 225.21 71.185 225.38 73.635 ;
      RECT 225.21 68.885 225.38 71.015 ;
      RECT 228.34 71.015 228.87 71.185 ;
      RECT 228.53 71.185 228.7 73.635 ;
      RECT 228.53 68.885 228.7 71.015 ;
      RECT 229.2 71.415 229.76 72.305 ;
      RECT 229.31 72.305 229.76 74.515 ;
      RECT 229.31 68.885 229.76 71.415 ;
      RECT 229.59 74.515 229.76 74.525 ;
      RECT 230.17 74.255 236.61 74.505 ;
      RECT 233.755 71.415 234.65 72.305 ;
      RECT 233.99 72.305 234.65 74.255 ;
      RECT 233.99 68.635 234.65 71.415 ;
      RECT 230.87 68.885 231.04 74.255 ;
      RECT 232.43 68.885 232.6 74.255 ;
      RECT 229.93 71.015 230.46 71.185 ;
      RECT 230.09 71.185 230.26 73.635 ;
      RECT 230.09 68.885 230.26 71.015 ;
      RECT 122.13 72.55 122.695 75.51 ;
      RECT 122.13 75.51 122.795 82.88 ;
      RECT 121.215 72.31 121.585 73.155 ;
      RECT 121.1 72.14 121.77 72.31 ;
      RECT 121.44 69.905 121.97 70.075 ;
      RECT 121.79 70.075 121.96 71.66 ;
      RECT 121.79 68.95 121.96 69.905 ;
      RECT 120.84 70.675 121.37 70.845 ;
      RECT 121.01 70.845 121.18 71.66 ;
      RECT 121.01 68.95 121.18 70.675 ;
      RECT 125.835 71.35 129.565 71.52 ;
      RECT 125.835 70.985 129.56 71.35 ;
      RECT 125.75 68.23 129.52 68.385 ;
      RECT 125.79 68.4 129.56 68.555 ;
      RECT 125.75 68.385 129.56 68.4 ;
      RECT 129.73 68.62 129.9 71.13 ;
      RECT 125.45 70.12 125.62 71.945 ;
      RECT 125.45 68.725 126.38 69.905 ;
      RECT 125.85 69.905 126.38 70.075 ;
      RECT 125.45 68.62 125.62 68.725 ;
      RECT 124.54 70.305 125.07 70.475 ;
      RECT 124.9 70.475 125.07 71.33 ;
      RECT 124.9 68.62 125.07 70.305 ;
      RECT 125.07 75.57 125.6 75.74 ;
      RECT 125.355 75.74 125.525 77.23 ;
      RECT 125.355 72.25 125.525 75.57 ;
      RECT 126.305 71.775 126.475 74.96 ;
      RECT 127.845 74 128.375 74.17 ;
      RECT 125.85 75.88 128.375 76.05 ;
      RECT 128.205 72.25 128.375 74 ;
      RECT 128.205 74.17 128.375 75.88 ;
      RECT 127.255 76.05 127.425 77.23 ;
      RECT 125.85 75.18 126.18 75.88 ;
      RECT 130.6 71.44 131.49 72.33 ;
      RECT 130.6 68.46 131.45 71.44 ;
      RECT 130.6 72.33 131.45 72.45 ;
      RECT 129.61 72.45 131.45 73.365 ;
      RECT 128.785 71.775 128.955 74.94 ;
      RECT 133.57 70.2 134.1 70.37 ;
      RECT 133.835 70.37 134.005 73.215 ;
      RECT 133.835 69.485 134.005 70.2 ;
      RECT 134.355 69.125 135.405 69.295 ;
      RECT 132.15 68.81 133.4 69.7 ;
      RECT 132.21 69.7 133.4 73.365 ;
      RECT 137.025 74 137.615 74.17 ;
      RECT 137.265 68.925 137.615 74 ;
      RECT 136.155 71.415 137.045 72.305 ;
      RECT 136.515 72.305 137.045 72.365 ;
      RECT 136.515 69.125 137.045 71.415 ;
      RECT 136.155 72.305 136.325 73.575 ;
      RECT 136.155 68.635 136.325 71.415 ;
      RECT 138.01 70.655 138.885 71.185 ;
      RECT 138.375 71.185 138.885 72.25 ;
      RECT 137.415 68.205 138.085 68.545 ;
      RECT 138.035 72.6 138.255 73.61 ;
      RECT 138.035 71.38 138.205 72.6 ;
      RECT 139.565 71.415 140.455 72.305 ;
      RECT 139.645 72.305 140.455 72.365 ;
      RECT 139.645 70.86 140.455 71.415 ;
      RECT 139.645 72.365 140.305 73.61 ;
      RECT 139.645 68.925 140.305 70.86 ;
      RECT 140.135 68.635 140.305 68.925 ;
      RECT 140.68 68.205 141.35 68.555 ;
      RECT 139.095 68.375 139.845 68.545 ;
      RECT 139.175 68.205 139.845 68.375 ;
      RECT 141.405 68.885 141.575 73.635 ;
      RECT 140.625 68.885 140.795 73.635 ;
      RECT 138.865 73.49 139.475 73.66 ;
      RECT 138.505 72.935 139.035 73.105 ;
      RECT 139.305 73.66 139.475 73.93 ;
      RECT 138.865 73.105 139.035 73.49 ;
      RECT 138.865 72.6 139.035 72.935 ;
      RECT 139.305 74 139.98 74.17 ;
      RECT 139.305 74.17 139.56 74.2 ;
      RECT 139.305 73.93 139.56 74 ;
      RECT 139.275 74.76 139.56 75.77 ;
      RECT 139.39 74.2 139.56 74.76 ;
      RECT 141.715 68.205 148.77 68.385 ;
      RECT 141.715 68.385 147.485 68.555 ;
      RECT 148.6 68.385 148.77 68.885 ;
      RECT 148.625 73.345 148.795 73.635 ;
      RECT 148.6 71.015 149.16 71.185 ;
      RECT 148.6 71.185 148.795 73.345 ;
      RECT 148.6 68.885 148.795 71.015 ;
      RECT 142.185 68.555 142.355 73.635 ;
      RECT 145.305 68.555 145.475 73.635 ;
      RECT 143.745 68.555 143.915 73.635 ;
      RECT 146.865 68.555 147.035 73.635 ;
      RECT 146.085 68.885 146.255 73.635 ;
      RECT 144.525 68.885 144.695 73.635 ;
      RECT 142.965 68.885 143.135 73.635 ;
      RECT 147.385 71.24 148.305 72.305 ;
      RECT 147.645 72.305 148.305 73.635 ;
      RECT 147.645 68.635 148.305 71.04 ;
      RECT 147.315 71.04 148.305 71.24 ;
      RECT 149.235 72.535 149.765 72.705 ;
      RECT 150.795 72.535 151.325 72.705 ;
      RECT 152.355 72.535 152.885 72.705 ;
      RECT 153.915 72.535 154.445 72.705 ;
      RECT 149.405 72.705 149.575 73.635 ;
      RECT 150.965 72.705 151.135 73.635 ;
      RECT 152.525 72.705 152.695 73.635 ;
      RECT 154.085 72.705 154.255 73.635 ;
      RECT 148.94 68.205 154.71 68.555 ;
      RECT 149.405 68.555 149.575 72.535 ;
      RECT 150.965 68.555 151.135 72.535 ;
      RECT 152.525 68.555 152.695 72.535 ;
      RECT 154.085 68.555 154.255 72.535 ;
      RECT 151.58 71.015 152.11 71.185 ;
      RECT 151.745 71.185 151.915 73.635 ;
      RECT 151.745 68.885 151.915 71.015 ;
      RECT 153.14 71.015 153.67 71.185 ;
      RECT 153.305 71.185 153.475 73.635 ;
      RECT 153.305 68.885 153.475 71.015 ;
      RECT 150.02 71.015 150.55 71.185 ;
      RECT 150.185 71.185 150.355 73.635 ;
      RECT 150.185 68.885 150.355 71.015 ;
      RECT 156.16 68.205 161.93 68.525 ;
      RECT 153.395 74.255 159.835 74.505 ;
      RECT 155.355 71.415 156.25 72.305 ;
      RECT 155.355 72.305 156.015 74.255 ;
      RECT 155.355 68.635 156.015 71.415 ;
      RECT 157.405 68.885 157.575 74.255 ;
      RECT 158.965 68.885 159.135 74.255 ;
      RECT 154.51 71.015 155.04 71.185 ;
      RECT 154.865 71.185 155.035 73.635 ;
      RECT 154.865 68.885 155.035 71.015 ;
      RECT 468.85 69.675 471.42 69.925 ;
      RECT 469.045 64.31 469.215 68.14 ;
      RECT 466.925 57.59 467.455 57.76 ;
      RECT 466.845 61.385 467.375 61.555 ;
      RECT 467.205 57.76 467.455 61.14 ;
      RECT 467.205 61.14 467.375 61.385 ;
      RECT 469.045 57.31 469.215 61.14 ;
      RECT 470.2 64.605 470.76 64.925 ;
      RECT 470.43 64.925 470.6 69.325 ;
      RECT 470.43 64.575 470.6 64.605 ;
      RECT 470.655 63.895 471.325 64.065 ;
      RECT 470.735 62.855 471.265 63.895 ;
      RECT 470.655 61.385 471.325 61.555 ;
      RECT 470.735 61.555 471.265 62.595 ;
      RECT 469.705 63.895 470.375 64.065 ;
      RECT 469.705 61.385 470.375 61.555 ;
      RECT 9.35 65.275 9.68 65.865 ;
      RECT 8.455 65.275 8.87 65.865 ;
      RECT 17.65 70.255 25.215 70.425 ;
      RECT 17.65 56.835 17.82 70.255 ;
      RECT 25.045 56.835 25.215 70.255 ;
      RECT 17.65 56.665 25.215 56.835 ;
      RECT 21.415 69.34 22.085 69.51 ;
      RECT 20.135 69.34 20.805 69.51 ;
      RECT 46.92 67.005 47.63 67.255 ;
      RECT 47.38 67.255 47.55 67.295 ;
      RECT 47.38 66.965 47.55 67.005 ;
      RECT 61.685 65.805 62.395 66.055 ;
      RECT 61.765 66.055 61.94 66.095 ;
      RECT 61.765 65.765 61.94 65.805 ;
      RECT 70.455 69.085 71.125 69.255 ;
      RECT 71.635 69.085 72.305 69.255 ;
      RECT 72.815 69.085 73.485 69.255 ;
      RECT 73.995 69.085 74.665 69.255 ;
      RECT 81.95 65.155 82.12 67.865 ;
      RECT 83.23 65.155 83.4 67.865 ;
      RECT 88.19 71.685 90.21 72.435 ;
      RECT 84.51 65.155 84.68 67.865 ;
      RECT 85.79 65.155 85.96 67.865 ;
      RECT 87.07 65.155 87.24 67.865 ;
      RECT 88.35 65.155 88.52 67.865 ;
      RECT 89.63 65.155 89.8 67.865 ;
      RECT 90.91 65.155 91.08 67.865 ;
      RECT 92.19 65.155 92.36 67.865 ;
      RECT 102.815 68.255 102.985 73.625 ;
      RECT 109.255 68.255 109.425 73.625 ;
      RECT 115.695 68.255 115.865 73.625 ;
      RECT 103.395 68.255 103.565 73.355 ;
      RECT 108.675 68.255 108.845 73.355 ;
      RECT 106.915 68.255 107.085 73.355 ;
      RECT 105.155 68.255 105.325 73.355 ;
      RECT 102.815 68.085 115.865 68.255 ;
      RECT 112.475 68.255 112.645 73.355 ;
      RECT 110.715 68.255 110.885 73.355 ;
      RECT 114.235 68.255 114.405 73.355 ;
      RECT 104.275 69.905 104.81 70.075 ;
      RECT 104.275 68.605 104.445 69.905 ;
      RECT 104.275 70.075 104.445 73.355 ;
      RECT 105.855 69.905 106.385 70.075 ;
      RECT 106.035 68.605 106.205 69.905 ;
      RECT 106.035 70.075 106.205 74.765 ;
      RECT 105.765 74.765 106.205 74.935 ;
      RECT 105.765 74.935 105.935 77.475 ;
      RECT 107.435 69.905 107.965 70.075 ;
      RECT 107.795 70.075 107.965 73.355 ;
      RECT 107.795 68.605 107.965 69.905 ;
      RECT 109.835 69.905 110.365 70.075 ;
      RECT 113.355 74.34 115.835 74.595 ;
      RECT 111.415 69.905 111.945 70.075 ;
      RECT 113.175 69.905 113.705 70.075 ;
      RECT 114.755 69.905 115.285 70.075 ;
      RECT 109.835 68.605 110.005 69.905 ;
      RECT 109.835 70.075 110.005 73.815 ;
      RECT 113.355 73.985 113.525 74.34 ;
      RECT 109.835 73.815 113.525 73.985 ;
      RECT 111.595 68.605 111.765 69.905 ;
      RECT 113.355 68.605 113.525 69.905 ;
      RECT 111.595 70.075 111.765 73.815 ;
      RECT 115.115 68.605 115.285 69.905 ;
      RECT 115.115 70.075 115.285 74.34 ;
      RECT 113.355 70.075 113.525 73.815 ;
      RECT 113.905 74.595 114.075 77.475 ;
      RECT 115.665 74.595 115.835 77.475 ;
      RECT 118.235 73.325 118.765 73.495 ;
      RECT 118.315 71.96 118.92 72.25 ;
      RECT 118.315 72.25 118.525 72.82 ;
      RECT 118.235 73.495 118.525 77.57 ;
      RECT 118.235 72.82 118.525 73.325 ;
      RECT 118.63 69.905 119.2 70.075 ;
      RECT 118.63 70.075 118.92 71.96 ;
      RECT 118.63 68.95 118.92 69.905 ;
      RECT 117.975 68.49 118.145 72.305 ;
      RECT 117.12 72.545 117.835 78.155 ;
      RECT 117.12 78.57 117.835 82.85 ;
      RECT 102.545 74.4 102.715 78.155 ;
      RECT 110.715 74.4 110.885 78.155 ;
      RECT 108.955 74.4 109.125 78.155 ;
      RECT 112.475 74.4 112.645 78.155 ;
      RECT 102.545 78.155 117.835 78.57 ;
      RECT 107.195 74.4 107.365 78.155 ;
      RECT 118.965 68.23 121.68 68.555 ;
      RECT 122.555 68.23 124.855 68.4 ;
      RECT 123.96 70.675 124.55 70.845 ;
      RECT 123.96 68.4 124.37 70.675 ;
      RECT 122.13 70.675 122.66 70.845 ;
      RECT 122.34 70.845 122.51 71.33 ;
      RECT 122.34 68.62 122.51 70.675 ;
      RECT 122.9 72.49 124.795 74.94 ;
      RECT 122.9 71.415 124.74 72.49 ;
      RECT 123.62 68.62 123.79 71.415 ;
      RECT 119.12 72.14 120.81 72.31 ;
      RECT 119.455 72.31 119.825 73.155 ;
      RECT 120.335 72.31 120.705 73.155 ;
      RECT 120.055 69.905 120.585 70.075 ;
      RECT 120.23 70.075 120.4 71.66 ;
      RECT 120.23 68.95 120.4 69.905 ;
      RECT 119.28 70.305 119.81 70.475 ;
      RECT 119.45 70.475 119.62 71.66 ;
      RECT 119.45 68.95 119.62 70.305 ;
      RECT 119.115 72.82 119.285 77.57 ;
      RECT 119.805 73.325 120.335 73.495 ;
      RECT 119.995 73.495 120.165 77.57 ;
      RECT 119.995 72.82 120.165 73.325 ;
      RECT 121.395 73.325 121.925 73.495 ;
      RECT 121.755 73.495 121.925 77.57 ;
      RECT 121.755 72.82 121.925 73.325 ;
      RECT 120.875 72.82 121.045 77.57 ;
      RECT 398.15 86.51 398.33 97.43 ;
      RECT 412.235 75.415 412.415 86.33 ;
      RECT 423.64 86.33 424.78 86.51 ;
      RECT 424.6 75.415 424.78 86.33 ;
      RECT 424.6 97.61 424.78 108.715 ;
      RECT 423.64 97.43 424.78 97.61 ;
      RECT 424.6 86.51 424.78 97.43 ;
      RECT 412.235 86.51 412.415 97.43 ;
      RECT 412.235 97.61 412.415 108.715 ;
      RECT 424.6 64.13 424.78 75.235 ;
      RECT 398.15 108.715 424.78 108.895 ;
      RECT 410.82 63.95 413.945 64.13 ;
      RECT 401.43 63.95 405.34 64.13 ;
      RECT 407.66 64.38 411.39 64.55 ;
      RECT 410.12 63.505 410.65 64.38 ;
      RECT 403.38 64.38 407.11 64.55 ;
      RECT 405.51 63.505 406.04 64.38 ;
      RECT 406.21 63.95 409.95 64.13 ;
      RECT 408.98 61.405 416.99 61.81 ;
      RECT 413.26 64.38 416.99 64.55 ;
      RECT 414.185 63.505 414.715 64.38 ;
      RECT 417.56 64.38 419.25 64.55 ;
      RECT 417.56 63.505 418.09 64.38 ;
      RECT 414.99 63.95 417.39 64.13 ;
      RECT 418.26 63.95 419.67 64.13 ;
      RECT 419.84 64.38 421.53 64.55 ;
      RECT 419.84 63.505 420.37 64.38 ;
      RECT 421.85 64.38 423.81 64.55 ;
      RECT 421.85 63.505 422.38 64.38 ;
      RECT 420.54 63.95 421.68 64.13 ;
      RECT 430.48 63.64 430.81 64.33 ;
      RECT 429.71 63.64 430.04 64.33 ;
      RECT 436.31 63.64 436.64 64.33 ;
      RECT 434.33 63.64 434.66 64.33 ;
      RECT 431.25 63.64 431.58 64.33 ;
      RECT 432.02 63.64 432.35 64.33 ;
      RECT 432.79 63.64 433.12 64.33 ;
      RECT 433.56 63.64 433.89 64.33 ;
      RECT 435.1 63.64 435.43 64.33 ;
      RECT 437.08 63.64 437.41 64.33 ;
      RECT 440.16 63.64 440.49 64.33 ;
      RECT 439.39 63.64 439.72 64.33 ;
      RECT 440.93 63.64 441.26 64.33 ;
      RECT 441.7 63.64 442.03 64.33 ;
      RECT 438.62 63.64 438.95 64.33 ;
      RECT 437.85 63.64 438.18 64.33 ;
      RECT 444.03 59.42 446.83 59.59 ;
      RECT 444.12 58.64 446.83 58.81 ;
      RECT 444.03 57.86 446.83 58.03 ;
      RECT 453.17 64.575 453.34 69.325 ;
      RECT 453.755 64.605 454.315 64.925 ;
      RECT 453.95 64.925 454.12 69.325 ;
      RECT 453.95 64.575 454.12 64.605 ;
      RECT 453.395 63.56 453.765 63.895 ;
      RECT 453.24 63.895 453.91 64.065 ;
      RECT 458.635 66.28 459.145 66.61 ;
      RECT 458.725 63.56 459.095 66.28 ;
      RECT 453.395 63.19 459.095 63.56 ;
      RECT 453.395 61.555 453.765 61.89 ;
      RECT 453.24 61.385 453.91 61.555 ;
      RECT 458.635 58.84 459.145 59.17 ;
      RECT 458.725 59.17 459.095 61.89 ;
      RECT 453.395 61.89 459.095 62.26 ;
      RECT 457.755 58.84 458.265 59.17 ;
      RECT 457.825 57.365 458.195 58.84 ;
      RECT 457.825 57.195 458.355 57.365 ;
      RECT 457.485 57.62 457.655 58.67 ;
      RECT 458.365 57.66 458.535 58.67 ;
      RECT 459.245 57.365 459.415 58.67 ;
      RECT 458.885 57.195 459.415 57.365 ;
      RECT 455.145 64.605 455.705 64.925 ;
      RECT 455.35 64.925 455.52 69.325 ;
      RECT 455.35 64.575 455.52 64.605 ;
      RECT 455.94 65.185 456.475 65.505 ;
      RECT 456.13 65.505 456.3 69.325 ;
      RECT 456.13 64.575 456.3 65.185 ;
      RECT 454.415 65.765 454.98 66.085 ;
      RECT 454.57 66.085 454.74 69.325 ;
      RECT 454.57 64.575 454.74 65.765 ;
      RECT 457.03 63.895 457.655 64.065 ;
      RECT 457.03 63.865 457.2 63.895 ;
      RECT 457.03 69.045 457.655 70.055 ;
      RECT 457.03 64.065 457.2 69.045 ;
      RECT 459.645 63.365 460.175 63.535 ;
      RECT 459.805 63.535 460.175 70.225 ;
      RECT 459.805 63.36 460.175 63.365 ;
      RECT 458.635 70.225 460.175 70.555 ;
      RECT 455.575 63.895 456.245 64.065 ;
      RECT 455.575 61.385 456.245 61.555 ;
      RECT 454.625 63.895 455.295 64.065 ;
      RECT 454.625 61.385 455.295 61.555 ;
      RECT 462.425 63.895 462.955 64.065 ;
      RECT 462.425 64.065 462.935 64.145 ;
      RECT 462.425 63.815 462.935 63.895 ;
      RECT 461.545 63.815 462.055 64.145 ;
      RECT 461.615 68.48 462.145 68.65 ;
      RECT 461.615 64.145 461.985 68.48 ;
      RECT 462.425 61.385 462.955 61.555 ;
      RECT 462.425 61.555 462.935 61.635 ;
      RECT 462.425 61.305 462.935 61.385 ;
      RECT 463.035 68.48 463.565 68.65 ;
      RECT 463.035 64.31 463.205 68.48 ;
      RECT 462.155 64.615 462.325 67.325 ;
      RECT 461.18 64.31 461.445 67.325 ;
      RECT 461.18 63.795 461.35 64.31 ;
      RECT 462.155 58.125 462.325 60.835 ;
      RECT 461.18 58.125 461.445 61.14 ;
      RECT 461.18 61.14 461.35 61.655 ;
      RECT 467.555 63.815 468.065 64.145 ;
      RECT 467.625 64.145 467.995 68.14 ;
      RECT 468.435 63.895 468.945 64.145 ;
      RECT 468.415 62.855 468.945 63.895 ;
      RECT 467.555 61.305 468.065 61.635 ;
      RECT 467.625 57.31 467.995 61.305 ;
      RECT 468.435 61.305 468.945 61.555 ;
      RECT 468.415 61.555 468.945 62.595 ;
      RECT 469.485 65.185 470.045 65.505 ;
      RECT 469.65 65.505 469.82 69.325 ;
      RECT 469.65 64.575 469.82 65.185 ;
      RECT 471.21 64.575 471.38 69.325 ;
      RECT 466.925 67.69 467.455 67.86 ;
      RECT 466.845 63.895 467.375 64.065 ;
      RECT 467.205 64.31 467.455 67.69 ;
      RECT 467.205 64.065 467.375 64.31 ;
      RECT 468.165 64.425 468.615 68.415 ;
      RECT 467.245 68.415 469.1 68.665 ;
      RECT 468.85 68.665 469.1 69.675 ;
      RECT 280.395 62.955 281.115 63.285 ;
      RECT 282.235 61.505 282.605 67.585 ;
      RECT 282.165 67.585 282.675 67.915 ;
      RECT 282.145 61.175 282.675 61.345 ;
      RECT 282.165 61.345 282.675 61.505 ;
      RECT 283.255 61.505 283.625 67.585 ;
      RECT 283.185 61.175 283.695 61.505 ;
      RECT 283.185 67.585 283.695 67.915 ;
      RECT 281.355 61.505 281.725 67.585 ;
      RECT 281.285 61.175 281.795 61.505 ;
      RECT 281.285 67.585 281.795 67.915 ;
      RECT 284.065 61.175 284.575 61.505 ;
      RECT 284.065 67.585 284.575 67.915 ;
      RECT 283.975 66.375 284.505 66.545 ;
      RECT 284.135 66.545 284.505 67.585 ;
      RECT 284.135 61.505 284.505 66.375 ;
      RECT 285.295 61.675 285.465 67.42 ;
      RECT 285.635 61.505 286.005 67.585 ;
      RECT 285.565 61.175 286.075 61.505 ;
      RECT 285.565 67.585 286.075 67.915 ;
      RECT 281.895 61.675 282.065 66.145 ;
      RECT 282.845 61.675 283.015 62.725 ;
      RECT 284.745 61.675 284.915 62.725 ;
      RECT 283.795 61.675 283.965 66.145 ;
      RECT 286.175 61.675 286.345 62.725 ;
      RECT 280.945 64.405 281.115 67.42 ;
      RECT 282.845 64.405 283.015 67.115 ;
      RECT 282.845 62.955 283.015 63.285 ;
      RECT 282.845 63.905 283.015 64.235 ;
      RECT 284.745 64.405 284.915 67.42 ;
      RECT 284.745 63.905 284.915 64.235 ;
      RECT 284.745 62.955 284.915 63.285 ;
      RECT 286.175 64.405 286.345 67.115 ;
      RECT 286.175 63.905 286.345 64.235 ;
      RECT 286.175 62.955 286.345 63.285 ;
      RECT 287.055 61.675 287.225 67.415 ;
      RECT 288.63 61.675 288.8 62.955 ;
      RECT 287.935 62.955 288.8 63.285 ;
      RECT 286.445 61.175 286.955 61.505 ;
      RECT 286.515 61.505 286.885 67.585 ;
      RECT 286.445 67.585 286.955 67.915 ;
      RECT 287.325 61.175 287.835 61.505 ;
      RECT 287.395 61.505 287.765 67.585 ;
      RECT 287.325 67.585 287.835 67.915 ;
      RECT 287.935 61.675 288.105 62.725 ;
      RECT 296.805 57.44 296.975 62.29 ;
      RECT 296.025 64.435 297.59 64.605 ;
      RECT 296.025 64.605 296.535 67.865 ;
      RECT 303.58 59.195 303.75 61.905 ;
      RECT 299.365 57.44 299.535 62.29 ;
      RECT 300.735 57.44 300.905 62.29 ;
      RECT 299.955 57.44 300.125 62.29 ;
      RECT 303.58 58.695 303.75 59.025 ;
      RECT 303.58 57.745 303.75 58.075 ;
      RECT 298.085 57.44 298.255 62.29 ;
      RECT 307.93 59.195 308.1 61.905 ;
      RECT 306.81 59.195 306.98 61.905 ;
      RECT 305.05 59.195 305.22 61.905 ;
      RECT 307.93 58.695 308.1 59.025 ;
      RECT 307.93 57.745 308.1 58.075 ;
      RECT 305.05 58.695 305.22 59.025 ;
      RECT 306.81 58.695 306.98 59.025 ;
      RECT 305.05 57.745 305.22 58.075 ;
      RECT 306.81 57.745 306.98 58.075 ;
      RECT 309.165 64.605 309.675 67.865 ;
      RECT 308.11 64.435 309.675 64.605 ;
      RECT 311.45 59.195 311.62 61.905 ;
      RECT 309.69 59.195 309.86 61.905 ;
      RECT 309.69 58.695 309.86 59.025 ;
      RECT 311.45 58.695 311.62 59.025 ;
      RECT 309.69 57.745 309.86 58.075 ;
      RECT 311.45 57.745 311.62 58.075 ;
      RECT 316.52 58.375 317.19 58.545 ;
      RECT 315.34 58.375 316.01 58.545 ;
      RECT 317.7 58.375 318.37 58.545 ;
      RECT 318.88 58.375 319.55 58.545 ;
      RECT 320.79 57.285 320.96 59.995 ;
      RECT 320.955 61.64 321.125 64.35 ;
      RECT 321.345 61.25 322.015 61.42 ;
      RECT 321.415 61.235 321.945 61.25 ;
      RECT 322.625 61.25 323.295 61.42 ;
      RECT 322.695 61.235 323.225 61.25 ;
      RECT 323.35 57.285 323.52 59.995 ;
      RECT 323.515 61.64 323.685 64.35 ;
      RECT 322.07 57.285 322.24 59.995 ;
      RECT 322.235 61.64 322.405 64.35 ;
      RECT 343.925 65.035 344.635 65.285 ;
      RECT 344.005 65.285 344.175 65.325 ;
      RECT 344.005 64.995 344.175 65.035 ;
      RECT 360.43 57.4 361.1 57.57 ;
      RECT 360.5 57.39 361.03 57.4 ;
      RECT 359.15 57.4 359.82 57.57 ;
      RECT 359.22 57.39 359.75 57.4 ;
      RECT 361.32 57.98 361.49 62.83 ;
      RECT 358.76 57.98 358.93 62.83 ;
      RECT 360.04 58.08 360.21 62.83 ;
      RECT 366.62 63.27 367.29 63.44 ;
      RECT 366.25 64.05 366.42 68.9 ;
      RECT 366.25 57.685 366.42 62.535 ;
      RECT 367.9 63.27 369.85 63.44 ;
      RECT 367.92 57.265 368.59 57.435 ;
      RECT 369.2 57.265 369.87 57.435 ;
      RECT 370.46 63.27 371.13 63.44 ;
      RECT 371.37 64.05 371.54 68.9 ;
      RECT 371.37 57.685 371.54 62.535 ;
      RECT 370.09 64.05 370.26 68.9 ;
      RECT 368.81 64.05 368.98 68.9 ;
      RECT 367.53 64.05 367.7 68.9 ;
      RECT 370.09 57.685 370.26 62.535 ;
      RECT 368.81 57.685 368.98 62.535 ;
      RECT 367.53 57.685 367.7 62.535 ;
      RECT 399.1 61.405 407.11 61.81 ;
      RECT 399.1 64.38 402.83 64.55 ;
      RECT 400.73 63.505 401.26 64.38 ;
      RECT 398.15 63.95 400.56 64.13 ;
      RECT 422.55 63.95 424.78 64.13 ;
      RECT 398.15 64.13 398.33 75.235 ;
      RECT 398.15 75.235 400.29 75.415 ;
      RECT 412.235 64.13 412.415 75.235 ;
      RECT 410.2 75.235 414.45 75.415 ;
      RECT 410.2 86.33 414.45 86.51 ;
      RECT 410.2 97.43 414.45 97.61 ;
      RECT 423.64 75.235 424.78 75.415 ;
      RECT 398.15 86.33 400.29 86.51 ;
      RECT 398.15 75.415 398.33 86.33 ;
      RECT 398.15 97.61 398.33 108.715 ;
      RECT 398.15 97.43 400.29 97.61 ;
      RECT 259.775 61.505 260.145 67.585 ;
      RECT 259.705 61.175 260.215 61.505 ;
      RECT 259.705 67.585 260.215 67.915 ;
      RECT 260.655 61.505 261.025 67.585 ;
      RECT 260.585 61.175 261.095 61.505 ;
      RECT 260.585 67.585 261.095 67.915 ;
      RECT 259.855 59.125 264.365 60.315 ;
      RECT 260.09 59.115 264.22 59.125 ;
      RECT 257.605 61.675 257.775 63.495 ;
      RECT 261.265 61.675 261.985 62.725 ;
      RECT 259.365 61.675 259.535 62.74 ;
      RECT 260.315 61.675 260.485 66.145 ;
      RECT 262.765 61.675 262.935 66.145 ;
      RECT 257.605 64.405 257.775 67.115 ;
      RECT 261.265 62.955 261.985 63.285 ;
      RECT 261.265 63.905 261.985 64.235 ;
      RECT 259.365 62.91 259.535 63.285 ;
      RECT 259.365 64.405 259.535 67.115 ;
      RECT 259.365 63.905 259.535 64.235 ;
      RECT 261.265 64.405 261.435 67.42 ;
      RECT 261.815 64.405 261.985 67.42 ;
      RECT 267.645 61.505 268.015 67.585 ;
      RECT 267.575 61.175 268.085 61.505 ;
      RECT 268.455 61.175 268.965 61.505 ;
      RECT 268.365 66.745 268.895 66.915 ;
      RECT 268.525 66.915 268.895 67.585 ;
      RECT 268.525 61.505 268.895 66.745 ;
      RECT 267.575 67.585 268.965 67.915 ;
      RECT 264.055 61.505 264.425 67.585 ;
      RECT 263.985 61.175 264.495 61.505 ;
      RECT 263.985 67.585 264.495 67.915 ;
      RECT 265.815 61.505 266.185 67.585 ;
      RECT 265.745 61.175 266.255 61.505 ;
      RECT 265.745 67.585 266.255 67.915 ;
      RECT 264.595 61.675 264.765 67.415 ;
      RECT 266.355 61.675 266.525 67.415 ;
      RECT 264.935 61.505 265.305 67.585 ;
      RECT 264.865 61.175 265.375 61.505 ;
      RECT 264.865 67.585 265.375 67.915 ;
      RECT 266.695 61.505 267.065 67.585 ;
      RECT 266.625 61.175 267.135 61.505 ;
      RECT 266.625 67.585 267.135 67.915 ;
      RECT 263.715 61.675 263.885 62.725 ;
      RECT 265.475 61.675 265.645 62.725 ;
      RECT 267.235 61.675 267.405 62.725 ;
      RECT 268.185 61.675 268.355 66.145 ;
      RECT 263.715 64.405 263.885 67.115 ;
      RECT 263.715 62.955 263.885 63.285 ;
      RECT 263.715 63.905 263.885 64.235 ;
      RECT 265.475 64.405 265.645 67.115 ;
      RECT 265.475 63.905 265.645 64.235 ;
      RECT 265.475 62.955 265.645 63.285 ;
      RECT 267.235 64.405 267.405 67.115 ;
      RECT 267.235 62.955 267.405 63.285 ;
      RECT 267.235 63.905 267.405 64.235 ;
      RECT 273.17 61.8 273.34 67.42 ;
      RECT 272.63 61.505 273 67.585 ;
      RECT 272.56 61.175 273.07 61.505 ;
      RECT 272.56 67.59 273.95 67.92 ;
      RECT 273.44 61.175 273.95 61.505 ;
      RECT 272.56 67.585 273.07 67.59 ;
      RECT 273.44 67.585 273.95 67.59 ;
      RECT 273.51 64.235 273.88 67.585 ;
      RECT 273.51 61.505 273.88 64.025 ;
      RECT 273.51 64.025 274.77 64.235 ;
      RECT 274.6 64.235 274.77 67.42 ;
      RECT 274.6 61.675 274.77 64.025 ;
      RECT 270.87 61.505 271.24 67.585 ;
      RECT 270.8 61.175 271.31 61.505 ;
      RECT 270.8 67.585 271.31 67.915 ;
      RECT 271.41 61.675 271.58 67.415 ;
      RECT 271.75 61.505 272.12 67.585 ;
      RECT 271.68 61.175 272.19 61.505 ;
      RECT 271.68 67.585 272.19 67.915 ;
      RECT 269.135 61.675 269.305 62.725 ;
      RECT 270.53 61.675 270.7 62.725 ;
      RECT 269.72 61.675 269.89 62.955 ;
      RECT 269.135 62.955 270.7 63.285 ;
      RECT 274.05 61.675 274.22 63.855 ;
      RECT 272.29 61.675 272.46 62.74 ;
      RECT 274.095 57.325 274.265 60.405 ;
      RECT 269.72 67.115 269.89 67.415 ;
      RECT 269.135 63.905 270.7 64.235 ;
      RECT 269.72 64.235 270.7 67.115 ;
      RECT 269.135 64.405 269.305 67.42 ;
      RECT 274.05 64.405 274.22 67.115 ;
      RECT 272.29 62.91 272.46 63.285 ;
      RECT 272.29 64.405 272.46 67.115 ;
      RECT 272.29 63.905 272.46 64.235 ;
      RECT 276.36 61.8 276.53 67.42 ;
      RECT 275.75 67.585 276.26 67.915 ;
      RECT 275.82 61.605 276.19 67.585 ;
      RECT 275.82 61.505 276.35 61.605 ;
      RECT 275.75 61.175 276.26 61.435 ;
      RECT 275.75 61.435 276.35 61.505 ;
      RECT 276.7 61.505 277.07 67.585 ;
      RECT 276.63 67.585 277.14 67.915 ;
      RECT 276.565 61.065 277.095 61.175 ;
      RECT 276.63 61.235 277.14 61.505 ;
      RECT 276.565 61.175 277.14 61.235 ;
      RECT 278.975 61.505 279.345 67.585 ;
      RECT 278.905 61.175 279.415 61.505 ;
      RECT 278.905 67.585 279.415 67.915 ;
      RECT 279.515 61.675 279.685 67.415 ;
      RECT 279.785 61.175 280.295 61.505 ;
      RECT 279.855 61.505 280.225 67.515 ;
      RECT 279.855 67.515 280.385 67.585 ;
      RECT 279.785 67.685 280.295 67.915 ;
      RECT 279.785 67.585 280.385 67.685 ;
      RECT 274.94 61.505 275.31 67.585 ;
      RECT 274.87 61.175 275.38 61.505 ;
      RECT 274.87 67.585 275.38 67.915 ;
      RECT 275.48 61.675 275.65 62.74 ;
      RECT 275.555 57.305 275.725 60.405 ;
      RECT 277.24 61.675 277.41 63.495 ;
      RECT 277.825 61.675 277.995 62.955 ;
      RECT 277.825 62.955 278.805 63.285 ;
      RECT 280.395 61.675 281.115 62.725 ;
      RECT 278.635 61.675 278.805 62.725 ;
      RECT 275.48 62.91 275.65 63.285 ;
      RECT 275.48 64.405 275.65 67.115 ;
      RECT 275.48 63.905 275.65 64.235 ;
      RECT 277.825 67.115 277.995 67.415 ;
      RECT 277.825 63.905 278.805 67.115 ;
      RECT 277.24 64.405 277.41 67.115 ;
      RECT 280.395 64.235 280.565 67.115 ;
      RECT 280.395 63.905 281.115 64.235 ;
      RECT 237.26 60.665 237.79 60.835 ;
      RECT 237.445 64.405 237.615 67.115 ;
      RECT 245.725 61.8 245.895 67.42 ;
      RECT 243.415 61.8 243.585 67.42 ;
      RECT 242.875 61.505 243.245 67.585 ;
      RECT 242.805 61.175 243.315 61.505 ;
      RECT 243.685 61.175 244.195 61.505 ;
      RECT 243.755 63.695 244.285 63.865 ;
      RECT 242.805 67.585 243.315 67.59 ;
      RECT 242.805 67.59 244.195 67.915 ;
      RECT 243.685 67.585 244.195 67.59 ;
      RECT 243.755 63.865 244.125 67.585 ;
      RECT 243.755 61.505 244.125 63.695 ;
      RECT 245.185 61.505 245.555 67.585 ;
      RECT 245.115 61.175 245.625 61.505 ;
      RECT 245.115 67.585 245.625 67.915 ;
      RECT 245.185 61.075 245.355 61.175 ;
      RECT 240.165 61.505 240.535 67.585 ;
      RECT 240.095 67.585 240.605 67.915 ;
      RECT 240.075 61.285 240.605 61.455 ;
      RECT 240.095 61.455 240.605 61.505 ;
      RECT 240.095 61.175 240.605 61.285 ;
      RECT 241.115 61.505 241.485 67.585 ;
      RECT 241.045 61.175 241.555 61.505 ;
      RECT 241.045 67.585 241.555 67.915 ;
      RECT 241.655 61.675 241.825 67.415 ;
      RECT 241.995 61.505 242.365 67.585 ;
      RECT 241.925 67.585 242.435 67.915 ;
      RECT 241.91 61.26 242.44 61.43 ;
      RECT 241.925 61.43 242.435 61.505 ;
      RECT 241.925 61.175 242.435 61.26 ;
      RECT 240.775 61.675 240.945 62.725 ;
      RECT 242.535 61.675 242.705 62.74 ;
      RECT 244.295 61.645 244.675 61.815 ;
      RECT 244.365 61.26 244.895 61.43 ;
      RECT 244.505 61.43 244.675 61.645 ;
      RECT 244.295 61.815 244.465 63.495 ;
      RECT 244.845 61.675 245.015 63.495 ;
      RECT 246.065 61.505 246.435 67.585 ;
      RECT 245.995 67.585 246.505 67.915 ;
      RECT 245.995 61.345 246.505 61.505 ;
      RECT 245.83 61.175 246.505 61.345 ;
      RECT 240.775 64.405 240.945 67.115 ;
      RECT 240.775 63.905 240.945 64.235 ;
      RECT 240.775 62.955 240.945 63.285 ;
      RECT 242.535 62.91 242.705 63.285 ;
      RECT 242.535 64.405 242.705 67.115 ;
      RECT 242.535 63.905 242.705 64.235 ;
      RECT 244.845 64.405 245.015 67.115 ;
      RECT 244.295 64.405 244.465 67.115 ;
      RECT 248.915 61.8 249.085 67.42 ;
      RECT 249.255 61.505 249.625 67.585 ;
      RECT 249.185 61.175 249.695 61.505 ;
      RECT 248.305 61.175 248.815 61.505 ;
      RECT 249.185 67.585 249.695 67.59 ;
      RECT 248.305 67.59 249.695 67.915 ;
      RECT 248.305 67.585 248.815 67.59 ;
      RECT 248.375 63.865 248.745 67.585 ;
      RECT 248.375 61.505 248.745 63.695 ;
      RECT 247.485 63.695 248.745 63.865 ;
      RECT 247.485 63.865 247.655 67.42 ;
      RECT 247.485 61.675 247.655 63.695 ;
      RECT 250.065 61.175 250.575 61.505 ;
      RECT 250.065 67.585 250.575 67.915 ;
      RECT 249.885 63.455 250.505 63.625 ;
      RECT 250.135 63.625 250.505 67.585 ;
      RECT 250.135 61.505 250.505 63.455 ;
      RECT 250.675 61.675 250.845 67.415 ;
      RECT 251.015 61.505 251.385 67.585 ;
      RECT 250.945 61.175 251.455 61.505 ;
      RECT 250.945 67.585 251.455 67.915 ;
      RECT 246.875 61.175 247.385 61.505 ;
      RECT 246.785 63.455 247.315 63.625 ;
      RECT 246.875 67.585 247.385 67.915 ;
      RECT 246.945 63.625 247.315 67.585 ;
      RECT 246.945 61.505 247.315 63.455 ;
      RECT 246.605 61.675 246.775 62.74 ;
      RECT 248.035 61.675 248.205 63.495 ;
      RECT 248.495 57.305 248.665 60.405 ;
      RECT 249.795 61.675 249.965 62.74 ;
      RECT 249.955 57.325 250.125 60.405 ;
      RECT 251.555 61.675 251.725 62.725 ;
      RECT 246.605 62.91 246.775 63.285 ;
      RECT 246.605 64.405 246.775 67.115 ;
      RECT 246.605 63.905 246.775 64.235 ;
      RECT 248.035 64.405 248.205 67.115 ;
      RECT 249.795 62.91 249.965 63.285 ;
      RECT 249.795 64.405 249.965 67.115 ;
      RECT 249.795 63.905 249.965 64.235 ;
      RECT 251.555 64.405 251.725 67.115 ;
      RECT 251.555 63.905 251.725 64.235 ;
      RECT 251.555 62.955 251.725 63.285 ;
      RECT 253.255 61.175 253.765 61.505 ;
      RECT 253.325 61.505 253.695 67.585 ;
      RECT 253.255 67.585 253.765 67.915 ;
      RECT 252.375 61.175 252.885 61.505 ;
      RECT 252.445 61.505 252.815 67.585 ;
      RECT 252.375 67.585 252.885 67.915 ;
      RECT 256.445 61.175 256.955 61.505 ;
      RECT 256.515 61.505 256.885 67.585 ;
      RECT 256.445 67.585 256.955 67.915 ;
      RECT 252.105 64.405 252.275 67.115 ;
      RECT 253.865 62.91 254.035 63.285 ;
      RECT 253.865 64.405 254.035 67.115 ;
      RECT 252.985 61.8 253.155 67.42 ;
      RECT 252.105 61.675 252.275 63.495 ;
      RECT 253.865 61.675 254.035 62.74 ;
      RECT 253.865 63.905 254.035 64.235 ;
      RECT 257.055 61.675 257.225 67.42 ;
      RECT 256.175 61.675 256.345 62.725 ;
      RECT 256.175 64.405 256.345 67.115 ;
      RECT 256.175 63.905 256.345 64.235 ;
      RECT 256.175 62.955 256.345 63.285 ;
      RECT 258.485 61.8 258.655 67.42 ;
      RECT 258.825 61.505 259.195 67.585 ;
      RECT 258.755 61.175 259.265 61.505 ;
      RECT 258.755 67.585 259.265 67.915 ;
      RECT 257.945 61.505 258.315 67.585 ;
      RECT 257.875 61.175 258.385 61.505 ;
      RECT 257.875 67.585 258.385 67.915 ;
      RECT 263.105 61.505 263.475 67.585 ;
      RECT 263.035 61.175 263.545 61.505 ;
      RECT 262.225 61.505 262.595 67.585 ;
      RECT 262.155 61.175 262.665 61.505 ;
      RECT 262.14 67.915 262.67 68.055 ;
      RECT 262.14 67.885 263.545 67.915 ;
      RECT 262.155 67.585 263.545 67.885 ;
      RECT 224.295 67.585 224.805 67.915 ;
      RECT 224.365 63.455 224.985 63.625 ;
      RECT 224.365 63.625 224.735 67.585 ;
      RECT 224.365 61.505 224.735 63.455 ;
      RECT 226.055 61.175 226.565 61.505 ;
      RECT 226.125 61.505 226.495 67.515 ;
      RECT 226.125 67.515 226.655 67.585 ;
      RECT 226.055 67.685 226.565 67.915 ;
      RECT 226.055 67.585 226.655 67.685 ;
      RECT 223.415 61.175 223.925 61.505 ;
      RECT 223.325 63.695 223.855 63.865 ;
      RECT 223.415 67.585 223.925 67.915 ;
      RECT 223.485 63.865 223.855 67.585 ;
      RECT 223.485 61.505 223.855 63.695 ;
      RECT 228.355 61.255 228.885 61.425 ;
      RECT 228.35 67.585 228.86 67.915 ;
      RECT 228.435 61.425 228.805 67.585 ;
      RECT 228.435 61.175 228.805 61.255 ;
      RECT 223.145 61.675 223.315 63.495 ;
      RECT 224.905 61.675 225.075 62.74 ;
      RECT 224.035 58.45 225.565 59.2 ;
      RECT 224.275 59.2 225.325 60.405 ;
      RECT 224.275 57.305 225.325 58.45 ;
      RECT 226.665 61.675 226.835 63.495 ;
      RECT 227.555 61.505 227.925 61.885 ;
      RECT 227.465 61.255 227.995 61.425 ;
      RECT 227.485 61.425 227.995 61.505 ;
      RECT 227.485 61.175 227.995 61.255 ;
      RECT 227.215 63.695 227.745 63.865 ;
      RECT 227.215 61.675 227.385 63.695 ;
      RECT 227.215 63.865 227.385 67.115 ;
      RECT 226.925 57.305 227.095 60.405 ;
      RECT 228.095 61.675 228.265 62.685 ;
      RECT 228.385 57.325 228.555 60.405 ;
      RECT 223.145 64.405 223.315 67.115 ;
      RECT 224.905 62.91 225.075 63.285 ;
      RECT 224.905 64.405 225.075 67.115 ;
      RECT 224.905 63.905 225.075 64.235 ;
      RECT 226.665 64.405 226.835 67.115 ;
      RECT 228.095 63.905 228.265 64.235 ;
      RECT 228.095 62.955 228.265 63.285 ;
      RECT 228.095 64.405 228.265 67.115 ;
      RECT 229.73 57.3 229.9 60.3 ;
      RECT 230.535 60.665 232.565 60.835 ;
      RECT 230.195 63.695 230.725 63.865 ;
      RECT 230.195 63.865 230.525 63.965 ;
      RECT 230.195 63.455 230.525 63.695 ;
      RECT 230.115 61.255 230.645 61.425 ;
      RECT 230.195 61.505 230.565 61.88 ;
      RECT 230.125 61.425 230.635 61.505 ;
      RECT 230.125 61.175 230.635 61.255 ;
      RECT 231.005 61.285 231.535 61.455 ;
      RECT 231.02 67.585 231.53 67.915 ;
      RECT 231.005 61.455 231.515 61.505 ;
      RECT 231.005 61.175 231.515 61.285 ;
      RECT 231.075 61.505 231.445 67.585 ;
      RECT 232.135 63.415 232.665 63.585 ;
      RECT 232.495 61.675 232.665 63.415 ;
      RECT 232.495 63.585 232.665 67.115 ;
      RECT 232.775 60.665 233.445 60.835 ;
      RECT 231.615 62.955 231.785 63.285 ;
      RECT 229.855 65.585 230.385 65.755 ;
      RECT 229.855 65.755 230.025 67.42 ;
      RECT 229.855 61.675 230.025 65.585 ;
      RECT 231.615 63.905 231.785 64.235 ;
      RECT 229.155 63.415 229.685 63.585 ;
      RECT 229.24 67.585 229.75 67.915 ;
      RECT 229.315 63.585 229.685 67.585 ;
      RECT 231.615 61.675 231.785 62.725 ;
      RECT 228.975 64.405 229.145 67.115 ;
      RECT 230.735 64.405 230.905 67.115 ;
      RECT 231.615 64.405 231.785 67.115 ;
      RECT 233.725 60.665 236.835 60.835 ;
      RECT 234.18 67.585 234.69 67.915 ;
      RECT 234.17 61.285 234.705 61.455 ;
      RECT 234.195 61.455 234.705 61.505 ;
      RECT 234.195 61.175 234.705 61.285 ;
      RECT 234.265 61.505 234.635 67.585 ;
      RECT 233.045 63.415 233.575 63.585 ;
      RECT 233.045 61.675 233.215 63.415 ;
      RECT 233.045 63.585 233.215 67.115 ;
      RECT 233.925 62.955 234.095 63.285 ;
      RECT 233.925 63.905 234.095 64.235 ;
      RECT 233.925 61.675 234.095 62.725 ;
      RECT 233.925 64.405 234.095 67.115 ;
      RECT 234.985 63.695 235.515 63.865 ;
      RECT 235.185 63.865 235.515 63.965 ;
      RECT 235.185 63.455 235.515 63.695 ;
      RECT 235.065 61.255 235.595 61.425 ;
      RECT 235.145 61.505 235.515 61.88 ;
      RECT 235.075 61.425 235.585 61.505 ;
      RECT 235.075 61.175 235.585 61.255 ;
      RECT 236.825 61.255 237.355 61.425 ;
      RECT 236.905 61.175 237.275 61.255 ;
      RECT 236.85 67.685 237.36 67.915 ;
      RECT 236.85 67.585 237.535 67.685 ;
      RECT 236.905 67.515 237.535 67.585 ;
      RECT 236.905 61.425 237.275 67.515 ;
      RECT 235.325 65.585 235.855 65.755 ;
      RECT 235.685 65.755 235.855 67.42 ;
      RECT 235.685 61.675 235.855 65.585 ;
      RECT 236.025 63.415 236.555 63.585 ;
      RECT 235.96 67.585 236.47 67.915 ;
      RECT 236.025 63.585 236.395 67.585 ;
      RECT 236.565 64.405 236.735 67.115 ;
      RECT 234.805 64.405 234.975 67.115 ;
      RECT 239.215 61.175 239.725 61.505 ;
      RECT 239.215 67.585 239.725 67.915 ;
      RECT 239.215 67.115 239.745 67.285 ;
      RECT 239.285 67.285 239.655 67.585 ;
      RECT 239.285 61.505 239.655 67.115 ;
      RECT 237.785 61.505 238.155 61.885 ;
      RECT 237.715 61.255 238.245 61.425 ;
      RECT 237.715 61.425 238.225 61.505 ;
      RECT 237.715 61.175 238.225 61.255 ;
      RECT 238.875 61.675 239.045 62.725 ;
      RECT 237.965 63.695 238.495 63.865 ;
      RECT 238.325 61.675 238.495 63.695 ;
      RECT 238.325 63.865 238.495 67.115 ;
      RECT 238.875 64.405 239.045 67.42 ;
      RECT 237.445 63.905 237.615 64.235 ;
      RECT 237.445 62.955 237.615 63.285 ;
      RECT 239.825 61.675 239.995 66.135 ;
      RECT 238.875 63.905 239.045 64.235 ;
      RECT 238.875 62.955 239.045 63.285 ;
      RECT 238.115 60.665 240.085 60.835 ;
      RECT 237.445 61.675 237.615 62.685 ;
      RECT 172.6 61.175 173.11 61.505 ;
      RECT 172.6 67.585 173.11 67.915 ;
      RECT 173.48 67.585 173.99 67.915 ;
      RECT 173.55 61.585 173.92 67.585 ;
      RECT 173.55 61.505 174.08 61.585 ;
      RECT 173.48 61.175 173.99 61.415 ;
      RECT 173.48 61.415 174.08 61.505 ;
      RECT 170.94 60.665 172.97 60.835 ;
      RECT 171.45 61.675 171.62 63.495 ;
      RECT 170.9 61.675 171.07 63.495 ;
      RECT 174.13 60.665 174.8 60.835 ;
      RECT 173.21 62.91 173.38 63.285 ;
      RECT 174.97 61.675 175.14 63.855 ;
      RECT 173.21 61.675 173.38 62.74 ;
      RECT 173.18 60.665 173.85 60.835 ;
      RECT 173.25 60.835 173.78 60.885 ;
      RECT 171.45 64.405 171.62 67.115 ;
      RECT 170.9 64.405 171.07 67.115 ;
      RECT 174.97 64.405 175.14 67.115 ;
      RECT 173.21 64.405 173.38 67.115 ;
      RECT 173.21 63.905 173.38 64.235 ;
      RECT 264.475 91.72 290.58 92.265 ;
      RECT 244.49 91.465 290.58 91.72 ;
      RECT 244.49 90.92 265.275 91.465 ;
      RECT 289.78 87.885 290.58 91.465 ;
      RECT 244.49 87.885 245.29 90.92 ;
      RECT 214.205 87.87 278.02 87.885 ;
      RECT 289.07 87.87 290.955 87.885 ;
      RECT 279.02 87.87 287.225 87.885 ;
      RECT 214.205 87.7 290.955 87.87 ;
      RECT 214.205 87.07 237.66 87.7 ;
      RECT 214.205 86.38 234.265 87.07 ;
      RECT 214.205 86.375 234.28 86.38 ;
      RECT 219.275 86.32 234.28 86.375 ;
      RECT 253.455 86.315 256.43 87.7 ;
      RECT 219.3 86.21 234.28 86.32 ;
      RECT 253.455 85.785 256.565 86.315 ;
      RECT 214.205 85.65 218.345 86.375 ;
      RECT 253.455 85.555 256.43 85.785 ;
      RECT 231.855 85.025 234.225 86.21 ;
      RECT 222.42 84.555 222.59 86.21 ;
      RECT 237.48 81.95 237.65 87.07 ;
      RECT 216.11 82.17 216.28 85.65 ;
      RECT 217.87 82.17 218.04 85.65 ;
      RECT 219.3 82.05 219.47 86.21 ;
      RECT 288.63 76.345 289.32 77.785 ;
      RECT 290.785 76.195 290.955 87.7 ;
      RECT 288.525 76.195 289.32 76.345 ;
      RECT 288.525 76.025 290.955 76.195 ;
      RECT 214.205 73.615 215.275 85.65 ;
      RECT 214.205 71.225 218.11 73.615 ;
      RECT 288.525 68.505 289.375 76.025 ;
      RECT 214.205 68.615 218.11 70.285 ;
      RECT 214.205 70.285 218.125 71.225 ;
      RECT 288.63 67.115 289.375 68.505 ;
      RECT 214.205 64.235 214.375 68.615 ;
      RECT 287.935 63.905 288.8 63.975 ;
      RECT 287.935 63.975 289.375 67.115 ;
      RECT 214.205 64.065 214.735 64.235 ;
      RECT 214.205 63.905 214.375 64.065 ;
      RECT 215.205 60.665 215.875 60.835 ;
      RECT 214.865 64.405 215.035 67.115 ;
      RECT 215.745 61.8 215.915 67.42 ;
      RECT 214.865 61.675 215.035 63.855 ;
      RECT 216.015 67.585 216.525 67.915 ;
      RECT 216.085 61.585 216.455 67.585 ;
      RECT 215.925 61.505 216.455 61.585 ;
      RECT 216.015 61.175 216.525 61.415 ;
      RECT 215.925 61.415 216.525 61.505 ;
      RECT 215.205 61.505 215.575 67.585 ;
      RECT 215.135 61.175 215.645 61.505 ;
      RECT 215.135 67.585 215.645 67.915 ;
      RECT 216.155 60.665 216.825 60.835 ;
      RECT 216.225 60.835 216.755 60.885 ;
      RECT 216.625 62.91 216.795 63.285 ;
      RECT 216.625 64.405 216.795 67.115 ;
      RECT 216.625 61.675 216.795 62.74 ;
      RECT 216.625 63.905 216.795 64.235 ;
      RECT 219.7 57.3 219.87 60.3 ;
      RECT 221.045 57.325 221.215 60.405 ;
      RECT 222.505 57.305 222.675 60.405 ;
      RECT 217.035 60.665 219.065 60.835 ;
      RECT 218.385 64.405 218.555 67.115 ;
      RECT 217.505 61.8 217.675 67.42 ;
      RECT 218.385 61.675 218.555 63.495 ;
      RECT 216.965 61.505 217.335 67.585 ;
      RECT 216.895 61.175 217.405 61.505 ;
      RECT 216.895 67.585 217.405 67.915 ;
      RECT 217.775 61.175 218.285 61.505 ;
      RECT 217.845 63.695 218.375 63.865 ;
      RECT 217.775 67.585 218.285 67.915 ;
      RECT 217.845 63.865 218.215 67.585 ;
      RECT 217.845 61.505 218.215 63.695 ;
      RECT 218.935 64.405 219.105 67.115 ;
      RECT 220.695 62.91 220.865 63.285 ;
      RECT 220.695 64.405 220.865 67.115 ;
      RECT 219.815 61.8 219.985 67.42 ;
      RECT 218.935 61.675 219.105 63.495 ;
      RECT 220.155 61.505 220.525 67.585 ;
      RECT 220.085 61.175 220.595 61.505 ;
      RECT 220.085 67.585 220.595 67.915 ;
      RECT 219.275 61.505 219.645 67.585 ;
      RECT 219.205 61.175 219.715 61.505 ;
      RECT 219.205 67.585 219.715 67.915 ;
      RECT 220.695 61.675 220.865 62.74 ;
      RECT 220.695 63.905 220.865 64.235 ;
      RECT 221.035 67.585 221.545 67.915 ;
      RECT 220.99 61.505 221.52 61.555 ;
      RECT 221.035 61.175 221.545 61.385 ;
      RECT 220.99 61.385 221.545 61.505 ;
      RECT 221.105 61.555 221.475 67.585 ;
      RECT 221.915 61.175 222.425 61.505 ;
      RECT 221.915 67.585 222.425 67.915 ;
      RECT 221.895 67.115 222.425 67.285 ;
      RECT 221.985 67.285 222.355 67.585 ;
      RECT 221.985 61.505 222.355 67.115 ;
      RECT 222.595 61.675 222.765 62.725 ;
      RECT 222.595 64.405 222.765 67.42 ;
      RECT 221.645 61.675 221.815 66.145 ;
      RECT 222.595 63.905 222.765 64.235 ;
      RECT 222.595 62.955 222.765 63.285 ;
      RECT 225.785 61.8 225.955 67.42 ;
      RECT 224.025 61.8 224.195 67.42 ;
      RECT 225.245 61.505 225.615 67.585 ;
      RECT 225.175 61.175 225.685 61.505 ;
      RECT 225.175 67.585 225.685 67.915 ;
      RECT 224.295 61.175 224.805 61.505 ;
      RECT 153.27 64.405 153.44 67.115 ;
      RECT 155.03 64.405 155.2 67.115 ;
      RECT 157.44 60.665 159.47 60.835 ;
      RECT 158.47 61.285 159 61.455 ;
      RECT 158.475 67.585 158.985 67.915 ;
      RECT 158.49 61.455 159 61.505 ;
      RECT 158.49 61.175 159 61.285 ;
      RECT 158.56 61.505 158.93 67.585 ;
      RECT 157.34 63.415 157.87 63.585 ;
      RECT 157.34 61.675 157.51 63.415 ;
      RECT 157.34 63.585 157.51 67.115 ;
      RECT 156.43 63.415 156.96 63.585 ;
      RECT 156.79 61.675 156.96 63.415 ;
      RECT 156.79 63.585 156.96 67.115 ;
      RECT 156.56 60.665 157.23 60.835 ;
      RECT 155.91 62.955 156.08 63.285 ;
      RECT 158.22 63.905 158.39 64.235 ;
      RECT 155.91 63.905 156.08 64.235 ;
      RECT 158.22 62.955 158.39 63.285 ;
      RECT 158.22 61.675 158.39 62.725 ;
      RECT 155.91 61.675 156.08 62.725 ;
      RECT 158.22 64.405 158.39 67.115 ;
      RECT 155.91 64.405 156.08 67.115 ;
      RECT 160.105 57.3 160.275 60.3 ;
      RECT 161.45 57.325 161.62 60.405 ;
      RECT 162.91 57.305 163.08 60.405 ;
      RECT 164.44 58.45 165.97 59.2 ;
      RECT 164.68 59.2 165.73 60.405 ;
      RECT 164.68 57.305 165.73 58.45 ;
      RECT 159.28 63.695 159.81 63.865 ;
      RECT 159.48 63.865 159.81 63.965 ;
      RECT 159.48 63.455 159.81 63.695 ;
      RECT 159.36 61.255 159.89 61.425 ;
      RECT 159.44 61.505 159.81 61.88 ;
      RECT 159.37 61.425 159.88 61.505 ;
      RECT 159.37 61.175 159.88 61.255 ;
      RECT 159.1 64.405 159.27 67.115 ;
      RECT 162.08 61.505 162.45 61.885 ;
      RECT 162.01 61.255 162.54 61.425 ;
      RECT 162.01 61.425 162.52 61.505 ;
      RECT 162.01 61.175 162.52 61.255 ;
      RECT 161.12 61.255 161.65 61.425 ;
      RECT 161.145 67.585 161.655 67.915 ;
      RECT 161.2 61.425 161.57 67.585 ;
      RECT 161.2 61.175 161.57 61.255 ;
      RECT 159.62 65.585 160.15 65.755 ;
      RECT 159.98 65.755 160.15 67.42 ;
      RECT 159.98 61.675 160.15 65.585 ;
      RECT 160.32 63.415 160.85 63.585 ;
      RECT 160.255 67.585 160.765 67.915 ;
      RECT 160.32 63.585 160.69 67.585 ;
      RECT 161.74 63.905 161.91 64.235 ;
      RECT 161.74 62.955 161.91 63.285 ;
      RECT 162.26 63.695 162.79 63.865 ;
      RECT 162.62 61.675 162.79 63.695 ;
      RECT 162.62 63.865 162.79 67.115 ;
      RECT 161.74 61.675 161.91 62.685 ;
      RECT 161.74 64.405 161.91 67.115 ;
      RECT 160.86 64.405 161.03 67.115 ;
      RECT 163.17 64.405 163.34 67.115 ;
      RECT 164.05 61.8 164.22 67.42 ;
      RECT 163.17 61.675 163.34 63.495 ;
      RECT 163.44 61.175 163.95 61.505 ;
      RECT 163.51 61.505 163.88 67.515 ;
      RECT 163.35 67.515 163.88 67.585 ;
      RECT 163.44 67.685 163.95 67.915 ;
      RECT 163.35 67.585 163.95 67.685 ;
      RECT 164.39 61.505 164.76 67.585 ;
      RECT 164.32 61.175 164.83 61.505 ;
      RECT 164.32 67.585 164.83 67.915 ;
      RECT 165.81 61.8 165.98 67.42 ;
      RECT 170.02 61.8 170.19 67.42 ;
      RECT 169.48 61.505 169.85 67.585 ;
      RECT 169.41 61.175 169.92 61.505 ;
      RECT 169.41 67.585 169.92 67.915 ;
      RECT 166.08 61.175 166.59 61.505 ;
      RECT 166.15 63.695 166.68 63.865 ;
      RECT 166.08 67.585 166.59 67.915 ;
      RECT 166.15 63.865 166.52 67.585 ;
      RECT 166.15 61.505 166.52 63.695 ;
      RECT 170.36 61.505 170.73 67.585 ;
      RECT 170.29 61.175 170.8 61.505 ;
      RECT 170.29 67.585 170.8 67.915 ;
      RECT 165.2 61.175 165.71 61.505 ;
      RECT 165.2 67.585 165.71 67.915 ;
      RECT 165.02 63.455 165.64 63.625 ;
      RECT 165.27 63.625 165.64 67.585 ;
      RECT 165.27 61.505 165.64 63.455 ;
      RECT 167.58 61.175 168.09 61.505 ;
      RECT 167.58 67.585 168.09 67.915 ;
      RECT 167.58 67.115 168.11 67.285 ;
      RECT 167.65 67.285 168.02 67.585 ;
      RECT 167.65 61.505 168.02 67.115 ;
      RECT 168.46 67.585 168.97 67.915 ;
      RECT 168.53 61.555 168.9 67.585 ;
      RECT 168.485 61.505 169.015 61.555 ;
      RECT 168.46 61.175 168.97 61.385 ;
      RECT 168.46 61.385 169.015 61.505 ;
      RECT 167.33 57.305 167.5 60.405 ;
      RECT 170.135 57.3 170.305 60.3 ;
      RECT 168.79 57.325 168.96 60.405 ;
      RECT 164.93 61.675 165.1 62.74 ;
      RECT 166.69 61.675 166.86 63.495 ;
      RECT 167.24 61.675 167.41 62.725 ;
      RECT 169.14 61.675 169.31 62.74 ;
      RECT 168.19 61.675 168.36 66.145 ;
      RECT 164.93 64.405 165.1 67.115 ;
      RECT 164.93 62.91 165.1 63.285 ;
      RECT 164.93 63.905 165.1 64.235 ;
      RECT 166.69 64.405 166.86 67.115 ;
      RECT 167.24 64.405 167.41 67.42 ;
      RECT 167.24 63.905 167.41 64.235 ;
      RECT 167.24 62.955 167.41 63.285 ;
      RECT 169.14 64.405 169.31 67.115 ;
      RECT 169.14 62.91 169.31 63.285 ;
      RECT 169.14 63.905 169.31 64.235 ;
      RECT 172.33 61.8 172.5 67.42 ;
      RECT 174.09 61.8 174.26 67.42 ;
      RECT 171.72 61.175 172.23 61.505 ;
      RECT 171.63 63.695 172.16 63.865 ;
      RECT 171.72 67.585 172.23 67.915 ;
      RECT 171.79 63.865 172.16 67.585 ;
      RECT 171.79 61.505 172.16 63.695 ;
      RECT 174.43 61.505 174.8 67.585 ;
      RECT 174.36 61.175 174.87 61.505 ;
      RECT 174.36 67.585 174.87 67.915 ;
      RECT 172.67 61.505 173.04 67.585 ;
      RECT 139.16 61.675 139.33 67.415 ;
      RECT 138.62 61.505 138.99 67.585 ;
      RECT 138.55 61.175 139.06 61.505 ;
      RECT 138.55 67.585 139.06 67.915 ;
      RECT 137.73 61.675 137.9 63.495 ;
      RECT 135.97 61.675 136.14 62.74 ;
      RECT 140.04 61.675 140.21 62.74 ;
      RECT 138.28 61.675 138.45 62.725 ;
      RECT 139.88 57.325 140.05 60.405 ;
      RECT 141.34 57.305 141.51 60.405 ;
      RECT 137.73 64.405 137.9 67.115 ;
      RECT 135.97 64.405 136.14 67.115 ;
      RECT 135.97 62.91 136.14 63.285 ;
      RECT 135.97 63.905 136.14 64.235 ;
      RECT 140.04 64.405 140.21 67.115 ;
      RECT 140.04 62.91 140.21 63.285 ;
      RECT 140.04 63.905 140.21 64.235 ;
      RECT 138.28 64.405 138.45 67.115 ;
      RECT 138.28 63.905 138.45 64.235 ;
      RECT 138.28 62.955 138.45 63.285 ;
      RECT 144.11 61.8 144.28 67.42 ;
      RECT 146.42 61.8 146.59 67.42 ;
      RECT 143.57 61.505 143.94 67.585 ;
      RECT 143.5 67.585 144.01 67.915 ;
      RECT 143.5 61.175 144.175 61.345 ;
      RECT 143.5 61.345 144.01 61.505 ;
      RECT 146.76 61.505 147.13 67.585 ;
      RECT 146.69 61.175 147.2 61.505 ;
      RECT 145.81 61.175 146.32 61.505 ;
      RECT 145.72 63.695 146.25 63.865 ;
      RECT 146.69 67.585 147.2 67.59 ;
      RECT 145.81 67.59 147.2 67.915 ;
      RECT 145.81 67.585 146.32 67.59 ;
      RECT 145.88 63.865 146.25 67.585 ;
      RECT 145.88 61.505 146.25 63.695 ;
      RECT 144.45 61.505 144.82 67.585 ;
      RECT 144.38 61.175 144.89 61.505 ;
      RECT 144.38 67.585 144.89 67.915 ;
      RECT 144.65 61.075 144.82 61.175 ;
      RECT 142.62 61.175 143.13 61.505 ;
      RECT 142.69 63.455 143.22 63.625 ;
      RECT 142.62 67.585 143.13 67.915 ;
      RECT 142.69 63.625 143.06 67.585 ;
      RECT 142.69 61.505 143.06 63.455 ;
      RECT 141.8 61.675 141.97 63.495 ;
      RECT 143.23 61.675 143.4 62.74 ;
      RECT 145.33 61.645 145.71 61.815 ;
      RECT 145.11 61.26 145.64 61.43 ;
      RECT 145.33 61.43 145.5 61.645 ;
      RECT 145.54 61.815 145.71 63.495 ;
      RECT 144.99 61.675 145.16 63.495 ;
      RECT 147.3 61.675 147.47 62.74 ;
      RECT 141.8 64.405 141.97 67.115 ;
      RECT 143.23 64.405 143.4 67.115 ;
      RECT 143.23 62.91 143.4 63.285 ;
      RECT 143.23 63.905 143.4 64.235 ;
      RECT 144.99 64.405 145.16 67.115 ;
      RECT 145.54 64.405 145.71 67.115 ;
      RECT 147.3 64.405 147.47 67.115 ;
      RECT 147.3 62.91 147.47 63.285 ;
      RECT 147.3 63.905 147.47 64.235 ;
      RECT 152.65 61.255 153.18 61.425 ;
      RECT 152.73 61.175 153.1 61.255 ;
      RECT 152.645 67.685 153.155 67.915 ;
      RECT 152.47 67.585 153.155 67.685 ;
      RECT 152.47 67.515 153.1 67.585 ;
      RECT 152.73 61.425 153.1 67.515 ;
      RECT 149.47 61.505 149.84 67.585 ;
      RECT 149.4 67.585 149.91 67.915 ;
      RECT 149.4 61.285 149.93 61.455 ;
      RECT 149.4 61.455 149.91 61.505 ;
      RECT 149.4 61.175 149.91 61.285 ;
      RECT 150.28 61.175 150.79 61.505 ;
      RECT 150.28 67.585 150.79 67.915 ;
      RECT 150.26 67.115 150.79 67.285 ;
      RECT 150.35 67.285 150.72 67.585 ;
      RECT 150.35 61.505 150.72 67.115 ;
      RECT 148.52 61.505 148.89 67.585 ;
      RECT 148.45 61.175 148.96 61.505 ;
      RECT 148.45 67.585 148.96 67.915 ;
      RECT 148.18 61.675 148.35 67.415 ;
      RECT 147.64 61.505 148.01 67.585 ;
      RECT 147.57 67.585 148.08 67.915 ;
      RECT 147.565 61.26 148.095 61.43 ;
      RECT 147.57 61.43 148.08 61.505 ;
      RECT 147.57 61.175 148.08 61.26 ;
      RECT 149.06 61.675 149.23 62.725 ;
      RECT 150.01 61.675 150.18 66.135 ;
      RECT 149.92 60.665 151.89 60.835 ;
      RECT 151.85 61.505 152.22 61.885 ;
      RECT 151.76 61.255 152.29 61.425 ;
      RECT 151.78 61.425 152.29 61.505 ;
      RECT 151.78 61.175 152.29 61.255 ;
      RECT 150.96 61.675 151.13 62.725 ;
      RECT 151.51 63.695 152.04 63.865 ;
      RECT 151.51 61.675 151.68 63.695 ;
      RECT 151.51 63.865 151.68 67.115 ;
      RECT 152.215 60.665 152.745 60.835 ;
      RECT 152.39 61.675 152.56 62.685 ;
      RECT 149.06 64.405 149.23 67.115 ;
      RECT 149.06 63.905 149.23 64.235 ;
      RECT 149.06 62.955 149.23 63.285 ;
      RECT 150.96 64.405 151.13 67.42 ;
      RECT 152.39 63.905 152.56 64.235 ;
      RECT 152.39 62.955 152.56 63.285 ;
      RECT 150.96 63.905 151.13 64.235 ;
      RECT 150.96 62.955 151.13 63.285 ;
      RECT 152.39 64.405 152.56 67.115 ;
      RECT 153.17 60.665 156.28 60.835 ;
      RECT 154.41 61.255 154.94 61.425 ;
      RECT 154.49 61.505 154.86 61.88 ;
      RECT 154.42 61.425 154.93 61.505 ;
      RECT 154.42 61.175 154.93 61.255 ;
      RECT 155.315 67.585 155.825 67.915 ;
      RECT 155.3 61.285 155.835 61.455 ;
      RECT 155.3 61.455 155.81 61.505 ;
      RECT 155.3 61.175 155.81 61.285 ;
      RECT 155.37 61.505 155.74 67.585 ;
      RECT 154.49 63.695 155.02 63.865 ;
      RECT 154.49 63.865 154.82 63.965 ;
      RECT 154.49 63.455 154.82 63.695 ;
      RECT 154.15 65.585 154.68 65.755 ;
      RECT 154.15 65.755 154.32 67.42 ;
      RECT 154.15 61.675 154.32 65.585 ;
      RECT 153.45 63.415 153.98 63.585 ;
      RECT 153.535 67.585 154.045 67.915 ;
      RECT 153.61 63.585 153.98 67.585 ;
      RECT 114.625 61.175 115.135 61.505 ;
      RECT 114.695 61.505 115.065 67.585 ;
      RECT 114.625 67.585 115.135 67.915 ;
      RECT 115.785 64.405 115.955 67.115 ;
      RECT 117.545 64.405 117.715 67.115 ;
      RECT 116.665 61.8 116.835 67.42 ;
      RECT 117.545 62.91 117.715 63.285 ;
      RECT 115.785 61.675 115.955 63.855 ;
      RECT 117.545 61.675 117.715 62.74 ;
      RECT 117.545 63.905 117.715 64.235 ;
      RECT 117.815 61.175 118.325 61.505 ;
      RECT 117.885 61.505 118.255 67.585 ;
      RECT 117.815 67.585 118.325 67.915 ;
      RECT 115.74 57.325 115.91 60.405 ;
      RECT 121.04 61.175 121.55 61.505 ;
      RECT 121.11 66.745 121.64 66.915 ;
      RECT 121.99 61.505 122.36 67.585 ;
      RECT 121.92 61.175 122.43 61.505 ;
      RECT 121.11 66.915 121.48 67.585 ;
      RECT 121.11 61.505 121.48 66.745 ;
      RECT 121.04 67.585 122.43 67.915 ;
      RECT 123.82 61.505 124.19 67.585 ;
      RECT 123.75 61.175 124.26 61.505 ;
      RECT 123.75 67.585 124.26 67.915 ;
      RECT 118.765 61.505 119.135 67.585 ;
      RECT 118.695 61.175 119.205 61.505 ;
      RECT 118.695 67.585 119.205 67.915 ;
      RECT 122.94 61.505 123.31 67.585 ;
      RECT 122.87 61.175 123.38 61.505 ;
      RECT 122.87 67.585 123.38 67.915 ;
      RECT 119.305 64.235 120.285 67.115 ;
      RECT 119.305 63.905 120.87 64.235 ;
      RECT 120.115 67.115 120.285 67.415 ;
      RECT 120.115 61.675 120.285 62.955 ;
      RECT 119.305 62.955 120.87 63.285 ;
      RECT 119.305 61.675 119.475 62.725 ;
      RECT 118.425 61.675 118.595 67.415 ;
      RECT 122.6 61.675 122.77 62.725 ;
      RECT 120.7 61.675 120.87 62.725 ;
      RECT 122.6 64.405 122.77 67.115 ;
      RECT 120.7 64.405 120.87 67.42 ;
      RECT 121.65 61.675 121.82 66.145 ;
      RECT 122.6 62.955 122.77 63.285 ;
      RECT 122.6 63.905 122.77 64.235 ;
      RECT 123.48 61.675 123.65 67.415 ;
      RECT 127.41 61.505 127.78 67.585 ;
      RECT 127.34 61.175 127.85 61.505 ;
      RECT 126.53 61.505 126.9 67.585 ;
      RECT 126.46 61.175 126.97 61.505 ;
      RECT 127.335 67.915 127.865 68.055 ;
      RECT 126.46 67.585 127.85 67.885 ;
      RECT 126.46 67.885 127.865 67.915 ;
      RECT 128.98 61.505 129.35 67.585 ;
      RECT 128.91 61.175 129.42 61.505 ;
      RECT 128.91 67.585 129.42 67.915 ;
      RECT 129.86 61.505 130.23 67.585 ;
      RECT 129.79 61.175 130.3 61.505 ;
      RECT 129.79 67.585 130.3 67.915 ;
      RECT 125.64 59.125 130.15 60.315 ;
      RECT 125.785 59.115 129.915 59.125 ;
      RECT 125.58 61.505 125.95 67.585 ;
      RECT 125.51 61.175 126.02 61.505 ;
      RECT 125.51 67.585 126.02 67.915 ;
      RECT 125.24 61.675 125.41 67.415 ;
      RECT 124.7 61.505 125.07 67.585 ;
      RECT 124.63 61.175 125.14 61.505 ;
      RECT 124.63 67.585 125.14 67.915 ;
      RECT 124.36 61.675 124.53 62.725 ;
      RECT 126.12 61.675 126.29 62.725 ;
      RECT 127.07 61.675 127.24 66.145 ;
      RECT 128.02 61.675 128.74 62.725 ;
      RECT 129.52 61.675 129.69 66.145 ;
      RECT 124.36 64.405 124.53 67.115 ;
      RECT 124.36 63.905 124.53 64.235 ;
      RECT 124.36 62.955 124.53 63.285 ;
      RECT 126.12 64.405 126.29 67.115 ;
      RECT 126.12 62.955 126.29 63.285 ;
      RECT 126.12 63.905 126.29 64.235 ;
      RECT 128.02 62.955 128.74 63.285 ;
      RECT 128.02 63.905 128.74 64.235 ;
      RECT 128.57 64.405 128.74 67.42 ;
      RECT 128.02 64.405 128.19 67.42 ;
      RECT 130.81 61.505 131.18 67.585 ;
      RECT 130.74 61.175 131.25 61.505 ;
      RECT 130.74 67.585 131.25 67.915 ;
      RECT 131.69 61.505 132.06 67.585 ;
      RECT 131.62 61.175 132.13 61.505 ;
      RECT 131.62 67.585 132.13 67.915 ;
      RECT 133.12 61.505 133.49 67.585 ;
      RECT 133.05 61.175 133.56 61.505 ;
      RECT 133.05 67.585 133.56 67.915 ;
      RECT 131.35 61.8 131.52 67.42 ;
      RECT 130.47 64.405 130.64 67.115 ;
      RECT 130.47 62.91 130.64 63.285 ;
      RECT 130.47 63.905 130.64 64.235 ;
      RECT 130.47 61.675 130.64 62.74 ;
      RECT 132.23 64.405 132.4 67.115 ;
      RECT 132.23 61.675 132.4 63.495 ;
      RECT 132.78 61.675 132.95 67.42 ;
      RECT 133.66 61.675 133.83 62.725 ;
      RECT 133.66 64.405 133.83 67.115 ;
      RECT 133.66 63.905 133.83 64.235 ;
      RECT 133.66 62.955 133.83 63.285 ;
      RECT 136.85 61.8 137.02 67.42 ;
      RECT 140.92 61.8 141.09 67.42 ;
      RECT 137.19 61.505 137.56 67.585 ;
      RECT 137.12 61.175 137.63 61.505 ;
      RECT 137.12 67.585 137.63 67.915 ;
      RECT 141.19 61.175 141.7 61.505 ;
      RECT 140.38 61.505 140.75 67.585 ;
      RECT 140.31 61.175 140.82 61.505 ;
      RECT 141.26 63.865 141.63 67.585 ;
      RECT 141.26 61.505 141.63 63.695 ;
      RECT 141.19 67.585 141.7 67.59 ;
      RECT 141.26 63.695 142.52 63.865 ;
      RECT 142.35 63.865 142.52 67.42 ;
      RECT 142.35 61.675 142.52 63.695 ;
      RECT 140.31 67.59 141.7 67.915 ;
      RECT 140.31 67.585 140.82 67.59 ;
      RECT 136.31 61.505 136.68 67.585 ;
      RECT 136.24 61.175 136.75 61.505 ;
      RECT 136.24 67.585 136.75 67.915 ;
      RECT 139.43 61.175 139.94 61.505 ;
      RECT 139.43 67.585 139.94 67.915 ;
      RECT 139.5 63.455 140.12 63.625 ;
      RECT 139.5 63.625 139.87 67.585 ;
      RECT 139.5 61.505 139.87 63.455 ;
      RECT 99.425 87.885 100.225 91.465 ;
      RECT 144.715 87.885 145.515 90.92 ;
      RECT 99.05 87.87 100.935 87.885 ;
      RECT 102.78 87.87 110.985 87.885 ;
      RECT 111.985 87.87 175.8 87.885 ;
      RECT 99.05 87.7 175.8 87.87 ;
      RECT 152.345 87.07 175.8 87.7 ;
      RECT 155.74 86.38 175.8 87.07 ;
      RECT 155.725 86.375 175.8 86.38 ;
      RECT 155.725 86.32 170.73 86.375 ;
      RECT 133.575 86.315 136.55 87.7 ;
      RECT 155.725 86.21 170.705 86.32 ;
      RECT 133.44 85.785 136.55 86.315 ;
      RECT 171.66 85.65 175.8 86.375 ;
      RECT 133.575 85.555 136.55 85.785 ;
      RECT 155.78 85.025 158.15 86.21 ;
      RECT 167.415 84.555 167.585 86.21 ;
      RECT 152.355 81.95 152.525 87.07 ;
      RECT 173.725 82.17 173.895 85.65 ;
      RECT 171.965 82.17 172.135 85.65 ;
      RECT 170.535 82.05 170.705 86.21 ;
      RECT 100.685 76.345 101.375 77.785 ;
      RECT 99.05 76.195 99.22 87.7 ;
      RECT 100.685 76.195 101.48 76.345 ;
      RECT 99.05 76.025 101.48 76.195 ;
      RECT 174.73 73.615 175.8 85.65 ;
      RECT 171.895 71.225 175.8 73.615 ;
      RECT 100.63 68.505 101.48 76.025 ;
      RECT 171.895 68.615 175.8 70.285 ;
      RECT 171.88 70.285 175.8 71.225 ;
      RECT 100.63 67.115 101.375 68.505 ;
      RECT 175.63 64.235 175.8 68.615 ;
      RECT 101.205 63.905 102.07 63.975 ;
      RECT 100.63 63.975 102.07 67.115 ;
      RECT 175.27 64.065 175.8 64.235 ;
      RECT 175.63 63.905 175.8 64.065 ;
      RECT 105.43 61.175 105.94 61.505 ;
      RECT 105.43 67.585 105.94 67.915 ;
      RECT 105.5 66.375 106.03 66.545 ;
      RECT 105.5 66.545 105.87 67.585 ;
      RECT 105.5 61.505 105.87 66.375 ;
      RECT 106.38 61.505 106.75 67.585 ;
      RECT 106.31 61.175 106.82 61.505 ;
      RECT 106.31 67.585 106.82 67.915 ;
      RECT 102.24 61.505 102.61 67.585 ;
      RECT 102.17 61.175 102.68 61.505 ;
      RECT 102.17 67.585 102.68 67.915 ;
      RECT 102.78 61.675 102.95 67.415 ;
      RECT 103.12 61.505 103.49 67.585 ;
      RECT 103.05 61.175 103.56 61.505 ;
      RECT 103.05 67.585 103.56 67.915 ;
      RECT 104.54 61.675 104.71 67.42 ;
      RECT 104 61.505 104.37 67.585 ;
      RECT 103.93 61.175 104.44 61.505 ;
      RECT 103.93 67.585 104.44 67.915 ;
      RECT 101.205 61.675 101.375 62.955 ;
      RECT 101.205 62.955 102.07 63.285 ;
      RECT 103.66 61.675 103.83 62.725 ;
      RECT 101.9 61.675 102.07 62.725 ;
      RECT 105.09 61.675 105.26 62.725 ;
      RECT 106.04 61.675 106.21 66.145 ;
      RECT 103.66 64.405 103.83 67.115 ;
      RECT 103.66 63.905 103.83 64.235 ;
      RECT 103.66 62.955 103.83 63.285 ;
      RECT 105.09 64.405 105.26 67.42 ;
      RECT 105.09 63.905 105.26 64.235 ;
      RECT 105.09 62.955 105.26 63.285 ;
      RECT 108.28 61.505 108.65 67.585 ;
      RECT 108.21 61.175 108.72 61.505 ;
      RECT 108.21 67.585 108.72 67.915 ;
      RECT 107.4 61.505 107.77 67.585 ;
      RECT 107.33 67.585 107.84 67.915 ;
      RECT 107.33 61.175 107.86 61.345 ;
      RECT 107.33 61.345 107.84 61.505 ;
      RECT 110.66 61.505 111.03 67.585 ;
      RECT 110.59 61.175 111.1 61.505 ;
      RECT 110.59 67.585 111.1 67.915 ;
      RECT 110.32 61.675 110.49 67.415 ;
      RECT 109.71 61.175 110.22 61.505 ;
      RECT 109.78 61.505 110.15 67.515 ;
      RECT 109.62 67.515 110.15 67.585 ;
      RECT 109.71 67.685 110.22 67.915 ;
      RECT 109.62 67.585 110.22 67.685 ;
      RECT 108.89 61.675 109.61 62.725 ;
      RECT 106.99 61.675 107.16 62.725 ;
      RECT 107.94 61.675 108.11 66.145 ;
      RECT 111.2 61.675 111.37 62.725 ;
      RECT 112.595 61.675 112.765 63.495 ;
      RECT 112.01 61.675 112.18 62.955 ;
      RECT 111.2 62.955 112.18 63.285 ;
      RECT 108.89 63.905 109.61 64.235 ;
      RECT 109.44 64.235 109.61 67.115 ;
      RECT 108.89 62.955 109.61 63.285 ;
      RECT 108.89 64.405 109.06 67.42 ;
      RECT 106.99 64.405 107.16 67.115 ;
      RECT 106.99 62.955 107.16 63.285 ;
      RECT 106.99 63.905 107.16 64.235 ;
      RECT 112.01 67.115 112.18 67.415 ;
      RECT 111.2 63.905 112.18 67.115 ;
      RECT 112.595 64.405 112.765 67.115 ;
      RECT 114.28 57.305 114.45 60.405 ;
      RECT 116.055 61.175 116.565 61.505 ;
      RECT 116.055 67.59 117.445 67.92 ;
      RECT 117.005 61.505 117.375 67.585 ;
      RECT 116.935 61.175 117.445 61.505 ;
      RECT 115.235 64.235 115.405 67.42 ;
      RECT 115.235 61.675 115.405 64.025 ;
      RECT 115.235 64.025 116.495 64.235 ;
      RECT 116.125 64.235 116.495 67.585 ;
      RECT 116.125 61.505 116.495 64.025 ;
      RECT 116.055 67.585 116.565 67.59 ;
      RECT 116.935 67.585 117.445 67.59 ;
      RECT 114.355 64.405 114.525 67.115 ;
      RECT 113.475 61.8 113.645 67.42 ;
      RECT 114.355 62.91 114.525 63.285 ;
      RECT 113.745 67.585 114.255 67.915 ;
      RECT 113.815 61.605 114.185 67.585 ;
      RECT 113.655 61.505 114.185 61.605 ;
      RECT 113.745 61.175 114.255 61.435 ;
      RECT 113.655 61.435 114.255 61.505 ;
      RECT 112.935 61.505 113.305 67.585 ;
      RECT 112.865 67.585 113.375 67.915 ;
      RECT 112.91 61.065 113.44 61.175 ;
      RECT 112.865 61.235 113.375 61.505 ;
      RECT 112.865 61.175 113.44 61.235 ;
      RECT 114.355 61.675 114.525 62.74 ;
      RECT 114.355 63.905 114.525 64.235 ;
      RECT 453.17 56.125 453.34 60.875 ;
      RECT 453.755 60.525 454.315 60.845 ;
      RECT 453.95 60.845 454.12 60.875 ;
      RECT 453.95 56.125 454.12 60.525 ;
      RECT 453.22 55.605 456.36 55.775 ;
      RECT 453.22 53.485 456.36 53.655 ;
      RECT 459.645 61.915 460.175 62.085 ;
      RECT 458.635 54.895 460.175 55.225 ;
      RECT 459.805 62.085 460.175 62.09 ;
      RECT 459.805 55.225 460.175 61.915 ;
      RECT 457.755 54.895 458.265 55.225 ;
      RECT 457.825 55.225 458.195 56.8 ;
      RECT 457.825 56.8 458.355 56.97 ;
      RECT 457.755 50.09 458.265 50.42 ;
      RECT 457.825 50.42 458.195 51.895 ;
      RECT 457.825 51.895 458.355 52.065 ;
      RECT 457.755 54.035 458.265 54.365 ;
      RECT 457.825 52.46 458.195 54.035 ;
      RECT 457.825 52.29 458.355 52.46 ;
      RECT 459.245 55.395 459.415 56.8 ;
      RECT 458.885 56.8 459.415 56.97 ;
      RECT 458.365 55.395 458.535 56.445 ;
      RECT 457.03 61.385 457.655 61.555 ;
      RECT 457.03 61.555 457.2 61.585 ;
      RECT 457.03 56.405 457.2 61.385 ;
      RECT 457.03 55.395 457.655 56.405 ;
      RECT 457.485 50.59 457.655 51.64 ;
      RECT 458.365 50.59 458.535 51.6 ;
      RECT 459.245 52.46 459.415 53.865 ;
      RECT 458.885 52.29 459.415 52.46 ;
      RECT 458.365 52.815 458.535 53.865 ;
      RECT 459.245 50.59 459.415 51.895 ;
      RECT 458.885 51.895 459.415 52.065 ;
      RECT 455.145 60.525 455.705 60.845 ;
      RECT 455.35 60.845 455.52 60.875 ;
      RECT 455.35 56.125 455.52 60.525 ;
      RECT 455.94 59.945 456.475 60.265 ;
      RECT 456.13 60.265 456.3 60.875 ;
      RECT 456.13 56.125 456.3 59.945 ;
      RECT 454.415 59.365 454.98 59.685 ;
      RECT 454.57 59.685 454.74 60.875 ;
      RECT 454.57 56.125 454.74 59.365 ;
      RECT 461.615 56.8 462.145 56.97 ;
      RECT 461.545 61.305 462.055 61.635 ;
      RECT 461.615 56.97 461.985 61.305 ;
      RECT 463.035 56.8 463.565 56.97 ;
      RECT 463.035 56.97 463.205 61.14 ;
      RECT 469.485 59.945 470.045 60.265 ;
      RECT 469.65 60.265 469.82 60.875 ;
      RECT 469.65 56.125 469.82 59.945 ;
      RECT 471.21 56.125 471.38 60.875 ;
      RECT 467.245 56.785 469.1 57.035 ;
      RECT 468.85 55.775 469.1 56.785 ;
      RECT 468.165 57.035 468.615 61.025 ;
      RECT 468.85 55.525 471.42 55.775 ;
      RECT 470.2 60.525 470.76 60.845 ;
      RECT 470.43 60.845 470.6 60.875 ;
      RECT 470.43 56.125 470.6 60.525 ;
      RECT 18.875 63.27 19.545 63.44 ;
      RECT 18.465 64.05 18.635 68.9 ;
      RECT 18.465 57.685 18.635 62.535 ;
      RECT 19.745 64.05 19.915 68.9 ;
      RECT 19.745 57.685 19.915 62.535 ;
      RECT 22.715 63.27 23.385 63.44 ;
      RECT 20.155 63.27 22.105 63.44 ;
      RECT 21.415 57.265 22.085 57.435 ;
      RECT 20.135 57.265 20.805 57.435 ;
      RECT 23.585 64.05 23.755 68.9 ;
      RECT 23.585 57.685 23.755 62.535 ;
      RECT 21.025 64.05 21.195 68.9 ;
      RECT 22.305 64.05 22.475 68.9 ;
      RECT 21.025 57.685 21.195 62.535 ;
      RECT 22.305 57.685 22.475 62.535 ;
      RECT 30.185 57.4 30.855 57.57 ;
      RECT 30.255 57.39 30.785 57.4 ;
      RECT 28.905 57.4 29.575 57.57 ;
      RECT 28.975 57.39 29.505 57.4 ;
      RECT 28.515 57.98 28.685 62.83 ;
      RECT 31.075 57.98 31.245 62.83 ;
      RECT 29.795 58.08 29.965 62.83 ;
      RECT 45.37 65.035 46.08 65.285 ;
      RECT 45.83 65.285 46 65.325 ;
      RECT 45.83 64.995 46 65.035 ;
      RECT 71.635 58.375 72.305 58.545 ;
      RECT 70.455 58.375 71.125 58.545 ;
      RECT 67.99 61.25 68.66 61.42 ;
      RECT 68.06 61.235 68.59 61.25 ;
      RECT 66.71 61.25 67.38 61.42 ;
      RECT 66.78 61.235 67.31 61.25 ;
      RECT 66.32 61.64 66.49 64.35 ;
      RECT 68.88 61.64 69.05 64.35 ;
      RECT 66.485 57.285 66.655 59.995 ;
      RECT 69.045 57.285 69.215 59.995 ;
      RECT 67.765 57.285 67.935 59.995 ;
      RECT 67.6 61.64 67.77 64.35 ;
      RECT 72.815 58.375 73.485 58.545 ;
      RECT 73.995 58.375 74.665 58.545 ;
      RECT 78.385 59.195 78.555 61.905 ;
      RECT 81.905 59.195 82.075 61.905 ;
      RECT 83.025 59.195 83.195 61.905 ;
      RECT 80.145 59.195 80.315 61.905 ;
      RECT 81.905 58.695 82.075 59.025 ;
      RECT 80.145 58.695 80.315 59.025 ;
      RECT 78.385 58.695 78.555 59.025 ;
      RECT 80.145 57.745 80.315 58.075 ;
      RECT 81.905 57.745 82.075 58.075 ;
      RECT 78.385 57.745 78.555 58.075 ;
      RECT 83.025 58.695 83.195 59.025 ;
      RECT 83.025 57.745 83.195 58.075 ;
      RECT 80.33 64.605 80.84 67.865 ;
      RECT 80.33 64.435 81.895 64.605 ;
      RECT 84.785 59.195 84.955 61.905 ;
      RECT 86.255 59.195 86.425 61.905 ;
      RECT 89.1 57.44 89.27 62.29 ;
      RECT 84.785 58.695 84.955 59.025 ;
      RECT 84.785 57.745 84.955 58.075 ;
      RECT 86.255 58.695 86.425 59.025 ;
      RECT 86.255 57.745 86.425 58.075 ;
      RECT 90.47 57.44 90.64 62.29 ;
      RECT 93.03 57.44 93.2 62.29 ;
      RECT 89.88 57.44 90.05 62.29 ;
      RECT 91.75 57.44 91.92 62.29 ;
      RECT 92.415 64.435 93.98 64.605 ;
      RECT 93.47 64.605 93.98 67.865 ;
      RECT 99.425 91.72 125.53 92.265 ;
      RECT 99.425 91.465 145.515 91.72 ;
      RECT 124.73 90.92 145.515 91.465 ;
      RECT 310.91 56.295 311.28 62.375 ;
      RECT 311.45 56.465 311.62 57.515 ;
      RECT 312.5 51 317.25 51.17 ;
      RECT 312.845 51.81 313.375 51.98 ;
      RECT 313.015 51.98 313.185 54.43 ;
      RECT 313.015 51.72 313.185 51.81 ;
      RECT 314.6 51.81 315.13 51.98 ;
      RECT 314.775 51.98 314.945 54.43 ;
      RECT 314.775 51.72 314.945 51.81 ;
      RECT 311.085 53.37 311.615 53.54 ;
      RECT 311.255 53.54 311.425 54.43 ;
      RECT 311.255 51.72 311.425 53.37 ;
      RECT 309.69 56.465 309.86 57.515 ;
      RECT 310.57 56.465 310.74 62.21 ;
      RECT 318.76 50.25 321.45 50.265 ;
      RECT 318.7 50.08 321.41 50.095 ;
      RECT 318.7 50.095 321.45 50.25 ;
      RECT 319.455 50.265 320.805 51.17 ;
      RECT 317.695 50.66 319.045 51.17 ;
      RECT 317.695 50.265 318.4 50.66 ;
      RECT 311.355 50.25 318.4 50.265 ;
      RECT 311.2 50.095 318.365 50.25 ;
      RECT 311.2 50.08 318.33 50.095 ;
      RECT 316.365 51.81 316.895 51.98 ;
      RECT 316.535 51.98 316.705 54.43 ;
      RECT 316.535 51.72 316.705 51.81 ;
      RECT 318.125 52.18 318.655 52.35 ;
      RECT 318.295 52.35 318.465 54.43 ;
      RECT 318.295 51.72 318.465 52.18 ;
      RECT 319.885 52.18 320.415 52.35 ;
      RECT 320.055 52.35 320.225 54.43 ;
      RECT 320.055 51.72 320.225 52.18 ;
      RECT 321.88 50.08 324.59 50.25 ;
      RECT 321.88 50.25 322.73 51 ;
      RECT 321.215 51 322.73 51.17 ;
      RECT 322.43 56.5 323.1 56.67 ;
      RECT 321.15 56.5 321.82 56.67 ;
      RECT 321.645 52.18 322.175 52.35 ;
      RECT 321.815 52.35 321.985 54.43 ;
      RECT 321.815 51.72 321.985 52.18 ;
      RECT 327.365 50.955 344.7 53.665 ;
      RECT 327.365 55.34 353.22 58.05 ;
      RECT 348.79 49.475 353.54 49.645 ;
      RECT 348.79 49.465 353.495 49.475 ;
      RECT 360.665 52.4 360.995 52.845 ;
      RECT 360.665 52.195 360.995 52.23 ;
      RECT 360.385 52.23 360.995 52.4 ;
      RECT 361.445 52.195 361.775 52.845 ;
      RECT 361.155 51.925 361.325 52.025 ;
      RECT 361.135 50.575 361.305 51.135 ;
      RECT 361.135 51.135 361.325 51.925 ;
      RECT 360.355 50.575 360.525 51.925 ;
      RECT 361.575 50.005 363.42 50.175 ;
      RECT 361.635 50 363.34 50.005 ;
      RECT 358.28 56.945 362.11 57.175 ;
      RECT 361.88 57.175 362.11 63.485 ;
      RECT 358.25 57.92 358.48 63.485 ;
      RECT 358.25 63.685 359.44 63.715 ;
      RECT 358.25 63.485 359.44 63.515 ;
      RECT 358.25 63.515 362.11 63.685 ;
      RECT 361.29 63.685 362.11 63.715 ;
      RECT 361.29 63.485 362.11 63.515 ;
      RECT 358.28 57.175 358.45 57.92 ;
      RECT 357.34 56.03 363.035 56.2 ;
      RECT 362.865 56.2 363.035 64.455 ;
      RECT 357.34 64.455 363.035 64.625 ;
      RECT 357.34 56.2 357.51 64.455 ;
      RECT 364.255 50.575 364.425 51.925 ;
      RECT 363.785 52.335 364.115 52.845 ;
      RECT 363.815 50.175 364.08 52.335 ;
      RECT 363.7 50.005 364.37 50.175 ;
      RECT 363.005 52.195 363.335 52.845 ;
      RECT 362.225 52.4 362.555 52.845 ;
      RECT 362.225 52.195 362.555 52.23 ;
      RECT 361.945 52.23 362.555 52.4 ;
      RECT 361.915 50.575 362.085 51.925 ;
      RECT 362.715 51.925 362.885 52.025 ;
      RECT 362.695 50.575 362.865 51.14 ;
      RECT 362.695 51.14 362.885 51.925 ;
      RECT 363.475 50.575 363.645 51.925 ;
      RECT 366.63 52.675 367.415 52.845 ;
      RECT 373.525 56.71 373.855 58.3 ;
      RECT 374.335 56.71 374.865 58.05 ;
      RECT 374.215 54.165 374.865 56.71 ;
      RECT 430.48 56.485 430.81 57.175 ;
      RECT 430.48 49.85 431.58 50.02 ;
      RECT 429.71 56.485 430.04 57.175 ;
      RECT 429.595 49.85 430.125 50.02 ;
      RECT 436.31 56.485 436.64 57.175 ;
      RECT 436.31 49.785 437.41 50.295 ;
      RECT 434.33 49.785 435.43 50.295 ;
      RECT 434.33 56.485 434.66 57.175 ;
      RECT 431.25 56.485 431.58 57.175 ;
      RECT 431.915 49.85 432.445 50.02 ;
      RECT 432.02 56.485 432.35 57.175 ;
      RECT 432.79 56.485 433.12 57.175 ;
      RECT 432.79 49.79 433.89 50.3 ;
      RECT 433.56 56.485 433.89 57.175 ;
      RECT 435.1 56.485 435.43 57.175 ;
      RECT 437.08 56.485 437.41 57.175 ;
      RECT 440.16 56.485 440.49 57.175 ;
      RECT 440.16 49.85 441.26 50.02 ;
      RECT 439.295 49.85 439.825 50.02 ;
      RECT 439.39 56.485 439.72 57.175 ;
      RECT 440.93 56.485 441.26 57.175 ;
      RECT 441.7 56.485 442.03 57.175 ;
      RECT 441.615 49.85 442.145 50.02 ;
      RECT 438.62 56.485 438.95 57.175 ;
      RECT 437.85 49.79 438.95 50.3 ;
      RECT 437.85 56.485 438.18 57.175 ;
      RECT 444.12 53.96 446.83 54.13 ;
      RECT 445.2 54.13 446.81 54.23 ;
      RECT 447.01 54.185 447.18 59.445 ;
      RECT 443.225 53.585 443.485 56.94 ;
      RECT 443.225 58.505 443.485 59.97 ;
      RECT 447.425 53.54 447.595 60.015 ;
      RECT 443.225 53.37 447.595 53.54 ;
      RECT 443.225 53.54 444.35 53.585 ;
      RECT 443.225 53.325 444.35 53.37 ;
      RECT 443.225 60.185 444.35 60.23 ;
      RECT 443.225 60.015 447.595 60.185 ;
      RECT 443.225 59.97 444.35 60.015 ;
      RECT 443.27 56.94 443.44 58.505 ;
      RECT 444.12 57.08 446.83 57.25 ;
      RECT 444.03 56.3 446.83 56.47 ;
      RECT 444.12 55.52 446.83 55.69 ;
      RECT 444.03 54.74 446.83 54.91 ;
      RECT 271.35 49.955 271.52 50.845 ;
      RECT 272.015 54.705 272.185 55.895 ;
      RECT 269.025 55.085 271.555 55.285 ;
      RECT 270.57 49.955 270.74 55.085 ;
      RECT 269.025 55.285 269.195 60.365 ;
      RECT 271.385 55.285 271.555 60.365 ;
      RECT 273.415 53.37 273.945 53.54 ;
      RECT 273.775 56.265 274.305 56.435 ;
      RECT 273.775 50.845 273.945 53.37 ;
      RECT 273.775 53.54 273.945 56.265 ;
      RECT 272.895 50.845 273.065 55.525 ;
      RECT 272.165 58.725 273.055 59.255 ;
      RECT 272.165 59.255 273.015 60.485 ;
      RECT 272.165 56.755 273.015 58.725 ;
      RECT 272.31 56.265 272.84 56.435 ;
      RECT 272.51 55.785 272.84 56.265 ;
      RECT 270.205 55.455 270.375 60.365 ;
      RECT 273.245 53.995 273.575 54.325 ;
      RECT 273.055 55.895 273.585 56.065 ;
      RECT 273.255 56.065 273.585 56.295 ;
      RECT 273.255 55.785 273.585 55.895 ;
      RECT 274.47 52.23 275 52.4 ;
      RECT 274.47 52.4 274.8 52.605 ;
      RECT 274.47 52.095 274.8 52.23 ;
      RECT 274.775 57.005 275.44 57.175 ;
      RECT 274.91 55.525 275.44 57.005 ;
      RECT 274.775 57.175 274.945 60.015 ;
      RECT 275.08 49.415 275.75 50.365 ;
      RECT 275.645 52.355 276.155 52.685 ;
      RECT 274.855 50.535 275.945 50.705 ;
      RECT 275.775 52.685 275.945 52.84 ;
      RECT 275.775 50.705 275.945 52.355 ;
      RECT 274.855 50.705 275.025 51.885 ;
      RECT 274.855 52.875 275.025 53.885 ;
      RECT 275.355 54.905 275.885 55.075 ;
      RECT 275.61 56.87 276.505 57.04 ;
      RECT 275.61 55.565 275.78 56.87 ;
      RECT 275.61 55.075 275.885 55.565 ;
      RECT 275.61 54.555 275.885 54.905 ;
      RECT 276.335 57.04 276.505 60.015 ;
      RECT 277.115 55.495 277.645 55.665 ;
      RECT 277.475 54.555 277.645 55.495 ;
      RECT 275.95 56.515 277.155 56.7 ;
      RECT 275.95 55.735 276.46 56.265 ;
      RECT 275.95 56.265 276.48 56.515 ;
      RECT 276.985 56.7 277.155 57.68 ;
      RECT 276.985 58.805 277.595 60.665 ;
      RECT 276.925 56.065 277.595 56.345 ;
      RECT 276.88 55.895 277.595 56.065 ;
      RECT 276.925 55.835 277.595 55.895 ;
      RECT 277.325 56.345 277.595 58.805 ;
      RECT 274.83 60.665 277.595 60.835 ;
      RECT 277.765 56.67 277.935 60.405 ;
      RECT 278.345 56.69 278.515 60.405 ;
      RECT 303.92 56.295 304.29 62.375 ;
      RECT 303.85 62.375 304.36 62.705 ;
      RECT 296.815 55.765 296.985 55.965 ;
      RECT 296.815 55.965 304.36 56.295 ;
      RECT 297.195 56.635 299.145 56.805 ;
      RECT 296.09 56.625 296.26 63.475 ;
      RECT 296.09 63.475 300.945 63.645 ;
      RECT 298.175 50.405 298.705 50.575 ;
      RECT 298.205 50.575 298.375 50.75 ;
      RECT 298.205 50.08 298.375 50.405 ;
      RECT 299.025 50.96 302.075 51.13 ;
      RECT 299.055 50.08 299.225 50.96 ;
      RECT 303.11 50.865 304.46 51.17 ;
      RECT 302.785 53.37 303.315 53.54 ;
      RECT 302.785 53.54 302.955 54.43 ;
      RECT 302.785 51.72 302.955 53.37 ;
      RECT 303.58 56.465 303.75 57.515 ;
      RECT 300.48 50 300.65 50.67 ;
      RECT 300.085 56.635 300.755 56.805 ;
      RECT 299.595 53 300.125 53.17 ;
      RECT 299.595 53.17 299.765 54.43 ;
      RECT 299.595 51.72 299.765 53 ;
      RECT 303.48 53 304.01 53.17 ;
      RECT 303.665 53.17 303.835 54.43 ;
      RECT 303.665 51.72 303.835 53 ;
      RECT 300.995 53 301.525 53.17 ;
      RECT 301.355 53.17 301.525 54.43 ;
      RECT 301.355 51.72 301.525 53 ;
      RECT 304.845 51 306.195 51.41 ;
      RECT 304.375 53.37 304.905 53.54 ;
      RECT 304.545 53.54 304.715 54.43 ;
      RECT 304.545 51.72 304.715 53.37 ;
      RECT 305.265 51.64 305.795 51.81 ;
      RECT 305.425 51.81 305.595 54.43 ;
      RECT 305.945 53.37 306.475 53.54 ;
      RECT 306.305 53.54 306.475 54.43 ;
      RECT 306.305 51.72 306.475 53.37 ;
      RECT 307.25 51.31 51.17 ;
      RECT 306.62 50.08 310.73 50.095 ;
      RECT 309.2 50.265 310.73 51 ;
      RECT 306.54 50.095 310.73 50.265 ;
      RECT 307.565 53.37 308.095 53.54 ;
      RECT 307.735 53.54 307.905 54.43 ;
      RECT 307.735 51.72 307.905 53.37 ;
      RECT 309.32 53.37 309.85 53.54 ;
      RECT 309.495 53.54 309.665 54.43 ;
      RECT 309.495 51.72 309.665 53.37 ;
      RECT 306.2 55.965 306.71 56.295 ;
      RECT 306.27 56.295 306.64 62.375 ;
      RECT 306.2 62.375 306.71 62.705 ;
      RECT 305.32 55.965 305.83 56.295 ;
      RECT 305.32 62.375 305.83 62.705 ;
      RECT 305.39 58.495 305.76 62.375 ;
      RECT 305.39 56.295 305.76 58.25 ;
      RECT 304.46 58.25 305.76 58.495 ;
      RECT 304.46 58.495 304.63 62.21 ;
      RECT 304.46 56.465 304.63 58.25 ;
      RECT 305.05 56.465 305.22 57.515 ;
      RECT 305.93 56.465 306.1 62.205 ;
      RECT 309.08 55.965 310.47 56.295 ;
      RECT 309.08 62.375 310.47 62.705 ;
      RECT 309.15 56.295 309.52 62.375 ;
      RECT 310.03 56.295 310.4 62.375 ;
      RECT 308.2 55.965 308.71 56.295 ;
      RECT 308.2 62.375 308.71 62.705 ;
      RECT 307.635 58.31 308.64 58.48 ;
      RECT 308.27 56.295 308.64 58.31 ;
      RECT 308.27 58.48 308.64 62.375 ;
      RECT 307.93 56.465 308.1 57.515 ;
      RECT 306.81 56.465 306.98 57.515 ;
      RECT 308.81 56.465 308.98 62.21 ;
      RECT 310.84 55.965 311.35 56.295 ;
      RECT 310.84 62.375 311.35 62.705 ;
      RECT 249.92 51.91 250.105 52.775 ;
      RECT 249.655 52.775 250.105 53.77 ;
      RECT 248.735 52.875 248.945 53.935 ;
      RECT 247.635 50.865 247.805 53.77 ;
      RECT 248.065 52.355 248.575 52.685 ;
      RECT 248.275 50.535 249.365 50.705 ;
      RECT 248.275 52.685 248.445 52.84 ;
      RECT 248.275 50.705 248.445 52.355 ;
      RECT 249.195 50.705 249.365 51.885 ;
      RECT 249.22 52.23 249.75 52.4 ;
      RECT 249.42 52.4 249.75 52.605 ;
      RECT 249.42 52.095 249.75 52.23 ;
      RECT 250.275 53.37 250.805 53.54 ;
      RECT 249.915 56.265 250.445 56.435 ;
      RECT 250.275 50.845 250.445 53.37 ;
      RECT 250.275 53.54 250.445 56.265 ;
      RECT 251.155 50.845 251.325 55.525 ;
      RECT 247.065 56.515 248.27 56.7 ;
      RECT 247.76 55.735 248.27 56.265 ;
      RECT 247.74 56.265 248.27 56.515 ;
      RECT 247.065 56.7 247.235 57.68 ;
      RECT 246.625 58.805 247.235 60.665 ;
      RECT 246.625 55.895 247.34 56.065 ;
      RECT 246.625 56.065 247.295 56.345 ;
      RECT 246.625 55.835 247.295 55.895 ;
      RECT 246.625 60.665 249.39 60.835 ;
      RECT 246.625 56.345 246.895 58.805 ;
      RECT 248.335 54.92 248.865 55.09 ;
      RECT 247.715 56.87 248.61 57.04 ;
      RECT 248.44 55.565 248.61 56.87 ;
      RECT 248.335 55.09 248.61 55.565 ;
      RECT 248.335 54.555 248.61 54.92 ;
      RECT 247.715 57.04 247.885 60.015 ;
      RECT 248.81 57.175 249.445 57.205 ;
      RECT 248.78 55.525 249.31 57.005 ;
      RECT 248.78 57.005 249.445 57.175 ;
      RECT 249.275 57.205 249.445 60.015 ;
      RECT 246.575 55.495 247.105 55.665 ;
      RECT 246.575 54.555 246.745 55.495 ;
      RECT 250.63 53.995 250.96 54.325 ;
      RECT 250.635 55.895 251.165 56.065 ;
      RECT 250.635 56.065 250.965 56.295 ;
      RECT 250.635 55.785 250.965 55.895 ;
      RECT 251.38 56.265 251.91 56.435 ;
      RECT 251.38 55.785 251.71 56.265 ;
      RECT 249.195 52.875 249.365 53.885 ;
      RECT 246.285 56.67 246.455 60.405 ;
      RECT 251.165 58.725 252.055 59.255 ;
      RECT 251.205 59.255 252.055 60.485 ;
      RECT 251.205 56.755 252.055 58.725 ;
      RECT 252.035 50.845 252.87 54.705 ;
      RECT 251.885 55.895 252.415 56.065 ;
      RECT 252.7 49.955 252.87 50.845 ;
      RECT 252.035 54.705 252.205 55.895 ;
      RECT 252.665 55.085 255.195 55.285 ;
      RECT 253.48 49.955 253.65 55.085 ;
      RECT 252.665 55.285 252.835 60.365 ;
      RECT 255.025 55.285 255.195 60.365 ;
      RECT 255.025 49.955 255.815 54.705 ;
      RECT 255.645 54.705 255.815 60.365 ;
      RECT 253.965 53.37 254.495 53.54 ;
      RECT 254.245 53.54 254.415 54.705 ;
      RECT 254.245 49.955 254.415 53.37 ;
      RECT 252.93 60.535 256.66 60.855 ;
      RECT 255.985 49.595 256.655 60.535 ;
      RECT 256.825 49.985 256.995 60.365 ;
      RECT 253.845 55.455 254.015 60.365 ;
      RECT 261.38 50.345 262.84 50.995 ;
      RECT 258.885 60.365 259.055 60.445 ;
      RECT 265.165 60.365 265.335 60.445 ;
      RECT 258.305 50.345 260.87 50.995 ;
      RECT 258.885 49.805 265.335 49.985 ;
      RECT 263.35 50.345 265.915 50.995 ;
      RECT 265.165 50.995 265.915 60.365 ;
      RECT 258.305 49.985 265.915 50.345 ;
      RECT 258.305 50.995 259.055 60.365 ;
      RECT 260.2 51.235 260.87 51.405 ;
      RECT 260.2 58.715 261.55 58.885 ;
      RECT 261.095 52.21 261.365 58.715 ;
      RECT 260.315 51.405 260.585 58.715 ;
      RECT 257.175 49.985 257.615 60.365 ;
      RECT 257.875 49.985 258.045 54.895 ;
      RECT 259.32 51.235 259.99 51.785 ;
      RECT 259.975 51.955 260.145 58.495 ;
      RECT 259.275 52.63 259.805 52.8 ;
      RECT 259.295 54.985 259.805 55.315 ;
      RECT 259.295 51.955 259.685 52.63 ;
      RECT 259.295 52.8 259.685 54.985 ;
      RECT 260.755 51.765 261.21 51.935 ;
      RECT 261.04 50.515 261.21 51.765 ;
      RECT 260.755 51.935 260.925 58.495 ;
      RECT 262.515 51.955 262.685 58.495 ;
      RECT 261.535 51.955 261.705 58.495 ;
      RECT 262.67 58.715 264.02 58.885 ;
      RECT 263.35 51.235 264.02 51.405 ;
      RECT 262.855 52.21 263.125 58.715 ;
      RECT 263.635 51.405 263.905 58.715 ;
      RECT 263.01 51.765 263.465 51.935 ;
      RECT 263.01 50.515 263.18 51.765 ;
      RECT 263.295 51.935 263.465 58.495 ;
      RECT 262.025 51.665 262.195 58.425 ;
      RECT 257.875 55.455 258.045 60.365 ;
      RECT 257.625 60.615 259.685 60.785 ;
      RECT 259.515 55.785 259.685 60.615 ;
      RECT 257.625 60.555 258.295 60.615 ;
      RECT 264.23 51.235 264.9 51.785 ;
      RECT 264.075 51.955 264.245 58.495 ;
      RECT 264.415 52.63 264.945 52.8 ;
      RECT 264.415 54.985 264.925 55.315 ;
      RECT 264.535 51.955 264.925 52.63 ;
      RECT 264.535 52.8 264.925 54.985 ;
      RECT 266.175 49.985 266.345 54.895 ;
      RECT 266.605 49.985 267.045 60.365 ;
      RECT 267.56 60.535 271.29 60.855 ;
      RECT 267.565 49.595 268.235 60.535 ;
      RECT 267.225 49.985 267.395 60.365 ;
      RECT 268.405 49.955 269.195 54.705 ;
      RECT 268.405 54.705 268.575 60.365 ;
      RECT 264.535 60.615 266.595 60.785 ;
      RECT 264.535 55.785 264.705 60.615 ;
      RECT 265.925 60.555 266.595 60.615 ;
      RECT 266.175 55.455 266.345 60.365 ;
      RECT 269.725 53.37 270.255 53.54 ;
      RECT 269.805 53.54 269.975 54.705 ;
      RECT 269.805 49.955 269.975 53.37 ;
      RECT 271.35 50.845 272.185 54.705 ;
      RECT 271.805 55.895 272.335 56.065 ;
      RECT 223.65 53.37 224.18 53.43 ;
      RECT 222.89 56.055 223.51 56.385 ;
      RECT 223.185 56.64 224.105 56.81 ;
      RECT 223.185 56.385 223.51 56.64 ;
      RECT 223.935 56.81 224.105 57.975 ;
      RECT 226.09 56.055 226.71 56.385 ;
      RECT 225.495 56.64 226.415 56.81 ;
      RECT 226.09 56.385 226.415 56.64 ;
      RECT 225.495 56.81 225.665 57.975 ;
      RECT 223.545 53.77 223.715 55.565 ;
      RECT 225.885 53.77 226.055 55.565 ;
      RECT 225.165 56 225.835 56.17 ;
      RECT 225.235 55.87 225.765 56 ;
      RECT 223.765 56 224.435 56.17 ;
      RECT 223.835 55.87 224.365 56 ;
      RECT 224.065 55.495 224.595 55.665 ;
      RECT 224.425 54.555 224.595 55.495 ;
      RECT 225.005 55.495 225.535 55.665 ;
      RECT 225.005 54.555 225.175 55.495 ;
      RECT 228.21 55.53 229.56 55.7 ;
      RECT 228.31 55.5 229.56 55.53 ;
      RECT 227.825 53.82 229.385 53.99 ;
      RECT 227.825 52.24 230.355 52.41 ;
      RECT 227.825 52.41 227.995 53.82 ;
      RECT 228.355 53.99 228.525 55.33 ;
      RECT 229.215 53.99 229.385 55.33 ;
      RECT 230.185 52.41 230.355 53.59 ;
      RECT 230.185 51.09 230.355 52.24 ;
      RECT 227.925 54.16 228.095 55.33 ;
      RECT 227.7 55.87 228.23 56.04 ;
      RECT 227.265 56.735 228.23 56.905 ;
      RECT 227.08 56.915 227.75 57.085 ;
      RECT 225.495 59.555 225.875 60.575 ;
      RECT 227.92 56.04 228.23 56.735 ;
      RECT 227.265 56.905 227.75 56.915 ;
      RECT 227.265 57.085 227.635 60.575 ;
      RECT 225.495 60.575 227.635 60.665 ;
      RECT 225.495 60.665 227.75 60.835 ;
      RECT 227.92 57.075 228.09 57.305 ;
      RECT 227.805 57.305 228.09 60.015 ;
      RECT 231.705 54.905 232.235 55.075 ;
      RECT 232.065 49.78 232.235 54.905 ;
      RECT 229.005 49.45 231.895 49.62 ;
      RECT 231.705 50.8 231.895 53.82 ;
      RECT 230.075 53.82 231.895 53.99 ;
      RECT 230.075 53.99 230.245 55.33 ;
      RECT 230.935 53.99 231.105 55.33 ;
      RECT 229.005 49.62 229.175 52.07 ;
      RECT 231.365 49.62 231.895 50.8 ;
      RECT 229.505 51.155 229.835 52.005 ;
      RECT 229.585 50.545 229.755 51.155 ;
      RECT 230.185 49.79 231.055 50.8 ;
      RECT 230.525 50.8 231.055 51.835 ;
      RECT 234.4 51.665 234.93 51.835 ;
      RECT 234.175 49.895 234.93 50.065 ;
      RECT 234.76 50.065 234.93 51.665 ;
      RECT 234.76 51.835 234.93 53.755 ;
      RECT 234.725 53.755 234.93 54.765 ;
      RECT 232.525 51.665 233.055 51.835 ;
      RECT 232.405 54.765 232.575 55.525 ;
      RECT 229.915 55.525 232.575 55.695 ;
      RECT 232.885 50.085 233.055 51.665 ;
      RECT 232.405 53.755 233.055 54.765 ;
      RECT 229.915 55.695 231.265 55.7 ;
      RECT 232.885 51.835 233.055 53.755 ;
      RECT 233.685 50.085 233.975 52.505 ;
      RECT 233.925 52.795 234.225 53.43 ;
      RECT 233.685 52.505 234.225 52.795 ;
      RECT 233.685 53.43 234.225 53.585 ;
      RECT 233.685 55.6 234.215 55.77 ;
      RECT 233.685 53.585 234.095 55.6 ;
      RECT 232.545 49.705 232.715 50.315 ;
      RECT 235.225 49.705 235.395 52 ;
      RECT 232.545 49.535 235.395 49.705 ;
      RECT 233.225 53 233.755 53.17 ;
      RECT 233.345 50.085 233.515 53 ;
      RECT 228.785 54.16 228.955 55.33 ;
      RECT 231.365 54.16 231.535 55.33 ;
      RECT 229.645 54.16 229.815 55.33 ;
      RECT 231.005 52.72 231.535 52.89 ;
      RECT 231.365 52.89 231.535 53.59 ;
      RECT 231.365 51.09 231.535 52.72 ;
      RECT 230.505 54.16 230.675 55.33 ;
      RECT 229.005 52.72 229.68 52.89 ;
      RECT 229.005 52.58 229.175 52.72 ;
      RECT 229.005 52.89 229.175 53.59 ;
      RECT 233.32 54.765 233.49 55.865 ;
      RECT 233.32 56.535 233.535 56.59 ;
      RECT 233.285 55.865 233.535 56.535 ;
      RECT 233.365 57.28 233.67 59.99 ;
      RECT 233.365 56.59 233.535 57.28 ;
      RECT 233.32 53.755 233.515 54.765 ;
      RECT 231.825 56.64 232.355 56.81 ;
      RECT 232.005 55.865 232.175 56.64 ;
      RECT 229.95 56.64 230.48 56.81 ;
      RECT 230.31 60.16 234.55 60.33 ;
      RECT 233.805 56.71 234.55 56.88 ;
      RECT 233.875 56.64 234.405 56.71 ;
      RECT 230.31 56.81 230.48 60.16 ;
      RECT 234.38 56.88 234.55 60.16 ;
      RECT 231.19 57.01 231.45 59.99 ;
      RECT 231.65 57.01 231.91 59.99 ;
      RECT 232.525 56.71 233.195 56.88 ;
      RECT 232.585 55.97 233.115 56.14 ;
      RECT 232.62 56.14 233.115 56.71 ;
      RECT 232.62 56.88 232.79 59.99 ;
      RECT 233.705 55.97 234.735 56.14 ;
      RECT 234.565 56.14 234.735 56.535 ;
      RECT 234.565 55.865 234.735 55.97 ;
      RECT 235.225 59.255 235.395 60.32 ;
      RECT 235.225 58.725 235.41 59.255 ;
      RECT 235.225 52.61 235.395 58.725 ;
      RECT 234.46 55.085 234.995 55.66 ;
      RECT 234.42 52.87 234.59 53.54 ;
      RECT 234.265 53.755 234.435 54.765 ;
      RECT 248.47 49.415 249.14 50.365 ;
      RECT 249.575 51.74 250.105 51.91 ;
      RECT 248.735 50.875 248.945 51.885 ;
      RECT 247.455 53.935 248.945 54.055 ;
      RECT 247.455 53.77 247.985 53.935 ;
      RECT 247.455 54.66 247.625 55.565 ;
      RECT 248.78 54.385 250.105 54.66 ;
      RECT 248.745 51.885 248.945 52.875 ;
      RECT 247.455 54.055 250.105 54.385 ;
      RECT 247.455 54.385 247.985 54.66 ;
      RECT 249.575 53.77 250.105 54.055 ;
      RECT 249.655 50.875 250.105 51.74 ;
      RECT 214.67 53.755 214.875 54.765 ;
      RECT 215.01 52.87 215.18 53.54 ;
      RECT 216.545 51.665 217.075 51.835 ;
      RECT 217.025 54.765 217.195 55.525 ;
      RECT 217.025 55.525 219.685 55.695 ;
      RECT 216.545 50.085 216.715 51.665 ;
      RECT 216.545 53.755 217.195 54.765 ;
      RECT 218.335 55.695 219.685 55.7 ;
      RECT 216.545 51.835 216.715 53.755 ;
      RECT 215.375 52.795 215.675 53.43 ;
      RECT 215.375 52.505 215.915 52.795 ;
      RECT 215.625 50.085 215.915 52.505 ;
      RECT 215.375 53.43 215.915 53.585 ;
      RECT 215.385 55.6 215.915 55.77 ;
      RECT 215.505 53.585 215.915 55.6 ;
      RECT 215.845 53 216.375 53.17 ;
      RECT 216.085 50.085 216.255 53 ;
      RECT 216.11 54.765 216.28 55.865 ;
      RECT 216.065 56.535 216.28 56.59 ;
      RECT 216.065 55.865 216.315 56.535 ;
      RECT 215.93 57.28 216.235 59.99 ;
      RECT 216.065 56.59 216.235 57.28 ;
      RECT 216.085 53.755 216.28 54.765 ;
      RECT 215.165 53.755 215.335 54.765 ;
      RECT 214.865 56.14 215.035 56.535 ;
      RECT 214.865 55.865 215.035 55.97 ;
      RECT 214.865 55.97 215.895 56.14 ;
      RECT 216.405 56.71 217.075 56.88 ;
      RECT 216.485 55.97 217.015 56.14 ;
      RECT 216.485 56.14 216.98 56.71 ;
      RECT 216.81 56.88 216.98 59.99 ;
      RECT 215.05 60.16 219.29 60.33 ;
      RECT 219.12 56.64 219.65 56.81 ;
      RECT 215.195 56.64 215.725 56.71 ;
      RECT 215.05 56.71 215.795 56.88 ;
      RECT 215.05 56.88 215.22 60.16 ;
      RECT 219.12 56.81 219.29 60.16 ;
      RECT 217.365 54.905 217.895 55.075 ;
      RECT 217.365 49.78 217.535 54.905 ;
      RECT 221.965 54.89 222.495 55.06 ;
      RECT 221.85 56.24 222.38 56.41 ;
      RECT 222.07 55.06 222.38 56.24 ;
      RECT 222.185 49.78 222.355 54.89 ;
      RECT 217.705 49.45 220.595 49.62 ;
      RECT 217.705 50.8 217.895 53.82 ;
      RECT 217.705 53.82 219.525 53.99 ;
      RECT 218.495 53.99 218.665 55.33 ;
      RECT 219.355 53.99 219.525 55.33 ;
      RECT 217.705 49.62 218.235 50.8 ;
      RECT 220.425 49.62 220.595 52.07 ;
      RECT 218.065 52.72 218.595 52.89 ;
      RECT 218.065 52.89 218.235 53.59 ;
      RECT 218.065 51.09 218.235 52.72 ;
      RECT 219.245 52.24 221.775 52.41 ;
      RECT 220.215 53.82 221.775 53.99 ;
      RECT 219.245 52.41 219.415 53.59 ;
      RECT 220.215 53.99 220.385 55.33 ;
      RECT 221.075 53.99 221.245 55.33 ;
      RECT 221.605 52.41 221.775 53.82 ;
      RECT 219.245 51.09 219.415 52.24 ;
      RECT 218.545 50.8 219.075 51.835 ;
      RECT 218.545 49.79 219.415 50.8 ;
      RECT 219.765 51.155 220.095 52.005 ;
      RECT 219.845 50.545 220.015 51.155 ;
      RECT 221.245 51.665 221.775 51.835 ;
      RECT 221.605 51.835 221.775 52.07 ;
      RECT 221.605 49.79 221.775 51.665 ;
      RECT 219.92 52.72 220.595 52.89 ;
      RECT 220.425 52.58 220.595 52.72 ;
      RECT 220.425 52.89 220.595 53.59 ;
      RECT 217.245 56.64 217.775 56.81 ;
      RECT 217.425 55.865 217.595 56.64 ;
      RECT 218.065 54.16 218.235 55.33 ;
      RECT 218.925 54.16 219.095 55.33 ;
      RECT 218.15 57.01 218.41 59.99 ;
      RECT 217.69 57.01 217.95 59.99 ;
      RECT 220.04 55.53 221.39 55.7 ;
      RECT 220.04 55.5 221.29 55.53 ;
      RECT 219.785 54.16 219.955 55.33 ;
      RECT 221.85 56.915 222.52 57.085 ;
      RECT 221.37 56.735 222.335 56.905 ;
      RECT 223.725 59.555 224.105 60.575 ;
      RECT 221.37 55.87 221.9 56.04 ;
      RECT 221.85 56.905 222.335 56.915 ;
      RECT 221.37 56.04 221.68 56.735 ;
      RECT 221.965 60.575 224.105 60.665 ;
      RECT 221.965 57.085 222.335 60.575 ;
      RECT 221.85 60.665 224.105 60.835 ;
      RECT 221.505 54.16 221.675 55.33 ;
      RECT 220.645 54.16 220.815 55.33 ;
      RECT 222.55 55.48 222.835 55.65 ;
      RECT 222.55 55.65 222.72 56.555 ;
      RECT 222.55 56.555 223.015 56.725 ;
      RECT 222.845 56.725 223.015 57.305 ;
      RECT 222.665 54.555 222.835 55.48 ;
      RECT 222.845 57.305 223.555 57.775 ;
      RECT 223.385 57.775 223.555 60.015 ;
      RECT 221.51 57.075 221.68 57.305 ;
      RECT 221.51 57.305 221.795 60.015 ;
      RECT 223.56 52.97 224.105 53.14 ;
      RECT 223.935 53.14 224.105 53.17 ;
      RECT 223.935 50.17 224.105 52.97 ;
      RECT 224.715 50.17 224.885 52.88 ;
      RECT 223.155 50.17 223.325 52.88 ;
      RECT 225.495 52.97 226.04 53.14 ;
      RECT 225.495 53.14 225.665 53.17 ;
      RECT 225.495 50.17 225.665 52.97 ;
      RECT 226.275 50.17 226.445 52.88 ;
      RECT 223.275 49.82 226.325 49.955 ;
      RECT 223.115 49.65 226.485 49.82 ;
      RECT 227.825 51.665 228.355 51.835 ;
      RECT 227.825 51.835 227.995 52.07 ;
      RECT 227.825 49.79 227.995 51.665 ;
      RECT 226.765 55.48 227.05 55.65 ;
      RECT 226.88 55.65 227.05 56.555 ;
      RECT 226.585 56.555 227.05 56.725 ;
      RECT 226.585 56.725 226.755 57.305 ;
      RECT 226.045 57.305 226.755 57.775 ;
      RECT 226.045 57.775 226.215 60.015 ;
      RECT 226.765 52.095 226.935 55.48 ;
      RECT 227.105 54.89 227.635 55.06 ;
      RECT 227.22 56.24 227.75 56.41 ;
      RECT 227.22 55.06 227.53 56.24 ;
      RECT 227.245 49.78 227.415 54.89 ;
      RECT 224.94 53.43 225.95 53.6 ;
      RECT 225.42 53.37 225.95 53.43 ;
      RECT 223.65 53.43 224.66 53.6 ;
      RECT 168.23 51.835 168.4 52.07 ;
      RECT 168.23 49.79 168.4 51.665 ;
      RECT 168.23 52.24 170.76 52.41 ;
      RECT 168.23 53.82 169.79 53.99 ;
      RECT 168.23 52.41 168.4 53.82 ;
      RECT 168.76 53.99 168.93 55.33 ;
      RECT 169.62 53.99 169.79 55.33 ;
      RECT 170.59 52.41 170.76 53.59 ;
      RECT 170.59 51.09 170.76 52.24 ;
      RECT 165.9 52.97 166.445 53.14 ;
      RECT 165.9 53.14 166.07 53.17 ;
      RECT 165.9 50.17 166.07 52.97 ;
      RECT 166.68 50.17 166.85 52.88 ;
      RECT 169.91 51.155 170.24 52.005 ;
      RECT 169.99 50.545 170.16 51.155 ;
      RECT 169.41 49.45 172.3 49.62 ;
      RECT 172.11 50.8 172.3 53.82 ;
      RECT 170.48 53.82 172.3 53.99 ;
      RECT 170.48 53.99 170.65 55.33 ;
      RECT 171.34 53.99 171.51 55.33 ;
      RECT 169.41 49.62 169.58 52.07 ;
      RECT 171.77 49.62 172.3 50.8 ;
      RECT 169.41 52.72 170.085 52.89 ;
      RECT 169.41 52.58 169.58 52.72 ;
      RECT 169.41 52.89 169.58 53.59 ;
      RECT 165.345 53.43 166.355 53.6 ;
      RECT 165.825 53.37 166.355 53.43 ;
      RECT 168.615 55.53 169.965 55.7 ;
      RECT 168.715 55.5 169.965 55.53 ;
      RECT 166.495 56.055 167.115 56.385 ;
      RECT 165.9 56.64 166.82 56.81 ;
      RECT 166.495 56.385 166.82 56.64 ;
      RECT 165.9 56.81 166.07 57.975 ;
      RECT 166.29 53.77 166.46 55.565 ;
      RECT 165.57 56 166.24 56.17 ;
      RECT 165.64 55.87 166.17 56 ;
      RECT 168.33 54.16 168.5 55.33 ;
      RECT 165.41 55.495 165.94 55.665 ;
      RECT 165.41 54.555 165.58 55.495 ;
      RECT 168.105 55.87 168.635 56.04 ;
      RECT 167.67 56.735 168.635 56.905 ;
      RECT 167.485 56.915 168.155 57.085 ;
      RECT 165.9 59.555 166.28 60.575 ;
      RECT 168.325 56.04 168.635 56.735 ;
      RECT 167.67 56.905 168.155 56.915 ;
      RECT 165.9 60.575 168.04 60.665 ;
      RECT 167.67 57.085 168.04 60.575 ;
      RECT 165.9 60.665 168.155 60.835 ;
      RECT 167.17 55.48 167.455 55.65 ;
      RECT 167.285 55.65 167.455 56.555 ;
      RECT 166.99 56.555 167.455 56.725 ;
      RECT 166.99 56.725 167.16 57.305 ;
      RECT 167.17 54.555 167.34 55.48 ;
      RECT 166.45 57.305 167.16 57.775 ;
      RECT 166.45 57.775 166.62 60.015 ;
      RECT 170.32 55.525 172.98 55.695 ;
      RECT 172.81 54.765 172.98 55.525 ;
      RECT 172.93 51.665 173.46 51.835 ;
      RECT 170.32 55.695 171.67 55.7 ;
      RECT 172.81 53.755 173.46 54.765 ;
      RECT 173.29 50.085 173.46 51.665 ;
      RECT 173.29 51.835 173.46 53.755 ;
      RECT 170.05 54.16 170.22 55.33 ;
      RECT 169.19 54.16 169.36 55.33 ;
      RECT 170.355 56.64 170.885 56.81 ;
      RECT 170.715 60.16 174.955 60.33 ;
      RECT 174.21 56.71 174.955 56.88 ;
      RECT 174.28 56.64 174.81 56.71 ;
      RECT 170.715 56.81 170.885 60.16 ;
      RECT 174.785 56.88 174.955 60.16 ;
      RECT 168.325 57.075 168.495 57.305 ;
      RECT 168.21 57.305 168.495 60.015 ;
      RECT 170.91 54.16 171.08 55.33 ;
      RECT 171.41 52.72 171.94 52.89 ;
      RECT 171.77 52.89 171.94 53.59 ;
      RECT 171.77 51.09 171.94 52.72 ;
      RECT 170.93 50.8 171.46 51.835 ;
      RECT 170.59 49.79 171.46 50.8 ;
      RECT 171.77 54.16 171.94 55.33 ;
      RECT 172.95 49.705 173.12 50.315 ;
      RECT 175.63 49.705 175.8 52 ;
      RECT 172.95 49.535 175.8 49.705 ;
      RECT 172.11 54.905 172.64 55.075 ;
      RECT 172.47 49.78 172.64 54.905 ;
      RECT 174.33 52.795 174.63 53.43 ;
      RECT 174.09 52.505 174.63 52.795 ;
      RECT 174.09 50.085 174.38 52.505 ;
      RECT 174.09 53.43 174.63 53.585 ;
      RECT 174.09 55.6 174.62 55.77 ;
      RECT 174.09 53.585 174.5 55.6 ;
      RECT 173.63 53 174.16 53.17 ;
      RECT 173.75 50.085 173.92 53 ;
      RECT 173.725 54.765 173.895 55.865 ;
      RECT 173.725 56.535 173.94 56.59 ;
      RECT 173.69 55.865 173.94 56.535 ;
      RECT 173.77 57.28 174.075 59.99 ;
      RECT 173.77 56.59 173.94 57.28 ;
      RECT 173.725 53.755 173.92 54.765 ;
      RECT 175.63 52.61 175.8 63.485 ;
      RECT 174.865 55.085 175.4 55.66 ;
      RECT 174.805 51.665 175.335 51.835 ;
      RECT 174.58 49.895 175.335 50.065 ;
      RECT 175.165 50.065 175.335 51.665 ;
      RECT 175.165 51.835 175.335 53.755 ;
      RECT 175.13 53.755 175.335 54.765 ;
      RECT 174.825 52.87 174.995 53.54 ;
      RECT 174.67 53.755 174.84 54.765 ;
      RECT 171.595 57.01 171.855 59.99 ;
      RECT 172.23 56.64 172.76 56.81 ;
      RECT 172.41 55.865 172.58 56.64 ;
      RECT 172.93 56.71 173.6 56.88 ;
      RECT 172.99 55.97 173.52 56.14 ;
      RECT 173.025 56.14 173.52 56.71 ;
      RECT 173.025 56.88 173.195 59.99 ;
      RECT 172.055 57.01 172.315 59.99 ;
      RECT 174.11 55.97 175.14 56.14 ;
      RECT 174.97 56.14 175.14 56.535 ;
      RECT 174.97 55.865 175.14 55.97 ;
      RECT 214.205 49.705 214.375 52 ;
      RECT 214.205 49.535 217.055 49.705 ;
      RECT 216.885 49.705 217.055 50.315 ;
      RECT 214.205 52.61 214.375 63.485 ;
      RECT 214.605 55.085 215.14 55.66 ;
      RECT 214.67 51.665 215.2 51.835 ;
      RECT 214.67 49.895 215.425 50.065 ;
      RECT 214.67 50.065 214.84 51.665 ;
      RECT 214.67 51.835 214.84 53.755 ;
      RECT 155.075 49.895 155.83 50.065 ;
      RECT 155.075 50.065 155.245 51.665 ;
      RECT 155.075 51.835 155.245 53.755 ;
      RECT 155.075 53.755 155.28 54.765 ;
      RECT 156.95 51.665 157.48 51.835 ;
      RECT 157.43 54.765 157.6 55.525 ;
      RECT 157.43 55.525 160.09 55.695 ;
      RECT 156.95 50.085 157.12 51.665 ;
      RECT 156.95 53.755 157.6 54.765 ;
      RECT 158.74 55.695 160.09 55.7 ;
      RECT 156.95 51.835 157.12 53.755 ;
      RECT 156.03 50.085 156.32 52.505 ;
      RECT 155.78 52.795 156.08 53.43 ;
      RECT 155.78 52.505 156.32 52.795 ;
      RECT 155.78 53.43 156.32 53.585 ;
      RECT 155.79 55.6 156.32 55.77 ;
      RECT 155.91 53.585 156.32 55.6 ;
      RECT 156.25 53 156.78 53.17 ;
      RECT 156.49 50.085 156.66 53 ;
      RECT 158.11 50.8 158.3 53.82 ;
      RECT 158.11 49.45 161 49.62 ;
      RECT 158.11 53.82 159.93 53.99 ;
      RECT 158.9 53.99 159.07 55.33 ;
      RECT 159.76 53.99 159.93 55.33 ;
      RECT 158.11 49.62 158.64 50.8 ;
      RECT 160.83 49.62 161 52.07 ;
      RECT 158.95 49.79 159.82 50.8 ;
      RECT 158.95 50.8 159.48 51.835 ;
      RECT 154.61 59.255 154.78 60.32 ;
      RECT 154.595 58.725 154.78 59.255 ;
      RECT 154.61 52.61 154.78 58.725 ;
      RECT 155.01 55.085 155.545 55.66 ;
      RECT 155.415 52.87 155.585 53.54 ;
      RECT 156.515 54.765 156.685 55.865 ;
      RECT 156.47 56.535 156.685 56.59 ;
      RECT 156.47 55.865 156.72 56.535 ;
      RECT 156.335 57.28 156.64 59.99 ;
      RECT 156.47 56.59 156.64 57.28 ;
      RECT 156.49 53.755 156.685 54.765 ;
      RECT 155.57 53.755 155.74 54.765 ;
      RECT 158.47 54.16 158.64 55.33 ;
      RECT 158.47 52.72 159 52.89 ;
      RECT 158.47 52.89 158.64 53.59 ;
      RECT 158.47 51.09 158.64 52.72 ;
      RECT 155.27 56.14 155.44 56.535 ;
      RECT 155.27 55.865 155.44 55.97 ;
      RECT 155.27 55.97 156.3 56.14 ;
      RECT 156.81 56.71 157.48 56.88 ;
      RECT 156.89 55.97 157.42 56.14 ;
      RECT 156.89 56.14 157.385 56.71 ;
      RECT 157.215 56.88 157.385 59.99 ;
      RECT 155.455 60.16 159.695 60.33 ;
      RECT 159.525 56.64 160.055 56.81 ;
      RECT 155.6 56.64 156.13 56.71 ;
      RECT 155.455 56.71 156.2 56.88 ;
      RECT 155.455 56.88 155.625 60.16 ;
      RECT 159.525 56.81 159.695 60.16 ;
      RECT 157.65 56.64 158.18 56.81 ;
      RECT 157.83 55.865 158 56.64 ;
      RECT 158.555 57.01 158.815 59.99 ;
      RECT 158.095 57.01 158.355 59.99 ;
      RECT 162.37 54.89 162.9 55.06 ;
      RECT 162.255 56.24 162.785 56.41 ;
      RECT 162.475 55.06 162.785 56.24 ;
      RECT 162.59 49.78 162.76 54.89 ;
      RECT 160.17 51.155 160.5 52.005 ;
      RECT 160.25 50.545 160.42 51.155 ;
      RECT 161.65 51.665 162.18 51.835 ;
      RECT 162.01 51.835 162.18 52.07 ;
      RECT 162.01 49.79 162.18 51.665 ;
      RECT 159.65 52.24 162.18 52.41 ;
      RECT 160.62 53.82 162.18 53.99 ;
      RECT 159.65 52.41 159.82 53.59 ;
      RECT 160.62 53.99 160.79 55.33 ;
      RECT 161.48 53.99 161.65 55.33 ;
      RECT 162.01 52.41 162.18 53.82 ;
      RECT 159.65 51.09 159.82 52.24 ;
      RECT 160.325 52.72 161 52.89 ;
      RECT 160.83 52.58 161 52.72 ;
      RECT 160.83 52.89 161 53.59 ;
      RECT 162.955 55.48 163.24 55.65 ;
      RECT 162.955 55.65 163.125 56.555 ;
      RECT 162.955 56.555 163.42 56.725 ;
      RECT 163.25 56.725 163.42 57.305 ;
      RECT 163.25 57.305 163.96 57.775 ;
      RECT 163.79 57.775 163.96 60.015 ;
      RECT 163.07 52.095 163.24 55.48 ;
      RECT 163.965 52.97 164.51 53.14 ;
      RECT 164.34 53.14 164.51 53.17 ;
      RECT 164.34 50.17 164.51 52.97 ;
      RECT 163.56 50.17 163.73 52.88 ;
      RECT 163.68 49.82 166.73 49.955 ;
      RECT 163.52 49.65 166.89 49.82 ;
      RECT 160.445 55.53 161.795 55.7 ;
      RECT 160.445 55.5 161.695 55.53 ;
      RECT 160.19 54.16 160.36 55.33 ;
      RECT 161.91 54.16 162.08 55.33 ;
      RECT 161.05 54.16 161.22 55.33 ;
      RECT 159.33 54.16 159.5 55.33 ;
      RECT 161.775 55.87 162.305 56.04 ;
      RECT 161.775 56.735 162.74 56.905 ;
      RECT 162.255 56.915 162.925 57.085 ;
      RECT 164.13 59.555 164.51 60.575 ;
      RECT 161.775 56.04 162.085 56.735 ;
      RECT 162.255 56.905 162.74 56.915 ;
      RECT 162.37 60.575 164.51 60.665 ;
      RECT 162.37 57.085 162.74 60.575 ;
      RECT 162.255 60.665 164.51 60.835 ;
      RECT 164.055 53.43 165.065 53.6 ;
      RECT 164.055 53.37 164.585 53.43 ;
      RECT 163.295 56.055 163.915 56.385 ;
      RECT 163.59 56.64 164.51 56.81 ;
      RECT 163.59 56.385 163.915 56.64 ;
      RECT 164.34 56.81 164.51 57.975 ;
      RECT 163.95 53.77 164.12 55.565 ;
      RECT 164.17 56 164.84 56.17 ;
      RECT 164.24 55.87 164.77 56 ;
      RECT 164.47 55.495 165 55.665 ;
      RECT 164.83 54.555 165 55.495 ;
      RECT 161.915 57.075 162.085 57.305 ;
      RECT 161.915 57.305 162.2 60.015 ;
      RECT 167.51 54.89 168.04 55.06 ;
      RECT 167.625 56.24 168.155 56.41 ;
      RECT 167.625 55.06 167.935 56.24 ;
      RECT 167.65 49.78 167.82 54.89 ;
      RECT 165.12 50.17 165.29 52.88 ;
      RECT 168.23 51.665 168.76 51.835 ;
      RECT 124.09 50.995 124.84 60.365 ;
      RECT 123.66 49.985 123.83 54.895 ;
      RECT 119.63 55.455 119.8 60.365 ;
      RECT 123.66 55.455 123.83 60.365 ;
      RECT 125.08 54.985 125.59 55.315 ;
      RECT 125.06 52.63 125.59 52.8 ;
      RECT 125.08 52.8 125.47 54.985 ;
      RECT 125.08 51.955 125.47 52.63 ;
      RECT 125.985 51.235 126.655 51.405 ;
      RECT 125.985 58.715 127.335 58.885 ;
      RECT 126.88 52.21 127.15 58.715 ;
      RECT 126.1 51.405 126.37 58.715 ;
      RECT 125.105 51.235 125.775 51.785 ;
      RECT 125.76 51.955 125.93 58.495 ;
      RECT 123.41 60.615 125.47 60.785 ;
      RECT 125.3 55.785 125.47 60.615 ;
      RECT 123.41 60.555 124.08 60.615 ;
      RECT 127.32 51.955 127.49 58.495 ;
      RECT 126.54 51.765 126.995 51.935 ;
      RECT 126.825 50.515 126.995 51.765 ;
      RECT 126.54 51.935 126.71 58.495 ;
      RECT 129.135 51.235 129.805 51.405 ;
      RECT 128.455 58.715 129.805 58.885 ;
      RECT 128.64 52.21 128.91 58.715 ;
      RECT 129.42 51.405 129.69 58.715 ;
      RECT 128.3 51.955 128.47 58.495 ;
      RECT 127.81 51.665 127.98 58.425 ;
      RECT 128.795 51.765 129.25 51.935 ;
      RECT 128.795 50.515 128.965 51.765 ;
      RECT 129.08 51.935 129.25 58.495 ;
      RECT 129.86 51.955 130.03 58.495 ;
      RECT 130.015 51.235 130.685 51.785 ;
      RECT 132.39 49.985 132.83 60.365 ;
      RECT 133.345 60.535 137.075 60.855 ;
      RECT 133.35 49.595 134.02 60.535 ;
      RECT 133.01 49.985 133.18 60.365 ;
      RECT 134.19 49.955 134.98 54.705 ;
      RECT 134.19 54.705 134.36 60.365 ;
      RECT 131.96 49.985 132.13 54.895 ;
      RECT 135.51 53.37 136.04 53.54 ;
      RECT 135.59 53.54 135.76 54.705 ;
      RECT 135.59 49.955 135.76 53.37 ;
      RECT 130.2 54.985 130.71 55.315 ;
      RECT 130.2 52.63 130.73 52.8 ;
      RECT 130.32 52.8 130.71 54.985 ;
      RECT 130.32 51.955 130.71 52.63 ;
      RECT 130.32 60.615 132.38 60.785 ;
      RECT 130.32 55.785 130.49 60.615 ;
      RECT 131.71 60.555 132.38 60.615 ;
      RECT 131.96 55.455 132.13 60.365 ;
      RECT 134.81 55.085 137.34 55.285 ;
      RECT 136.355 49.955 136.525 55.085 ;
      RECT 134.81 55.285 134.98 60.365 ;
      RECT 137.17 55.285 137.34 60.365 ;
      RECT 137.135 50.845 137.97 54.705 ;
      RECT 137.59 55.895 138.12 56.065 ;
      RECT 137.135 49.955 137.305 50.845 ;
      RECT 137.8 54.705 137.97 55.895 ;
      RECT 139.045 53.995 139.375 54.325 ;
      RECT 141.43 52.355 141.94 52.685 ;
      RECT 140.64 50.535 141.73 50.705 ;
      RECT 141.56 52.685 141.73 52.84 ;
      RECT 141.56 50.705 141.73 52.355 ;
      RECT 140.64 50.705 140.81 51.885 ;
      RECT 140.255 52.23 140.785 52.4 ;
      RECT 140.255 52.4 140.585 52.605 ;
      RECT 140.255 52.095 140.585 52.23 ;
      RECT 139.2 53.37 139.73 53.54 ;
      RECT 139.56 56.265 140.09 56.435 ;
      RECT 139.56 50.845 139.73 53.37 ;
      RECT 139.56 53.54 139.73 56.265 ;
      RECT 140.865 49.415 141.535 50.365 ;
      RECT 139.9 51.74 140.43 51.91 ;
      RECT 141.06 50.875 141.27 51.885 ;
      RECT 141.06 53.935 142.55 54.055 ;
      RECT 142.02 53.77 142.55 53.935 ;
      RECT 139.9 53.77 140.43 54.055 ;
      RECT 139.9 54.385 141.225 54.66 ;
      RECT 142.38 54.66 142.55 55.565 ;
      RECT 139.9 51.91 140.085 52.775 ;
      RECT 141.06 51.885 141.26 52.875 ;
      RECT 139.9 54.055 142.55 54.385 ;
      RECT 142.02 54.385 142.55 54.66 ;
      RECT 139.9 52.775 140.35 53.77 ;
      RECT 139.9 50.875 140.35 51.74 ;
      RECT 141.06 52.875 141.27 53.935 ;
      RECT 142.2 50.865 142.37 53.77 ;
      RECT 140.64 52.875 140.81 53.885 ;
      RECT 138.68 50.845 138.85 55.525 ;
      RECT 137.95 58.725 138.84 59.255 ;
      RECT 137.95 59.255 138.8 60.485 ;
      RECT 137.95 56.755 138.8 58.725 ;
      RECT 138.095 56.265 138.625 56.435 ;
      RECT 138.295 55.785 138.625 56.265 ;
      RECT 135.99 55.455 136.16 60.365 ;
      RECT 138.84 55.895 139.37 56.065 ;
      RECT 139.04 56.065 139.37 56.295 ;
      RECT 139.04 55.785 139.37 55.895 ;
      RECT 140.56 57.175 141.195 57.205 ;
      RECT 140.695 55.525 141.225 57.005 ;
      RECT 140.56 57.205 140.73 60.015 ;
      RECT 140.56 57.005 141.225 57.175 ;
      RECT 141.14 54.92 141.67 55.09 ;
      RECT 141.395 56.87 142.29 57.04 ;
      RECT 141.395 55.565 141.565 56.87 ;
      RECT 141.395 55.09 141.67 55.565 ;
      RECT 141.395 54.555 141.67 54.92 ;
      RECT 142.12 57.04 142.29 60.015 ;
      RECT 141.735 56.515 142.94 56.7 ;
      RECT 141.735 55.735 142.245 56.265 ;
      RECT 141.735 56.265 142.265 56.515 ;
      RECT 142.77 56.7 142.94 57.68 ;
      RECT 142.77 58.805 143.38 60.665 ;
      RECT 142.665 55.895 143.38 56.065 ;
      RECT 142.71 56.065 143.38 56.345 ;
      RECT 142.71 55.835 143.38 55.895 ;
      RECT 140.615 60.665 143.38 60.835 ;
      RECT 143.11 56.345 143.38 58.805 ;
      RECT 143.55 56.67 143.72 60.405 ;
      RECT 142.9 55.495 143.43 55.665 ;
      RECT 143.26 54.555 143.43 55.495 ;
      RECT 157.77 54.905 158.3 55.075 ;
      RECT 157.77 49.78 157.94 54.905 ;
      RECT 154.61 49.705 154.78 52 ;
      RECT 154.61 49.535 157.46 49.705 ;
      RECT 157.29 49.705 157.46 50.315 ;
      RECT 155.075 51.665 155.605 51.835 ;
      RECT 81.365 58.31 82.37 58.48 ;
      RECT 81.365 56.295 81.735 58.31 ;
      RECT 81.365 58.48 81.735 62.375 ;
      RECT 83.295 55.965 83.805 56.295 ;
      RECT 83.365 56.295 83.735 62.375 ;
      RECT 83.295 62.375 83.805 62.705 ;
      RECT 78.385 56.465 78.555 57.515 ;
      RECT 81.905 56.465 82.075 57.515 ;
      RECT 83.025 56.465 83.195 57.515 ;
      RECT 80.145 56.465 80.315 57.515 ;
      RECT 79.265 56.465 79.435 62.21 ;
      RECT 81.025 56.465 81.195 62.21 ;
      RECT 83.81 51 85.16 51.41 ;
      RECT 85.545 50.865 86.895 51.17 ;
      RECT 87.93 50.96 90.98 51.13 ;
      RECT 90.78 50.08 90.95 50.96 ;
      RECT 84.175 55.965 84.685 56.295 ;
      RECT 84.175 62.375 84.685 62.705 ;
      RECT 84.245 58.495 84.615 62.375 ;
      RECT 84.245 56.295 84.615 58.25 ;
      RECT 84.245 58.25 85.545 58.495 ;
      RECT 85.375 58.495 85.545 62.21 ;
      RECT 85.375 56.465 85.545 58.25 ;
      RECT 85.715 56.295 86.085 62.375 ;
      RECT 85.645 62.375 86.155 62.705 ;
      RECT 85.645 55.965 93.19 56.295 ;
      RECT 93.02 55.765 93.19 55.965 ;
      RECT 85.1 53.37 85.63 53.54 ;
      RECT 85.29 53.54 85.46 54.43 ;
      RECT 85.29 51.72 85.46 53.37 ;
      RECT 86.69 53.37 87.22 53.54 ;
      RECT 87.05 53.54 87.22 54.43 ;
      RECT 87.05 51.72 87.22 53.37 ;
      RECT 84.785 56.465 84.955 57.515 ;
      RECT 86.255 56.465 86.425 57.515 ;
      RECT 89.355 50 89.525 50.67 ;
      RECT 89.25 56.635 89.92 56.805 ;
      RECT 88.48 53 89.01 53.17 ;
      RECT 88.48 53.17 88.65 54.43 ;
      RECT 88.48 51.72 88.65 53 ;
      RECT 85.995 53 86.525 53.17 ;
      RECT 86.17 53.17 86.34 54.43 ;
      RECT 86.17 51.72 86.34 53 ;
      RECT 84.21 51.64 84.74 51.81 ;
      RECT 84.41 51.81 84.58 54.43 ;
      RECT 83.905 56.465 84.075 62.205 ;
      RECT 91.3 50.405 91.83 50.575 ;
      RECT 91.63 50.575 91.8 50.75 ;
      RECT 91.63 50.08 91.8 50.405 ;
      RECT 90.86 56.635 92.81 56.805 ;
      RECT 89.88 53 90.41 53.17 ;
      RECT 90.24 53.17 90.41 54.43 ;
      RECT 90.24 51.72 90.41 53 ;
      RECT 93.745 56.625 93.915 63.475 ;
      RECT 89.06 63.475 93.915 63.645 ;
      RECT 112.41 58.805 113.02 60.665 ;
      RECT 112.41 55.895 113.125 56.065 ;
      RECT 112.41 56.065 113.08 56.345 ;
      RECT 112.41 55.835 113.08 55.895 ;
      RECT 112.41 60.665 115.175 60.835 ;
      RECT 112.41 56.345 112.68 58.805 ;
      RECT 112.07 56.67 112.24 60.405 ;
      RECT 112.36 55.495 112.89 55.665 ;
      RECT 112.36 54.555 112.53 55.495 ;
      RECT 111.49 56.69 111.66 60.405 ;
      RECT 114.255 49.415 114.925 50.365 ;
      RECT 114.06 50.535 115.15 50.705 ;
      RECT 113.85 52.355 114.36 52.685 ;
      RECT 114.98 50.705 115.15 51.885 ;
      RECT 114.06 52.685 114.23 52.84 ;
      RECT 114.06 50.705 114.23 52.355 ;
      RECT 116.06 53.37 116.59 53.54 ;
      RECT 115.7 56.265 116.23 56.435 ;
      RECT 116.06 50.845 116.23 53.37 ;
      RECT 116.06 53.54 116.23 56.265 ;
      RECT 117.82 50.845 118.655 54.705 ;
      RECT 117.67 55.895 118.2 56.065 ;
      RECT 118.485 49.955 118.655 50.845 ;
      RECT 117.82 54.705 117.99 55.895 ;
      RECT 116.94 50.845 117.11 55.525 ;
      RECT 112.85 56.515 114.055 56.7 ;
      RECT 113.545 55.735 114.055 56.265 ;
      RECT 113.525 56.265 114.055 56.515 ;
      RECT 112.85 56.7 113.02 57.68 ;
      RECT 115.005 52.23 115.535 52.4 ;
      RECT 115.205 52.4 115.535 52.605 ;
      RECT 115.205 52.095 115.535 52.23 ;
      RECT 114.98 52.875 115.15 53.885 ;
      RECT 114.12 54.905 114.65 55.075 ;
      RECT 113.5 56.87 114.395 57.04 ;
      RECT 114.12 54.555 114.395 54.905 ;
      RECT 114.225 55.565 114.395 56.87 ;
      RECT 114.12 55.075 114.395 55.565 ;
      RECT 113.5 57.04 113.67 60.015 ;
      RECT 114.565 55.525 115.095 57.005 ;
      RECT 114.565 57.005 115.23 57.175 ;
      RECT 115.06 57.175 115.23 60.015 ;
      RECT 116.43 53.995 116.76 54.325 ;
      RECT 116.42 55.895 116.95 56.065 ;
      RECT 116.42 56.065 116.75 56.295 ;
      RECT 116.42 55.785 116.75 55.895 ;
      RECT 117.165 56.265 117.695 56.435 ;
      RECT 117.165 55.785 117.495 56.265 ;
      RECT 116.95 58.725 117.84 59.255 ;
      RECT 116.99 59.255 117.84 60.485 ;
      RECT 116.99 56.755 117.84 58.725 ;
      RECT 118.45 55.085 120.98 55.285 ;
      RECT 119.265 49.955 119.435 55.085 ;
      RECT 118.45 55.285 118.62 60.365 ;
      RECT 120.81 55.285 120.98 60.365 ;
      RECT 119.75 53.37 120.28 53.54 ;
      RECT 120.03 53.54 120.2 54.705 ;
      RECT 120.03 49.955 120.2 53.37 ;
      RECT 120.81 49.955 121.6 54.705 ;
      RECT 121.43 54.705 121.6 60.365 ;
      RECT 118.715 60.535 122.445 60.855 ;
      RECT 121.77 49.595 122.44 60.535 ;
      RECT 122.61 49.985 122.78 60.365 ;
      RECT 122.96 49.985 123.4 60.365 ;
      RECT 127.165 50.345 128.625 50.995 ;
      RECT 130.95 60.365 131.12 60.445 ;
      RECT 124.67 60.365 124.84 60.445 ;
      RECT 129.135 50.345 131.7 50.995 ;
      RECT 124.67 49.805 131.12 49.985 ;
      RECT 124.09 50.345 126.655 50.995 ;
      RECT 124.09 49.985 131.7 50.345 ;
      RECT 130.95 50.995 131.7 60.365 ;
      RECT 461.18 48.12 461.445 51.135 ;
      RECT 461.18 47.605 461.35 48.12 ;
      RECT 467.555 47.625 468.065 47.955 ;
      RECT 467.625 47.955 467.995 51.95 ;
      RECT 468.435 47.705 468.945 47.955 ;
      RECT 468.415 46.665 468.945 47.705 ;
      RECT 469.485 48.995 470.045 49.315 ;
      RECT 469.65 49.315 469.82 53.135 ;
      RECT 469.65 48.385 469.82 48.995 ;
      RECT 471.21 48.385 471.38 53.135 ;
      RECT 466.925 51.5 467.455 51.67 ;
      RECT 466.845 47.705 467.375 47.875 ;
      RECT 467.205 48.12 467.455 51.5 ;
      RECT 467.205 47.875 467.375 48.12 ;
      RECT 468.165 48.235 468.615 52.225 ;
      RECT 467.245 52.225 469.1 52.475 ;
      RECT 468.85 52.475 469.1 53.485 ;
      RECT 468.85 53.485 471.42 53.735 ;
      RECT 469.045 48.12 469.215 51.95 ;
      RECT 470.2 48.415 470.76 48.735 ;
      RECT 470.43 48.735 470.6 53.135 ;
      RECT 470.43 48.385 470.6 48.415 ;
      RECT 470.655 47.705 471.325 47.875 ;
      RECT 470.735 46.665 471.265 47.705 ;
      RECT 469.705 47.705 470.375 47.875 ;
      RECT 16.15 56.71 16.48 58.3 ;
      RECT 15.14 56.71 15.67 58.05 ;
      RECT 15.14 54.165 15.79 56.71 ;
      RECT 25.58 50.575 25.75 51.925 ;
      RECT 25.635 50.005 26.305 50.175 ;
      RECT 25.925 50.175 26.19 52.335 ;
      RECT 25.89 52.335 26.22 52.845 ;
      RECT 22.59 52.675 23.375 52.845 ;
      RECT 29.01 52.4 29.34 52.845 ;
      RECT 29.01 52.195 29.34 52.23 ;
      RECT 29.01 52.23 29.62 52.4 ;
      RECT 26.67 52.195 27 52.845 ;
      RECT 27.45 52.4 27.78 52.845 ;
      RECT 27.45 52.195 27.78 52.23 ;
      RECT 27.45 52.23 28.06 52.4 ;
      RECT 28.23 52.195 28.56 52.845 ;
      RECT 26.36 50.575 26.53 51.925 ;
      RECT 27.92 50.575 28.09 51.925 ;
      RECT 27.12 51.925 27.29 52.025 ;
      RECT 27.14 50.575 27.31 51.14 ;
      RECT 27.12 51.14 27.31 51.925 ;
      RECT 28.68 51.925 28.85 52.025 ;
      RECT 28.7 50.575 28.87 51.135 ;
      RECT 28.68 51.135 28.87 51.925 ;
      RECT 29.48 50.575 29.65 51.925 ;
      RECT 26.585 50.005 28.43 50.175 ;
      RECT 26.665 50 28.37 50.005 ;
      RECT 27.895 57.175 28.125 63.485 ;
      RECT 27.895 56.945 31.725 57.175 ;
      RECT 31.525 57.92 31.755 63.485 ;
      RECT 27.895 63.685 28.715 63.715 ;
      RECT 27.895 63.485 28.715 63.515 ;
      RECT 27.895 63.515 31.755 63.685 ;
      RECT 30.565 63.685 31.755 63.715 ;
      RECT 30.565 63.485 31.755 63.515 ;
      RECT 31.555 57.175 31.725 57.92 ;
      RECT 26.97 56.03 32.665 56.2 ;
      RECT 26.97 56.2 27.14 64.455 ;
      RECT 26.97 64.455 32.665 64.625 ;
      RECT 32.495 56.2 32.665 64.455 ;
      RECT 36.465 49.475 41.215 49.645 ;
      RECT 36.51 49.465 41.215 49.475 ;
      RECT 36.785 55.34 62.64 58.05 ;
      RECT 45.305 50.955 62.64 53.665 ;
      RECT 65.415 50.08 68.125 50.25 ;
      RECT 67.275 50.25 68.125 51 ;
      RECT 67.275 51 68.79 51.17 ;
      RECT 68.555 50.25 71.245 50.265 ;
      RECT 68.595 50.08 71.305 50.095 ;
      RECT 68.555 50.095 71.305 50.25 ;
      RECT 69.2 50.265 70.55 51.17 ;
      RECT 70.96 50.66 72.31 51.17 ;
      RECT 71.605 50.265 72.31 50.66 ;
      RECT 71.605 50.25 78.65 50.265 ;
      RECT 71.64 50.095 78.805 50.25 ;
      RECT 71.675 50.08 78.805 50.095 ;
      RECT 66.905 56.5 67.575 56.67 ;
      RECT 68.185 56.5 68.855 56.67 ;
      RECT 71.35 52.18 71.88 52.35 ;
      RECT 71.54 52.35 71.71 54.43 ;
      RECT 71.54 51.72 71.71 52.18 ;
      RECT 69.59 52.18 70.12 52.35 ;
      RECT 69.78 52.35 69.95 54.43 ;
      RECT 69.78 51.72 69.95 52.18 ;
      RECT 67.83 52.18 68.36 52.35 ;
      RECT 68.02 52.35 68.19 54.43 ;
      RECT 68.02 51.72 68.19 52.18 ;
      RECT 72.755 51 77.505 51.17 ;
      RECT 76.63 51.81 77.16 51.98 ;
      RECT 76.82 51.98 76.99 54.43 ;
      RECT 76.82 51.72 76.99 51.81 ;
      RECT 74.875 51.81 75.405 51.98 ;
      RECT 75.06 51.98 75.23 54.43 ;
      RECT 75.06 51.72 75.23 51.81 ;
      RECT 73.11 51.81 73.64 51.98 ;
      RECT 73.3 51.98 73.47 54.43 ;
      RECT 73.3 51.72 73.47 51.81 ;
      RECT 78.005 51 82.755 51.17 ;
      RECT 79.275 50.265 80.805 51 ;
      RECT 79.275 50.08 83.385 50.095 ;
      RECT 79.275 50.095 83.465 50.265 ;
      RECT 83.53 53.37 84.06 53.54 ;
      RECT 83.53 53.54 83.7 54.43 ;
      RECT 83.53 51.72 83.7 53.37 ;
      RECT 81.91 53.37 82.44 53.54 ;
      RECT 82.1 53.54 82.27 54.43 ;
      RECT 82.1 51.72 82.27 53.37 ;
      RECT 80.155 53.37 80.685 53.54 ;
      RECT 80.34 53.54 80.51 54.43 ;
      RECT 80.34 51.72 80.51 53.37 ;
      RECT 78.39 53.37 78.92 53.54 ;
      RECT 78.58 53.54 78.75 54.43 ;
      RECT 78.58 51.72 78.75 53.37 ;
      RECT 78.655 55.965 79.165 56.295 ;
      RECT 78.655 62.375 79.165 62.705 ;
      RECT 78.725 56.295 79.095 62.375 ;
      RECT 79.535 55.965 80.925 56.295 ;
      RECT 80.485 56.295 80.855 62.375 ;
      RECT 79.535 62.375 80.925 62.705 ;
      RECT 79.605 56.295 79.975 62.375 ;
      RECT 81.295 55.965 81.805 56.295 ;
      RECT 81.295 62.375 81.805 62.705 ;
      RECT 362.13 48.245 362.3 49.595 ;
      RECT 363.475 48.245 363.645 49.595 ;
      RECT 366.63 42.025 367.415 42.195 ;
      RECT 366.805 42.195 367.355 42.495 ;
      RECT 367.585 42.025 368.71 42.195 ;
      RECT 367.585 52.675 368.71 52.845 ;
      RECT 367.585 42.195 367.755 52.675 ;
      RECT 372.225 42.025 373.35 42.195 ;
      RECT 372.225 52.675 373.35 52.845 ;
      RECT 372.225 42.195 372.395 52.675 ;
      RECT 368.99 42.025 370.115 42.195 ;
      RECT 368.99 52.675 370.115 52.845 ;
      RECT 369.945 42.195 370.115 52.675 ;
      RECT 375.465 43.425 375.795 44.015 ;
      RECT 386.27 47.58 386.6 48.23 ;
      RECT 387.53 47.58 387.86 48.23 ;
      RECT 386.9 47.58 387.23 48.23 ;
      RECT 388.79 47.58 389.12 48.23 ;
      RECT 388.16 47.58 388.49 48.23 ;
      RECT 390.05 47.58 390.38 48.23 ;
      RECT 389.42 47.58 389.75 48.23 ;
      RECT 386.27 48.61 386.6 49.26 ;
      RECT 386.9 48.61 387.23 49.26 ;
      RECT 387.53 48.61 387.86 49.26 ;
      RECT 388.79 48.61 389.12 49.26 ;
      RECT 388.16 48.61 388.49 49.26 ;
      RECT 389.42 48.61 389.75 49.26 ;
      RECT 390.05 48.61 390.38 49.26 ;
      RECT 393.83 47.17 394.16 48.23 ;
      RECT 390.68 47.58 391.01 48.23 ;
      RECT 391.31 47.58 391.64 48.23 ;
      RECT 391.94 47.58 392.27 48.23 ;
      RECT 393.2 47.72 393.53 49.26 ;
      RECT 392.57 47.58 392.9 48.23 ;
      RECT 390.68 48.61 391.01 49.26 ;
      RECT 391.31 48.61 391.64 49.26 ;
      RECT 391.94 48.61 392.27 49.26 ;
      RECT 393.83 48.61 394.16 49.26 ;
      RECT 394.46 48.61 394.79 49.26 ;
      RECT 392.57 48.61 392.9 49.26 ;
      RECT 421.065 47.58 445.335 47.75 ;
      RECT 421.065 43.2 421.815 43.73 ;
      RECT 421.065 43.73 421.235 47.58 ;
      RECT 445.165 47.075 445.335 47.58 ;
      RECT 444.585 43.4 445.335 43.73 ;
      RECT 445.16 43.73 445.335 47.075 ;
      RECT 421.645 43.9 421.815 46.61 ;
      RECT 423.075 43.9 423.245 46.61 ;
      RECT 424.835 43.9 425.005 46.61 ;
      RECT 424.835 43.2 425.005 43.73 ;
      RECT 424.835 42.405 425.005 42.78 ;
      RECT 426.595 43.9 426.765 46.61 ;
      RECT 427.145 43.9 427.315 46.61 ;
      RECT 428.905 43.9 429.075 46.61 ;
      RECT 430.805 43.9 430.975 46.915 ;
      RECT 428.905 43.2 429.075 43.73 ;
      RECT 428.905 42.405 429.075 42.78 ;
      RECT 430.805 43.4 431.525 43.73 ;
      RECT 430.805 42.45 431.525 42.78 ;
      RECT 431.355 43.9 431.525 46.915 ;
      RECT 433.255 43.9 433.425 46.61 ;
      RECT 433.255 42.405 433.425 42.78 ;
      RECT 433.255 43.4 433.425 43.73 ;
      RECT 435.565 43.9 435.735 46.61 ;
      RECT 435.015 43.9 435.185 46.61 ;
      RECT 437.325 42.405 437.495 42.78 ;
      RECT 439.085 42.45 439.255 42.78 ;
      RECT 439.085 43.4 439.255 43.73 ;
      RECT 437.325 43.2 437.495 43.73 ;
      RECT 440.515 43.2 440.685 43.73 ;
      RECT 440.515 42.405 440.685 42.78 ;
      RECT 439.085 43.9 439.255 46.61 ;
      RECT 437.325 43.9 437.495 46.61 ;
      RECT 442.275 43.9 442.445 46.61 ;
      RECT 440.515 43.9 440.685 46.61 ;
      RECT 442.825 43.9 442.995 46.61 ;
      RECT 444.585 43.9 444.755 46.61 ;
      RECT 453.445 44.355 457.145 44.525 ;
      RECT 453.445 43.955 454.925 44.355 ;
      RECT 453.17 48.385 453.34 53.135 ;
      RECT 453.755 48.415 454.315 48.735 ;
      RECT 453.95 48.735 454.12 53.135 ;
      RECT 453.95 48.385 454.12 48.415 ;
      RECT 453.395 47.37 453.765 47.705 ;
      RECT 453.24 47.705 453.91 47.875 ;
      RECT 458.635 50.09 459.145 50.42 ;
      RECT 458.725 47.37 459.095 50.09 ;
      RECT 453.395 47 459.095 47.37 ;
      RECT 454.925 45.78 456.875 46.13 ;
      RECT 456.34 45.1 456.875 45.78 ;
      RECT 455.65 45.065 455.82 45.595 ;
      RECT 457.1 45.18 458.515 45.48 ;
      RECT 454.615 44.88 455.07 45.43 ;
      RECT 454.615 44.71 456.545 44.88 ;
      RECT 455.205 43.955 456.685 44.125 ;
      RECT 455.145 48.415 455.705 48.735 ;
      RECT 455.35 48.735 455.52 53.135 ;
      RECT 455.35 48.385 455.52 48.415 ;
      RECT 455.94 48.995 456.475 49.315 ;
      RECT 456.13 49.315 456.3 53.135 ;
      RECT 456.13 48.385 456.3 48.995 ;
      RECT 454.415 49.575 454.98 49.895 ;
      RECT 454.57 49.895 454.74 53.135 ;
      RECT 454.57 48.385 454.74 49.575 ;
      RECT 457.03 47.705 457.655 47.875 ;
      RECT 457.03 47.675 457.2 47.705 ;
      RECT 457.03 52.855 457.655 53.865 ;
      RECT 457.03 47.875 457.2 52.855 ;
      RECT 459.645 47.175 460.175 47.345 ;
      RECT 459.805 47.345 460.175 54.035 ;
      RECT 459.805 47.17 460.175 47.175 ;
      RECT 458.635 54.035 460.175 54.365 ;
      RECT 455.575 47.705 456.245 47.875 ;
      RECT 454.625 47.705 455.295 47.875 ;
      RECT 462.415 42.435 464.1 42.605 ;
      RECT 461.62 44.615 462.57 45.865 ;
      RECT 462.055 43.095 462.565 44.615 ;
      RECT 463.275 43.155 463.445 45.865 ;
      RECT 462.425 47.705 462.955 47.875 ;
      RECT 462.425 47.875 462.935 47.955 ;
      RECT 462.425 47.625 462.935 47.705 ;
      RECT 461.545 47.625 462.055 47.955 ;
      RECT 461.615 52.29 462.145 52.46 ;
      RECT 461.615 47.955 461.985 52.29 ;
      RECT 463.035 52.29 463.565 52.46 ;
      RECT 463.035 48.12 463.205 52.29 ;
      RECT 462.155 48.425 462.325 51.135 ;
      RECT 308.525 44.82 308.695 47.57 ;
      RECT 305.235 48.37 305.765 48.54 ;
      RECT 305.405 48.54 305.575 49.57 ;
      RECT 305.405 44.82 305.575 48.37 ;
      RECT 309.815 42.65 327.825 42.98 ;
      RECT 309.725 47.57 310.255 47.74 ;
      RECT 310.085 47.74 310.255 49.57 ;
      RECT 310.085 44.82 310.255 47.57 ;
      RECT 315.075 47.555 315.605 47.725 ;
      RECT 315.265 47.725 315.435 49.57 ;
      RECT 315.265 44.82 315.435 47.555 ;
      RECT 313.315 47.555 313.845 47.725 ;
      RECT 313.505 47.725 313.675 49.57 ;
      RECT 313.505 44.82 313.675 47.555 ;
      RECT 311.555 47.555 312.085 47.725 ;
      RECT 311.745 47.725 311.915 49.57 ;
      RECT 311.745 44.82 311.915 47.555 ;
      RECT 318.455 48.355 318.985 48.525 ;
      RECT 318.455 48.525 318.625 49.57 ;
      RECT 318.455 44.82 318.625 48.355 ;
      RECT 319.825 48.355 320.355 48.525 ;
      RECT 320.015 48.525 320.185 49.57 ;
      RECT 320.015 44.82 320.185 48.355 ;
      RECT 319.045 47.555 319.575 47.725 ;
      RECT 319.235 47.725 319.405 49.57 ;
      RECT 319.235 44.82 319.405 47.555 ;
      RECT 320.605 47.555 321.135 47.725 ;
      RECT 320.795 47.725 320.965 49.57 ;
      RECT 320.795 44.82 320.965 47.555 ;
      RECT 316.835 47.555 317.365 47.725 ;
      RECT 317.025 47.725 317.195 49.57 ;
      RECT 317.025 44.82 317.195 47.555 ;
      RECT 321.385 48.355 321.915 48.525 ;
      RECT 321.575 48.525 321.745 49.57 ;
      RECT 321.575 44.82 321.745 48.355 ;
      RECT 324.335 48.355 324.865 48.525 ;
      RECT 324.695 48.525 324.865 49.57 ;
      RECT 324.695 44.82 324.865 48.355 ;
      RECT 322.95 48.355 323.48 48.525 ;
      RECT 323.135 48.525 323.305 49.57 ;
      RECT 323.135 44.82 323.305 48.355 ;
      RECT 322.185 47.97 322.715 48.14 ;
      RECT 322.355 48.14 322.525 49.57 ;
      RECT 322.355 44.82 322.525 47.97 ;
      RECT 323.745 47.97 324.275 48.14 ;
      RECT 323.915 48.14 324.085 49.57 ;
      RECT 323.915 44.82 324.085 47.97 ;
      RECT 327.365 47.305 344.7 50.015 ;
      RECT 332.38 45.27 332.91 45.44 ;
      RECT 332.39 45.44 332.9 45.535 ;
      RECT 332.39 45.205 332.9 45.27 ;
      RECT 328.095 45.245 328.885 45.495 ;
      RECT 328.495 45.495 328.885 45.535 ;
      RECT 328.495 45.205 328.885 45.245 ;
      RECT 328.095 43.945 333.41 44.275 ;
      RECT 328.095 44.575 333.41 44.905 ;
      RECT 328.095 44.275 328.765 44.575 ;
      RECT 330.695 42.755 331.225 42.925 ;
      RECT 336.89 45.27 337.42 45.44 ;
      RECT 336.9 45.44 337.41 45.535 ;
      RECT 336.9 45.205 337.41 45.27 ;
      RECT 335.52 42.02 337.545 42.35 ;
      RECT 335.515 42.65 336.31 42.98 ;
      RECT 336.875 42.65 337.545 43.61 ;
      RECT 335.105 44.64 335.635 44.81 ;
      RECT 335.115 44.81 335.625 44.905 ;
      RECT 335.115 44.575 335.625 44.64 ;
      RECT 335.105 44.02 335.635 44.19 ;
      RECT 335.115 44.19 335.625 44.275 ;
      RECT 335.115 43.945 335.625 44.02 ;
      RECT 341.4 45.27 341.93 45.44 ;
      RECT 341.41 45.44 341.92 45.535 ;
      RECT 341.41 45.205 341.92 45.27 ;
      RECT 341.4 44.025 341.93 44.195 ;
      RECT 341.41 44.195 341.92 44.275 ;
      RECT 341.41 43.945 341.92 44.025 ;
      RECT 341.4 44.64 341.93 44.81 ;
      RECT 341.41 44.81 341.92 44.905 ;
      RECT 341.41 44.575 341.92 44.64 ;
      RECT 348.79 48.415 353.54 48.585 ;
      RECT 347.695 44.64 348.225 44.81 ;
      RECT 347.705 44.81 348.215 44.905 ;
      RECT 347.705 44.575 348.215 44.64 ;
      RECT 347.695 44.015 348.225 44.185 ;
      RECT 347.705 44.185 348.215 44.275 ;
      RECT 347.705 43.945 348.215 44.015 ;
      RECT 347.695 45.27 348.225 45.44 ;
      RECT 347.705 45.44 348.215 45.535 ;
      RECT 347.705 45.205 348.215 45.27 ;
      RECT 348.79 48.945 353.54 49.115 ;
      RECT 348.08 48.105 348.25 48.825 ;
      RECT 348.08 49.185 348.25 49.955 ;
      RECT 348.79 47.905 354.305 47.935 ;
      RECT 354.13 48.105 354.305 49.955 ;
      RECT 348.195 50.125 354.305 50.135 ;
      RECT 348.08 47.935 354.305 48.105 ;
      RECT 348.08 49.955 354.305 50.125 ;
      RECT 353.92 44.575 354.59 45.535 ;
      RECT 353.91 43.61 354.59 44.275 ;
      RECT 353.91 43.28 363.37 43.61 ;
      RECT 353.76 48.64 353.93 49.42 ;
      RECT 357.51 48.245 357.68 49.74 ;
      RECT 360.795 47.675 361.465 47.845 ;
      RECT 360.96 47.845 361.13 48.78 ;
      RECT 359.79 48.245 359.96 49.74 ;
      RECT 360.57 48.245 360.74 49.595 ;
      RECT 361.35 48.1 361.52 49.595 ;
      RECT 356.885 50.37 360.03 50.54 ;
      RECT 362.995 45.925 364.905 46.095 ;
      RECT 356.885 46.8 363.165 46.97 ;
      RECT 362.995 46.095 363.165 46.8 ;
      RECT 356.885 53.265 364.875 53.345 ;
      RECT 359.86 53.095 364.905 53.175 ;
      RECT 356.885 53.175 364.905 53.265 ;
      RECT 364.735 46.095 364.905 53.095 ;
      RECT 359.86 52.535 360.03 53.095 ;
      RECT 359.705 51.305 360.03 52.535 ;
      RECT 359.86 50.82 360.03 51.305 ;
      RECT 356.885 46.97 357.055 50.37 ;
      RECT 359.045 50.54 360.03 50.82 ;
      RECT 356.885 50.54 357.055 53.175 ;
      RECT 357.735 47.675 360.515 47.845 ;
      RECT 364.255 48.245 364.425 49.595 ;
      RECT 362.695 48.245 362.865 49.595 ;
      RECT 363.475 46.445 363.645 47.795 ;
      RECT 364.255 46.445 364.425 47.795 ;
      RECT 362.7 42.02 363.37 42.98 ;
      RECT 276.215 48.105 276.97 48.275 ;
      RECT 276.8 46.505 276.97 48.105 ;
      RECT 276.8 44.415 276.97 46.335 ;
      RECT 280.425 43.095 280.955 43.265 ;
      RECT 280.425 43.265 280.595 48.39 ;
      RECT 280.085 42.645 280.255 43.405 ;
      RECT 280.085 42.475 282.745 42.645 ;
      RECT 279.605 46.335 280.135 46.505 ;
      RECT 281.395 42.47 282.745 42.475 ;
      RECT 279.605 46.505 279.775 48.085 ;
      RECT 279.605 44.415 279.775 46.335 ;
      RECT 279.605 43.405 280.255 44.415 ;
      RECT 276.46 44.63 276.63 45.3 ;
      RECT 275.265 45 275.795 45.17 ;
      RECT 275.385 45.17 275.555 48.085 ;
      RECT 278.905 45 279.435 45.17 ;
      RECT 279.145 45.17 279.315 48.085 ;
      RECT 285.025 43.11 285.555 43.28 ;
      RECT 284.91 41.76 285.44 41.93 ;
      RECT 285.13 41.93 285.44 43.11 ;
      RECT 285.245 43.28 285.415 48.39 ;
      RECT 280.765 44.35 280.955 47.37 ;
      RECT 280.765 44.18 282.585 44.35 ;
      RECT 280.765 48.55 283.655 48.72 ;
      RECT 281.555 42.84 281.725 44.18 ;
      RECT 282.415 42.84 282.585 44.18 ;
      RECT 280.765 47.37 281.295 48.55 ;
      RECT 283.485 46.1 283.655 48.55 ;
      RECT 283.1 42.47 284.45 42.64 ;
      RECT 283.1 42.64 284.35 42.67 ;
      RECT 281.125 42.84 281.295 44.01 ;
      RECT 282.845 42.84 283.015 44.01 ;
      RECT 281.125 45.28 281.655 45.45 ;
      RECT 281.125 44.58 281.295 45.28 ;
      RECT 281.125 45.45 281.295 47.08 ;
      RECT 283.275 44.18 284.835 44.35 ;
      RECT 282.305 45.76 284.835 45.93 ;
      RECT 283.275 42.84 283.445 44.18 ;
      RECT 284.135 42.84 284.305 44.18 ;
      RECT 282.305 44.58 282.475 45.76 ;
      RECT 284.665 44.35 284.835 45.76 ;
      RECT 282.305 45.93 282.475 47.08 ;
      RECT 283.705 42.84 283.875 44.01 ;
      RECT 281.985 42.84 282.155 44.01 ;
      RECT 282.98 45.28 283.655 45.45 ;
      RECT 283.485 45.45 283.655 45.59 ;
      RECT 283.485 44.58 283.655 45.28 ;
      RECT 284.565 42.84 284.735 44.01 ;
      RECT 282.825 46.165 283.155 47.015 ;
      RECT 282.905 47.015 283.075 47.625 ;
      RECT 281.605 47.37 282.475 48.38 ;
      RECT 281.605 46.335 282.135 47.37 ;
      RECT 284.305 46.335 284.835 46.505 ;
      RECT 284.665 46.1 284.835 46.335 ;
      RECT 284.665 46.505 284.835 48.38 ;
      RECT 286.215 45.29 286.385 48 ;
      RECT 286.335 48.215 287.945 48.35 ;
      RECT 286.175 48.385 287.86 48.52 ;
      RECT 286.175 48.35 287.945 48.385 ;
      RECT 286.605 44.57 287.72 44.74 ;
      RECT 286.605 44.74 287.24 44.8 ;
      RECT 286.605 42.605 286.775 44.57 ;
      RECT 286.825 42 287.495 42.17 ;
      RECT 286.895 42.17 287.425 42.3 ;
      RECT 286.62 45.03 287.165 45.2 ;
      RECT 286.995 45 287.165 45.03 ;
      RECT 286.995 45.2 287.165 48 ;
      RECT 287.775 45.29 287.945 48 ;
      RECT 287.125 42.505 287.655 42.675 ;
      RECT 287.485 42.675 287.655 43.615 ;
      RECT 290.115 46.99 294.245 47.125 ;
      RECT 290.035 46.5 294.285 46.99 ;
      RECT 289.205 43.51 289.375 44.4 ;
      RECT 322.92 50.61 324.53 50.665 ;
      RECT 322.92 50.44 325.445 50.61 ;
      RECT 295.045 44.3 325.445 44.47 ;
      RECT 325.275 44.47 325.445 50.44 ;
      RECT 317.905 44.47 318.075 49.57 ;
      RECT 316.145 44.47 316.315 49.57 ;
      RECT 310.865 44.47 311.035 49.57 ;
      RECT 312.625 44.47 312.795 49.57 ;
      RECT 314.385 44.47 314.555 49.57 ;
      RECT 298.615 44.47 298.785 49.57 ;
      RECT 300.175 44.47 300.345 49.57 ;
      RECT 296.405 44.47 296.575 49.57 ;
      RECT 309.305 44.47 309.475 49.57 ;
      RECT 304.625 44.47 304.795 49.57 ;
      RECT 306.185 44.47 306.355 49.57 ;
      RECT 307.745 44.47 307.915 49.57 ;
      RECT 301.505 44.47 301.675 49.57 ;
      RECT 303.065 44.47 303.235 49.57 ;
      RECT 295.045 44.47 295.215 49.84 ;
      RECT 297.715 49.74 299.955 49.91 ;
      RECT 297.715 51.24 298.245 51.41 ;
      RECT 297.715 44.82 298.005 49.74 ;
      RECT 297.715 51.41 298.005 54.43 ;
      RECT 297.715 49.91 298.005 51.24 ;
      RECT 299.785 49.91 299.955 50.67 ;
      RECT 296.485 50.035 297.015 50.205 ;
      RECT 295.525 50.84 296.955 51.14 ;
      RECT 295.525 51.14 295.795 54.43 ;
      RECT 295.525 44.82 295.795 50.84 ;
      RECT 296.785 50.015 296.955 50.035 ;
      RECT 296.785 50.205 296.955 50.84 ;
      RECT 296.925 49.665 297.455 49.835 ;
      RECT 297.185 49.835 297.455 54.43 ;
      RECT 297.185 44.82 297.455 49.665 ;
      RECT 295.965 45.575 296.235 50 ;
      RECT 295.965 50 296.255 50.67 ;
      RECT 299.225 48.845 299.755 49.015 ;
      RECT 299.395 49.015 299.565 49.57 ;
      RECT 299.395 44.82 299.565 48.845 ;
      RECT 300.595 48.845 301.125 49.015 ;
      RECT 300.955 44.82 301.125 48.845 ;
      RECT 300.955 49.015 301.125 50.08 ;
      RECT 300.955 50.08 306.01 50.265 ;
      RECT 302.095 48.355 302.625 48.525 ;
      RECT 302.285 48.525 302.455 49.57 ;
      RECT 302.285 44.82 302.455 48.355 ;
      RECT 303.675 48.355 304.205 48.525 ;
      RECT 303.845 48.525 304.015 49.57 ;
      RECT 303.845 44.82 304.015 48.355 ;
      RECT 306.785 47.57 307.315 47.74 ;
      RECT 306.965 47.74 307.135 49.57 ;
      RECT 306.965 44.82 307.135 47.57 ;
      RECT 308.345 47.57 308.875 47.74 ;
      RECT 308.525 47.74 308.695 49.57 ;
      RECT 262.465 44.58 262.635 45.28 ;
      RECT 257.625 49.045 258.295 49.765 ;
      RECT 261.805 46.165 262.135 47.015 ;
      RECT 261.885 47.015 262.055 47.625 ;
      RECT 260.585 46.335 261.115 47.37 ;
      RECT 260.585 47.37 261.455 48.38 ;
      RECT 263.545 42.84 263.715 44.01 ;
      RECT 265.585 42.605 265.755 44.4 ;
      RECT 265.805 42 266.475 42.17 ;
      RECT 265.875 42.17 266.405 42.3 ;
      RECT 263.89 41.76 264.42 41.93 ;
      RECT 264.11 41.93 264.42 43.11 ;
      RECT 264.005 43.11 264.535 48.39 ;
      RECT 266.105 42.505 266.635 42.675 ;
      RECT 266.465 42.675 266.635 43.615 ;
      RECT 267.925 42.605 268.095 44.4 ;
      RECT 267.205 42 267.875 42.17 ;
      RECT 267.275 42.17 267.805 42.3 ;
      RECT 267.045 42.505 267.575 42.675 ;
      RECT 267.045 42.675 267.215 43.615 ;
      RECT 263.285 46.335 263.815 46.505 ;
      RECT 263.645 46.1 263.815 46.335 ;
      RECT 263.645 46.505 263.815 48.38 ;
      RECT 265.69 44.57 266.7 44.74 ;
      RECT 265.69 44.74 266.22 44.8 ;
      RECT 265.6 45.03 266.145 45.2 ;
      RECT 265.975 45 266.145 45.03 ;
      RECT 265.975 45.2 266.145 48 ;
      RECT 265.195 45.29 265.365 48 ;
      RECT 265.925 49.045 266.595 49.765 ;
      RECT 265.315 48.215 268.365 48.35 ;
      RECT 265.155 48.35 268.525 48.52 ;
      RECT 266.98 44.57 267.99 44.74 ;
      RECT 267.46 44.74 267.99 44.8 ;
      RECT 266.755 45.29 266.925 48 ;
      RECT 267.535 45.03 268.08 45.2 ;
      RECT 267.535 45 267.705 45.03 ;
      RECT 267.535 45.2 267.705 48 ;
      RECT 268.315 45.29 268.485 48 ;
      RECT 273.745 43.095 274.275 43.265 ;
      RECT 274.05 49.785 274.905 49.955 ;
      RECT 274.05 49.015 274.58 49.785 ;
      RECT 274.105 43.265 274.275 49.015 ;
      RECT 269.26 41.76 269.79 41.93 ;
      RECT 269.26 41.93 269.57 43.11 ;
      RECT 269.145 43.11 269.675 48.39 ;
      RECT 270.25 42.47 271.6 42.64 ;
      RECT 270.35 42.64 271.6 42.67 ;
      RECT 269.965 42.84 270.135 44.01 ;
      RECT 269.865 44.18 271.425 44.35 ;
      RECT 269.865 45.76 272.395 45.93 ;
      RECT 270.395 42.84 270.565 44.18 ;
      RECT 271.255 42.84 271.425 44.18 ;
      RECT 272.225 44.58 272.395 45.76 ;
      RECT 269.865 44.35 270.035 45.76 ;
      RECT 272.225 45.93 272.395 47.08 ;
      RECT 270.825 42.84 270.995 44.01 ;
      RECT 271.955 42.475 274.615 42.645 ;
      RECT 274.445 42.645 274.615 43.405 ;
      RECT 274.565 46.335 275.095 46.505 ;
      RECT 271.955 42.47 273.305 42.475 ;
      RECT 274.445 43.405 275.095 44.415 ;
      RECT 274.925 46.505 275.095 48.085 ;
      RECT 274.925 44.415 275.095 46.335 ;
      RECT 273.405 42.84 273.575 44.01 ;
      RECT 271.685 42.84 271.855 44.01 ;
      RECT 272.115 44.18 273.935 44.35 ;
      RECT 273.745 44.35 273.935 47.37 ;
      RECT 271.045 48.55 273.935 48.72 ;
      RECT 272.115 42.84 272.285 44.18 ;
      RECT 272.975 42.84 273.145 44.18 ;
      RECT 273.405 47.37 273.935 48.55 ;
      RECT 271.045 46.1 271.215 48.55 ;
      RECT 272.545 42.84 272.715 44.01 ;
      RECT 271.545 46.165 271.875 47.015 ;
      RECT 271.625 47.015 271.795 47.625 ;
      RECT 269.865 46.335 270.395 46.505 ;
      RECT 269.865 46.1 270.035 46.335 ;
      RECT 269.865 46.505 270.035 48.38 ;
      RECT 271.045 45.28 271.72 45.45 ;
      RECT 271.045 44.58 271.215 45.28 ;
      RECT 271.045 45.45 271.215 45.59 ;
      RECT 273.045 45.28 273.575 45.45 ;
      RECT 273.405 44.58 273.575 45.28 ;
      RECT 273.405 45.45 273.575 47.08 ;
      RECT 272.565 46.335 273.095 47.37 ;
      RECT 272.225 47.37 273.095 48.38 ;
      RECT 269.255 49.595 271.285 49.765 ;
      RECT 269.695 48.99 270.225 49.595 ;
      RECT 274.585 47.855 274.755 48.465 ;
      RECT 277.265 47.855 277.435 48.465 ;
      RECT 279.945 47.855 280.115 48.465 ;
      RECT 274.585 48.465 280.115 48.635 ;
      RECT 272.355 50.625 272.725 55.42 ;
      RECT 272.17 49.085 272.84 50.625 ;
      RECT 273.12 49.09 273.79 50.625 ;
      RECT 276.605 42.2 276.775 42.305 ;
      RECT 276.605 41.635 276.775 42.03 ;
      RECT 275.745 42.03 276.775 42.2 ;
      RECT 277.925 42.2 278.095 42.305 ;
      RECT 277.925 41.635 278.095 42.03 ;
      RECT 277.925 42.03 278.955 42.2 ;
      RECT 277.665 42.51 278.2 43.085 ;
      RECT 276.5 42.51 277.035 43.085 ;
      RECT 278.445 42.4 278.975 42.57 ;
      RECT 278.485 44.585 278.975 44.74 ;
      RECT 278.485 44.74 278.735 45.375 ;
      RECT 278.485 45.375 278.975 45.665 ;
      RECT 278.685 45.665 278.975 48.085 ;
      RECT 278.565 42.57 278.975 44.585 ;
      RECT 277.73 46.335 278.26 46.505 ;
      RECT 277.73 43.405 277.935 44.415 ;
      RECT 277.73 48.105 278.485 48.275 ;
      RECT 277.73 46.505 277.9 48.105 ;
      RECT 277.73 44.415 277.9 46.335 ;
      RECT 275.725 42.4 276.255 42.57 ;
      RECT 275.725 44.585 276.265 44.74 ;
      RECT 275.965 44.74 276.265 45.375 ;
      RECT 275.725 45.375 276.265 45.665 ;
      RECT 275.725 45.665 276.015 48.085 ;
      RECT 275.725 42.57 276.135 44.585 ;
      RECT 278.105 43.405 278.395 44.415 ;
      RECT 278.105 44.415 278.275 44.52 ;
      RECT 278.07 44.52 278.275 45.3 ;
      RECT 276.305 43.405 276.475 44.415 ;
      RECT 276.44 46.335 276.97 46.505 ;
      RECT 276.765 43.405 276.97 44.415 ;
      RECT 253.425 43.405 254.075 44.415 ;
      RECT 253.905 46.505 254.075 48.085 ;
      RECT 253.905 44.415 254.075 46.335 ;
      RECT 245.96 44.57 246.97 44.74 ;
      RECT 246.44 44.74 246.97 44.8 ;
      RECT 246.025 42.505 246.555 42.675 ;
      RECT 246.025 42.675 246.195 43.615 ;
      RECT 246.905 42.605 247.075 44.4 ;
      RECT 248.845 46.335 249.375 46.505 ;
      RECT 248.845 46.1 249.015 46.335 ;
      RECT 248.845 46.505 249.015 48.38 ;
      RECT 248.845 44.18 250.405 44.35 ;
      RECT 248.845 45.76 251.375 45.93 ;
      RECT 248.845 44.35 249.015 45.76 ;
      RECT 249.375 42.84 249.545 44.18 ;
      RECT 250.235 42.84 250.405 44.18 ;
      RECT 251.205 44.58 251.375 45.76 ;
      RECT 251.205 45.93 251.375 47.08 ;
      RECT 246.515 45.03 247.06 45.2 ;
      RECT 246.515 45 246.685 45.03 ;
      RECT 246.515 45.2 246.685 48 ;
      RECT 247.295 45.29 247.465 48 ;
      RECT 248.945 42.84 249.115 44.01 ;
      RECT 249.805 42.84 249.975 44.01 ;
      RECT 250.525 46.165 250.855 47.015 ;
      RECT 250.605 47.015 250.775 47.625 ;
      RECT 250.665 42.84 250.835 44.01 ;
      RECT 250.025 48.55 252.915 48.72 ;
      RECT 252.725 44.35 252.915 47.37 ;
      RECT 251.095 44.18 252.915 44.35 ;
      RECT 251.095 42.84 251.265 44.18 ;
      RECT 251.955 42.84 252.125 44.18 ;
      RECT 250.025 46.1 250.195 48.55 ;
      RECT 252.385 47.37 252.915 48.55 ;
      RECT 251.525 42.84 251.695 44.01 ;
      RECT 251.545 46.335 252.075 47.37 ;
      RECT 251.205 47.37 252.075 48.38 ;
      RECT 250.025 45.28 250.7 45.45 ;
      RECT 250.025 44.58 250.195 45.28 ;
      RECT 250.025 45.45 250.195 45.59 ;
      RECT 251.38 49.005 252.58 49.175 ;
      RECT 251.38 49.175 252.05 50.625 ;
      RECT 250.43 49.09 251.1 50.625 ;
      RECT 252.725 43.095 253.255 43.265 ;
      RECT 253.085 43.265 253.255 48.39 ;
      RECT 256.71 46.335 257.24 46.505 ;
      RECT 256.71 43.405 256.915 44.415 ;
      RECT 256.71 48.105 257.465 48.275 ;
      RECT 256.71 46.505 256.88 48.105 ;
      RECT 256.71 44.415 256.88 46.335 ;
      RECT 255.42 46.335 255.95 46.505 ;
      RECT 255.745 43.405 255.95 44.415 ;
      RECT 255.195 48.105 255.95 48.275 ;
      RECT 255.78 46.505 255.95 48.105 ;
      RECT 255.78 44.415 255.95 46.335 ;
      RECT 253.565 47.855 253.735 48.465 ;
      RECT 258.925 47.855 259.095 48.465 ;
      RECT 256.245 45.065 256.415 48.465 ;
      RECT 253.565 48.465 259.095 48.635 ;
      RECT 252.385 42.84 252.555 44.01 ;
      RECT 252.025 45.28 252.555 45.45 ;
      RECT 252.385 44.58 252.555 45.28 ;
      RECT 252.385 45.45 252.555 47.08 ;
      RECT 254.245 45 254.775 45.17 ;
      RECT 254.365 45.17 254.535 48.085 ;
      RECT 254.725 42.03 255.755 42.2 ;
      RECT 255.585 42.2 255.755 42.305 ;
      RECT 255.585 41.635 255.755 42.03 ;
      RECT 254.705 42.4 255.235 42.57 ;
      RECT 254.705 44.585 255.245 44.74 ;
      RECT 254.945 44.74 255.245 45.375 ;
      RECT 254.705 45.375 255.245 45.665 ;
      RECT 254.705 45.665 254.995 48.085 ;
      RECT 254.705 42.57 255.115 44.585 ;
      RECT 255.48 42.51 256.015 43.085 ;
      RECT 255.44 44.63 255.61 45.3 ;
      RECT 255.285 43.405 255.455 44.415 ;
      RECT 256.905 42.2 257.075 42.305 ;
      RECT 256.905 41.635 257.075 42.03 ;
      RECT 256.905 42.03 257.935 42.2 ;
      RECT 256.645 42.51 257.18 43.085 ;
      RECT 257.05 44.63 257.22 45.3 ;
      RECT 257.205 43.405 257.375 44.415 ;
      RECT 257.415 44.74 257.715 45.375 ;
      RECT 257.415 44.585 257.955 44.74 ;
      RECT 257.415 45.375 257.955 45.665 ;
      RECT 257.665 45.665 257.955 48.085 ;
      RECT 257.425 42.4 257.955 42.57 ;
      RECT 257.545 42.57 257.955 44.585 ;
      RECT 252.935 49.595 255.815 49.765 ;
      RECT 255.285 49.045 255.815 49.595 ;
      RECT 259.405 43.095 259.935 43.265 ;
      RECT 259.405 43.265 259.575 48.39 ;
      RECT 259.745 48.55 262.635 48.72 ;
      RECT 259.745 44.35 259.935 47.37 ;
      RECT 259.745 44.18 261.565 44.35 ;
      RECT 260.535 42.84 260.705 44.18 ;
      RECT 261.395 42.84 261.565 44.18 ;
      RECT 259.745 47.37 260.275 48.55 ;
      RECT 262.465 46.1 262.635 48.55 ;
      RECT 261.285 45.76 263.815 45.93 ;
      RECT 262.255 44.18 263.815 44.35 ;
      RECT 261.285 44.58 261.455 45.76 ;
      RECT 262.255 42.84 262.425 44.18 ;
      RECT 263.115 42.84 263.285 44.18 ;
      RECT 263.645 44.35 263.815 45.76 ;
      RECT 261.285 45.93 261.455 47.08 ;
      RECT 259.065 42.475 261.725 42.645 ;
      RECT 259.065 42.645 259.235 43.405 ;
      RECT 258.585 46.335 259.115 46.505 ;
      RECT 260.375 42.47 261.725 42.475 ;
      RECT 258.585 43.405 259.235 44.415 ;
      RECT 258.585 46.505 258.755 48.085 ;
      RECT 258.585 44.415 258.755 46.335 ;
      RECT 257.885 45 258.415 45.17 ;
      RECT 258.125 45.17 258.295 48.085 ;
      RECT 260.105 42.84 260.275 44.01 ;
      RECT 260.105 45.28 260.635 45.45 ;
      RECT 260.105 44.58 260.275 45.28 ;
      RECT 260.105 45.45 260.275 47.08 ;
      RECT 261.825 42.84 261.995 44.01 ;
      RECT 260.965 42.84 261.135 44.01 ;
      RECT 262.08 42.47 263.43 42.64 ;
      RECT 262.08 42.64 263.33 42.67 ;
      RECT 262.685 42.84 262.855 44.01 ;
      RECT 261.96 45.28 262.635 45.45 ;
      RECT 262.465 45.45 262.635 45.59 ;
      RECT 232.545 47.855 232.715 48.465 ;
      RECT 237.905 47.855 238.075 48.465 ;
      RECT 235.225 45.065 235.395 48.465 ;
      RECT 232.545 48.465 238.075 48.635 ;
      RECT 229.645 42.84 229.815 44.01 ;
      RECT 228.785 42.84 228.955 44.01 ;
      RECT 231.365 42.84 231.535 44.01 ;
      RECT 230.505 42.84 230.675 44.01 ;
      RECT 233.705 42.03 234.735 42.2 ;
      RECT 234.565 42.2 234.735 42.305 ;
      RECT 234.565 41.635 234.735 42.03 ;
      RECT 233.685 42.4 234.215 42.57 ;
      RECT 233.685 44.585 234.225 44.74 ;
      RECT 233.925 44.74 234.225 45.375 ;
      RECT 233.685 45.375 234.225 45.665 ;
      RECT 233.685 45.665 233.975 48.085 ;
      RECT 233.685 42.57 234.095 44.585 ;
      RECT 229.505 46.165 229.835 47.015 ;
      RECT 229.585 47.015 229.755 47.625 ;
      RECT 229.005 45.28 229.68 45.45 ;
      RECT 229.005 44.58 229.175 45.28 ;
      RECT 229.005 45.45 229.175 45.59 ;
      RECT 231.005 45.28 231.535 45.45 ;
      RECT 231.365 44.58 231.535 45.28 ;
      RECT 231.365 45.45 231.535 47.08 ;
      RECT 230.525 46.335 231.055 47.37 ;
      RECT 230.185 47.37 231.055 48.38 ;
      RECT 234.4 46.335 234.93 46.505 ;
      RECT 234.175 48.105 234.93 48.275 ;
      RECT 234.76 46.505 234.93 48.105 ;
      RECT 234.76 44.415 234.93 46.335 ;
      RECT 234.725 43.405 234.93 44.415 ;
      RECT 233.225 45 233.755 45.17 ;
      RECT 233.345 45.17 233.515 48.085 ;
      RECT 238.725 48.55 241.615 48.72 ;
      RECT 238.725 44.35 238.915 47.37 ;
      RECT 238.725 44.18 240.545 44.35 ;
      RECT 239.515 42.84 239.685 44.18 ;
      RECT 240.375 42.84 240.545 44.18 ;
      RECT 238.725 47.37 239.255 48.55 ;
      RECT 241.445 46.1 241.615 48.55 ;
      RECT 235.885 42.2 236.055 42.305 ;
      RECT 235.885 41.635 236.055 42.03 ;
      RECT 235.885 42.03 236.915 42.2 ;
      RECT 236.405 42.4 236.935 42.57 ;
      RECT 236.395 44.585 236.935 44.74 ;
      RECT 236.395 44.74 236.695 45.375 ;
      RECT 236.395 45.375 236.935 45.665 ;
      RECT 236.645 45.665 236.935 48.085 ;
      RECT 236.525 42.57 236.935 44.585 ;
      RECT 238.045 42.475 240.705 42.645 ;
      RECT 238.045 42.645 238.215 43.405 ;
      RECT 237.565 46.335 238.095 46.505 ;
      RECT 239.355 42.47 240.705 42.475 ;
      RECT 237.565 43.405 238.215 44.415 ;
      RECT 237.565 46.505 237.735 48.085 ;
      RECT 237.565 44.415 237.735 46.335 ;
      RECT 235.625 42.51 236.16 43.085 ;
      RECT 234.46 42.51 234.995 43.085 ;
      RECT 235.69 46.335 236.22 46.505 ;
      RECT 235.69 48.105 236.445 48.275 ;
      RECT 235.69 46.505 235.86 48.105 ;
      RECT 235.69 44.415 235.86 46.335 ;
      RECT 235.69 43.405 235.895 44.415 ;
      RECT 234.42 44.63 234.59 45.3 ;
      RECT 234.265 43.405 234.435 44.415 ;
      RECT 236.03 44.63 236.2 45.3 ;
      RECT 238.385 43.095 238.915 43.265 ;
      RECT 238.385 43.265 238.555 48.39 ;
      RECT 236.865 45 237.395 45.17 ;
      RECT 237.105 45.17 237.275 48.085 ;
      RECT 236.185 43.405 236.355 44.415 ;
      RECT 239.085 42.84 239.255 44.01 ;
      RECT 239.085 45.28 239.615 45.45 ;
      RECT 239.085 44.58 239.255 45.28 ;
      RECT 239.085 45.45 239.255 47.08 ;
      RECT 239.945 42.84 240.115 44.01 ;
      RECT 239.565 46.335 240.095 47.37 ;
      RECT 239.565 47.37 240.435 48.38 ;
      RECT 242.87 41.76 243.4 41.93 ;
      RECT 243.09 41.93 243.4 43.11 ;
      RECT 242.985 43.11 243.515 48.39 ;
      RECT 241.06 42.47 242.41 42.64 ;
      RECT 241.06 42.64 242.31 42.67 ;
      RECT 240.805 42.84 240.975 44.01 ;
      RECT 242.525 42.84 242.695 44.01 ;
      RECT 241.665 42.84 241.835 44.01 ;
      RECT 241.235 44.18 242.795 44.35 ;
      RECT 240.265 45.76 242.795 45.93 ;
      RECT 242.095 42.84 242.265 44.18 ;
      RECT 241.235 42.84 241.405 44.18 ;
      RECT 240.265 44.58 240.435 45.76 ;
      RECT 242.625 44.35 242.795 45.76 ;
      RECT 240.265 45.93 240.435 47.08 ;
      RECT 244.565 42.605 244.735 44.4 ;
      RECT 244.785 42 245.455 42.17 ;
      RECT 244.855 42.17 245.385 42.3 ;
      RECT 245.085 42.505 245.615 42.675 ;
      RECT 245.445 42.675 245.615 43.615 ;
      RECT 240.785 46.165 241.115 47.015 ;
      RECT 240.865 47.015 241.035 47.625 ;
      RECT 242.265 46.335 242.795 46.505 ;
      RECT 242.625 46.1 242.795 46.335 ;
      RECT 242.625 46.505 242.795 48.38 ;
      RECT 240.94 45.28 241.615 45.45 ;
      RECT 241.445 44.58 241.615 45.28 ;
      RECT 241.445 45.45 241.615 45.59 ;
      RECT 244.67 44.57 245.68 44.74 ;
      RECT 244.67 44.74 245.2 44.8 ;
      RECT 245.735 45.29 245.905 48 ;
      RECT 244.58 45.03 245.125 45.2 ;
      RECT 244.955 45 245.125 45.03 ;
      RECT 244.955 45.2 245.125 48 ;
      RECT 244.175 45.29 244.345 48 ;
      RECT 244.295 48.215 247.345 48.35 ;
      RECT 244.135 48.35 247.505 48.52 ;
      RECT 248.24 41.76 248.77 41.93 ;
      RECT 248.24 41.93 248.55 43.11 ;
      RECT 248.125 43.11 248.655 48.39 ;
      RECT 246.185 42 246.855 42.17 ;
      RECT 246.255 42.17 246.785 42.3 ;
      RECT 249.23 42.47 250.58 42.64 ;
      RECT 249.33 42.64 250.58 42.67 ;
      RECT 250.935 42.475 253.595 42.645 ;
      RECT 253.425 42.645 253.595 43.405 ;
      RECT 253.545 46.335 254.075 46.505 ;
      RECT 250.935 42.47 252.285 42.475 ;
      RECT 214.865 41.635 215.035 42.03 ;
      RECT 214.865 42.03 215.895 42.2 ;
      RECT 214.605 42.51 215.14 43.085 ;
      RECT 215.01 44.63 215.18 45.3 ;
      RECT 214.67 46.335 215.2 46.505 ;
      RECT 214.67 48.105 215.425 48.275 ;
      RECT 214.67 46.505 214.84 48.105 ;
      RECT 214.67 44.415 214.84 46.335 ;
      RECT 214.67 43.405 214.875 44.415 ;
      RECT 216.545 46.335 217.075 46.505 ;
      RECT 217.025 42.645 217.195 43.405 ;
      RECT 217.025 42.475 219.685 42.645 ;
      RECT 216.545 46.505 216.715 48.085 ;
      RECT 216.545 43.405 217.195 44.415 ;
      RECT 218.335 42.47 219.685 42.475 ;
      RECT 216.545 44.415 216.715 46.335 ;
      RECT 215.625 45.665 215.915 48.085 ;
      RECT 215.375 45.375 215.915 45.665 ;
      RECT 215.375 44.74 215.675 45.375 ;
      RECT 215.375 44.585 215.915 44.74 ;
      RECT 215.385 42.4 215.915 42.57 ;
      RECT 215.505 42.57 215.915 44.585 ;
      RECT 214.205 45.065 214.375 48.465 ;
      RECT 214.205 48.635 214.66 48.655 ;
      RECT 215.585 48.635 216.755 48.655 ;
      RECT 214.205 48.465 217.055 48.635 ;
      RECT 216.885 47.855 217.055 48.465 ;
      RECT 215.845 45 216.375 45.17 ;
      RECT 216.085 45.17 216.255 48.085 ;
      RECT 215.165 43.405 215.335 44.415 ;
      RECT 217.365 43.095 217.895 43.265 ;
      RECT 217.365 43.265 217.535 48.39 ;
      RECT 217.705 48.55 220.595 48.72 ;
      RECT 217.705 44.35 217.895 47.37 ;
      RECT 217.705 44.18 219.525 44.35 ;
      RECT 218.495 42.84 218.665 44.18 ;
      RECT 219.355 42.84 219.525 44.18 ;
      RECT 217.705 47.37 218.235 48.55 ;
      RECT 220.425 46.1 220.595 48.55 ;
      RECT 219.245 45.76 221.775 45.93 ;
      RECT 220.215 44.18 221.775 44.35 ;
      RECT 219.245 44.58 219.415 45.76 ;
      RECT 220.215 42.84 220.385 44.18 ;
      RECT 221.075 42.84 221.245 44.18 ;
      RECT 221.605 44.35 221.775 45.76 ;
      RECT 219.245 45.93 219.415 47.08 ;
      RECT 221.965 43.11 222.495 43.28 ;
      RECT 221.85 41.76 222.38 41.93 ;
      RECT 222.07 41.93 222.38 43.11 ;
      RECT 222.185 43.28 222.355 48.39 ;
      RECT 218.065 42.84 218.235 44.01 ;
      RECT 218.065 45.28 218.595 45.45 ;
      RECT 218.065 44.58 218.235 45.28 ;
      RECT 218.065 45.45 218.235 47.08 ;
      RECT 218.925 42.84 219.095 44.01 ;
      RECT 220.04 42.47 221.39 42.64 ;
      RECT 220.04 42.64 221.29 42.67 ;
      RECT 219.785 42.84 219.955 44.01 ;
      RECT 220.645 42.84 220.815 44.01 ;
      RECT 219.92 45.28 220.595 45.45 ;
      RECT 220.425 45.45 220.595 45.59 ;
      RECT 220.425 44.58 220.595 45.28 ;
      RECT 221.505 42.84 221.675 44.01 ;
      RECT 218.545 46.335 219.075 47.37 ;
      RECT 218.545 47.37 219.415 48.38 ;
      RECT 219.765 46.165 220.095 47.015 ;
      RECT 219.845 47.015 220.015 47.625 ;
      RECT 221.245 46.335 221.775 46.505 ;
      RECT 221.605 46.1 221.775 46.335 ;
      RECT 221.605 46.505 221.775 48.38 ;
      RECT 227.825 45.76 230.355 45.93 ;
      RECT 227.825 44.18 229.385 44.35 ;
      RECT 230.185 44.58 230.355 45.76 ;
      RECT 228.355 42.84 228.525 44.18 ;
      RECT 229.215 42.84 229.385 44.18 ;
      RECT 227.825 44.35 227.995 45.76 ;
      RECT 230.185 45.93 230.355 47.08 ;
      RECT 227.22 41.76 227.75 41.93 ;
      RECT 227.22 41.93 227.53 43.11 ;
      RECT 227.105 43.11 227.635 48.39 ;
      RECT 223.545 42.605 223.715 44.4 ;
      RECT 223.765 42 224.435 42.17 ;
      RECT 223.835 42.17 224.365 42.3 ;
      RECT 224.065 42.505 224.595 42.675 ;
      RECT 224.425 42.675 224.595 43.615 ;
      RECT 225.885 42.605 226.055 44.4 ;
      RECT 225.165 42 225.835 42.17 ;
      RECT 225.235 42.17 225.765 42.3 ;
      RECT 225.005 42.505 225.535 42.675 ;
      RECT 225.005 42.675 225.175 43.615 ;
      RECT 228.21 42.47 229.56 42.64 ;
      RECT 228.31 42.64 229.56 42.67 ;
      RECT 227.925 42.84 228.095 44.01 ;
      RECT 223.65 44.57 224.66 44.74 ;
      RECT 223.65 44.74 224.18 44.8 ;
      RECT 223.56 45.03 224.105 45.2 ;
      RECT 223.935 45 224.105 45.03 ;
      RECT 223.935 45.2 224.105 48 ;
      RECT 223.155 45.29 223.325 48 ;
      RECT 223.275 48.215 226.325 48.35 ;
      RECT 223.115 48.35 226.485 48.52 ;
      RECT 224.94 44.57 225.95 44.74 ;
      RECT 225.42 44.74 225.95 44.8 ;
      RECT 224.715 45.29 224.885 48 ;
      RECT 225.495 45.03 226.04 45.2 ;
      RECT 225.495 45 225.665 45.03 ;
      RECT 225.495 45.2 225.665 48 ;
      RECT 226.275 45.29 226.445 48 ;
      RECT 227.825 46.335 228.355 46.505 ;
      RECT 227.825 46.1 227.995 46.335 ;
      RECT 227.825 46.505 227.995 48.38 ;
      RECT 231.705 43.095 232.235 43.265 ;
      RECT 232.065 43.265 232.235 48.39 ;
      RECT 229.005 48.55 231.895 48.72 ;
      RECT 231.705 44.35 231.895 47.37 ;
      RECT 230.075 44.18 231.895 44.35 ;
      RECT 230.075 42.84 230.245 44.18 ;
      RECT 230.935 42.84 231.105 44.18 ;
      RECT 229.005 46.1 229.175 48.55 ;
      RECT 231.365 47.37 231.895 48.55 ;
      RECT 229.915 42.475 232.575 42.645 ;
      RECT 232.405 42.645 232.575 43.405 ;
      RECT 232.525 46.335 233.055 46.505 ;
      RECT 229.915 42.47 231.265 42.475 ;
      RECT 232.405 43.405 233.055 44.415 ;
      RECT 232.885 46.505 233.055 48.085 ;
      RECT 232.885 44.415 233.055 46.335 ;
      RECT 158.47 42.84 158.64 44.01 ;
      RECT 158.47 45.28 159 45.45 ;
      RECT 158.47 44.58 158.64 45.28 ;
      RECT 158.47 45.45 158.64 47.08 ;
      RECT 158.95 46.335 159.48 47.37 ;
      RECT 158.95 47.37 159.82 48.38 ;
      RECT 163.68 48.215 166.73 48.35 ;
      RECT 163.52 48.35 166.89 48.52 ;
      RECT 159.65 45.76 162.18 45.93 ;
      RECT 160.62 44.18 162.18 44.35 ;
      RECT 159.65 44.58 159.82 45.76 ;
      RECT 160.62 42.84 160.79 44.18 ;
      RECT 161.48 42.84 161.65 44.18 ;
      RECT 162.01 44.35 162.18 45.76 ;
      RECT 159.65 45.93 159.82 47.08 ;
      RECT 162.255 41.76 162.785 41.93 ;
      RECT 162.475 41.93 162.785 43.11 ;
      RECT 162.37 43.11 162.9 48.39 ;
      RECT 160.445 42.47 161.795 42.64 ;
      RECT 160.445 42.64 161.695 42.67 ;
      RECT 160.19 42.84 160.36 44.01 ;
      RECT 159.33 42.84 159.5 44.01 ;
      RECT 161.91 42.84 162.08 44.01 ;
      RECT 161.05 42.84 161.22 44.01 ;
      RECT 163.95 42.605 164.12 44.4 ;
      RECT 164.17 42 164.84 42.17 ;
      RECT 164.24 42.17 164.77 42.3 ;
      RECT 164.47 42.505 165 42.675 ;
      RECT 164.83 42.675 165 43.615 ;
      RECT 160.17 46.165 160.5 47.015 ;
      RECT 160.25 47.015 160.42 47.625 ;
      RECT 160.325 45.28 161 45.45 ;
      RECT 160.83 44.58 161 45.28 ;
      RECT 160.83 45.45 161 45.59 ;
      RECT 161.65 46.335 162.18 46.505 ;
      RECT 162.01 46.1 162.18 46.335 ;
      RECT 162.01 46.505 162.18 48.38 ;
      RECT 163.56 45.29 163.73 48 ;
      RECT 164.055 44.57 165.065 44.74 ;
      RECT 164.055 44.74 164.585 44.8 ;
      RECT 163.965 45.03 164.51 45.2 ;
      RECT 164.34 45 164.51 45.03 ;
      RECT 164.34 45.2 164.51 48 ;
      RECT 167.51 43.11 168.04 43.28 ;
      RECT 167.625 41.76 168.155 41.93 ;
      RECT 167.625 41.93 167.935 43.11 ;
      RECT 167.65 43.28 167.82 48.39 ;
      RECT 168.615 42.47 169.965 42.64 ;
      RECT 168.715 42.64 169.965 42.67 ;
      RECT 165.345 44.57 166.355 44.74 ;
      RECT 165.825 44.74 166.355 44.8 ;
      RECT 166.29 42.605 166.46 44.4 ;
      RECT 168.23 44.18 169.79 44.35 ;
      RECT 168.23 45.76 170.76 45.93 ;
      RECT 168.23 44.35 168.4 45.76 ;
      RECT 168.76 42.84 168.93 44.18 ;
      RECT 169.62 42.84 169.79 44.18 ;
      RECT 170.59 44.58 170.76 45.76 ;
      RECT 170.59 45.93 170.76 47.08 ;
      RECT 165.57 42 166.24 42.17 ;
      RECT 165.64 42.17 166.17 42.3 ;
      RECT 168.33 42.84 168.5 44.01 ;
      RECT 165.41 42.505 165.94 42.675 ;
      RECT 165.41 42.675 165.58 43.615 ;
      RECT 170.32 42.475 172.98 42.645 ;
      RECT 172.81 42.645 172.98 43.405 ;
      RECT 172.93 46.335 173.46 46.505 ;
      RECT 170.32 42.47 171.67 42.475 ;
      RECT 172.81 43.405 173.46 44.415 ;
      RECT 173.29 46.505 173.46 48.085 ;
      RECT 173.29 44.415 173.46 46.335 ;
      RECT 170.05 42.84 170.22 44.01 ;
      RECT 169.19 42.84 169.36 44.01 ;
      RECT 170.48 44.18 172.3 44.35 ;
      RECT 172.11 44.35 172.3 47.37 ;
      RECT 169.41 48.55 172.3 48.72 ;
      RECT 170.48 42.84 170.65 44.18 ;
      RECT 171.34 42.84 171.51 44.18 ;
      RECT 171.77 47.37 172.3 48.55 ;
      RECT 169.41 46.1 169.58 48.55 ;
      RECT 169.41 45.28 170.085 45.45 ;
      RECT 169.41 45.45 169.58 45.59 ;
      RECT 169.41 44.58 169.58 45.28 ;
      RECT 168.23 46.335 168.76 46.505 ;
      RECT 168.23 46.1 168.4 46.335 ;
      RECT 168.23 46.505 168.4 48.38 ;
      RECT 165.12 45.29 165.29 48 ;
      RECT 165.9 45.03 166.445 45.2 ;
      RECT 165.9 45 166.07 45.03 ;
      RECT 165.9 45.2 166.07 48 ;
      RECT 166.68 45.29 166.85 48 ;
      RECT 169.91 46.165 170.24 47.015 ;
      RECT 169.99 47.015 170.16 47.625 ;
      RECT 174.97 42.2 175.14 42.305 ;
      RECT 174.97 41.635 175.14 42.03 ;
      RECT 174.11 42.03 175.14 42.2 ;
      RECT 171.77 42.84 171.94 44.01 ;
      RECT 171.41 45.28 171.94 45.45 ;
      RECT 171.77 44.58 171.94 45.28 ;
      RECT 171.77 45.45 171.94 47.08 ;
      RECT 170.91 42.84 171.08 44.01 ;
      RECT 172.95 47.855 173.12 48.465 ;
      RECT 173.25 48.635 174.42 48.655 ;
      RECT 175.345 48.635 175.8 48.655 ;
      RECT 175.63 45.065 175.8 48.465 ;
      RECT 172.95 48.465 175.8 48.635 ;
      RECT 170.93 46.335 171.46 47.37 ;
      RECT 170.59 47.37 171.46 48.38 ;
      RECT 172.11 43.095 172.64 43.265 ;
      RECT 172.47 43.265 172.64 48.39 ;
      RECT 174.865 42.51 175.4 43.085 ;
      RECT 174.805 46.335 175.335 46.505 ;
      RECT 174.58 48.105 175.335 48.275 ;
      RECT 175.165 46.505 175.335 48.105 ;
      RECT 175.165 44.415 175.335 46.335 ;
      RECT 175.13 43.405 175.335 44.415 ;
      RECT 174.825 44.63 174.995 45.3 ;
      RECT 174.09 45.665 174.38 48.085 ;
      RECT 174.09 45.375 174.63 45.665 ;
      RECT 174.33 44.74 174.63 45.375 ;
      RECT 174.09 44.585 174.63 44.74 ;
      RECT 174.09 42.4 174.62 42.57 ;
      RECT 174.09 42.57 174.5 44.585 ;
      RECT 173.63 45 174.16 45.17 ;
      RECT 173.75 45.17 173.92 48.085 ;
      RECT 174.67 43.405 174.84 44.415 ;
      RECT 214.865 42.2 215.035 42.305 ;
      RECT 144.55 42 145.22 42.17 ;
      RECT 144.62 42.17 145.15 42.3 ;
      RECT 146.605 41.76 147.135 41.93 ;
      RECT 146.605 41.93 146.915 43.11 ;
      RECT 146.49 43.11 147.02 48.39 ;
      RECT 143.035 44.57 144.045 44.74 ;
      RECT 143.035 44.74 143.565 44.8 ;
      RECT 142.93 42.605 143.1 44.4 ;
      RECT 144.1 45.29 144.27 48 ;
      RECT 142.945 45.03 143.49 45.2 ;
      RECT 143.32 45 143.49 45.03 ;
      RECT 143.32 45.2 143.49 48 ;
      RECT 142.54 45.29 142.71 48 ;
      RECT 143.45 42.505 143.98 42.675 ;
      RECT 143.81 42.675 143.98 43.615 ;
      RECT 142.66 48.215 145.71 48.35 ;
      RECT 142.5 48.35 145.87 48.52 ;
      RECT 144.325 44.57 145.335 44.74 ;
      RECT 144.805 44.74 145.335 44.8 ;
      RECT 145.27 42.605 145.44 44.4 ;
      RECT 144.88 45.03 145.425 45.2 ;
      RECT 144.88 45 145.05 45.03 ;
      RECT 144.88 45.2 145.05 48 ;
      RECT 145.66 45.29 145.83 48 ;
      RECT 144.39 42.505 144.92 42.675 ;
      RECT 144.39 42.675 144.56 43.615 ;
      RECT 147.21 46.335 147.74 46.505 ;
      RECT 147.21 46.1 147.38 46.335 ;
      RECT 147.21 46.505 147.38 48.38 ;
      RECT 147.21 45.76 149.74 45.93 ;
      RECT 147.21 44.18 148.77 44.35 ;
      RECT 147.21 44.35 147.38 45.76 ;
      RECT 147.74 42.84 147.91 44.18 ;
      RECT 148.6 42.84 148.77 44.18 ;
      RECT 149.57 44.58 149.74 45.76 ;
      RECT 149.57 45.93 149.74 47.08 ;
      RECT 147.31 42.84 147.48 44.01 ;
      RECT 151.09 43.095 151.62 43.265 ;
      RECT 151.45 43.265 151.62 48.39 ;
      RECT 148.39 48.55 151.28 48.72 ;
      RECT 151.09 44.35 151.28 47.37 ;
      RECT 149.46 44.18 151.28 44.35 ;
      RECT 149.46 42.84 149.63 44.18 ;
      RECT 150.32 42.84 150.49 44.18 ;
      RECT 148.39 46.1 148.56 48.55 ;
      RECT 150.75 47.37 151.28 48.55 ;
      RECT 149.3 42.475 151.96 42.645 ;
      RECT 151.79 42.645 151.96 43.405 ;
      RECT 151.91 46.335 152.44 46.505 ;
      RECT 149.3 42.47 150.65 42.475 ;
      RECT 151.79 43.405 152.44 44.415 ;
      RECT 152.27 46.505 152.44 48.085 ;
      RECT 152.27 44.415 152.44 46.335 ;
      RECT 147.595 42.47 148.945 42.64 ;
      RECT 147.695 42.64 148.945 42.67 ;
      RECT 148.17 42.84 148.34 44.01 ;
      RECT 149.03 42.84 149.2 44.01 ;
      RECT 149.89 42.84 150.06 44.01 ;
      RECT 150.75 42.84 150.92 44.01 ;
      RECT 153.09 42.03 154.12 42.2 ;
      RECT 153.95 42.2 154.12 42.305 ;
      RECT 153.95 41.635 154.12 42.03 ;
      RECT 153.07 42.4 153.6 42.57 ;
      RECT 153.07 44.585 153.61 44.74 ;
      RECT 153.31 44.74 153.61 45.375 ;
      RECT 153.07 45.375 153.61 45.665 ;
      RECT 153.07 45.665 153.36 48.085 ;
      RECT 153.07 42.57 153.48 44.585 ;
      RECT 148.39 45.28 149.065 45.45 ;
      RECT 148.39 44.58 148.56 45.28 ;
      RECT 148.39 45.45 148.56 45.59 ;
      RECT 148.89 46.165 149.22 47.015 ;
      RECT 148.97 47.015 149.14 47.625 ;
      RECT 149.91 46.335 150.44 47.37 ;
      RECT 149.57 47.37 150.44 48.38 ;
      RECT 150.39 45.28 150.92 45.45 ;
      RECT 150.75 44.58 150.92 45.28 ;
      RECT 150.75 45.45 150.92 47.08 ;
      RECT 151.93 47.855 152.1 48.465 ;
      RECT 157.29 47.855 157.46 48.465 ;
      RECT 151.93 48.465 157.46 48.635 ;
      RECT 154.61 45.065 154.78 48.465 ;
      RECT 152.61 45 153.14 45.17 ;
      RECT 152.73 45.17 152.9 48.085 ;
      RECT 158.11 48.55 161 48.72 ;
      RECT 158.11 44.35 158.3 47.37 ;
      RECT 158.11 44.18 159.93 44.35 ;
      RECT 158.9 42.84 159.07 44.18 ;
      RECT 159.76 42.84 159.93 44.18 ;
      RECT 158.11 47.37 158.64 48.55 ;
      RECT 160.83 46.1 161 48.55 ;
      RECT 155.27 42.2 155.44 42.305 ;
      RECT 155.27 41.635 155.44 42.03 ;
      RECT 155.27 42.03 156.3 42.2 ;
      RECT 155.79 42.4 156.32 42.57 ;
      RECT 155.78 44.585 156.32 44.74 ;
      RECT 155.78 44.74 156.08 45.375 ;
      RECT 155.78 45.375 156.32 45.665 ;
      RECT 156.03 45.665 156.32 48.085 ;
      RECT 155.91 42.57 156.32 44.585 ;
      RECT 153.845 42.51 154.38 43.085 ;
      RECT 155.01 42.51 155.545 43.085 ;
      RECT 153.785 46.335 154.315 46.505 ;
      RECT 153.56 48.105 154.315 48.275 ;
      RECT 154.145 46.505 154.315 48.105 ;
      RECT 154.145 44.415 154.315 46.335 ;
      RECT 154.11 43.405 154.315 44.415 ;
      RECT 153.805 44.63 153.975 45.3 ;
      RECT 155.075 46.335 155.605 46.505 ;
      RECT 155.075 48.105 155.83 48.275 ;
      RECT 155.075 46.505 155.245 48.105 ;
      RECT 155.075 44.415 155.245 46.335 ;
      RECT 155.075 43.405 155.28 44.415 ;
      RECT 153.65 43.405 153.82 44.415 ;
      RECT 155.415 44.63 155.585 45.3 ;
      RECT 156.95 46.335 157.48 46.505 ;
      RECT 157.43 42.645 157.6 43.405 ;
      RECT 157.43 42.475 160.09 42.645 ;
      RECT 156.95 46.505 157.12 48.085 ;
      RECT 156.95 43.405 157.6 44.415 ;
      RECT 158.74 42.47 160.09 42.475 ;
      RECT 156.95 44.415 157.12 46.335 ;
      RECT 156.25 45 156.78 45.17 ;
      RECT 156.49 45.17 156.66 48.085 ;
      RECT 157.77 43.095 158.3 43.265 ;
      RECT 157.77 43.265 157.94 48.39 ;
      RECT 155.57 43.405 155.74 44.415 ;
      RECT 128.28 42.475 130.94 42.645 ;
      RECT 130.77 42.645 130.94 43.405 ;
      RECT 130.89 46.335 131.42 46.505 ;
      RECT 128.28 42.47 129.63 42.475 ;
      RECT 130.77 43.405 131.42 44.415 ;
      RECT 131.25 46.505 131.42 48.085 ;
      RECT 131.25 44.415 131.42 46.335 ;
      RECT 124.25 42.605 124.42 44.4 ;
      RECT 126.575 42.47 127.925 42.64 ;
      RECT 126.675 42.64 127.925 42.67 ;
      RECT 126.29 42.84 126.46 44.01 ;
      RECT 127.15 42.84 127.32 44.01 ;
      RECT 127.37 45.28 128.045 45.45 ;
      RECT 127.37 45.45 127.54 45.59 ;
      RECT 127.37 44.58 127.54 45.28 ;
      RECT 128.01 42.84 128.18 44.01 ;
      RECT 128.87 42.84 129.04 44.01 ;
      RECT 129.73 42.84 129.9 44.01 ;
      RECT 129.37 45.28 129.9 45.45 ;
      RECT 129.73 44.58 129.9 45.28 ;
      RECT 129.73 45.45 129.9 47.08 ;
      RECT 124.64 45.29 124.81 48 ;
      RECT 126.19 46.335 126.72 46.505 ;
      RECT 126.19 46.1 126.36 46.335 ;
      RECT 126.19 46.505 126.36 48.38 ;
      RECT 127.87 46.165 128.2 47.015 ;
      RECT 127.95 47.015 128.12 47.625 ;
      RECT 128.89 46.335 129.42 47.37 ;
      RECT 128.55 47.37 129.42 48.38 ;
      RECT 130.91 47.855 131.08 48.465 ;
      RECT 136.27 47.855 136.44 48.465 ;
      RECT 133.59 45.065 133.76 48.465 ;
      RECT 130.91 48.465 136.44 48.635 ;
      RECT 130.07 43.095 130.6 43.265 ;
      RECT 130.43 43.265 130.6 48.39 ;
      RECT 132.07 42.03 133.1 42.2 ;
      RECT 132.93 42.2 133.1 42.305 ;
      RECT 132.93 41.635 133.1 42.03 ;
      RECT 132.05 42.4 132.58 42.57 ;
      RECT 132.05 44.585 132.59 44.74 ;
      RECT 132.29 44.74 132.59 45.375 ;
      RECT 132.05 45.375 132.59 45.665 ;
      RECT 132.05 45.665 132.34 48.085 ;
      RECT 132.05 42.57 132.46 44.585 ;
      RECT 132.825 42.51 133.36 43.085 ;
      RECT 133.99 42.51 134.525 43.085 ;
      RECT 132.63 43.405 132.8 44.415 ;
      RECT 132.765 46.335 133.295 46.505 ;
      RECT 133.09 43.405 133.295 44.415 ;
      RECT 132.54 48.105 133.295 48.275 ;
      RECT 133.125 46.505 133.295 48.105 ;
      RECT 133.125 44.415 133.295 46.335 ;
      RECT 134.055 46.335 134.585 46.505 ;
      RECT 134.055 43.405 134.26 44.415 ;
      RECT 134.055 48.105 134.81 48.275 ;
      RECT 134.055 46.505 134.225 48.105 ;
      RECT 134.055 44.415 134.225 46.335 ;
      RECT 134.25 42.2 134.42 42.305 ;
      RECT 134.25 41.635 134.42 42.03 ;
      RECT 134.25 42.03 135.28 42.2 ;
      RECT 134.77 42.4 135.3 42.57 ;
      RECT 134.76 44.585 135.3 44.74 ;
      RECT 134.76 44.74 135.06 45.375 ;
      RECT 134.76 45.375 135.3 45.665 ;
      RECT 135.01 45.665 135.3 48.085 ;
      RECT 134.89 42.57 135.3 44.585 ;
      RECT 134.55 43.405 134.72 44.415 ;
      RECT 131.71 49.045 132.38 49.765 ;
      RECT 131.59 45 132.12 45.17 ;
      RECT 131.71 45.17 131.88 48.085 ;
      RECT 132.785 44.63 132.955 45.3 ;
      RECT 134.19 49.595 137.07 49.765 ;
      RECT 134.19 49.045 134.72 49.595 ;
      RECT 134.395 44.63 134.565 45.3 ;
      RECT 135.23 45 135.76 45.17 ;
      RECT 135.47 45.17 135.64 48.085 ;
      RECT 136.75 43.095 137.28 43.265 ;
      RECT 136.75 43.265 136.92 48.39 ;
      RECT 141.235 41.76 141.765 41.93 ;
      RECT 141.455 41.93 141.765 43.11 ;
      RECT 141.35 43.11 141.88 48.39 ;
      RECT 135.93 46.335 136.46 46.505 ;
      RECT 136.41 42.645 136.58 43.405 ;
      RECT 136.41 42.475 139.07 42.645 ;
      RECT 135.93 43.405 136.58 44.415 ;
      RECT 135.93 46.505 136.1 48.085 ;
      RECT 137.72 42.47 139.07 42.475 ;
      RECT 135.93 44.415 136.1 46.335 ;
      RECT 137.45 42.84 137.62 44.01 ;
      RECT 137.45 45.28 137.98 45.45 ;
      RECT 137.45 44.58 137.62 45.28 ;
      RECT 137.45 45.45 137.62 47.08 ;
      RECT 138.31 42.84 138.48 44.01 ;
      RECT 137.09 44.18 138.91 44.35 ;
      RECT 137.09 44.35 137.28 47.37 ;
      RECT 137.09 48.55 139.98 48.72 ;
      RECT 137.88 42.84 138.05 44.18 ;
      RECT 138.74 42.84 138.91 44.18 ;
      RECT 137.09 47.37 137.62 48.55 ;
      RECT 139.81 46.1 139.98 48.55 ;
      RECT 139.425 42.47 140.775 42.64 ;
      RECT 139.425 42.64 140.675 42.67 ;
      RECT 139.15 46.165 139.48 47.015 ;
      RECT 139.23 47.015 139.4 47.625 ;
      RECT 139.17 42.84 139.34 44.01 ;
      RECT 140.63 46.335 141.16 46.505 ;
      RECT 140.99 46.1 141.16 46.335 ;
      RECT 140.99 46.505 141.16 48.38 ;
      RECT 138.63 45.76 141.16 45.93 ;
      RECT 139.6 44.18 141.16 44.35 ;
      RECT 138.63 44.58 138.8 45.76 ;
      RECT 139.6 42.84 139.77 44.18 ;
      RECT 140.46 42.84 140.63 44.18 ;
      RECT 140.99 44.35 141.16 45.76 ;
      RECT 138.63 45.93 138.8 47.08 ;
      RECT 140.89 42.84 141.06 44.01 ;
      RECT 140.03 42.84 140.2 44.01 ;
      RECT 139.305 45.28 139.98 45.45 ;
      RECT 139.81 44.58 139.98 45.28 ;
      RECT 139.81 45.45 139.98 45.59 ;
      RECT 137.425 49.005 138.625 49.175 ;
      RECT 137.955 49.175 138.625 50.625 ;
      RECT 137.93 46.335 138.46 47.37 ;
      RECT 137.93 47.37 138.8 48.38 ;
      RECT 138.905 49.09 139.575 50.625 ;
      RECT 143.15 42 143.82 42.17 ;
      RECT 143.22 42.17 143.75 42.3 ;
      RECT 111.03 45.375 111.52 45.665 ;
      RECT 111.03 45.665 111.32 48.085 ;
      RECT 111.03 42.4 111.56 42.57 ;
      RECT 111.03 42.57 111.44 44.585 ;
      RECT 106.85 46.165 107.18 47.015 ;
      RECT 106.93 47.015 107.1 47.625 ;
      RECT 107.53 47.37 108.4 48.38 ;
      RECT 107.87 46.335 108.4 47.37 ;
      RECT 109.89 47.855 110.06 48.465 ;
      RECT 112.57 47.855 112.74 48.465 ;
      RECT 115.25 47.855 115.42 48.465 ;
      RECT 109.89 48.465 115.42 48.635 ;
      RECT 110.57 45 111.1 45.17 ;
      RECT 110.69 45.17 110.86 48.085 ;
      RECT 115.73 43.095 116.26 43.265 ;
      RECT 115.1 49.785 115.955 49.955 ;
      RECT 115.425 49.015 115.955 49.785 ;
      RECT 115.73 43.265 115.9 49.015 ;
      RECT 113.035 46.335 113.565 46.505 ;
      RECT 113.035 43.405 113.24 44.415 ;
      RECT 113.035 48.105 113.79 48.275 ;
      RECT 113.035 46.505 113.205 48.105 ;
      RECT 113.035 44.415 113.205 46.335 ;
      RECT 113.23 42.2 113.4 42.305 ;
      RECT 113.23 41.635 113.4 42.03 ;
      RECT 113.23 42.03 114.26 42.2 ;
      RECT 112.97 42.51 113.505 43.085 ;
      RECT 116.43 42.84 116.6 44.01 ;
      RECT 116.43 45.28 116.96 45.45 ;
      RECT 116.43 44.58 116.6 45.28 ;
      RECT 116.43 45.45 116.6 47.08 ;
      RECT 113.375 44.63 113.545 45.3 ;
      RECT 114.91 46.335 115.44 46.505 ;
      RECT 115.39 42.645 115.56 43.405 ;
      RECT 115.39 42.475 118.05 42.645 ;
      RECT 114.91 46.505 115.08 48.085 ;
      RECT 114.91 43.405 115.56 44.415 ;
      RECT 116.7 42.47 118.05 42.475 ;
      RECT 114.91 44.415 115.08 46.335 ;
      RECT 113.99 45.665 114.28 48.085 ;
      RECT 113.74 45.375 114.28 45.665 ;
      RECT 113.74 44.74 114.04 45.375 ;
      RECT 113.74 44.585 114.28 44.74 ;
      RECT 113.75 42.4 114.28 42.57 ;
      RECT 113.87 42.57 114.28 44.585 ;
      RECT 114.21 45 114.74 45.17 ;
      RECT 114.45 45.17 114.62 48.085 ;
      RECT 113.53 43.405 113.7 44.415 ;
      RECT 116.07 44.35 116.26 47.37 ;
      RECT 116.07 44.18 117.89 44.35 ;
      RECT 116.07 48.55 118.96 48.72 ;
      RECT 116.86 42.84 117.03 44.18 ;
      RECT 117.72 42.84 117.89 44.18 ;
      RECT 116.07 47.37 116.6 48.55 ;
      RECT 118.79 46.1 118.96 48.55 ;
      RECT 118.405 42.47 119.755 42.64 ;
      RECT 118.405 42.64 119.655 42.67 ;
      RECT 118.15 42.84 118.32 44.01 ;
      RECT 117.29 42.84 117.46 44.01 ;
      RECT 118.285 45.28 118.96 45.45 ;
      RECT 118.79 44.58 118.96 45.28 ;
      RECT 118.79 45.45 118.96 45.59 ;
      RECT 117.61 45.76 120.14 45.93 ;
      RECT 118.58 44.18 120.14 44.35 ;
      RECT 117.61 44.58 117.78 45.76 ;
      RECT 118.58 42.84 118.75 44.18 ;
      RECT 119.44 42.84 119.61 44.18 ;
      RECT 119.97 44.35 120.14 45.76 ;
      RECT 117.61 45.93 117.78 47.08 ;
      RECT 116.215 49.09 116.885 50.625 ;
      RECT 118.13 46.165 118.46 47.015 ;
      RECT 118.21 47.015 118.38 47.625 ;
      RECT 116.91 46.335 117.44 47.37 ;
      RECT 116.91 47.37 117.78 48.38 ;
      RECT 117.28 50.625 117.65 55.42 ;
      RECT 117.165 49.085 117.835 50.625 ;
      RECT 120.215 41.76 120.745 41.93 ;
      RECT 120.435 41.93 120.745 43.11 ;
      RECT 120.33 43.11 120.86 48.39 ;
      RECT 119.01 42.84 119.18 44.01 ;
      RECT 119.87 42.84 120.04 44.01 ;
      RECT 122.015 44.57 123.025 44.74 ;
      RECT 122.015 44.74 122.545 44.8 ;
      RECT 121.91 42.605 122.08 44.4 ;
      RECT 122.13 42 122.8 42.17 ;
      RECT 122.2 42.17 122.73 42.3 ;
      RECT 121.925 45.03 122.47 45.2 ;
      RECT 122.3 45 122.47 45.03 ;
      RECT 122.3 45.2 122.47 48 ;
      RECT 122.43 42.505 122.96 42.675 ;
      RECT 122.79 42.675 122.96 43.615 ;
      RECT 123.305 44.57 124.315 44.74 ;
      RECT 123.785 44.74 124.315 44.8 ;
      RECT 123.53 42 124.2 42.17 ;
      RECT 123.6 42.17 124.13 42.3 ;
      RECT 123.86 45.03 124.405 45.2 ;
      RECT 123.86 45 124.03 45.03 ;
      RECT 123.86 45.2 124.03 48 ;
      RECT 123.37 42.505 123.9 42.675 ;
      RECT 123.37 42.675 123.54 43.615 ;
      RECT 119.61 46.335 120.14 46.505 ;
      RECT 119.97 46.1 120.14 46.335 ;
      RECT 119.97 46.505 120.14 48.38 ;
      RECT 118.72 49.595 120.75 49.765 ;
      RECT 119.78 48.99 120.31 49.595 ;
      RECT 123.08 45.29 123.25 48 ;
      RECT 121.52 45.29 121.69 48 ;
      RECT 121.64 48.215 124.69 48.35 ;
      RECT 121.48 48.35 124.85 48.52 ;
      RECT 123.41 49.045 124.08 49.765 ;
      RECT 127.37 48.55 130.26 48.72 ;
      RECT 130.07 44.35 130.26 47.37 ;
      RECT 128.44 44.18 130.26 44.35 ;
      RECT 128.44 42.84 128.61 44.18 ;
      RECT 129.3 42.84 129.47 44.18 ;
      RECT 127.37 46.1 127.54 48.55 ;
      RECT 129.73 47.37 130.26 48.55 ;
      RECT 126.19 45.76 128.72 45.93 ;
      RECT 126.19 44.18 127.75 44.35 ;
      RECT 128.55 44.58 128.72 45.76 ;
      RECT 126.72 42.84 126.89 44.18 ;
      RECT 127.58 42.84 127.75 44.18 ;
      RECT 126.19 44.35 126.36 45.76 ;
      RECT 128.55 45.93 128.72 47.08 ;
      RECT 125.585 41.76 126.115 41.93 ;
      RECT 125.585 41.93 125.895 43.11 ;
      RECT 125.47 43.11 126 48.39 ;
      RECT 72.81 44.82 72.98 47.555 ;
      RECT 74.4 47.555 74.93 47.725 ;
      RECT 74.57 47.725 74.74 49.57 ;
      RECT 74.57 44.82 74.74 47.555 ;
      RECT 76.16 47.555 76.69 47.725 ;
      RECT 76.33 47.725 76.5 49.57 ;
      RECT 76.33 44.82 76.5 47.555 ;
      RECT 77.92 47.555 78.45 47.725 ;
      RECT 78.09 47.725 78.26 49.57 ;
      RECT 78.09 44.82 78.26 47.555 ;
      RECT 82.69 47.57 83.22 47.74 ;
      RECT 82.87 47.74 83.04 49.57 ;
      RECT 82.87 44.82 83.04 47.57 ;
      RECT 79.75 47.57 80.28 47.74 ;
      RECT 79.75 47.74 79.92 49.57 ;
      RECT 79.75 44.82 79.92 47.57 ;
      RECT 81.13 47.57 81.66 47.74 ;
      RECT 81.31 47.74 81.48 49.57 ;
      RECT 81.31 44.82 81.48 47.57 ;
      RECT 88.88 48.845 89.41 49.015 ;
      RECT 88.88 44.82 89.05 48.845 ;
      RECT 88.88 49.015 89.05 50.08 ;
      RECT 83.995 50.08 89.05 50.265 ;
      RECT 87.38 48.355 87.91 48.525 ;
      RECT 87.55 48.525 87.72 49.57 ;
      RECT 87.55 44.82 87.72 48.355 ;
      RECT 85.8 48.355 86.33 48.525 ;
      RECT 85.99 48.525 86.16 49.57 ;
      RECT 85.99 44.82 86.16 48.355 ;
      RECT 84.24 48.37 84.77 48.54 ;
      RECT 84.43 48.54 84.6 49.57 ;
      RECT 84.43 44.82 84.6 48.37 ;
      RECT 90.05 49.74 92.29 49.91 ;
      RECT 91.76 51.24 92.29 51.41 ;
      RECT 92 44.82 92.29 49.74 ;
      RECT 92 51.41 92.29 54.43 ;
      RECT 92 49.91 92.29 51.24 ;
      RECT 90.05 49.91 90.22 50.67 ;
      RECT 90.25 48.845 90.78 49.015 ;
      RECT 90.44 49.015 90.61 49.57 ;
      RECT 90.44 44.82 90.61 48.845 ;
      RECT 92.99 50.035 93.52 50.205 ;
      RECT 93.05 50.84 94.48 51.14 ;
      RECT 94.21 51.14 94.48 54.43 ;
      RECT 94.21 44.82 94.48 50.84 ;
      RECT 93.05 50.015 93.22 50.035 ;
      RECT 93.05 50.205 93.22 50.84 ;
      RECT 92.55 49.665 93.08 49.835 ;
      RECT 92.55 49.835 92.82 54.43 ;
      RECT 92.55 44.82 92.82 49.665 ;
      RECT 93.77 45.575 94.04 50 ;
      RECT 93.75 50 94.04 50.67 ;
      RECT 95.76 46.99 99.89 47.125 ;
      RECT 95.72 46.5 99.97 46.99 ;
      RECT 100.63 43.51 100.8 44.4 ;
      RECT 104.45 43.11 104.98 43.28 ;
      RECT 104.565 41.76 105.095 41.93 ;
      RECT 104.565 41.93 104.875 43.11 ;
      RECT 104.59 43.28 104.76 48.39 ;
      RECT 105.17 45.76 107.7 45.93 ;
      RECT 105.17 44.18 106.73 44.35 ;
      RECT 107.53 44.58 107.7 45.76 ;
      RECT 105.7 42.84 105.87 44.18 ;
      RECT 106.56 42.84 106.73 44.18 ;
      RECT 105.17 44.35 105.34 45.76 ;
      RECT 107.53 45.93 107.7 47.08 ;
      RECT 106.35 48.55 109.24 48.72 ;
      RECT 109.05 44.35 109.24 47.37 ;
      RECT 107.42 44.18 109.24 44.35 ;
      RECT 107.42 42.84 107.59 44.18 ;
      RECT 108.28 42.84 108.45 44.18 ;
      RECT 106.35 46.1 106.52 48.55 ;
      RECT 108.71 47.37 109.24 48.55 ;
      RECT 102.285 44.57 103.4 44.74 ;
      RECT 102.765 44.74 103.4 44.8 ;
      RECT 103.23 42.605 103.4 44.57 ;
      RECT 102.51 42 103.18 42.17 ;
      RECT 102.58 42.17 103.11 42.3 ;
      RECT 102.35 42.505 102.88 42.675 ;
      RECT 102.35 42.675 102.52 43.615 ;
      RECT 105.555 42.47 106.905 42.64 ;
      RECT 105.655 42.64 106.905 42.67 ;
      RECT 105.27 42.84 105.44 44.01 ;
      RECT 106.13 42.84 106.3 44.01 ;
      RECT 106.35 45.28 107.025 45.45 ;
      RECT 106.35 45.45 106.52 45.59 ;
      RECT 106.35 44.58 106.52 45.28 ;
      RECT 102.84 45.03 103.385 45.2 ;
      RECT 102.84 45 103.01 45.03 ;
      RECT 102.84 45.2 103.01 48 ;
      RECT 102.06 45.29 102.23 48 ;
      RECT 103.62 45.29 103.79 48 ;
      RECT 102.06 48.215 103.67 48.35 ;
      RECT 102.145 48.385 103.83 48.52 ;
      RECT 102.06 48.35 103.83 48.385 ;
      RECT 105.17 46.335 105.7 46.505 ;
      RECT 105.17 46.1 105.34 46.335 ;
      RECT 105.17 46.505 105.34 48.38 ;
      RECT 109.05 43.095 109.58 43.265 ;
      RECT 109.41 43.265 109.58 48.39 ;
      RECT 107.26 42.475 109.92 42.645 ;
      RECT 109.75 42.645 109.92 43.405 ;
      RECT 109.87 46.335 110.4 46.505 ;
      RECT 107.26 42.47 108.61 42.475 ;
      RECT 110.23 46.505 110.4 48.085 ;
      RECT 110.23 44.415 110.4 46.335 ;
      RECT 109.75 43.405 110.4 44.415 ;
      RECT 111.745 46.335 112.275 46.505 ;
      RECT 112.07 43.405 112.275 44.415 ;
      RECT 111.52 48.105 112.275 48.275 ;
      RECT 112.105 46.505 112.275 48.105 ;
      RECT 112.105 44.415 112.275 46.335 ;
      RECT 106.99 42.84 107.16 44.01 ;
      RECT 108.71 42.84 108.88 44.01 ;
      RECT 108.35 45.28 108.88 45.45 ;
      RECT 108.71 44.58 108.88 45.28 ;
      RECT 108.71 45.45 108.88 47.08 ;
      RECT 107.85 42.84 108.02 44.01 ;
      RECT 111.91 42.2 112.08 42.305 ;
      RECT 111.91 41.635 112.08 42.03 ;
      RECT 111.05 42.03 112.08 42.2 ;
      RECT 111.805 42.51 112.34 43.085 ;
      RECT 111.73 44.415 111.9 44.52 ;
      RECT 111.61 43.405 111.9 44.415 ;
      RECT 111.73 44.52 111.935 45.3 ;
      RECT 111.27 44.74 111.52 45.375 ;
      RECT 111.03 44.585 111.52 44.74 ;
      RECT 29.975 51.305 30.3 52.535 ;
      RECT 29.975 50.82 30.145 51.305 ;
      RECT 32.95 46.97 33.12 50.37 ;
      RECT 26.84 46.8 33.12 46.97 ;
      RECT 25.1 53.175 33.12 53.265 ;
      RECT 29.975 50.54 30.96 50.82 ;
      RECT 32.95 50.54 33.12 53.175 ;
      RECT 22.59 42.025 23.375 42.195 ;
      RECT 22.65 42.195 23.2 42.495 ;
      RECT 21.295 42.025 22.42 42.195 ;
      RECT 21.295 52.675 22.42 52.845 ;
      RECT 22.25 42.195 22.42 52.675 ;
      RECT 27.14 48.245 27.31 49.595 ;
      RECT 28.54 47.675 29.21 47.845 ;
      RECT 28.875 47.845 29.045 48.78 ;
      RECT 26.36 46.445 26.53 47.795 ;
      RECT 26.635 42.02 27.305 42.98 ;
      RECT 35.415 43.61 36.095 44.275 ;
      RECT 26.635 43.28 36.095 43.61 ;
      RECT 30.045 48.245 30.215 49.74 ;
      RECT 26.36 48.245 26.53 49.595 ;
      RECT 29.265 48.245 29.435 49.595 ;
      RECT 28.485 48.1 28.655 49.595 ;
      RECT 27.705 48.245 27.875 49.595 ;
      RECT 29.49 47.675 32.27 47.845 ;
      RECT 32.325 48.245 32.495 49.74 ;
      RECT 36.465 48.415 41.215 48.585 ;
      RECT 35.415 44.575 36.085 45.535 ;
      RECT 36.465 48.945 41.215 49.115 ;
      RECT 36.075 48.64 36.245 49.42 ;
      RECT 41.755 49.185 41.925 49.955 ;
      RECT 41.755 48.105 41.925 48.825 ;
      RECT 35.7 48.105 35.875 49.955 ;
      RECT 35.7 47.905 41.215 47.935 ;
      RECT 35.7 50.125 41.81 50.135 ;
      RECT 35.7 47.935 41.925 48.105 ;
      RECT 35.7 49.955 41.925 50.125 ;
      RECT 41.78 45.27 42.31 45.44 ;
      RECT 41.79 45.44 42.3 45.535 ;
      RECT 41.79 45.205 42.3 45.27 ;
      RECT 41.78 44.64 42.31 44.81 ;
      RECT 41.79 44.81 42.3 44.905 ;
      RECT 41.79 44.575 42.3 44.64 ;
      RECT 41.78 44.015 42.31 44.185 ;
      RECT 41.79 44.185 42.3 44.275 ;
      RECT 41.79 43.945 42.3 44.015 ;
      RECT 45.305 47.305 62.64 50.015 ;
      RECT 48.075 45.27 48.605 45.44 ;
      RECT 48.085 45.44 48.595 45.535 ;
      RECT 48.085 45.205 48.595 45.27 ;
      RECT 48.075 44.025 48.605 44.195 ;
      RECT 48.085 44.195 48.595 44.275 ;
      RECT 48.085 43.945 48.595 44.025 ;
      RECT 48.075 44.64 48.605 44.81 ;
      RECT 48.085 44.81 48.595 44.905 ;
      RECT 48.085 44.575 48.595 44.64 ;
      RECT 52.585 45.27 53.115 45.44 ;
      RECT 52.595 45.44 53.105 45.535 ;
      RECT 52.595 45.205 53.105 45.27 ;
      RECT 53.695 42.65 54.49 42.98 ;
      RECT 52.46 42.65 53.13 43.61 ;
      RECT 52.46 42.02 54.485 42.35 ;
      RECT 54.37 44.64 54.9 44.81 ;
      RECT 54.38 44.81 54.89 44.905 ;
      RECT 54.38 44.575 54.89 44.64 ;
      RECT 54.37 44.02 54.9 44.19 ;
      RECT 54.38 44.19 54.89 44.275 ;
      RECT 54.38 43.945 54.89 44.02 ;
      RECT 57.095 45.27 57.625 45.44 ;
      RECT 57.105 45.44 57.615 45.535 ;
      RECT 57.105 45.205 57.615 45.27 ;
      RECT 58.78 42.755 59.31 42.925 ;
      RECT 56.595 44.575 61.91 44.905 ;
      RECT 56.595 43.945 61.91 44.275 ;
      RECT 61.24 44.275 61.91 44.575 ;
      RECT 65.475 50.61 67.085 50.665 ;
      RECT 64.56 50.44 67.085 50.61 ;
      RECT 64.56 44.3 94.96 44.47 ;
      RECT 91.22 44.47 91.39 49.57 ;
      RECT 89.66 44.47 89.83 49.57 ;
      RECT 93.43 44.47 93.6 49.57 ;
      RECT 80.53 44.47 80.7 49.57 ;
      RECT 83.65 44.47 83.82 49.57 ;
      RECT 82.09 44.47 82.26 49.57 ;
      RECT 85.21 44.47 85.38 49.57 ;
      RECT 86.77 44.47 86.94 49.57 ;
      RECT 88.33 44.47 88.5 49.57 ;
      RECT 94.79 44.47 94.96 49.84 ;
      RECT 64.56 44.47 64.73 50.44 ;
      RECT 71.93 44.47 72.1 49.57 ;
      RECT 73.69 44.47 73.86 49.57 ;
      RECT 77.21 44.47 77.38 49.57 ;
      RECT 75.45 44.47 75.62 49.57 ;
      RECT 78.97 44.47 79.14 49.57 ;
      RECT 65.14 48.355 65.67 48.525 ;
      RECT 65.14 48.525 65.31 49.57 ;
      RECT 65.14 44.82 65.31 48.355 ;
      RECT 61.12 45.245 61.91 45.495 ;
      RECT 61.12 45.495 61.51 45.535 ;
      RECT 61.12 45.205 61.51 45.245 ;
      RECT 65.73 47.97 66.26 48.14 ;
      RECT 65.92 48.14 66.09 49.57 ;
      RECT 65.92 44.82 66.09 47.97 ;
      RECT 62.18 42.65 80.19 42.98 ;
      RECT 68.09 48.355 68.62 48.525 ;
      RECT 68.26 48.525 68.43 49.57 ;
      RECT 68.26 44.82 68.43 48.355 ;
      RECT 71.02 48.355 71.55 48.525 ;
      RECT 71.38 48.525 71.55 49.57 ;
      RECT 71.38 44.82 71.55 48.355 ;
      RECT 66.525 48.355 67.055 48.525 ;
      RECT 66.7 48.525 66.87 49.57 ;
      RECT 66.7 44.82 66.87 48.355 ;
      RECT 67.29 47.97 67.82 48.14 ;
      RECT 67.48 48.14 67.65 49.57 ;
      RECT 67.48 44.82 67.65 47.97 ;
      RECT 69.65 48.355 70.18 48.525 ;
      RECT 69.82 48.525 69.99 49.57 ;
      RECT 69.82 44.82 69.99 48.355 ;
      RECT 70.43 47.555 70.96 47.725 ;
      RECT 70.6 47.725 70.77 49.57 ;
      RECT 70.6 44.82 70.77 47.555 ;
      RECT 68.87 47.555 69.4 47.725 ;
      RECT 69.04 47.725 69.21 49.57 ;
      RECT 69.04 44.82 69.21 47.555 ;
      RECT 72.64 47.555 73.17 47.725 ;
      RECT 72.81 47.725 72.98 49.57 ;
      RECT 422.525 41.17 422.695 46.915 ;
      RECT 421.645 41.17 421.815 42.22 ;
      RECT 424.835 41.17 425.005 42.235 ;
      RECT 423.075 41.17 423.245 42.99 ;
      RECT 423.955 41.295 424.125 46.915 ;
      RECT 421.065 40.2 423.165 40.37 ;
      RECT 421.065 40.37 421.235 42.45 ;
      RECT 421.065 42.45 421.815 42.78 ;
      RECT 424.035 40.2 424.925 40.37 ;
      RECT 426.055 41 426.425 47.08 ;
      RECT 425.975 38.175 426.505 41 ;
      RECT 425.985 47.08 426.495 47.41 ;
      RECT 427.485 41 427.855 47.08 ;
      RECT 427.405 39.375 427.935 41 ;
      RECT 427.415 47.08 427.925 47.41 ;
      RECT 428.295 40.67 428.805 41 ;
      RECT 428.365 41 428.735 47.08 ;
      RECT 428.295 47.08 428.805 47.41 ;
      RECT 429.315 41 429.685 47.08 ;
      RECT 429.235 38.575 429.765 41 ;
      RECT 429.245 47.08 429.755 47.41 ;
      RECT 430.195 41 430.565 47.08 ;
      RECT 430.115 38.575 430.645 41 ;
      RECT 430.125 47.08 430.635 47.41 ;
      RECT 426.595 41.17 426.765 42.99 ;
      RECT 427.145 41.17 427.315 42.99 ;
      RECT 428.905 41.17 429.075 42.235 ;
      RECT 430.805 41.17 430.975 42.22 ;
      RECT 425.715 41.295 425.885 46.915 ;
      RECT 428.025 41.295 428.195 46.915 ;
      RECT 426.69 40.2 427.22 40.37 ;
      RECT 429.855 41.17 430.025 45.64 ;
      RECT 430.815 40.17 432.385 40.37 ;
      RECT 428.135 40.2 429.025 40.37 ;
      RECT 432.645 41 433.015 47.08 ;
      RECT 432.565 37.775 433.095 41 ;
      RECT 432.575 47.08 433.085 47.41 ;
      RECT 431.695 40.67 432.205 41 ;
      RECT 431.765 41 432.135 47.08 ;
      RECT 431.695 47.08 432.205 47.41 ;
      RECT 435.905 41 436.275 47.08 ;
      RECT 435.825 38.145 436.355 41 ;
      RECT 435.835 47.08 436.345 47.41 ;
      RECT 436.785 41 437.155 47.08 ;
      RECT 436.705 38.575 437.235 41 ;
      RECT 436.715 47.08 437.225 47.41 ;
      RECT 434.475 41 434.845 47.08 ;
      RECT 434.395 39.375 434.925 41 ;
      RECT 434.405 47.08 434.915 47.41 ;
      RECT 433.525 40.67 434.035 41 ;
      RECT 433.595 41 433.965 47.08 ;
      RECT 433.525 47.08 434.035 47.41 ;
      RECT 435.565 41.17 435.735 43.35 ;
      RECT 435.015 41.17 435.185 42.99 ;
      RECT 433.255 41.17 433.425 42.235 ;
      RECT 431.355 41.17 431.525 42.22 ;
      RECT 436.445 41.295 436.615 46.915 ;
      RECT 434.135 41.295 434.305 46.915 ;
      RECT 435.095 40.2 435.655 40.37 ;
      RECT 433.265 40.2 434.225 40.37 ;
      RECT 432.305 41.17 432.475 45.64 ;
      RECT 437.325 41.17 437.495 42.235 ;
      RECT 437.405 40.2 440.605 40.37 ;
      RECT 439.355 40.67 439.865 41 ;
      RECT 439.425 41 439.795 47.08 ;
      RECT 439.355 47.08 439.865 47.41 ;
      RECT 439.525 40.57 439.695 40.67 ;
      RECT 438.475 40.67 438.985 41 ;
      RECT 438.545 41 438.915 47.08 ;
      RECT 438.475 47.08 438.985 47.41 ;
      RECT 437.595 40.67 438.105 41 ;
      RECT 437.665 41 438.035 47.08 ;
      RECT 437.595 47.08 438.105 47.41 ;
      RECT 441.735 41 442.105 47.08 ;
      RECT 441.655 38.565 442.185 41 ;
      RECT 441.665 47.08 442.175 47.41 ;
      RECT 440.855 41 441.225 47.08 ;
      RECT 440.775 36.975 441.305 41 ;
      RECT 440.785 47.08 441.295 47.41 ;
      RECT 439.085 41.17 439.255 42.22 ;
      RECT 442.275 41.17 442.445 43.35 ;
      RECT 440.515 41.17 440.685 42.235 ;
      RECT 439.965 41.17 440.135 46.915 ;
      RECT 438.205 41.17 438.375 46.91 ;
      RECT 441.395 41.295 441.565 46.915 ;
      RECT 442.355 40.2 442.915 40.37 ;
      RECT 443.165 41 443.535 47.08 ;
      RECT 443.085 38.965 443.615 41 ;
      RECT 443.095 47.08 443.605 47.41 ;
      RECT 443.975 40.67 444.485 41 ;
      RECT 444.045 41 444.415 47.08 ;
      RECT 443.975 47.08 444.485 47.41 ;
      RECT 442.825 41.17 442.995 42.99 ;
      RECT 444.585 41.17 444.755 42.235 ;
      RECT 443.705 41.295 443.875 46.915 ;
      RECT 443.785 40.17 445.335 40.37 ;
      RECT 444.955 40.37 445.335 41.74 ;
      RECT 444.955 41.74 446.35 42.405 ;
      RECT 444.585 42.405 446.35 42.78 ;
      RECT 454.1 38.695 454.27 43.445 ;
      RECT 453.22 38.695 453.39 43.445 ;
      RECT 455.86 38.695 456.03 43.445 ;
      RECT 456.74 38.695 457.25 43.505 ;
      RECT 454.98 38.695 455.15 43.445 ;
      RECT 463.275 37.215 463.445 39.925 ;
      RECT 461.845 38.695 462.565 39.945 ;
      RECT 462.055 39.945 462.565 39.985 ;
      RECT 462.055 37.215 462.565 38.695 ;
      RECT 463.275 33.955 463.445 36.665 ;
      RECT 461.845 35.415 462.565 36.665 ;
      RECT 462.055 33.895 462.565 35.415 ;
      RECT 14.21 43.425 14.54 44.015 ;
      RECT 16.655 42.025 17.78 42.195 ;
      RECT 16.655 52.675 17.78 52.845 ;
      RECT 17.61 42.195 17.78 52.675 ;
      RECT 19.89 42.025 21.015 42.195 ;
      RECT 19.89 52.675 21.015 52.845 ;
      RECT 19.89 42.195 20.06 52.675 ;
      RECT 25.58 48.245 25.75 49.595 ;
      RECT 25.58 46.445 25.75 47.795 ;
      RECT 25.1 45.925 27.01 46.095 ;
      RECT 29.975 50.37 33.12 50.54 ;
      RECT 26.84 46.095 27.01 46.8 ;
      RECT 25.1 46.095 25.27 53.095 ;
      RECT 25.1 53.095 30.145 53.175 ;
      RECT 25.13 53.265 33.12 53.345 ;
      RECT 29.975 52.535 30.145 53.095 ;
      RECT 292.755 38.09 292.925 38.73 ;
      RECT 296.845 36.955 297.38 37.125 ;
      RECT 296.845 37.125 297.015 37.41 ;
      RECT 296.845 35.93 297.015 36.955 ;
      RECT 292.755 40.575 293.29 40.745 ;
      RECT 292.755 40.745 292.925 40.93 ;
      RECT 292.755 39.65 292.925 40.575 ;
      RECT 296.845 40.575 297.38 40.745 ;
      RECT 296.845 40.745 297.015 40.93 ;
      RECT 296.845 37.69 297.015 40.575 ;
      RECT 297.235 40.985 299.945 41.155 ;
      RECT 297.235 37.465 299.945 37.635 ;
      RECT 293.585 40.985 296.295 41.155 ;
      RECT 293.585 37.465 296.295 37.635 ;
      RECT 297.235 35.705 299.945 35.875 ;
      RECT 293.585 35.705 296.295 35.875 ;
      RECT 297.235 40.105 299.945 40.275 ;
      RECT 297.235 39.225 299.945 39.395 ;
      RECT 297.235 38.345 299.945 38.515 ;
      RECT 293.585 40.105 296.295 40.275 ;
      RECT 293.585 39.225 296.295 39.395 ;
      RECT 293.585 38.345 296.295 38.515 ;
      RECT 297.235 36.585 299.945 36.755 ;
      RECT 293.585 36.585 296.295 36.755 ;
      RECT 301.835 35.125 306.195 35.295 ;
      RECT 306.025 35.295 306.195 41.565 ;
      RECT 301.835 41.565 306.195 41.735 ;
      RECT 301.92 35.04 306.11 35.125 ;
      RECT 301.445 39.185 302.005 39.355 ;
      RECT 301.835 39.355 302.005 41.565 ;
      RECT 301.835 35.295 302.005 39.185 ;
      RECT 302.245 39.78 302.415 40.93 ;
      RECT 302.245 39.61 302.83 39.78 ;
      RECT 302.245 37.69 302.415 39.61 ;
      RECT 300.495 40.745 300.665 40.93 ;
      RECT 300.095 40.575 300.665 40.745 ;
      RECT 300.495 37.69 300.665 40.575 ;
      RECT 302.245 36.955 302.78 37.125 ;
      RECT 302.245 37.125 302.415 37.41 ;
      RECT 302.245 35.93 302.415 36.955 ;
      RECT 300.495 35.93 300.665 37.52 ;
      RECT 302.635 37.465 305.345 37.635 ;
      RECT 302.635 40.985 305.345 41.155 ;
      RECT 302.635 35.705 305.345 35.875 ;
      RECT 302.635 38.345 305.345 38.515 ;
      RECT 302.635 39.225 305.345 39.395 ;
      RECT 302.635 40.105 305.345 40.275 ;
      RECT 302.635 36.585 305.345 36.755 ;
      RECT 306.665 41.355 308.685 42.105 ;
      RECT 309.815 37.61 331.93 37.94 ;
      RECT 309.815 38.24 331.93 38.57 ;
      RECT 309.815 37.94 310.485 38.24 ;
      RECT 309.815 38.87 331.93 39.2 ;
      RECT 309.815 39.5 331.93 39.83 ;
      RECT 309.815 39.2 310.485 39.5 ;
      RECT 309.815 40.76 331.93 41.09 ;
      RECT 309.815 40.13 331.93 40.46 ;
      RECT 309.815 40.46 310.485 40.76 ;
      RECT 309.815 36.98 327.76 37.31 ;
      RECT 309.815 41.39 331.93 41.72 ;
      RECT 309.815 42.02 331.93 42.35 ;
      RECT 309.815 41.72 310.485 42.02 ;
      RECT 330.695 37.055 331.225 37.225 ;
      RECT 335.5 36.98 336.31 37.31 ;
      RECT 335.52 38.24 336.31 39.2 ;
      RECT 335.52 37.61 336.31 37.94 ;
      RECT 335.52 40.76 337.545 41.09 ;
      RECT 336.875 40.13 363.37 40.46 ;
      RECT 335.52 39.5 336.31 40.46 ;
      RECT 335.52 41.39 337.545 41.72 ;
      RECT 339.435 35.025 339.605 35.695 ;
      RECT 339.435 33.845 339.605 34.515 ;
      RECT 350.145 33.845 350.315 34.515 ;
      RECT 350.145 35.025 350.315 35.695 ;
      RECT 351.025 35.025 351.195 35.695 ;
      RECT 351.025 33.845 351.195 34.515 ;
      RECT 366.265 38.545 366.435 41.255 ;
      RECT 361.735 35.025 361.905 35.695 ;
      RECT 361.735 33.845 361.905 34.515 ;
      RECT 362.7 40.76 363.37 41.72 ;
      RECT 366.345 34.025 366.515 36.775 ;
      RECT 366.57 37.285 367.57 37.455 ;
      RECT 367.37 37.825 368.85 37.995 ;
      RECT 366.42 37.825 367.09 37.995 ;
      RECT 371.275 34.325 372.285 34.345 ;
      RECT 372.865 34.325 373.535 34.345 ;
      RECT 371.275 34.345 373.96 34.515 ;
      RECT 371.275 37.105 372.285 37.125 ;
      RECT 372.865 37.105 373.535 37.125 ;
      RECT 371.275 36.935 373.96 37.105 ;
      RECT 370.915 37.675 371.085 40.385 ;
      RECT 372.475 37.675 372.645 40.385 ;
      RECT 367.625 34.025 367.795 36.735 ;
      RECT 368.025 38.385 368.29 41.255 ;
      RECT 371.695 37.675 371.865 40.385 ;
      RECT 370.49 40.635 374.405 40.805 ;
      RECT 374.235 37.365 374.405 40.635 ;
      RECT 367.85 37.285 368.85 37.455 ;
      RECT 373.755 37.675 373.925 40.385 ;
      RECT 399.1 40.34 407.11 40.745 ;
      RECT 399.1 40.33 402.83 40.34 ;
      RECT 403.38 40.33 407.11 40.34 ;
      RECT 407.955 40.09 408.135 62.06 ;
      RECT 398.15 40.09 398.33 62.06 ;
      RECT 417.76 40.09 417.94 62.06 ;
      RECT 398.15 39.91 417.94 40.09 ;
      RECT 398.15 62.06 417.94 62.24 ;
      RECT 403 35.08 408.77 35.25 ;
      RECT 409.21 35.08 410.56 35.25 ;
      RECT 410.905 35.08 411.915 35.25 ;
      RECT 411.705 37.585 412.295 37.755 ;
      RECT 411.705 35.25 411.915 37.585 ;
      RECT 408.98 40.34 416.99 40.745 ;
      RECT 408.98 40.33 412.71 40.34 ;
      RECT 413.26 40.33 416.99 40.34 ;
      RECT 421.915 40.67 422.425 41 ;
      RECT 421.985 41 422.355 47.08 ;
      RECT 421.915 47.08 422.425 47.41 ;
      RECT 425.175 41 425.545 47.08 ;
      RECT 425.095 36.975 425.625 40.67 ;
      RECT 425.105 47.08 425.615 47.41 ;
      RECT 424.295 41 424.665 47.08 ;
      RECT 424.225 47.08 424.735 47.41 ;
      RECT 424.225 40.67 425.625 41 ;
      RECT 423.415 41 423.785 47.08 ;
      RECT 423.335 39.345 423.865 41 ;
      RECT 423.345 47.08 423.855 47.41 ;
      RECT 269.12 41.085 269.79 41.255 ;
      RECT 269.305 41.265 270.27 41.435 ;
      RECT 269.74 42.13 270.27 42.3 ;
      RECT 267.535 37.505 269.675 37.595 ;
      RECT 269.305 37.595 269.675 41.085 ;
      RECT 269.305 41.255 269.79 41.265 ;
      RECT 269.96 41.435 270.27 42.13 ;
      RECT 267.535 37.335 269.79 37.505 ;
      RECT 268.965 37.765 269.135 40.865 ;
      RECT 268.625 40.865 268.795 41.445 ;
      RECT 268.625 41.445 269.09 41.615 ;
      RECT 268.92 41.615 269.09 42.52 ;
      RECT 268.805 42.52 269.09 42.69 ;
      RECT 268.085 40.395 268.795 40.865 ;
      RECT 268.805 42.69 268.975 43.615 ;
      RECT 268.085 38.155 268.255 40.395 ;
      RECT 272.575 37.045 274.605 37.505 ;
      RECT 273.69 38.18 273.95 41.16 ;
      RECT 274.565 41.29 275.235 41.46 ;
      RECT 274.625 42.03 275.155 42.2 ;
      RECT 274.66 41.46 275.155 42.03 ;
      RECT 274.66 38.18 274.83 41.29 ;
      RECT 271.99 41.36 272.52 41.53 ;
      RECT 272.35 37.84 276.59 38.01 ;
      RECT 275.845 41.29 276.59 41.46 ;
      RECT 275.915 41.46 276.445 41.53 ;
      RECT 272.35 38.01 272.52 41.36 ;
      RECT 276.42 38.01 276.59 41.29 ;
      RECT 273.23 38.18 273.49 41.16 ;
      RECT 269.96 40.865 270.13 41.095 ;
      RECT 269.845 38.155 270.13 40.865 ;
      RECT 271.77 37.87 271.94 40.87 ;
      RECT 273.865 41.36 274.395 41.53 ;
      RECT 274.045 41.53 274.215 42.305 ;
      RECT 270.425 37.765 270.595 40.845 ;
      RECT 280.095 37.335 282.125 37.505 ;
      RECT 278.11 37.84 282.35 38.01 ;
      RECT 282.18 41.36 282.71 41.53 ;
      RECT 278.11 41.29 278.855 41.46 ;
      RECT 278.255 41.46 278.785 41.53 ;
      RECT 278.11 38.01 278.28 41.29 ;
      RECT 282.18 38.01 282.35 41.36 ;
      RECT 279.465 41.29 280.135 41.46 ;
      RECT 279.545 42.03 280.075 42.2 ;
      RECT 279.545 41.46 280.04 42.03 ;
      RECT 279.87 38.18 280.04 41.29 ;
      RECT 277.62 37.505 277.79 39.51 ;
      RECT 277.62 37.335 279.885 37.505 ;
      RECT 274.815 37.335 275.485 37.505 ;
      RECT 275.765 37.335 276.435 37.505 ;
      RECT 275.865 37.505 276.035 37.51 ;
      RECT 275.865 36.98 276.035 37.335 ;
      RECT 280.305 41.36 280.835 41.53 ;
      RECT 280.485 41.53 280.655 42.305 ;
      RECT 278.99 38.18 279.295 40.89 ;
      RECT 279.125 40.89 279.295 41.58 ;
      RECT 279.125 41.635 279.375 42.305 ;
      RECT 279.125 41.58 279.34 41.635 ;
      RECT 279.17 42.305 279.34 43.405 ;
      RECT 279.145 43.405 279.34 44.415 ;
      RECT 275.18 39.675 275.71 39.845 ;
      RECT 275.405 40.89 275.575 41.58 ;
      RECT 275.405 39.845 275.71 40.89 ;
      RECT 275.405 38.18 275.71 39.675 ;
      RECT 275.325 41.635 275.575 42.305 ;
      RECT 275.36 41.58 275.575 41.635 ;
      RECT 275.36 42.305 275.53 43.405 ;
      RECT 275.36 43.405 275.555 44.415 ;
      RECT 277.265 40.87 277.435 44.425 ;
      RECT 277 37.87 277.435 40.87 ;
      RECT 278.615 34.015 281.615 34.325 ;
      RECT 280.75 38.18 281.01 41.16 ;
      RECT 281.21 38.18 281.47 41.16 ;
      RECT 284.91 41.085 285.58 41.255 ;
      RECT 284.43 41.265 285.395 41.435 ;
      RECT 286.785 37.595 287.165 38.615 ;
      RECT 284.43 42.13 284.96 42.3 ;
      RECT 284.91 41.255 285.395 41.265 ;
      RECT 284.43 41.435 284.74 42.13 ;
      RECT 285.025 37.505 287.165 37.595 ;
      RECT 285.025 37.595 285.395 41.085 ;
      RECT 284.91 37.335 287.165 37.505 ;
      RECT 285.565 37.765 285.735 40.865 ;
      RECT 284.57 40.865 284.74 41.095 ;
      RECT 284.57 38.155 284.855 40.865 ;
      RECT 282.76 37.87 282.93 40.87 ;
      RECT 285.61 41.445 286.075 41.615 ;
      RECT 285.905 40.865 286.075 41.445 ;
      RECT 285.61 41.615 285.78 42.52 ;
      RECT 285.61 42.52 285.895 42.69 ;
      RECT 285.905 40.395 286.615 40.865 ;
      RECT 285.725 42.69 285.895 43.615 ;
      RECT 286.445 38.155 286.615 40.395 ;
      RECT 286.245 41.53 286.57 41.785 ;
      RECT 285.95 41.785 286.57 42.115 ;
      RECT 286.245 41.36 287.165 41.53 ;
      RECT 286.995 40.195 287.165 41.36 ;
      RECT 284.105 37.765 284.275 40.845 ;
      RECT 289.205 37.87 289.375 42.475 ;
      RECT 290.445 41.465 301.075 41.635 ;
      RECT 300.905 35.395 301.075 41.465 ;
      RECT 290.445 34.845 290.615 41.465 ;
      RECT 294.605 34.845 294.775 35.04 ;
      RECT 290.445 34.64 294.775 34.845 ;
      RECT 294.605 35.04 301.075 35.395 ;
      RECT 292.075 36.46 292.325 37.26 ;
      RECT 292.075 35.325 292.245 36.46 ;
      RECT 290.895 35.155 292.245 35.325 ;
      RECT 288.755 34.32 288.925 35.6 ;
      RECT 287.525 34.095 288.535 34.265 ;
      RECT 287.525 35.655 288.535 35.825 ;
      RECT 292.415 39.595 292.585 40.985 ;
      RECT 292.415 38.035 292.585 39.425 ;
      RECT 290.895 40.985 292.585 41.155 ;
      RECT 290.895 39.425 292.585 39.595 ;
      RECT 290.895 37.865 292.585 38.035 ;
      RECT 290.895 37.315 291.905 37.485 ;
      RECT 290.895 36.235 291.905 36.405 ;
      RECT 287.095 38.97 287.945 39.72 ;
      RECT 287.335 39.72 287.945 40.865 ;
      RECT 287.335 37.765 287.945 38.97 ;
      RECT 287.525 34.875 288.535 35.045 ;
      RECT 290.895 38.645 292.245 38.815 ;
      RECT 290.895 40.205 292.245 40.375 ;
      RECT 292.48 35.38 292.65 36.37 ;
      RECT 292.755 38.73 293.29 38.9 ;
      RECT 292.755 38.9 292.925 39.37 ;
      RECT 242.985 37.505 245.125 37.595 ;
      RECT 242.985 37.595 243.355 41.085 ;
      RECT 242.87 37.335 245.125 37.505 ;
      RECT 242.53 40.865 242.7 41.095 ;
      RECT 242.53 38.155 242.815 40.865 ;
      RECT 240.72 37.87 240.89 40.87 ;
      RECT 242.065 37.765 242.235 40.845 ;
      RECT 245.055 38.97 246.585 39.72 ;
      RECT 245.295 39.72 246.345 40.865 ;
      RECT 245.295 37.765 246.345 38.97 ;
      RECT 243.91 41.785 244.53 42.115 ;
      RECT 244.205 41.53 244.53 41.785 ;
      RECT 244.205 41.36 245.125 41.53 ;
      RECT 244.955 40.195 245.125 41.36 ;
      RECT 243.525 37.765 243.695 40.865 ;
      RECT 243.865 40.865 244.035 41.445 ;
      RECT 243.57 41.445 244.035 41.615 ;
      RECT 243.57 41.615 243.74 42.52 ;
      RECT 243.57 42.52 243.855 42.69 ;
      RECT 243.865 40.395 244.575 40.865 ;
      RECT 243.685 42.69 243.855 43.615 ;
      RECT 244.405 38.155 244.575 40.395 ;
      RECT 246.515 37.595 246.895 38.615 ;
      RECT 248.1 41.085 248.77 41.255 ;
      RECT 248.285 41.265 249.25 41.435 ;
      RECT 248.72 42.13 249.25 42.3 ;
      RECT 248.285 41.255 248.77 41.265 ;
      RECT 248.94 41.435 249.25 42.13 ;
      RECT 248.285 37.595 248.655 41.085 ;
      RECT 246.515 37.505 248.655 37.595 ;
      RECT 246.515 37.335 248.77 37.505 ;
      RECT 247.11 41.785 247.73 42.115 ;
      RECT 247.11 41.53 247.435 41.785 ;
      RECT 246.515 41.36 247.435 41.53 ;
      RECT 246.515 40.195 246.685 41.36 ;
      RECT 247.945 37.765 248.115 40.865 ;
      RECT 248.94 40.865 249.11 41.095 ;
      RECT 248.825 38.155 249.11 40.865 ;
      RECT 247.605 40.865 247.775 41.445 ;
      RECT 247.605 41.445 248.07 41.615 ;
      RECT 247.9 41.615 248.07 42.52 ;
      RECT 247.785 42.52 248.07 42.69 ;
      RECT 247.065 40.395 247.775 40.865 ;
      RECT 247.785 42.69 247.955 43.615 ;
      RECT 247.065 38.155 247.235 40.395 ;
      RECT 250.75 37.87 250.92 40.87 ;
      RECT 249.405 37.765 249.575 40.845 ;
      RECT 251.555 37.335 253.585 37.505 ;
      RECT 250.97 41.36 251.5 41.53 ;
      RECT 251.33 37.84 255.57 38.01 ;
      RECT 254.825 41.29 255.57 41.46 ;
      RECT 254.895 41.46 255.425 41.53 ;
      RECT 251.33 38.01 251.5 41.36 ;
      RECT 255.4 38.01 255.57 41.29 ;
      RECT 252.21 38.18 252.47 41.16 ;
      RECT 252.67 38.18 252.93 41.16 ;
      RECT 253.545 41.29 254.215 41.46 ;
      RECT 253.605 42.03 254.135 42.2 ;
      RECT 253.64 41.46 254.135 42.03 ;
      RECT 253.64 38.18 253.81 41.29 ;
      RECT 253.795 37.335 254.465 37.505 ;
      RECT 254.745 37.335 255.415 37.505 ;
      RECT 254.385 40.89 254.555 41.58 ;
      RECT 254.385 38.18 254.69 40.89 ;
      RECT 254.305 41.635 254.555 42.305 ;
      RECT 254.34 41.58 254.555 41.635 ;
      RECT 254.34 42.305 254.51 43.405 ;
      RECT 254.34 43.405 254.535 44.415 ;
      RECT 256.245 37.87 256.415 44.425 ;
      RECT 252.845 41.36 253.375 41.53 ;
      RECT 253.025 41.53 253.195 42.305 ;
      RECT 257.09 37.84 261.33 38.01 ;
      RECT 261.16 41.36 261.69 41.53 ;
      RECT 257.09 41.29 257.835 41.46 ;
      RECT 257.235 41.46 257.765 41.53 ;
      RECT 257.09 38.01 257.26 41.29 ;
      RECT 261.16 38.01 261.33 41.36 ;
      RECT 257.245 37.335 257.915 37.505 ;
      RECT 259.075 37.335 261.105 37.505 ;
      RECT 259.73 38.18 259.99 41.16 ;
      RECT 258.445 41.29 259.115 41.46 ;
      RECT 258.525 42.03 259.055 42.2 ;
      RECT 258.525 41.46 259.02 42.03 ;
      RECT 258.85 38.18 259.02 41.29 ;
      RECT 260.19 38.18 260.45 41.16 ;
      RECT 258.195 37.335 258.865 37.505 ;
      RECT 258.105 40.89 258.275 41.58 ;
      RECT 257.97 38.18 258.275 40.89 ;
      RECT 258.105 41.635 258.355 42.305 ;
      RECT 258.105 41.58 258.32 41.635 ;
      RECT 258.15 42.305 258.32 43.405 ;
      RECT 258.125 43.405 258.32 44.415 ;
      RECT 261.74 37.87 261.91 40.87 ;
      RECT 259.285 41.36 259.815 41.53 ;
      RECT 259.465 41.53 259.635 42.305 ;
      RECT 263.085 37.765 263.255 40.845 ;
      RECT 263.89 41.085 264.56 41.255 ;
      RECT 263.41 41.265 264.375 41.435 ;
      RECT 265.765 37.595 266.145 38.615 ;
      RECT 263.41 42.13 263.94 42.3 ;
      RECT 263.89 41.255 264.375 41.265 ;
      RECT 263.41 41.435 263.72 42.13 ;
      RECT 264.005 37.505 266.145 37.595 ;
      RECT 264.005 37.595 264.375 41.085 ;
      RECT 263.89 37.335 266.145 37.505 ;
      RECT 264.545 37.765 264.715 40.865 ;
      RECT 263.55 40.865 263.72 41.095 ;
      RECT 263.55 38.155 263.835 40.865 ;
      RECT 264.885 40.865 265.055 41.445 ;
      RECT 264.59 41.445 265.055 41.615 ;
      RECT 264.59 41.615 264.76 42.52 ;
      RECT 264.59 42.52 264.875 42.69 ;
      RECT 264.885 40.395 265.595 40.865 ;
      RECT 265.425 38.155 265.595 40.395 ;
      RECT 264.705 42.69 264.875 43.615 ;
      RECT 266.075 38.97 267.605 39.72 ;
      RECT 266.315 39.72 267.365 40.865 ;
      RECT 266.315 37.765 267.365 38.97 ;
      RECT 264.93 41.785 265.55 42.115 ;
      RECT 265.225 41.53 265.55 41.785 ;
      RECT 265.225 41.36 266.145 41.53 ;
      RECT 265.975 40.195 266.145 41.36 ;
      RECT 268.13 41.785 268.75 42.115 ;
      RECT 268.13 41.53 268.455 41.785 ;
      RECT 267.535 41.36 268.455 41.53 ;
      RECT 267.535 40.195 267.705 41.36 ;
      RECT 267.535 37.595 267.915 38.615 ;
      RECT 216.715 34.145 216.885 35.165 ;
      RECT 216.715 33.815 217.435 34.145 ;
      RECT 214.205 37.87 214.375 44.425 ;
      RECT 218.685 33.815 218.855 34.145 ;
      RECT 217.265 34.315 217.435 35.325 ;
      RECT 218.685 34.315 218.855 35.325 ;
      RECT 220.655 35.165 221.185 35.335 ;
      RECT 220.655 34.145 220.825 35.165 ;
      RECT 220.105 33.815 220.825 34.145 ;
      RECT 220.105 34.315 220.275 35.325 ;
      RECT 217.035 37.335 219.065 37.505 ;
      RECT 217.69 38.18 217.95 41.16 ;
      RECT 218.15 38.18 218.41 41.16 ;
      RECT 217.245 41.36 217.775 41.53 ;
      RECT 217.425 41.53 217.595 42.305 ;
      RECT 221.85 41.085 222.52 41.255 ;
      RECT 221.37 41.265 222.335 41.435 ;
      RECT 223.725 37.595 224.105 38.615 ;
      RECT 221.37 42.13 221.9 42.3 ;
      RECT 221.85 41.255 222.335 41.265 ;
      RECT 221.37 41.435 221.68 42.13 ;
      RECT 221.965 37.505 224.105 37.595 ;
      RECT 221.965 37.595 222.335 41.085 ;
      RECT 221.85 37.335 224.105 37.505 ;
      RECT 222.505 37.765 222.675 40.865 ;
      RECT 221.51 40.865 221.68 41.095 ;
      RECT 221.51 38.155 221.795 40.865 ;
      RECT 219.7 37.87 219.87 40.87 ;
      RECT 221.045 37.765 221.215 40.845 ;
      RECT 222.55 41.445 223.015 41.615 ;
      RECT 222.845 40.865 223.015 41.445 ;
      RECT 222.55 41.615 222.72 42.52 ;
      RECT 222.55 42.52 222.835 42.69 ;
      RECT 222.845 40.395 223.555 40.865 ;
      RECT 222.665 42.69 222.835 43.615 ;
      RECT 223.385 38.155 223.555 40.395 ;
      RECT 223.305 33.86 223.475 34.915 ;
      RECT 224.035 38.97 225.565 39.72 ;
      RECT 224.275 39.72 225.325 40.865 ;
      RECT 224.275 37.765 225.325 38.97 ;
      RECT 222.89 41.785 223.51 42.115 ;
      RECT 223.185 41.53 223.51 41.785 ;
      RECT 223.185 41.36 224.105 41.53 ;
      RECT 223.935 40.195 224.105 41.36 ;
      RECT 225.495 37.595 225.875 38.615 ;
      RECT 227.08 41.085 227.75 41.255 ;
      RECT 227.265 41.265 228.23 41.435 ;
      RECT 227.7 42.13 228.23 42.3 ;
      RECT 225.495 37.505 227.635 37.595 ;
      RECT 227.265 37.595 227.635 41.085 ;
      RECT 227.265 41.255 227.75 41.265 ;
      RECT 227.92 41.435 228.23 42.13 ;
      RECT 225.495 37.335 227.75 37.505 ;
      RECT 226.09 41.785 226.71 42.115 ;
      RECT 226.09 41.53 226.415 41.785 ;
      RECT 225.495 41.36 226.415 41.53 ;
      RECT 225.495 40.195 225.665 41.36 ;
      RECT 223.21 35.165 231.785 35.335 ;
      RECT 225.865 33.86 226.035 34.915 ;
      RECT 226.925 37.765 227.095 40.865 ;
      RECT 227.92 40.865 228.09 41.095 ;
      RECT 227.805 38.155 228.09 40.865 ;
      RECT 226.585 40.865 226.755 41.445 ;
      RECT 226.585 41.445 227.05 41.615 ;
      RECT 226.88 41.615 227.05 42.52 ;
      RECT 226.765 42.52 227.05 42.69 ;
      RECT 226.045 40.395 226.755 40.865 ;
      RECT 226.765 42.69 226.935 43.615 ;
      RECT 226.045 38.155 226.215 40.395 ;
      RECT 228.385 37.765 228.555 40.845 ;
      RECT 230.535 37.335 232.565 37.505 ;
      RECT 231.65 38.18 231.91 41.16 ;
      RECT 232.525 41.29 233.195 41.46 ;
      RECT 232.585 42.03 233.115 42.2 ;
      RECT 232.62 41.46 233.115 42.03 ;
      RECT 232.62 38.18 232.79 41.29 ;
      RECT 229.95 41.36 230.48 41.53 ;
      RECT 230.31 37.84 234.55 38.01 ;
      RECT 233.805 41.29 234.55 41.46 ;
      RECT 233.875 41.46 234.405 41.53 ;
      RECT 230.31 38.01 230.48 41.36 ;
      RECT 234.38 38.01 234.55 41.29 ;
      RECT 231.19 38.18 231.45 41.16 ;
      RECT 228.975 33.86 229.145 34.915 ;
      RECT 231.535 33.86 231.705 34.915 ;
      RECT 232.775 37.335 233.445 37.505 ;
      RECT 233.725 37.335 234.395 37.505 ;
      RECT 233.365 40.89 233.535 41.58 ;
      RECT 233.365 38.18 233.67 40.89 ;
      RECT 233.285 41.635 233.535 42.305 ;
      RECT 233.32 41.58 233.535 41.635 ;
      RECT 233.32 42.305 233.49 43.405 ;
      RECT 233.32 43.405 233.515 44.415 ;
      RECT 229.73 37.87 229.9 40.87 ;
      RECT 231.825 41.36 232.355 41.53 ;
      RECT 232.005 41.53 232.175 42.305 ;
      RECT 236.07 37.84 240.31 38.01 ;
      RECT 240.14 41.36 240.67 41.53 ;
      RECT 236.07 41.29 236.815 41.46 ;
      RECT 236.215 41.46 236.745 41.53 ;
      RECT 236.07 38.01 236.24 41.29 ;
      RECT 240.14 38.01 240.31 41.36 ;
      RECT 235.225 37.87 235.395 44.425 ;
      RECT 238.055 37.335 240.085 37.505 ;
      RECT 239.17 38.18 239.43 41.16 ;
      RECT 238.71 38.18 238.97 41.16 ;
      RECT 237.425 41.29 238.095 41.46 ;
      RECT 237.505 42.03 238.035 42.2 ;
      RECT 237.505 41.46 238 42.03 ;
      RECT 237.83 38.18 238 41.29 ;
      RECT 237.175 37.335 237.845 37.505 ;
      RECT 237.585 36.975 237.755 37.335 ;
      RECT 236.225 37.335 236.895 37.505 ;
      RECT 237.085 40.89 237.255 41.58 ;
      RECT 236.95 38.18 237.255 40.89 ;
      RECT 237.085 41.635 237.335 42.305 ;
      RECT 237.085 41.58 237.3 41.635 ;
      RECT 237.13 42.305 237.3 43.405 ;
      RECT 237.105 43.405 237.3 44.415 ;
      RECT 238.265 41.36 238.795 41.53 ;
      RECT 238.445 41.53 238.615 42.305 ;
      RECT 242.87 41.085 243.54 41.255 ;
      RECT 242.39 41.265 243.355 41.435 ;
      RECT 244.745 37.595 245.125 38.615 ;
      RECT 242.39 42.13 242.92 42.3 ;
      RECT 242.87 41.255 243.355 41.265 ;
      RECT 242.39 41.435 242.7 42.13 ;
      RECT 156.89 42.03 157.42 42.2 ;
      RECT 156.89 41.46 157.385 42.03 ;
      RECT 157.215 38.18 157.385 41.29 ;
      RECT 158.555 38.18 158.815 41.16 ;
      RECT 156.56 37.335 157.23 37.505 ;
      RECT 155.61 37.335 156.28 37.505 ;
      RECT 156.47 40.89 156.64 41.58 ;
      RECT 156.335 38.18 156.64 40.89 ;
      RECT 156.47 41.635 156.72 42.305 ;
      RECT 156.47 41.58 156.685 41.635 ;
      RECT 156.515 42.305 156.685 43.405 ;
      RECT 156.49 43.405 156.685 44.415 ;
      RECT 157.65 41.36 158.18 41.53 ;
      RECT 157.83 41.53 158 42.305 ;
      RECT 163.97 33.86 164.14 34.915 ;
      RECT 160.86 33.86 161.03 34.915 ;
      RECT 164.13 37.595 164.51 38.615 ;
      RECT 162.255 41.085 162.925 41.255 ;
      RECT 161.775 41.265 162.74 41.435 ;
      RECT 161.775 42.13 162.305 42.3 ;
      RECT 162.255 41.255 162.74 41.265 ;
      RECT 161.775 41.435 162.085 42.13 ;
      RECT 162.37 37.595 162.74 41.085 ;
      RECT 162.37 37.505 164.51 37.595 ;
      RECT 162.255 37.335 164.51 37.505 ;
      RECT 163.295 41.785 163.915 42.115 ;
      RECT 163.59 41.53 163.915 41.785 ;
      RECT 163.59 41.36 164.51 41.53 ;
      RECT 164.34 40.195 164.51 41.36 ;
      RECT 162.91 37.765 163.08 40.865 ;
      RECT 161.915 40.865 162.085 41.095 ;
      RECT 161.915 38.155 162.2 40.865 ;
      RECT 163.25 40.865 163.42 41.445 ;
      RECT 162.955 41.445 163.42 41.615 ;
      RECT 162.955 41.615 163.125 42.52 ;
      RECT 162.955 42.52 163.24 42.69 ;
      RECT 163.25 40.395 163.96 40.865 ;
      RECT 163.07 42.69 163.24 43.615 ;
      RECT 163.79 38.155 163.96 40.395 ;
      RECT 160.105 37.87 160.275 40.87 ;
      RECT 161.45 37.765 161.62 40.845 ;
      RECT 164.44 38.97 165.97 39.72 ;
      RECT 164.68 39.72 165.73 40.865 ;
      RECT 164.68 37.765 165.73 38.97 ;
      RECT 166.53 33.86 166.7 34.915 ;
      RECT 168.82 35.165 169.35 35.335 ;
      RECT 169.18 34.145 169.35 35.165 ;
      RECT 169.18 33.815 169.9 34.145 ;
      RECT 169.73 34.315 169.9 35.325 ;
      RECT 165.9 37.595 166.28 38.615 ;
      RECT 167.485 41.085 168.155 41.255 ;
      RECT 167.67 41.265 168.635 41.435 ;
      RECT 168.105 42.13 168.635 42.3 ;
      RECT 167.67 41.255 168.155 41.265 ;
      RECT 168.325 41.435 168.635 42.13 ;
      RECT 167.67 37.595 168.04 41.085 ;
      RECT 165.9 37.505 168.04 37.595 ;
      RECT 165.9 37.335 168.155 37.505 ;
      RECT 166.495 41.785 167.115 42.115 ;
      RECT 166.495 41.53 166.82 41.785 ;
      RECT 165.9 41.36 166.82 41.53 ;
      RECT 165.9 40.195 166.07 41.36 ;
      RECT 167.33 37.765 167.5 40.865 ;
      RECT 166.99 40.865 167.16 41.445 ;
      RECT 166.99 41.445 167.455 41.615 ;
      RECT 167.285 41.615 167.455 42.52 ;
      RECT 167.17 42.52 167.455 42.69 ;
      RECT 166.45 40.395 167.16 40.865 ;
      RECT 167.17 42.69 167.34 43.615 ;
      RECT 166.45 38.155 166.62 40.395 ;
      RECT 168.325 40.865 168.495 41.095 ;
      RECT 168.21 38.155 168.495 40.865 ;
      RECT 170.355 41.36 170.885 41.53 ;
      RECT 170.715 37.84 174.955 38.01 ;
      RECT 174.21 41.29 174.955 41.46 ;
      RECT 174.28 41.46 174.81 41.53 ;
      RECT 170.715 38.01 170.885 41.36 ;
      RECT 174.785 38.01 174.955 41.29 ;
      RECT 170.135 37.87 170.305 40.87 ;
      RECT 168.79 37.765 168.96 40.845 ;
      RECT 171.15 33.815 171.32 34.145 ;
      RECT 171.15 34.315 171.32 35.325 ;
      RECT 172.91 35.165 173.44 35.335 ;
      RECT 173.12 34.145 173.29 35.165 ;
      RECT 172.57 33.815 173.29 34.145 ;
      RECT 172.57 34.315 172.74 35.325 ;
      RECT 170.94 37.335 172.97 37.505 ;
      RECT 172.055 38.18 172.315 41.16 ;
      RECT 172.93 41.29 173.6 41.46 ;
      RECT 172.99 42.03 173.52 42.2 ;
      RECT 173.025 41.46 173.52 42.03 ;
      RECT 173.025 38.18 173.195 41.29 ;
      RECT 171.595 38.18 171.855 41.16 ;
      RECT 173.18 37.335 173.85 37.505 ;
      RECT 173.27 36.975 173.44 37.335 ;
      RECT 174.13 37.335 174.8 37.505 ;
      RECT 173.77 40.89 173.94 41.58 ;
      RECT 173.77 38.18 174.075 40.89 ;
      RECT 173.69 41.635 173.94 42.305 ;
      RECT 173.725 41.58 173.94 41.635 ;
      RECT 173.725 42.305 173.895 43.405 ;
      RECT 173.725 43.405 173.92 44.415 ;
      RECT 175.63 37.87 175.8 44.425 ;
      RECT 172.23 41.36 172.76 41.53 ;
      RECT 172.41 41.53 172.58 42.305 ;
      RECT 176.975 34.245 178.995 34.995 ;
      RECT 211.01 34.245 213.03 34.995 ;
      RECT 215.05 37.84 219.29 38.01 ;
      RECT 219.12 41.36 219.65 41.53 ;
      RECT 215.05 41.29 215.795 41.46 ;
      RECT 215.195 41.46 215.725 41.53 ;
      RECT 215.05 38.01 215.22 41.29 ;
      RECT 219.12 38.01 219.29 41.36 ;
      RECT 216.405 41.29 217.075 41.46 ;
      RECT 216.485 42.03 217.015 42.2 ;
      RECT 216.485 41.46 216.98 42.03 ;
      RECT 216.81 38.18 216.98 41.29 ;
      RECT 216.155 37.335 216.825 37.505 ;
      RECT 216.565 36.975 216.735 37.335 ;
      RECT 215.205 37.335 215.875 37.505 ;
      RECT 216.065 40.89 216.235 41.58 ;
      RECT 215.93 38.18 216.235 40.89 ;
      RECT 216.065 41.635 216.315 42.305 ;
      RECT 216.065 41.58 216.28 41.635 ;
      RECT 216.11 42.305 216.28 43.405 ;
      RECT 216.085 43.405 216.28 44.415 ;
      RECT 216.565 35.165 217.095 35.335 ;
      RECT 138.505 41.36 139.035 41.53 ;
      RECT 134.435 41.29 135.18 41.46 ;
      RECT 134.58 41.46 135.11 41.53 ;
      RECT 134.435 38.01 134.605 41.29 ;
      RECT 138.505 38.01 138.675 41.36 ;
      RECT 130.015 38.18 130.275 41.16 ;
      RECT 130.19 41.36 130.72 41.53 ;
      RECT 130.37 41.53 130.54 42.305 ;
      RECT 130.89 41.29 131.56 41.46 ;
      RECT 130.95 42.03 131.48 42.2 ;
      RECT 130.985 41.46 131.48 42.03 ;
      RECT 130.985 38.18 131.155 41.29 ;
      RECT 131.14 37.335 131.81 37.505 ;
      RECT 132.09 37.335 132.76 37.505 ;
      RECT 131.73 40.89 131.9 41.58 ;
      RECT 131.73 38.18 132.035 40.89 ;
      RECT 131.65 41.635 131.9 42.305 ;
      RECT 131.685 41.58 131.9 41.635 ;
      RECT 131.685 42.305 131.855 43.405 ;
      RECT 131.685 43.405 131.88 44.415 ;
      RECT 133.59 37.87 133.76 44.425 ;
      RECT 135.54 37.335 136.21 37.505 ;
      RECT 134.59 37.335 135.26 37.505 ;
      RECT 135.45 40.89 135.62 41.58 ;
      RECT 135.315 38.18 135.62 40.89 ;
      RECT 135.45 41.635 135.7 42.305 ;
      RECT 135.45 41.58 135.665 41.635 ;
      RECT 135.495 42.305 135.665 43.405 ;
      RECT 135.47 43.405 135.665 44.415 ;
      RECT 136.42 37.335 138.45 37.505 ;
      RECT 137.075 38.18 137.335 41.16 ;
      RECT 135.79 41.29 136.46 41.46 ;
      RECT 135.87 42.03 136.4 42.2 ;
      RECT 135.87 41.46 136.365 42.03 ;
      RECT 136.195 38.18 136.365 41.29 ;
      RECT 137.535 38.18 137.795 41.16 ;
      RECT 141.235 41.085 141.905 41.255 ;
      RECT 140.755 41.265 141.72 41.435 ;
      RECT 143.11 37.595 143.49 38.615 ;
      RECT 140.755 42.13 141.285 42.3 ;
      RECT 141.235 41.255 141.72 41.265 ;
      RECT 140.755 41.435 141.065 42.13 ;
      RECT 141.35 37.505 143.49 37.595 ;
      RECT 141.35 37.595 141.72 41.085 ;
      RECT 141.235 37.335 143.49 37.505 ;
      RECT 140.895 40.865 141.065 41.095 ;
      RECT 140.895 38.155 141.18 40.865 ;
      RECT 139.085 37.87 139.255 40.87 ;
      RECT 136.63 41.36 137.16 41.53 ;
      RECT 136.81 41.53 136.98 42.305 ;
      RECT 140.43 37.765 140.6 40.845 ;
      RECT 142.275 41.785 142.895 42.115 ;
      RECT 142.57 41.53 142.895 41.785 ;
      RECT 142.57 41.36 143.49 41.53 ;
      RECT 143.32 40.195 143.49 41.36 ;
      RECT 141.89 37.765 142.06 40.865 ;
      RECT 142.23 40.865 142.4 41.445 ;
      RECT 141.935 41.445 142.4 41.615 ;
      RECT 141.935 41.615 142.105 42.52 ;
      RECT 141.935 42.52 142.22 42.69 ;
      RECT 142.23 40.395 142.94 40.865 ;
      RECT 142.05 42.69 142.22 43.615 ;
      RECT 142.77 38.155 142.94 40.395 ;
      RECT 143.42 38.97 144.95 39.72 ;
      RECT 143.66 39.72 144.71 40.865 ;
      RECT 143.66 37.765 144.71 38.97 ;
      RECT 144.88 37.595 145.26 38.615 ;
      RECT 146.465 41.085 147.135 41.255 ;
      RECT 146.65 41.265 147.615 41.435 ;
      RECT 147.085 42.13 147.615 42.3 ;
      RECT 144.88 37.505 147.02 37.595 ;
      RECT 146.65 37.595 147.02 41.085 ;
      RECT 146.65 41.255 147.135 41.265 ;
      RECT 147.305 41.435 147.615 42.13 ;
      RECT 144.88 37.335 147.135 37.505 ;
      RECT 145.475 41.785 146.095 42.115 ;
      RECT 145.475 41.53 145.8 41.785 ;
      RECT 144.88 41.36 145.8 41.53 ;
      RECT 144.88 40.195 145.05 41.36 ;
      RECT 145.97 40.865 146.14 41.445 ;
      RECT 145.97 41.445 146.435 41.615 ;
      RECT 146.265 41.615 146.435 42.52 ;
      RECT 146.15 42.52 146.435 42.69 ;
      RECT 145.43 40.395 146.14 40.865 ;
      RECT 146.15 42.69 146.32 43.615 ;
      RECT 145.43 38.155 145.6 40.395 ;
      RECT 146.31 37.765 146.48 40.865 ;
      RECT 147.305 40.865 147.475 41.095 ;
      RECT 147.19 38.155 147.475 40.865 ;
      RECT 149.695 37.84 153.935 38.01 ;
      RECT 149.335 41.36 149.865 41.53 ;
      RECT 153.19 41.29 153.935 41.46 ;
      RECT 153.26 41.46 153.79 41.53 ;
      RECT 149.695 38.01 149.865 41.36 ;
      RECT 153.765 38.01 153.935 41.29 ;
      RECT 149.115 37.87 149.285 40.87 ;
      RECT 147.77 37.765 147.94 40.845 ;
      RECT 149.92 37.335 151.95 37.505 ;
      RECT 151.035 38.18 151.295 41.16 ;
      RECT 150.575 38.18 150.835 41.16 ;
      RECT 151.21 41.36 151.74 41.53 ;
      RECT 151.39 41.53 151.56 42.305 ;
      RECT 151.91 41.29 152.58 41.46 ;
      RECT 151.97 42.03 152.5 42.2 ;
      RECT 152.005 41.46 152.5 42.03 ;
      RECT 152.005 38.18 152.175 41.29 ;
      RECT 152.16 37.335 152.83 37.505 ;
      RECT 152.25 36.975 152.42 37.335 ;
      RECT 153.11 37.335 153.78 37.505 ;
      RECT 152.75 40.89 152.92 41.58 ;
      RECT 152.75 38.18 153.055 40.89 ;
      RECT 152.67 41.635 152.92 42.305 ;
      RECT 152.705 41.58 152.92 41.635 ;
      RECT 152.705 42.305 152.875 43.405 ;
      RECT 152.705 43.405 152.9 44.415 ;
      RECT 158.3 33.86 158.47 34.915 ;
      RECT 158.22 35.165 166.795 35.335 ;
      RECT 154.61 37.87 154.78 44.425 ;
      RECT 157.44 37.335 159.47 37.505 ;
      RECT 155.455 37.84 159.695 38.01 ;
      RECT 159.525 41.36 160.055 41.53 ;
      RECT 155.455 41.29 156.2 41.46 ;
      RECT 155.6 41.46 156.13 41.53 ;
      RECT 155.455 38.01 155.625 41.29 ;
      RECT 159.525 38.01 159.695 41.36 ;
      RECT 158.095 38.18 158.355 41.16 ;
      RECT 156.81 41.29 157.48 41.46 ;
      RECT 105.265 40.865 105.435 41.095 ;
      RECT 105.15 38.155 105.435 40.865 ;
      RECT 103.93 40.865 104.1 41.445 ;
      RECT 103.93 41.445 104.395 41.615 ;
      RECT 104.225 41.615 104.395 42.52 ;
      RECT 104.11 42.52 104.395 42.69 ;
      RECT 103.39 40.395 104.1 40.865 ;
      RECT 103.39 38.155 103.56 40.395 ;
      RECT 104.11 42.69 104.28 43.615 ;
      RECT 105.73 37.765 105.9 40.845 ;
      RECT 101.47 34.875 102.48 35.045 ;
      RECT 107.88 37.335 109.91 37.505 ;
      RECT 107.655 37.84 111.895 38.01 ;
      RECT 107.295 41.36 107.825 41.53 ;
      RECT 111.15 41.29 111.895 41.46 ;
      RECT 111.22 41.46 111.75 41.53 ;
      RECT 111.725 38.01 111.895 41.29 ;
      RECT 107.655 38.01 107.825 41.36 ;
      RECT 108.995 38.18 109.255 41.16 ;
      RECT 109.87 41.29 110.54 41.46 ;
      RECT 109.93 42.03 110.46 42.2 ;
      RECT 109.965 41.46 110.46 42.03 ;
      RECT 109.965 38.18 110.135 41.29 ;
      RECT 108.535 38.18 108.795 41.16 ;
      RECT 112.215 37.505 112.385 39.51 ;
      RECT 110.12 37.335 112.385 37.505 ;
      RECT 109.17 41.36 109.7 41.53 ;
      RECT 109.35 41.53 109.52 42.305 ;
      RECT 107.075 37.87 107.245 40.87 ;
      RECT 110.71 38.18 111.015 40.89 ;
      RECT 110.71 40.89 110.88 41.58 ;
      RECT 110.63 41.635 110.88 42.305 ;
      RECT 110.665 41.58 110.88 41.635 ;
      RECT 110.665 42.305 110.835 43.405 ;
      RECT 110.665 43.405 110.86 44.415 ;
      RECT 112.57 40.87 112.74 44.425 ;
      RECT 112.57 37.87 113.005 40.87 ;
      RECT 108.39 34.015 111.39 34.325 ;
      RECT 115.4 37.045 117.43 37.505 ;
      RECT 113.415 37.84 117.655 38.01 ;
      RECT 117.485 41.36 118.015 41.53 ;
      RECT 113.415 41.29 114.16 41.46 ;
      RECT 113.56 41.46 114.09 41.53 ;
      RECT 113.415 38.01 113.585 41.29 ;
      RECT 117.485 38.01 117.655 41.36 ;
      RECT 116.055 38.18 116.315 41.16 ;
      RECT 114.77 41.29 115.44 41.46 ;
      RECT 114.85 42.03 115.38 42.2 ;
      RECT 114.85 41.46 115.345 42.03 ;
      RECT 115.175 38.18 115.345 41.29 ;
      RECT 116.515 38.18 116.775 41.16 ;
      RECT 114.52 37.335 115.19 37.505 ;
      RECT 113.57 37.335 114.24 37.505 ;
      RECT 113.97 37.505 114.14 37.51 ;
      RECT 113.97 36.98 114.14 37.335 ;
      RECT 114.295 39.675 114.825 39.845 ;
      RECT 114.43 40.89 114.6 41.58 ;
      RECT 114.295 39.845 114.6 40.89 ;
      RECT 114.295 38.18 114.6 39.675 ;
      RECT 114.43 41.635 114.68 42.305 ;
      RECT 114.43 41.58 114.645 41.635 ;
      RECT 114.475 42.305 114.645 43.405 ;
      RECT 114.45 43.405 114.645 44.415 ;
      RECT 118.065 37.87 118.235 40.87 ;
      RECT 115.61 41.36 116.14 41.53 ;
      RECT 115.79 41.53 115.96 42.305 ;
      RECT 120.215 41.085 120.885 41.255 ;
      RECT 119.735 41.265 120.7 41.435 ;
      RECT 122.09 37.595 122.47 38.615 ;
      RECT 119.735 42.13 120.265 42.3 ;
      RECT 120.215 41.255 120.7 41.265 ;
      RECT 119.735 41.435 120.045 42.13 ;
      RECT 120.33 37.505 122.47 37.595 ;
      RECT 120.33 37.595 120.7 41.085 ;
      RECT 120.215 37.335 122.47 37.505 ;
      RECT 120.87 37.765 121.04 40.865 ;
      RECT 119.875 40.865 120.045 41.095 ;
      RECT 119.875 38.155 120.16 40.865 ;
      RECT 119.41 37.765 119.58 40.845 ;
      RECT 120.915 41.445 121.38 41.615 ;
      RECT 121.21 40.865 121.38 41.445 ;
      RECT 120.915 41.615 121.085 42.52 ;
      RECT 120.915 42.52 121.2 42.69 ;
      RECT 121.21 40.395 121.92 40.865 ;
      RECT 121.03 42.69 121.2 43.615 ;
      RECT 121.75 38.155 121.92 40.395 ;
      RECT 122.4 38.97 123.93 39.72 ;
      RECT 122.64 39.72 123.69 40.865 ;
      RECT 122.64 37.765 123.69 38.97 ;
      RECT 121.255 41.785 121.875 42.115 ;
      RECT 121.55 41.53 121.875 41.785 ;
      RECT 121.55 41.36 122.47 41.53 ;
      RECT 122.3 40.195 122.47 41.36 ;
      RECT 123.86 37.595 124.24 38.615 ;
      RECT 125.445 41.085 126.115 41.255 ;
      RECT 125.63 41.265 126.595 41.435 ;
      RECT 126.065 42.13 126.595 42.3 ;
      RECT 123.86 37.505 126 37.595 ;
      RECT 125.63 37.595 126 41.085 ;
      RECT 125.63 41.255 126.115 41.265 ;
      RECT 126.285 41.435 126.595 42.13 ;
      RECT 123.86 37.335 126.115 37.505 ;
      RECT 124.455 41.785 125.075 42.115 ;
      RECT 124.455 41.53 124.78 41.785 ;
      RECT 123.86 41.36 124.78 41.53 ;
      RECT 123.86 40.195 124.03 41.36 ;
      RECT 125.29 37.765 125.46 40.865 ;
      RECT 126.285 40.865 126.455 41.095 ;
      RECT 126.17 38.155 126.455 40.865 ;
      RECT 124.95 40.865 125.12 41.445 ;
      RECT 124.95 41.445 125.415 41.615 ;
      RECT 125.245 41.615 125.415 42.52 ;
      RECT 125.13 42.52 125.415 42.69 ;
      RECT 124.41 40.395 125.12 40.865 ;
      RECT 125.13 42.69 125.3 43.615 ;
      RECT 124.41 38.155 124.58 40.395 ;
      RECT 128.095 37.87 128.265 40.87 ;
      RECT 128.315 41.36 128.845 41.53 ;
      RECT 128.675 37.84 132.915 38.01 ;
      RECT 132.17 41.29 132.915 41.46 ;
      RECT 132.24 41.46 132.77 41.53 ;
      RECT 128.675 38.01 128.845 41.36 ;
      RECT 132.745 38.01 132.915 41.29 ;
      RECT 126.75 37.765 126.92 40.845 ;
      RECT 128.9 37.335 130.93 37.505 ;
      RECT 129.555 38.18 129.815 41.16 ;
      RECT 134.435 37.84 138.675 38.01 ;
      RECT 22.21 34.025 22.38 36.735 ;
      RECT 21.715 38.385 21.98 41.255 ;
      RECT 21.155 37.285 22.155 37.455 ;
      RECT 22.435 37.285 23.435 37.455 ;
      RECT 21.155 37.825 22.635 37.995 ;
      RECT 22.915 37.825 23.585 37.995 ;
      RECT 28.1 33.845 28.27 34.515 ;
      RECT 28.1 35.025 28.27 35.695 ;
      RECT 26.635 40.76 27.305 41.72 ;
      RECT 26.635 40.13 53.13 40.46 ;
      RECT 38.81 35.025 38.98 35.695 ;
      RECT 38.81 33.845 38.98 34.515 ;
      RECT 39.69 33.845 39.86 34.515 ;
      RECT 39.69 35.025 39.86 35.695 ;
      RECT 50.4 33.845 50.57 34.515 ;
      RECT 50.4 35.025 50.57 35.695 ;
      RECT 53.695 36.98 54.505 37.31 ;
      RECT 53.695 37.61 54.485 37.94 ;
      RECT 53.695 38.24 54.485 39.2 ;
      RECT 52.46 40.76 54.485 41.09 ;
      RECT 52.46 41.39 54.485 41.72 ;
      RECT 53.695 39.5 54.485 40.46 ;
      RECT 58.78 37.055 59.31 37.225 ;
      RECT 58.075 41.39 80.19 41.72 ;
      RECT 58.075 42.02 80.19 42.35 ;
      RECT 79.52 41.72 80.19 42.02 ;
      RECT 58.075 39.5 80.19 39.83 ;
      RECT 58.075 38.87 80.19 39.2 ;
      RECT 79.52 39.2 80.19 39.5 ;
      RECT 58.075 40.13 80.19 40.46 ;
      RECT 58.075 40.76 80.19 41.09 ;
      RECT 79.52 40.46 80.19 40.76 ;
      RECT 58.075 38.24 80.19 38.57 ;
      RECT 58.075 37.61 80.19 37.94 ;
      RECT 79.52 37.94 80.19 38.24 ;
      RECT 62.245 36.98 80.19 37.31 ;
      RECT 81.32 41.355 83.34 42.105 ;
      RECT 83.81 35.125 88.17 35.295 ;
      RECT 83.81 35.295 83.98 41.565 ;
      RECT 83.81 41.565 88.17 41.735 ;
      RECT 83.895 35.04 88.085 35.125 ;
      RECT 88 39.185 88.56 39.355 ;
      RECT 88 39.355 88.17 41.565 ;
      RECT 88 35.295 88.17 39.185 ;
      RECT 87.59 39.78 87.76 40.93 ;
      RECT 87.175 39.61 87.76 39.78 ;
      RECT 87.59 37.69 87.76 39.61 ;
      RECT 88.93 35.395 89.1 41.465 ;
      RECT 88.93 41.465 99.56 41.635 ;
      RECT 99.39 34.845 99.56 41.465 ;
      RECT 95.23 34.845 95.4 35.04 ;
      RECT 88.93 35.04 95.4 35.395 ;
      RECT 95.23 34.64 99.56 34.845 ;
      RECT 89.34 40.745 89.51 40.93 ;
      RECT 89.34 40.575 89.91 40.745 ;
      RECT 89.34 37.69 89.51 40.575 ;
      RECT 87.225 36.955 87.76 37.125 ;
      RECT 87.59 37.125 87.76 37.41 ;
      RECT 87.59 35.93 87.76 36.955 ;
      RECT 89.34 35.93 89.51 37.52 ;
      RECT 84.66 37.465 87.37 37.635 ;
      RECT 84.66 40.985 87.37 41.155 ;
      RECT 84.66 35.705 87.37 35.875 ;
      RECT 84.66 38.345 87.37 38.515 ;
      RECT 84.66 39.225 87.37 39.395 ;
      RECT 84.66 40.105 87.37 40.275 ;
      RECT 84.66 36.585 87.37 36.755 ;
      RECT 92.625 36.955 93.16 37.125 ;
      RECT 92.99 37.125 93.16 37.41 ;
      RECT 92.99 35.93 93.16 36.955 ;
      RECT 92.625 40.575 93.16 40.745 ;
      RECT 92.99 40.745 93.16 40.93 ;
      RECT 92.99 37.69 93.16 40.575 ;
      RECT 90.06 40.985 92.77 41.155 ;
      RECT 90.06 37.465 92.77 37.635 ;
      RECT 93.71 40.985 96.42 41.155 ;
      RECT 93.71 37.465 96.42 37.635 ;
      RECT 90.06 35.705 92.77 35.875 ;
      RECT 93.71 35.705 96.42 35.875 ;
      RECT 90.06 40.105 92.77 40.275 ;
      RECT 90.06 39.225 92.77 39.395 ;
      RECT 90.06 38.345 92.77 38.515 ;
      RECT 93.71 40.105 96.42 40.275 ;
      RECT 93.71 39.225 96.42 39.395 ;
      RECT 93.71 38.345 96.42 38.515 ;
      RECT 90.06 36.585 92.77 36.755 ;
      RECT 93.71 36.585 96.42 36.755 ;
      RECT 100.63 37.87 100.8 42.475 ;
      RECT 97.355 35.38 97.525 36.37 ;
      RECT 97.68 36.46 97.93 37.26 ;
      RECT 97.76 35.325 97.93 36.46 ;
      RECT 97.76 35.155 99.11 35.325 ;
      RECT 96.715 40.575 97.25 40.745 ;
      RECT 97.08 40.745 97.25 40.93 ;
      RECT 97.08 39.65 97.25 40.575 ;
      RECT 96.715 38.73 97.25 38.9 ;
      RECT 97.08 38.9 97.25 39.37 ;
      RECT 97.08 38.09 97.25 38.73 ;
      RECT 97.42 39.595 97.59 40.985 ;
      RECT 97.42 38.035 97.59 39.425 ;
      RECT 97.42 40.985 99.11 41.155 ;
      RECT 97.42 39.425 99.11 39.595 ;
      RECT 97.42 37.865 99.11 38.035 ;
      RECT 98.1 37.315 99.11 37.485 ;
      RECT 98.1 36.235 99.11 36.405 ;
      RECT 97.76 38.645 99.11 38.815 ;
      RECT 97.76 40.205 99.11 40.375 ;
      RECT 101.08 34.32 101.25 35.6 ;
      RECT 101.47 34.095 102.48 34.265 ;
      RECT 101.47 35.655 102.48 35.825 ;
      RECT 102.84 37.595 103.22 38.615 ;
      RECT 104.425 41.085 105.095 41.255 ;
      RECT 104.61 41.265 105.575 41.435 ;
      RECT 105.045 42.13 105.575 42.3 ;
      RECT 104.61 41.255 105.095 41.265 ;
      RECT 105.265 41.435 105.575 42.13 ;
      RECT 104.61 37.595 104.98 41.085 ;
      RECT 102.84 37.505 104.98 37.595 ;
      RECT 102.84 37.335 105.095 37.505 ;
      RECT 102.06 38.97 102.91 39.72 ;
      RECT 102.06 39.72 102.67 40.865 ;
      RECT 102.06 37.765 102.67 38.97 ;
      RECT 103.435 41.785 104.055 42.115 ;
      RECT 103.435 41.53 103.76 41.785 ;
      RECT 102.84 41.36 103.76 41.53 ;
      RECT 102.84 40.195 103.01 41.36 ;
      RECT 104.27 37.765 104.44 40.865 ;
      RECT 413.855 31.215 414.385 31.385 ;
      RECT 414.155 31.385 414.325 31.755 ;
      RECT 414.155 31.085 414.325 31.215 ;
      RECT 417.295 30.475 417.465 30.805 ;
      RECT 417.295 31.425 417.465 31.755 ;
      RECT 416.57 35.185 417.395 35.355 ;
      RECT 417.225 34.635 417.395 35.185 ;
      RECT 416.415 31.925 417.465 34.635 ;
      RECT 413.855 31.925 414.385 35.28 ;
      RECT 416.075 28.895 416.605 31.045 ;
      RECT 414.075 28.895 414.725 30.175 ;
      RECT 415.635 31.925 415.805 34.635 ;
      RECT 414.495 30.845 415.025 31.015 ;
      RECT 414.555 31.015 415.025 34.635 ;
      RECT 414.555 30.815 415.025 30.845 ;
      RECT 415.195 29.165 415.805 31.3 ;
      RECT 415.195 31.3 416.245 31.755 ;
      RECT 415.195 31.755 415.465 35.08 ;
      RECT 415.975 31.755 416.245 35.08 ;
      RECT 415.195 35.08 416.245 36.06 ;
      RECT 418.995 28.995 420.265 29.025 ;
      RECT 419.065 29.025 419.435 35.09 ;
      RECT 418.995 28.695 422.71 28.995 ;
      RECT 419.945 29.025 420.265 35.09 ;
      RECT 418.995 35.09 420.265 35.435 ;
      RECT 418.725 29.195 418.895 34.94 ;
      RECT 418.175 29.195 418.345 34.94 ;
      RECT 426.935 29.025 427.305 35.105 ;
      RECT 423.66 28.695 427.375 28.995 ;
      RECT 426.105 28.995 427.375 29.025 ;
      RECT 426.105 29.025 426.425 35.105 ;
      RECT 426.105 35.105 427.375 35.435 ;
      RECT 419.605 29.195 419.775 30.245 ;
      RECT 419.605 30.475 419.775 30.805 ;
      RECT 419.605 31.425 419.775 31.755 ;
      RECT 419.605 31.925 419.775 34.635 ;
      RECT 420.465 29.165 420.995 35.69 ;
      RECT 422.685 30.85 422.855 31.755 ;
      RECT 421.03 27.735 421.7 27.905 ;
      RECT 421.98 27.735 422.65 27.905 ;
      RECT 422.685 31.925 423.685 36.06 ;
      RECT 421.985 29.165 422.995 30.175 ;
      RECT 421.985 30.175 422.515 35.69 ;
      RECT 423.1 30.43 423.27 30.805 ;
      RECT 421.265 29.165 421.815 36.06 ;
      RECT 423.515 30.85 423.685 31.755 ;
      RECT 424.48 27.735 425.15 27.905 ;
      RECT 423.375 29.165 424.385 30.175 ;
      RECT 423.855 30.175 424.385 35.69 ;
      RECT 424.555 29.165 425.105 36.06 ;
      RECT 425.375 29.165 425.905 35.69 ;
      RECT 428.295 28.695 432.01 28.995 ;
      RECT 428.295 28.995 429.565 29.025 ;
      RECT 428.365 29.025 428.735 35.09 ;
      RECT 428.295 35.105 429.565 35.435 ;
      RECT 429.245 29.025 429.565 35.09 ;
      RECT 428.365 35.09 429.565 35.105 ;
      RECT 425.43 27.735 426.1 27.905 ;
      RECT 428.025 29.195 428.195 34.94 ;
      RECT 428.905 29.195 429.075 30.245 ;
      RECT 427.475 29.195 427.645 34.94 ;
      RECT 426.595 29.195 426.765 30.245 ;
      RECT 428.905 30.475 429.075 30.805 ;
      RECT 426.595 30.475 426.765 30.805 ;
      RECT 428.905 31.425 429.075 31.755 ;
      RECT 426.595 31.425 426.765 31.755 ;
      RECT 428.905 31.925 429.075 34.635 ;
      RECT 426.595 31.925 426.765 34.635 ;
      RECT 429.765 29.165 430.295 34.635 ;
      RECT 430.565 29.165 431.115 36.06 ;
      RECT 436.125 29.165 436.295 30.245 ;
      RECT 431.985 30.85 432.155 31.755 ;
      RECT 438.525 29.165 439.075 30.6 ;
      RECT 438.525 30.77 439.075 32.635 ;
      RECT 438.105 32.635 439.075 33.305 ;
      RECT 438.525 33.305 439.075 33.985 ;
      RECT 438.525 33.985 439.535 34.155 ;
      RECT 436.925 30.6 439.075 30.77 ;
      RECT 431.985 31.925 432.515 36.06 ;
      RECT 436.125 32.255 436.295 34.965 ;
      RECT 431.285 29.165 432.295 30.175 ;
      RECT 431.285 30.175 431.815 34.635 ;
      RECT 436.585 29.165 436.755 34.965 ;
      RECT 435.645 35.315 441.255 35.485 ;
      RECT 435.645 31.945 435.815 35.315 ;
      RECT 437.525 31.945 437.695 35.315 ;
      RECT 441.085 31.945 441.255 35.315 ;
      RECT 437.745 29.165 437.915 30.245 ;
      RECT 437.045 29.165 437.215 30.245 ;
      RECT 439.305 29.165 439.475 30.245 ;
      RECT 440.865 29.165 441.035 30.245 ;
      RECT 442.01 27.735 442.72 27.905 ;
      RECT 439.245 33.445 440.255 33.615 ;
      RECT 439.705 34.295 440.675 34.965 ;
      RECT 439.705 33.615 440.255 34.295 ;
      RECT 439.705 29.165 440.255 33.445 ;
      RECT 437.945 30.94 438.355 31.47 ;
      RECT 437.045 32.255 437.215 34.965 ;
      RECT 438.025 33.575 438.335 34.965 ;
      RECT 440.445 32.555 440.765 34.025 ;
      RECT 440.425 30.94 440.755 31.47 ;
      RECT 443 27.735 443.67 27.905 ;
      RECT 453.22 31.915 453.39 36.665 ;
      RECT 454.1 31.915 454.27 36.665 ;
      RECT 453.445 30.785 456.74 30.955 ;
      RECT 453.445 30.955 454.925 31.405 ;
      RECT 454.98 31.915 455.15 36.665 ;
      RECT 456.74 31.855 457.25 36.665 ;
      RECT 455.205 31.235 456.685 31.405 ;
      RECT 455.86 31.915 456.03 36.665 ;
      RECT 460.84 33.235 463.23 33.405 ;
      RECT 460.84 33.405 461.01 33.515 ;
      RECT 460.84 32.985 461.01 33.235 ;
      RECT 17.72 34.325 18.73 34.345 ;
      RECT 16.47 34.325 17.14 34.345 ;
      RECT 16.045 34.345 18.73 34.515 ;
      RECT 17.72 37.105 18.73 37.125 ;
      RECT 16.47 37.105 17.14 37.125 ;
      RECT 16.045 36.935 18.73 37.105 ;
      RECT 18.92 37.675 19.09 40.385 ;
      RECT 17.36 37.675 17.53 40.385 ;
      RECT 16.08 37.675 16.25 40.385 ;
      RECT 18.14 37.675 18.31 40.385 ;
      RECT 15.6 40.635 19.515 40.805 ;
      RECT 15.6 37.365 15.77 40.635 ;
      RECT 23.57 38.545 23.74 41.255 ;
      RECT 23.49 34.025 23.66 36.775 ;
      RECT 339.435 32.665 339.605 33.335 ;
      RECT 339.435 31.485 339.605 32.155 ;
      RECT 341.195 25.785 341.845 26.115 ;
      RECT 341.195 27.045 341.845 27.375 ;
      RECT 341.195 26.415 341.845 26.745 ;
      RECT 341.195 27.675 341.845 28.005 ;
      RECT 338.535 30.425 338.705 36.59 ;
      RECT 362.36 30.425 362.53 36.58 ;
      RECT 338.535 36.75 340.015 36.76 ;
      RECT 338.535 30.255 362.53 30.425 ;
      RECT 339.905 36.58 362.53 36.59 ;
      RECT 338.535 36.59 362.53 36.75 ;
      RECT 344.795 27.4 345.465 27.9 ;
      RECT 347.875 27.305 350.585 27.475 ;
      RECT 355.175 27.305 357.885 27.475 ;
      RECT 350.145 32.665 350.315 33.335 ;
      RECT 350.145 31.485 350.315 32.155 ;
      RECT 351.025 32.665 351.195 33.335 ;
      RECT 351.025 31.485 351.195 32.155 ;
      RECT 366.265 30.195 366.435 32.905 ;
      RECT 367.145 30.195 367.315 32.905 ;
      RECT 365.3 29.49 365.47 30.665 ;
      RECT 363.855 30.665 365.47 30.835 ;
      RECT 365.3 29.32 367.46 29.49 ;
      RECT 363.855 30.295 365.11 30.465 ;
      RECT 364.94 29.15 365.11 30.295 ;
      RECT 364.94 28.98 368.25 29.15 ;
      RECT 367.72 29.15 368.25 29.49 ;
      RECT 361.735 32.665 361.905 33.335 ;
      RECT 361.735 31.485 361.905 32.155 ;
      RECT 365.67 53.095 374.155 53.265 ;
      RECT 365.67 52.565 365.965 53.095 ;
      RECT 365.67 51.935 365.84 52.565 ;
      RECT 373.985 42.71 374.155 53.095 ;
      RECT 373.985 41.775 374.32 42.71 ;
      RECT 370.665 41.775 371.675 53.095 ;
      RECT 365.67 41.775 365.965 51.935 ;
      RECT 365.67 41.605 375.34 41.775 ;
      RECT 368.905 41.57 375.34 41.605 ;
      RECT 365.67 39.135 365.965 41.605 ;
      RECT 368.905 38.545 369.67 41.57 ;
      RECT 367.145 41.13 367.315 41.605 ;
      RECT 367.145 38.545 367.315 39.04 ;
      RECT 367.145 39.04 367.32 41.13 ;
      RECT 365.67 37.025 365.84 39.135 ;
      RECT 369.5 36.775 369.67 38.545 ;
      RECT 375.17 36.4 375.34 41.57 ;
      RECT 368.905 36.4 369.67 36.775 ;
      RECT 368.905 35.05 375.34 36.4 ;
      RECT 368.905 34.025 369.67 35.05 ;
      RECT 369.5 32.905 369.67 34.025 ;
      RECT 365.67 30.35 365.965 37.025 ;
      RECT 365.67 29.845 365.84 30.35 ;
      RECT 375.17 29.88 375.34 35.05 ;
      RECT 368.905 29.88 369.67 32.905 ;
      RECT 368.905 29.845 375.34 29.88 ;
      RECT 365.67 29.675 375.34 29.845 ;
      RECT 366.42 33.455 367.09 33.625 ;
      RECT 367.37 33.455 368.85 33.625 ;
      RECT 370.915 31.065 371.085 33.775 ;
      RECT 372.475 31.065 372.645 33.775 ;
      RECT 368.025 30.195 368.26 33.065 ;
      RECT 371.695 31.065 371.865 33.775 ;
      RECT 370.435 30.645 374.405 30.815 ;
      RECT 374.235 30.815 374.405 34.085 ;
      RECT 370.435 30.815 370.605 34.085 ;
      RECT 373.755 31.065 373.925 33.775 ;
      RECT 375.285 27.93 377.305 28.68 ;
      RECT 388.79 27.735 389.12 29.785 ;
      RECT 388.16 27.735 388.49 29.785 ;
      RECT 387.53 27.735 387.86 29.785 ;
      RECT 386.27 27.735 386.6 29.785 ;
      RECT 386.9 27.735 387.23 29.785 ;
      RECT 389.42 27.735 389.75 29.785 ;
      RECT 390.05 27.735 390.38 29.785 ;
      RECT 390.68 27.735 391.01 31.07 ;
      RECT 391.31 27.735 391.64 29.885 ;
      RECT 393.2 27.735 393.53 29.885 ;
      RECT 393.83 27.56 394.16 29.885 ;
      RECT 391.94 27.735 392.27 29.885 ;
      RECT 392.57 27.735 392.9 29.885 ;
      RECT 395.72 27.735 396.05 29.855 ;
      RECT 395.09 27.56 395.42 29.855 ;
      RECT 394.46 27.735 394.79 29.855 ;
      RECT 396.35 27.56 396.68 29.855 ;
      RECT 393.83 33.58 394.16 35.64 ;
      RECT 394.46 33.58 394.79 35.64 ;
      RECT 395.72 33.58 396.05 35.075 ;
      RECT 395.09 33.58 395.42 35.075 ;
      RECT 396.35 35.89 396.91 36.06 ;
      RECT 396.35 33.58 396.68 35.89 ;
      RECT 402.09 35.49 411.535 35.67 ;
      RECT 402.09 29.29 412.72 29.47 ;
      RECT 412.54 29.47 412.72 35.49 ;
      RECT 412.085 35.49 412.72 35.67 ;
      RECT 402.09 29.47 402.27 35.49 ;
      RECT 398.87 27.295 399.2 29.855 ;
      RECT 398.24 27.735 398.57 29.855 ;
      RECT 397.61 27.56 397.94 29.855 ;
      RECT 396.98 27.735 397.31 29.855 ;
      RECT 399.5 27.735 399.83 29.855 ;
      RECT 399.5 33.58 399.83 35.075 ;
      RECT 398.87 33.58 399.2 35.075 ;
      RECT 398.24 33.58 398.57 35.075 ;
      RECT 397.61 33.58 397.94 35.075 ;
      RECT 396.98 33.58 397.31 35.075 ;
      RECT 402.68 29.82 402.85 34.57 ;
      RECT 404.41 27.735 405.08 27.905 ;
      RECT 403.46 27.735 404.13 27.905 ;
      RECT 407.36 29.82 407.53 34.57 ;
      RECT 405.8 29.82 405.97 34.57 ;
      RECT 404.24 29.82 404.41 34.57 ;
      RECT 406.58 29.82 406.75 34.57 ;
      RECT 405.02 29.82 405.19 34.57 ;
      RECT 403.46 29.82 403.63 34.57 ;
      RECT 408.92 29.82 409.09 34.57 ;
      RECT 410.68 29.82 410.85 34.57 ;
      RECT 411.96 29.82 412.13 34.57 ;
      RECT 413.485 31.495 413.665 36.23 ;
      RECT 413.485 36.23 432.885 36.41 ;
      RECT 432.705 31.495 432.885 36.23 ;
      RECT 409.8 29.82 409.97 34.57 ;
      RECT 408.14 29.82 408.31 34.57 ;
      RECT 417.635 29.025 418.005 35.105 ;
      RECT 417.565 35.105 418.075 35.435 ;
      RECT 416.805 28.695 418.075 29.025 ;
      RECT 417.295 29.195 417.465 30.245 ;
      RECT 268.785 30.285 268.955 31.335 ;
      RECT 266.885 30.285 267.055 31.335 ;
      RECT 266.265 33.015 266.435 36.03 ;
      RECT 268.785 33.015 268.955 36.03 ;
      RECT 266.885 33.015 267.055 35.725 ;
      RECT 267.835 30.285 268.005 34.755 ;
      RECT 266.885 31.565 267.055 31.895 ;
      RECT 266.265 32.515 266.435 32.845 ;
      RECT 268.785 32.515 268.955 32.845 ;
      RECT 266.885 32.515 267.055 32.845 ;
      RECT 266.265 31.565 266.435 31.895 ;
      RECT 268.785 31.565 268.955 31.895 ;
      RECT 269.48 30.285 269.65 31.795 ;
      RECT 269.48 32.515 269.65 36.025 ;
      RECT 278.7 30.555 281.61 30.725 ;
      RECT 278.9 29.275 281.61 29.445 ;
      RECT 278.595 31.87 281.305 32.04 ;
      RECT 279.81 32.04 280.45 32.08 ;
      RECT 279.81 31.82 280.45 31.87 ;
      RECT 278.595 33.43 281.305 33.6 ;
      RECT 279.81 33.6 280.45 33.645 ;
      RECT 279.81 33.385 280.45 33.43 ;
      RECT 278.205 32.095 278.375 33.375 ;
      RECT 278.18 30.03 278.35 30.5 ;
      RECT 278.175 29.5 278.35 30.03 ;
      RECT 278.595 32.65 281.305 32.82 ;
      RECT 278.685 32.82 279.325 32.865 ;
      RECT 278.685 32.605 279.325 32.65 ;
      RECT 293.715 28.765 293.885 31.995 ;
      RECT 290.545 31.995 293.885 32.165 ;
      RECT 290.545 28.765 290.715 31.785 ;
      RECT 290.545 31.785 290.8 31.995 ;
      RECT 290.545 28.41 293.885 28.765 ;
      RECT 291.345 29.095 292.035 29.405 ;
      RECT 288.755 32.69 288.925 33.49 ;
      RECT 288.285 32.08 288.925 32.25 ;
      RECT 288.755 32.25 288.925 32.41 ;
      RECT 288.755 31.61 288.925 32.08 ;
      RECT 291.345 31.435 292.035 31.665 ;
      RECT 290.955 29.755 291.54 29.925 ;
      RECT 290.955 29.925 291.125 31.38 ;
      RECT 290.955 29.38 291.125 29.755 ;
      RECT 288.755 28.9 288.925 30.78 ;
      RECT 288.395 27.225 288.925 27.395 ;
      RECT 288.755 27.395 288.925 28.62 ;
      RECT 288.755 26.74 288.925 27.225 ;
      RECT 287.525 32.465 288.535 32.635 ;
      RECT 287.525 26.515 288.535 26.685 ;
      RECT 287.525 28.675 288.535 28.845 ;
      RECT 287.525 30.835 288.535 31.005 ;
      RECT 287.525 31.385 288.535 31.555 ;
      RECT 287.525 33.545 288.535 33.715 ;
      RECT 287.525 29.755 288.535 29.925 ;
      RECT 287.525 27.595 288.535 27.765 ;
      RECT 296.83 27.97 297 29.905 ;
      RECT 296.83 26.145 297 26.815 ;
      RECT 293.285 29.04 293.475 31.38 ;
      RECT 292.365 31.435 293.055 31.665 ;
      RECT 292.365 29.095 293.055 29.955 ;
      RECT 297.42 27.65 298.09 27.82 ;
      RECT 297.42 26.87 298.09 27.04 ;
      RECT 297.42 26.09 298.09 26.26 ;
      RECT 297.3 29.96 298.31 30.13 ;
      RECT 297.3 28.2 298.31 28.37 ;
      RECT 297.3 33.48 298.31 33.65 ;
      RECT 297.3 29.08 298.31 29.25 ;
      RECT 297.3 32.6 298.31 32.77 ;
      RECT 297.3 31.72 298.31 31.89 ;
      RECT 297.3 30.84 298.31 31.01 ;
      RECT 300.415 30.405 301.855 30.575 ;
      RECT 301.185 30.1 301.855 30.405 ;
      RECT 300.415 30.575 300.585 31.665 ;
      RECT 300.415 31.84 300.585 33.425 ;
      RECT 298.62 30.185 298.79 33.425 ;
      RECT 298.62 26.87 298.79 27.595 ;
      RECT 300.415 27.955 300.615 28.955 ;
      RECT 300.6 29.235 300.955 30.235 ;
      RECT 300.785 28.885 300.955 29.235 ;
      RECT 300.845 30.84 301.855 31.01 ;
      RECT 300.845 31.72 301.855 31.89 ;
      RECT 300.845 33.48 301.855 33.65 ;
      RECT 300.845 27.18 301.855 27.35 ;
      RECT 301.185 27.73 301.855 27.9 ;
      RECT 301.185 29.01 301.855 29.18 ;
      RECT 300.845 32.6 301.855 32.77 ;
      RECT 300.845 26 301.855 26.17 ;
      RECT 308.155 27.875 309.505 28.045 ;
      RECT 304.315 28.025 307.025 28.195 ;
      RECT 306.665 30.775 308.685 31.525 ;
      RECT 314.415 27.78 315.545 27.95 ;
      RECT 314.415 26.925 314.585 27.78 ;
      RECT 314.875 26.7 315.545 26.87 ;
      RECT 320.06 31.575 321.07 31.745 ;
      RECT 320.06 32.755 321.07 32.925 ;
      RECT 320.025 25.785 320.675 26.115 ;
      RECT 320.025 26.415 320.675 26.745 ;
      RECT 320.025 27.675 320.705 28.005 ;
      RECT 320.025 27.045 320.675 27.375 ;
      RECT 319.45 33.355 322.02 33.525 ;
      RECT 319.45 31.05 319.62 33.355 ;
      RECT 321.85 31.05 322.02 33.355 ;
      RECT 319.45 30.88 322.02 31.05 ;
      RECT 325.735 31.89 325.905 32.56 ;
      RECT 321.32 31.89 321.49 32.56 ;
      RECT 324.475 32.755 325.485 32.925 ;
      RECT 324.475 31.575 325.485 31.745 ;
      RECT 323.85 33.355 326.42 33.525 ;
      RECT 323.85 31.05 324.02 33.355 ;
      RECT 326.25 31.05 326.42 33.355 ;
      RECT 323.85 30.88 326.42 31.05 ;
      RECT 330.025 31.89 330.195 32.56 ;
      RECT 328.765 32.755 329.775 32.925 ;
      RECT 328.765 31.575 329.775 31.745 ;
      RECT 328.425 25.785 329.075 26.115 ;
      RECT 327.395 25.785 328.045 26.115 ;
      RECT 328.16 33.355 330.73 33.525 ;
      RECT 328.16 31.05 328.33 33.355 ;
      RECT 330.56 31.05 330.73 33.355 ;
      RECT 328.16 30.88 330.78 31.05 ;
      RECT 335.705 31.89 335.875 32.56 ;
      RECT 334.445 32.755 335.455 32.925 ;
      RECT 334.445 31.575 335.455 31.745 ;
      RECT 336.21 31.05 336.38 33.355 ;
      RECT 333.81 33.355 336.38 33.525 ;
      RECT 333.81 30.88 336.38 31.05 ;
      RECT 333.81 31.05 333.98 33.355 ;
      RECT 343.615 27.4 344.285 27.9 ;
      RECT 246.745 30.085 247.255 30.115 ;
      RECT 246.745 36.225 248.135 36.525 ;
      RECT 246.745 36.195 247.255 36.225 ;
      RECT 248.575 30.115 248.945 36.195 ;
      RECT 248.505 29.785 249.015 30.115 ;
      RECT 248.505 36.195 249.015 36.525 ;
      RECT 249.995 30.285 250.165 36.045 ;
      RECT 249.385 29.785 249.895 30.115 ;
      RECT 249.385 36.195 249.895 36.525 ;
      RECT 249.455 30.115 249.825 36.195 ;
      RECT 250.265 36.195 251.655 36.525 ;
      RECT 250.265 29.785 251.655 30.115 ;
      RECT 250.335 30.115 250.705 36.195 ;
      RECT 251.215 30.115 251.585 36.195 ;
      RECT 247.355 30.285 247.525 31.895 ;
      RECT 250.875 30.285 251.045 31.895 ;
      RECT 249.115 30.285 249.285 31.895 ;
      RECT 247.355 32.515 247.525 35.725 ;
      RECT 250.875 32.515 251.045 35.725 ;
      RECT 249.115 32.515 249.285 35.725 ;
      RECT 256.8 26.165 256.97 26.835 ;
      RECT 255.24 26.165 255.41 26.835 ;
      RECT 252.005 29.945 252.535 30.115 ;
      RECT 252.025 36.195 252.535 36.525 ;
      RECT 252.025 29.785 252.535 29.945 ;
      RECT 252.095 30.115 252.465 36.195 ;
      RECT 251.755 30.285 251.925 36.03 ;
      RECT 252.635 30.285 252.805 31.895 ;
      RECT 252.635 32.515 252.805 35.725 ;
      RECT 254.065 33.015 254.235 35.725 ;
      RECT 254.945 30.41 255.115 36.045 ;
      RECT 254.065 30.285 254.235 32.105 ;
      RECT 254.405 30.115 254.775 36.195 ;
      RECT 254.335 29.785 254.845 30.115 ;
      RECT 254.325 36.195 254.855 36.845 ;
      RECT 252.975 30.115 253.345 36.195 ;
      RECT 252.905 36.195 253.415 36.525 ;
      RECT 252.885 29.575 253.415 30.115 ;
      RECT 253.585 29.945 254.115 30.115 ;
      RECT 253.585 30.115 253.895 30.26 ;
      RECT 253.515 30.26 253.895 36.03 ;
      RECT 255.825 32.515 255.995 35.725 ;
      RECT 255.825 31.52 255.995 31.895 ;
      RECT 255.285 30.115 255.655 36.195 ;
      RECT 255.215 29.785 255.725 30.115 ;
      RECT 257.925 30.115 258.295 36.195 ;
      RECT 258.805 30.115 259.175 36.195 ;
      RECT 257.71 29.785 259.24 30.115 ;
      RECT 255.215 36.195 259.325 36.525 ;
      RECT 255.825 30.285 255.995 31.35 ;
      RECT 256.705 33.015 256.875 35.725 ;
      RECT 255.47 27.175 256.75 28.305 ;
      RECT 258.325 27.35 262.765 27.52 ;
      RECT 262.04 26.315 262.57 27.35 ;
      RECT 263.755 36.195 264.265 36.22 ;
      RECT 261.115 36.195 261.625 36.22 ;
      RECT 261.185 32.31 261.555 36.195 ;
      RECT 260.92 32.14 261.555 32.31 ;
      RECT 262.945 30.115 263.315 36.195 ;
      RECT 263.825 30.115 264.195 36.195 ;
      RECT 262.065 30.115 262.435 36.195 ;
      RECT 261.995 36.195 263.385 36.22 ;
      RECT 261.115 36.22 264.265 36.525 ;
      RECT 261.185 30.115 261.555 32.14 ;
      RECT 261.115 29.785 264.265 30.115 ;
      RECT 260.305 30.115 260.675 36.195 ;
      RECT 260.235 29.785 260.745 30.115 ;
      RECT 260.235 36.195 260.745 36.525 ;
      RECT 258.1 26.78 258.74 27.04 ;
      RECT 258.1 27.04 258.27 27.1 ;
      RECT 258.1 26.09 258.27 26.78 ;
      RECT 257.585 30.285 257.755 31.335 ;
      RECT 260.225 26.78 260.865 27.04 ;
      RECT 260.46 27.04 260.63 27.1 ;
      RECT 260.46 26.09 260.63 26.78 ;
      RECT 259.345 30.285 259.515 31.335 ;
      RECT 260.845 30.285 261.015 31.335 ;
      RECT 259.605 32.14 260.135 32.31 ;
      RECT 259.965 32.31 260.135 36.03 ;
      RECT 259.965 30.285 260.135 32.14 ;
      RECT 258.465 30.285 258.635 35.725 ;
      RECT 261.11 26.145 261.81 26.405 ;
      RECT 261.64 26.09 261.81 26.145 ;
      RECT 261.64 26.405 261.81 27.1 ;
      RECT 262.82 26.78 263.475 27.04 ;
      RECT 262.82 27.04 262.99 27.1 ;
      RECT 262.82 26.09 262.99 26.78 ;
      RECT 262.605 30.285 262.775 31.335 ;
      RECT 261.725 30.285 261.895 36.03 ;
      RECT 263.045 27.35 263.945 27.52 ;
      RECT 257.585 33.015 257.755 35.725 ;
      RECT 260.845 33.015 261.015 35.725 ;
      RECT 259.345 33.015 259.515 35.725 ;
      RECT 260.845 32.515 261.015 32.845 ;
      RECT 260.845 31.565 261.015 31.895 ;
      RECT 262.605 33.015 262.775 35.725 ;
      RECT 262.605 32.515 262.775 32.845 ;
      RECT 262.605 31.565 262.775 31.895 ;
      RECT 264 26.06 264.53 27.1 ;
      RECT 265.585 29.785 266.095 30.115 ;
      RECT 265.585 36.195 266.095 36.525 ;
      RECT 265.5 35.11 266.03 35.28 ;
      RECT 265.655 35.28 266.025 36.195 ;
      RECT 265.655 30.115 266.025 35.11 ;
      RECT 264.705 29.785 265.215 30.115 ;
      RECT 264.615 32.14 265.145 32.31 ;
      RECT 264.705 36.195 265.215 36.525 ;
      RECT 264.775 32.31 265.145 36.195 ;
      RECT 264.775 30.115 265.145 32.14 ;
      RECT 264.365 30.285 264.535 31.335 ;
      RECT 264.365 33.015 264.535 35.725 ;
      RECT 265.315 30.285 265.485 34.755 ;
      RECT 264.365 31.565 264.535 31.895 ;
      RECT 264.365 32.515 264.535 32.845 ;
      RECT 263.485 30.285 263.655 36.03 ;
      RECT 268.175 30.115 268.545 36.195 ;
      RECT 268.105 29.785 268.615 30.115 ;
      RECT 268.09 36.265 268.62 36.435 ;
      RECT 268.105 36.435 268.615 36.525 ;
      RECT 268.105 36.195 268.615 36.265 ;
      RECT 267.225 36.195 267.735 36.525 ;
      RECT 267.205 29.575 267.735 29.745 ;
      RECT 267.225 29.745 267.735 30.115 ;
      RECT 267.075 32.075 267.665 32.245 ;
      RECT 267.295 32.245 267.665 36.195 ;
      RECT 267.295 30.115 267.665 32.075 ;
      RECT 266.265 30.285 266.435 31.335 ;
      RECT 221.56 32.785 222.45 33.6 ;
      RECT 221.56 32.71 223.475 32.785 ;
      RECT 221.58 31.765 223.475 32.71 ;
      RECT 225.865 31.735 226.035 32.855 ;
      RECT 228.975 31.735 229.145 32.855 ;
      RECT 231.535 31.735 232.945 32.785 ;
      RECT 221.56 31.595 224.175 31.765 ;
      RECT 230.835 31.535 232.945 31.735 ;
      RECT 228.975 31.535 230.085 31.735 ;
      RECT 221.58 31.485 224.175 31.595 ;
      RECT 224.925 31.485 226.035 31.735 ;
      RECT 221.58 30.145 226.035 31.485 ;
      RECT 228.975 30.145 232.945 31.535 ;
      RECT 229.555 29.405 232.945 30.145 ;
      RECT 221.58 29.19 225.455 30.145 ;
      RECT 229.555 29.19 270.96 29.405 ;
      RECT 221.58 28.555 270.96 29.19 ;
      RECT 220.655 32.125 220.825 32.135 ;
      RECT 220.105 32.135 220.825 33.645 ;
      RECT 218.685 32.135 218.855 33.645 ;
      RECT 219.765 31.635 219.935 35.825 ;
      RECT 218.345 31.965 218.515 35.495 ;
      RECT 218.345 31.635 219.195 31.965 ;
      RECT 218.345 35.495 219.195 35.825 ;
      RECT 219.025 31.965 219.195 35.495 ;
      RECT 217.975 31.635 218.145 35.995 ;
      RECT 217.945 35.995 219.565 36.165 ;
      RECT 219.395 31.635 219.565 35.995 ;
      RECT 217.605 31.635 217.775 35.825 ;
      RECT 228.055 33.255 230.085 33.425 ;
      RECT 224.925 33.255 226.615 33.425 ;
      RECT 226.965 33.255 227.495 33.425 ;
      RECT 227.145 30.145 227.315 33.255 ;
      RECT 227.145 33.425 227.315 34.915 ;
      RECT 227.485 32.885 228.015 33.055 ;
      RECT 227.695 33.055 227.865 34.915 ;
      RECT 227.695 30.145 227.865 32.885 ;
      RECT 224.175 32.165 224.755 32.335 ;
      RECT 224.585 31.775 224.755 32.165 ;
      RECT 224.585 32.335 224.755 34.915 ;
      RECT 228.06 29.42 228.73 29.59 ;
      RECT 228.14 29.59 228.67 30.115 ;
      RECT 226.3 29.425 226.97 29.595 ;
      RECT 226.38 29.595 226.91 29.745 ;
      RECT 230.255 31.775 230.425 34.915 ;
      RECT 233.98 31.565 235.205 31.735 ;
      RECT 234.34 31.735 235.205 31.795 ;
      RECT 234.34 30.285 235.205 31.565 ;
      RECT 235.035 31.795 235.205 31.895 ;
      RECT 234.34 35.725 234.51 36.025 ;
      RECT 234.34 32.515 235.205 35.725 ;
      RECT 236.795 30.285 236.965 31.895 ;
      RECT 236.795 32.515 236.965 35.725 ;
      RECT 237.135 30.115 237.505 36.195 ;
      RECT 236.255 30.115 236.625 36.195 ;
      RECT 237.065 30.085 237.575 30.115 ;
      RECT 236.185 29.785 237.575 30.085 ;
      RECT 236.185 30.085 236.695 30.115 ;
      RECT 237.07 36.195 237.58 36.225 ;
      RECT 236.185 36.225 237.58 36.525 ;
      RECT 236.185 36.195 236.695 36.225 ;
      RECT 235.305 29.785 235.815 30.115 ;
      RECT 235.375 30.115 235.745 36.195 ;
      RECT 235.305 36.195 235.815 36.525 ;
      RECT 235.915 30.285 236.085 36.025 ;
      RECT 238.555 30.285 238.725 31.895 ;
      RECT 238.555 32.515 238.725 35.725 ;
      RECT 238.015 30.115 238.385 36.195 ;
      RECT 238.895 30.115 239.265 36.195 ;
      RECT 237.945 30.085 238.455 30.115 ;
      RECT 237.945 29.785 239.335 30.085 ;
      RECT 238.825 30.085 239.335 30.115 ;
      RECT 237.945 36.195 238.455 36.225 ;
      RECT 237.945 36.225 239.335 36.525 ;
      RECT 238.825 36.195 239.335 36.225 ;
      RECT 239.775 30.115 240.145 36.195 ;
      RECT 240.655 30.115 241.025 36.195 ;
      RECT 239.705 30.085 240.215 30.115 ;
      RECT 239.705 36.195 240.215 36.225 ;
      RECT 239.705 29.785 241.095 30.085 ;
      RECT 240.585 30.085 241.095 30.115 ;
      RECT 239.705 36.225 241.095 36.525 ;
      RECT 240.585 36.195 241.095 36.225 ;
      RECT 239.435 30.285 239.605 36.025 ;
      RECT 237.675 30.285 237.845 36.025 ;
      RECT 240.285 27.55 245.035 27.72 ;
      RECT 240.285 26.47 245.035 26.64 ;
      RECT 242.415 30.115 242.785 36.195 ;
      RECT 242.345 29.785 242.855 30.115 ;
      RECT 242.345 36.195 242.855 36.525 ;
      RECT 242.955 30.285 243.125 36.025 ;
      RECT 241.195 30.285 241.365 36.025 ;
      RECT 244.715 30.285 244.885 36.025 ;
      RECT 243.295 30.115 243.665 36.195 ;
      RECT 244.175 30.115 244.545 36.195 ;
      RECT 243.225 30.085 243.735 30.115 ;
      RECT 243.225 36.195 243.735 36.225 ;
      RECT 243.225 29.785 244.615 30.085 ;
      RECT 244.105 30.085 244.615 30.115 ;
      RECT 243.225 36.225 244.62 36.525 ;
      RECT 244.11 36.195 244.62 36.225 ;
      RECT 241.535 30.115 241.905 36.195 ;
      RECT 241.465 29.785 241.975 30.115 ;
      RECT 241.465 36.195 241.975 36.525 ;
      RECT 245.055 30.115 245.425 36.195 ;
      RECT 245.935 30.115 246.305 36.195 ;
      RECT 244.985 30.085 245.495 30.115 ;
      RECT 244.985 36.195 245.495 36.225 ;
      RECT 244.985 29.785 246.375 30.085 ;
      RECT 245.865 30.085 246.375 30.115 ;
      RECT 244.985 36.225 246.375 36.525 ;
      RECT 245.865 36.195 246.375 36.225 ;
      RECT 242.075 30.285 242.245 31.895 ;
      RECT 240.315 30.285 240.485 31.895 ;
      RECT 245.595 30.285 245.765 31.895 ;
      RECT 243.835 30.285 244.005 31.895 ;
      RECT 242.075 32.515 242.245 35.725 ;
      RECT 240.315 32.515 240.485 35.725 ;
      RECT 245.595 32.515 245.765 35.725 ;
      RECT 243.835 32.515 244.005 35.725 ;
      RECT 246.475 30.285 246.645 36.025 ;
      RECT 248.235 30.285 248.405 36.025 ;
      RECT 247.695 30.115 248.065 36.195 ;
      RECT 246.815 30.115 247.185 36.195 ;
      RECT 247.625 30.085 248.135 30.115 ;
      RECT 247.625 36.195 248.135 36.225 ;
      RECT 246.745 29.785 248.135 30.085 ;
      RECT 142.75 36.195 143.26 36.225 ;
      RECT 141.87 36.225 143.26 36.525 ;
      RECT 141.87 36.195 142.38 36.225 ;
      RECT 141.6 30.285 141.77 36.025 ;
      RECT 143.36 30.285 143.53 36.025 ;
      RECT 144.24 30.285 144.41 31.895 ;
      RECT 144.24 32.515 144.41 35.725 ;
      RECT 146 30.285 146.17 31.895 ;
      RECT 146 32.515 146.17 35.725 ;
      RECT 145.46 30.115 145.83 36.195 ;
      RECT 146.34 30.115 146.71 36.195 ;
      RECT 145.39 30.085 145.9 30.115 ;
      RECT 145.39 29.785 146.78 30.085 ;
      RECT 146.27 30.085 146.78 30.115 ;
      RECT 145.385 36.195 145.895 36.225 ;
      RECT 145.385 36.225 146.78 36.525 ;
      RECT 146.27 36.195 146.78 36.225 ;
      RECT 145.12 30.285 145.29 36.025 ;
      RECT 147.15 29.785 147.66 30.115 ;
      RECT 147.22 30.115 147.59 36.195 ;
      RECT 147.15 36.195 147.66 36.525 ;
      RECT 146.88 30.285 147.05 36.025 ;
      RECT 147.76 30.285 147.93 31.895 ;
      RECT 147.76 32.515 147.93 35.725 ;
      RECT 148.03 29.785 148.54 30.115 ;
      RECT 148.1 30.115 148.47 36.195 ;
      RECT 148.03 36.195 148.54 36.525 ;
      RECT 149.52 30.285 149.69 31.895 ;
      RECT 149.52 32.515 149.69 35.725 ;
      RECT 150.74 30.115 151.11 36.195 ;
      RECT 151.62 30.115 151.99 36.195 ;
      RECT 150.67 30.085 151.18 30.115 ;
      RECT 150.67 36.195 151.18 36.225 ;
      RECT 150.67 29.785 152.06 30.085 ;
      RECT 151.55 30.085 152.06 30.115 ;
      RECT 150.67 36.225 152.06 36.525 ;
      RECT 151.55 36.195 152.06 36.225 ;
      RECT 149.86 30.115 150.23 36.195 ;
      RECT 148.98 30.115 149.35 36.195 ;
      RECT 149.79 30.085 150.3 30.115 ;
      RECT 148.91 29.785 150.3 30.085 ;
      RECT 148.91 30.085 149.42 30.115 ;
      RECT 149.79 36.195 150.3 36.225 ;
      RECT 148.91 36.225 150.3 36.525 ;
      RECT 148.91 36.195 149.42 36.225 ;
      RECT 148.64 30.285 148.81 36.025 ;
      RECT 150.4 30.285 150.57 36.025 ;
      RECT 151.28 30.285 151.45 31.895 ;
      RECT 151.28 32.515 151.45 35.725 ;
      RECT 153.04 30.285 153.21 31.895 ;
      RECT 153.04 32.515 153.21 35.725 ;
      RECT 152.5 30.115 152.87 36.195 ;
      RECT 153.38 30.115 153.75 36.195 ;
      RECT 152.43 30.085 152.94 30.115 ;
      RECT 152.43 29.785 153.82 30.085 ;
      RECT 153.31 30.085 153.82 30.115 ;
      RECT 152.425 36.195 152.935 36.225 ;
      RECT 152.425 36.225 153.82 36.525 ;
      RECT 153.31 36.195 153.82 36.225 ;
      RECT 152.16 30.285 152.33 36.025 ;
      RECT 157.06 35.945 168.445 36.455 ;
      RECT 167.555 35.565 168.445 35.945 ;
      RECT 167.575 33.6 168.425 35.565 ;
      RECT 157.06 32.785 157.57 35.945 ;
      RECT 167.555 32.785 168.445 33.6 ;
      RECT 166.53 32.71 168.445 32.785 ;
      RECT 166.53 31.765 168.425 32.71 ;
      RECT 160.86 31.735 161.03 32.855 ;
      RECT 163.97 31.735 164.14 32.855 ;
      RECT 157.06 31.735 158.47 32.785 ;
      RECT 165.83 31.595 168.445 31.765 ;
      RECT 157.06 31.535 159.17 31.735 ;
      RECT 159.92 31.535 161.03 31.735 ;
      RECT 163.97 31.485 165.08 31.735 ;
      RECT 165.83 31.485 168.425 31.595 ;
      RECT 163.97 30.145 168.425 31.485 ;
      RECT 157.06 30.145 161.03 31.535 ;
      RECT 157.06 29.405 160.45 30.145 ;
      RECT 164.55 29.19 168.425 30.145 ;
      RECT 119.045 29.19 160.45 29.405 ;
      RECT 119.045 28.555 168.425 29.19 ;
      RECT 154.8 31.565 156.025 31.735 ;
      RECT 154.8 31.795 154.97 31.895 ;
      RECT 154.8 31.735 155.665 31.795 ;
      RECT 154.8 30.285 155.665 31.565 ;
      RECT 155.495 35.725 155.665 36.025 ;
      RECT 154.8 32.515 155.665 35.725 ;
      RECT 154.19 29.785 154.7 30.115 ;
      RECT 154.26 30.115 154.63 36.195 ;
      RECT 154.19 36.195 154.7 36.525 ;
      RECT 153.92 30.285 154.09 36.025 ;
      RECT 159.92 33.255 161.95 33.425 ;
      RECT 163.39 33.255 165.08 33.425 ;
      RECT 162.51 33.255 163.04 33.425 ;
      RECT 162.69 30.145 162.86 33.255 ;
      RECT 162.69 33.425 162.86 34.915 ;
      RECT 161.99 32.885 162.52 33.055 ;
      RECT 162.14 33.055 162.31 34.915 ;
      RECT 162.14 30.145 162.31 32.885 ;
      RECT 159.58 31.775 159.75 34.915 ;
      RECT 161.275 29.42 161.945 29.59 ;
      RECT 161.335 29.59 161.865 30.115 ;
      RECT 163.035 29.425 163.705 29.595 ;
      RECT 163.095 29.595 163.625 29.745 ;
      RECT 169.18 32.125 169.35 32.135 ;
      RECT 169.18 32.135 169.9 33.645 ;
      RECT 165.25 32.165 165.83 32.335 ;
      RECT 165.25 31.775 165.42 32.165 ;
      RECT 165.25 32.335 165.42 34.915 ;
      RECT 170.07 31.635 170.24 35.825 ;
      RECT 170.44 31.635 170.61 35.995 ;
      RECT 170.44 35.995 172.06 36.165 ;
      RECT 171.86 31.635 172.03 35.995 ;
      RECT 171.15 32.135 171.32 33.645 ;
      RECT 173.12 32.125 173.29 32.135 ;
      RECT 172.57 32.135 173.29 33.645 ;
      RECT 170.81 31.965 170.98 35.495 ;
      RECT 170.81 31.635 171.66 31.965 ;
      RECT 170.81 35.495 171.66 35.825 ;
      RECT 171.49 31.965 171.66 35.495 ;
      RECT 172.23 31.635 172.4 35.825 ;
      RECT 216.715 32.125 216.885 32.135 ;
      RECT 216.715 32.135 217.435 33.645 ;
      RECT 221.56 35.945 232.945 36.455 ;
      RECT 221.56 35.565 222.45 35.945 ;
      RECT 221.58 33.6 222.43 35.565 ;
      RECT 232.435 32.785 232.945 35.945 ;
      RECT 122.95 32.515 123.12 32.845 ;
      RECT 123.57 31.565 123.74 31.895 ;
      RECT 121.05 31.565 121.22 31.895 ;
      RECT 120.355 30.285 120.525 31.795 ;
      RECT 120.355 32.515 120.525 36.025 ;
      RECT 124.79 29.785 125.3 30.115 ;
      RECT 124.86 32.14 125.39 32.31 ;
      RECT 124.79 36.195 125.3 36.525 ;
      RECT 124.86 32.31 125.23 36.195 ;
      RECT 124.86 30.115 125.23 32.14 ;
      RECT 127.24 27.35 131.68 27.52 ;
      RECT 127.435 26.315 127.965 27.35 ;
      RECT 126.35 30.285 126.52 36.03 ;
      RECT 128.11 30.285 128.28 36.03 ;
      RECT 125.74 36.195 126.25 36.22 ;
      RECT 128.38 36.195 128.89 36.22 ;
      RECT 128.45 32.14 129.085 32.31 ;
      RECT 128.45 30.115 128.82 32.14 ;
      RECT 125.81 30.115 126.18 36.195 ;
      RECT 126.69 30.115 127.06 36.195 ;
      RECT 127.57 30.115 127.94 36.195 ;
      RECT 126.62 36.195 128.01 36.22 ;
      RECT 125.74 29.785 128.89 30.115 ;
      RECT 125.74 36.22 128.89 36.525 ;
      RECT 128.45 32.31 128.82 36.195 ;
      RECT 129.87 32.14 130.4 32.31 ;
      RECT 129.87 32.31 130.04 36.03 ;
      RECT 129.87 30.285 130.04 32.14 ;
      RECT 129.33 30.115 129.7 36.195 ;
      RECT 129.26 29.785 129.77 30.115 ;
      RECT 129.26 36.195 129.77 36.525 ;
      RECT 125.47 30.285 125.64 31.335 ;
      RECT 124.52 30.285 124.69 34.755 ;
      RECT 125.475 26.06 126.005 27.1 ;
      RECT 126.06 27.35 126.96 27.52 ;
      RECT 126.53 26.78 127.185 27.04 ;
      RECT 127.015 27.04 127.185 27.1 ;
      RECT 127.015 26.09 127.185 26.78 ;
      RECT 128.195 26.145 128.895 26.405 ;
      RECT 128.195 26.405 128.365 27.1 ;
      RECT 128.195 26.09 128.365 26.145 ;
      RECT 127.23 30.285 127.4 31.335 ;
      RECT 129.14 26.78 129.78 27.04 ;
      RECT 129.375 27.04 129.545 27.1 ;
      RECT 129.375 26.09 129.545 26.78 ;
      RECT 128.99 30.285 129.16 31.335 ;
      RECT 125.47 33.015 125.64 35.725 ;
      RECT 125.47 31.565 125.64 31.895 ;
      RECT 125.47 32.515 125.64 32.845 ;
      RECT 127.23 33.015 127.4 35.725 ;
      RECT 127.23 32.515 127.4 32.845 ;
      RECT 127.23 31.565 127.4 31.895 ;
      RECT 128.99 33.015 129.16 35.725 ;
      RECT 128.99 32.515 129.16 32.845 ;
      RECT 128.99 31.565 129.16 31.895 ;
      RECT 131.265 26.78 131.905 27.04 ;
      RECT 131.735 27.04 131.905 27.1 ;
      RECT 131.735 26.09 131.905 26.78 ;
      RECT 133.035 26.165 133.205 26.835 ;
      RECT 130.83 30.115 131.2 36.195 ;
      RECT 130.765 29.785 132.295 30.115 ;
      RECT 131.71 30.115 132.08 36.195 ;
      RECT 134.35 30.115 134.72 36.195 ;
      RECT 134.28 29.785 134.79 30.115 ;
      RECT 130.68 36.195 134.79 36.525 ;
      RECT 132.25 30.285 132.42 31.335 ;
      RECT 130.49 30.285 130.66 31.335 ;
      RECT 130.49 33.015 130.66 35.725 ;
      RECT 131.37 30.285 131.54 35.725 ;
      RECT 132.25 33.015 132.42 35.725 ;
      RECT 133.13 33.015 133.3 35.725 ;
      RECT 134.01 32.515 134.18 35.725 ;
      RECT 134.595 26.165 134.765 26.835 ;
      RECT 135.77 33.015 135.94 35.725 ;
      RECT 134.01 31.52 134.18 31.895 ;
      RECT 135.77 30.285 135.94 32.105 ;
      RECT 134.89 30.41 135.06 36.045 ;
      RECT 135.23 30.115 135.6 36.195 ;
      RECT 135.16 29.785 135.67 30.115 ;
      RECT 135.15 36.195 135.68 36.845 ;
      RECT 134.01 30.285 134.18 31.35 ;
      RECT 133.255 27.175 134.535 28.305 ;
      RECT 141.06 30.115 141.43 36.195 ;
      RECT 140.99 29.785 141.5 30.115 ;
      RECT 140.99 36.195 141.5 36.525 ;
      RECT 139.84 30.285 140.01 36.045 ;
      RECT 138.08 30.285 138.25 36.03 ;
      RECT 140.11 29.785 140.62 30.115 ;
      RECT 140.11 36.195 140.62 36.525 ;
      RECT 140.18 30.115 140.55 36.195 ;
      RECT 138.35 36.195 139.74 36.525 ;
      RECT 138.35 29.785 139.74 30.115 ;
      RECT 139.3 30.115 139.67 36.195 ;
      RECT 138.42 30.115 138.79 36.195 ;
      RECT 137.47 29.945 138 30.115 ;
      RECT 137.47 36.195 137.98 36.525 ;
      RECT 137.47 29.785 137.98 29.945 ;
      RECT 137.54 30.115 137.91 36.195 ;
      RECT 135.89 29.945 136.42 30.115 ;
      RECT 136.11 30.115 136.42 30.26 ;
      RECT 136.11 30.26 136.49 36.03 ;
      RECT 136.66 30.115 137.03 36.195 ;
      RECT 136.59 36.195 137.1 36.525 ;
      RECT 136.59 29.575 137.12 30.115 ;
      RECT 137.2 30.285 137.37 31.895 ;
      RECT 138.96 30.285 139.13 31.895 ;
      RECT 140.72 30.285 140.89 31.895 ;
      RECT 137.2 32.515 137.37 35.725 ;
      RECT 138.96 32.515 139.13 35.725 ;
      RECT 140.72 32.515 140.89 35.725 ;
      RECT 144.97 27.55 149.72 27.72 ;
      RECT 144.97 26.47 149.72 26.64 ;
      RECT 142.48 30.285 142.65 31.895 ;
      RECT 142.48 32.515 142.65 35.725 ;
      RECT 143.7 30.115 144.07 36.195 ;
      RECT 144.58 30.115 144.95 36.195 ;
      RECT 143.63 30.085 144.14 30.115 ;
      RECT 143.63 36.195 144.14 36.225 ;
      RECT 143.63 29.785 145.02 30.085 ;
      RECT 144.51 30.085 145.02 30.115 ;
      RECT 143.63 36.225 145.02 36.525 ;
      RECT 144.51 36.195 145.02 36.225 ;
      RECT 142.82 30.115 143.19 36.195 ;
      RECT 141.94 30.115 142.31 36.195 ;
      RECT 142.75 30.085 143.26 30.115 ;
      RECT 141.87 29.785 143.26 30.085 ;
      RECT 141.87 30.085 142.38 30.115 ;
      RECT 59.275 31.05 59.445 33.355 ;
      RECT 61.675 31.05 61.845 33.355 ;
      RECT 59.225 30.88 61.845 31.05 ;
      RECT 64.1 31.89 64.27 32.56 ;
      RECT 64.52 32.755 65.53 32.925 ;
      RECT 64.52 31.575 65.53 31.745 ;
      RECT 60.93 25.785 61.58 26.115 ;
      RECT 61.96 25.785 62.61 26.115 ;
      RECT 63.585 33.355 66.155 33.525 ;
      RECT 63.585 31.05 63.755 33.355 ;
      RECT 65.985 31.05 66.155 33.355 ;
      RECT 63.585 30.88 66.155 31.05 ;
      RECT 68.515 31.89 68.685 32.56 ;
      RECT 68.935 32.755 69.945 32.925 ;
      RECT 68.935 31.575 69.945 31.745 ;
      RECT 69.33 25.785 69.98 26.115 ;
      RECT 69.33 26.415 69.98 26.745 ;
      RECT 69.3 27.675 69.98 28.005 ;
      RECT 69.33 27.045 69.98 27.375 ;
      RECT 67.985 33.355 70.555 33.525 ;
      RECT 67.985 31.05 68.155 33.355 ;
      RECT 70.385 31.05 70.555 33.355 ;
      RECT 67.985 30.88 70.555 31.05 ;
      RECT 74.46 27.78 75.59 27.95 ;
      RECT 75.42 26.925 75.59 27.78 ;
      RECT 74.46 26.7 75.13 26.87 ;
      RECT 80.5 27.875 81.85 28.045 ;
      RECT 82.98 28.025 85.69 28.195 ;
      RECT 81.32 30.775 83.34 31.525 ;
      RECT 88.15 30.405 89.59 30.575 ;
      RECT 88.15 30.1 88.82 30.405 ;
      RECT 89.42 30.575 89.59 31.665 ;
      RECT 89.42 31.84 89.59 33.425 ;
      RECT 89.39 27.955 89.59 28.955 ;
      RECT 89.05 29.235 89.405 30.235 ;
      RECT 89.05 28.885 89.22 29.235 ;
      RECT 88.15 30.84 89.16 31.01 ;
      RECT 88.15 31.72 89.16 31.89 ;
      RECT 88.15 33.48 89.16 33.65 ;
      RECT 88.15 27.18 89.16 27.35 ;
      RECT 88.15 27.73 88.82 27.9 ;
      RECT 88.15 29.01 88.82 29.18 ;
      RECT 88.15 32.6 89.16 32.77 ;
      RECT 88.15 26 89.16 26.17 ;
      RECT 91.215 30.185 91.385 33.425 ;
      RECT 93.005 27.97 93.175 29.905 ;
      RECT 91.215 26.87 91.385 27.595 ;
      RECT 93.005 26.145 93.175 26.815 ;
      RECT 91.915 27.65 92.585 27.82 ;
      RECT 91.915 26.87 92.585 27.04 ;
      RECT 91.915 26.09 92.585 26.26 ;
      RECT 91.695 33.48 92.705 33.65 ;
      RECT 91.695 29.96 92.705 30.13 ;
      RECT 91.695 28.2 92.705 28.37 ;
      RECT 91.695 29.08 92.705 29.25 ;
      RECT 91.695 32.6 92.705 32.77 ;
      RECT 91.695 31.72 92.705 31.89 ;
      RECT 91.695 30.84 92.705 31.01 ;
      RECT 96.53 29.04 96.72 31.38 ;
      RECT 96.12 28.765 96.29 31.995 ;
      RECT 96.12 31.995 99.46 32.165 ;
      RECT 99.29 28.765 99.46 31.785 ;
      RECT 99.205 31.785 99.46 31.995 ;
      RECT 96.12 28.41 99.46 28.765 ;
      RECT 97.97 29.095 98.66 29.405 ;
      RECT 96.95 31.435 97.64 31.665 ;
      RECT 97.97 31.435 98.66 31.665 ;
      RECT 98.465 29.755 99.05 29.925 ;
      RECT 98.88 29.925 99.05 31.38 ;
      RECT 98.88 29.38 99.05 29.755 ;
      RECT 96.95 29.095 97.64 29.955 ;
      RECT 101.08 32.69 101.25 33.49 ;
      RECT 101.08 32.08 101.72 32.25 ;
      RECT 101.08 32.25 101.25 32.41 ;
      RECT 101.08 31.61 101.25 32.08 ;
      RECT 101.08 28.9 101.25 30.78 ;
      RECT 101.08 27.225 101.61 27.395 ;
      RECT 101.08 27.395 101.25 28.62 ;
      RECT 101.08 26.74 101.25 27.225 ;
      RECT 101.47 28.675 102.48 28.845 ;
      RECT 101.47 30.835 102.48 31.005 ;
      RECT 101.47 31.385 102.48 31.555 ;
      RECT 101.47 32.465 102.48 32.635 ;
      RECT 101.47 33.545 102.48 33.715 ;
      RECT 101.47 26.515 102.48 26.685 ;
      RECT 101.47 29.755 102.48 29.925 ;
      RECT 101.47 27.595 102.48 27.765 ;
      RECT 108.395 30.555 111.305 30.725 ;
      RECT 108.395 29.275 111.105 29.445 ;
      RECT 108.7 33.43 111.41 33.6 ;
      RECT 109.555 33.6 110.195 33.645 ;
      RECT 109.555 33.385 110.195 33.43 ;
      RECT 108.7 31.87 111.41 32.04 ;
      RECT 109.555 32.04 110.195 32.08 ;
      RECT 109.555 31.82 110.195 31.87 ;
      RECT 111.63 32.095 111.8 33.375 ;
      RECT 111.655 30.03 111.825 30.5 ;
      RECT 111.655 29.5 111.83 30.03 ;
      RECT 108.7 32.65 111.41 32.82 ;
      RECT 110.68 32.82 111.32 32.865 ;
      RECT 110.68 32.605 111.32 32.65 ;
      RECT 123.91 29.785 124.42 30.115 ;
      RECT 123.91 36.195 124.42 36.525 ;
      RECT 123.975 35.11 124.505 35.28 ;
      RECT 123.98 35.28 124.35 36.195 ;
      RECT 123.98 30.115 124.35 35.11 ;
      RECT 121.46 30.115 121.83 36.195 ;
      RECT 121.39 29.785 121.9 30.115 ;
      RECT 121.385 36.265 121.915 36.435 ;
      RECT 121.39 36.435 121.9 36.525 ;
      RECT 121.39 36.195 121.9 36.265 ;
      RECT 122.27 36.195 122.78 36.525 ;
      RECT 122.27 29.575 122.8 29.745 ;
      RECT 122.27 29.745 122.78 30.115 ;
      RECT 122.34 32.075 122.93 32.245 ;
      RECT 122.34 32.245 122.71 36.195 ;
      RECT 122.34 30.115 122.71 32.075 ;
      RECT 123.57 30.285 123.74 31.335 ;
      RECT 121.05 30.285 121.22 31.335 ;
      RECT 122.95 30.285 123.12 31.335 ;
      RECT 123.57 33.015 123.74 36.03 ;
      RECT 121.05 33.015 121.22 36.03 ;
      RECT 122.95 33.015 123.12 35.725 ;
      RECT 122 30.285 122.17 34.755 ;
      RECT 122.95 31.565 123.12 31.895 ;
      RECT 123.57 32.515 123.74 32.845 ;
      RECT 121.05 32.515 121.22 32.845 ;
      RECT 442.595 21.835 442.765 22.935 ;
      RECT 442.595 23.605 442.81 23.66 ;
      RECT 442.56 22.935 442.81 23.605 ;
      RECT 442.64 24.35 442.945 27.06 ;
      RECT 442.64 23.66 442.81 24.35 ;
      RECT 442.595 20.825 442.79 21.835 ;
      RECT 437.195 24.145 437.365 24.375 ;
      RECT 437.08 24.375 437.365 27.085 ;
      RECT 437.485 22.6 438.835 22.77 ;
      RECT 437.585 22.57 438.835 22.6 ;
      RECT 439.225 23.71 439.755 23.88 ;
      RECT 439.585 27.23 443.825 27.4 ;
      RECT 443.08 23.78 443.825 23.95 ;
      RECT 443.15 23.71 443.68 23.78 ;
      RECT 439.585 23.88 439.755 27.23 ;
      RECT 443.655 23.95 443.825 27.23 ;
      RECT 438.305 27.655 441.84 27.905 ;
      RECT 438.305 25.395 438.835 27.655 ;
      RECT 439.005 24.37 439.175 27.37 ;
      RECT 437.66 24.395 437.83 27.475 ;
      RECT 441.1 23.71 441.63 23.88 ;
      RECT 441.28 22.935 441.45 23.71 ;
      RECT 440.925 24.08 441.185 27.06 ;
      RECT 441.8 23.78 442.47 23.95 ;
      RECT 441.86 23.04 442.39 23.21 ;
      RECT 441.895 23.21 442.39 23.78 ;
      RECT 441.895 23.95 442.065 27.06 ;
      RECT 440.465 24.08 440.725 27.06 ;
      RECT 443.84 23.21 444.01 23.605 ;
      RECT 443.84 22.935 444.01 23.04 ;
      RECT 442.98 23.04 444.01 23.21 ;
      RECT 443.735 22.155 444.27 22.73 ;
      RECT 443.695 19.94 443.865 20.61 ;
      RECT 443.67 19.075 443.84 19.77 ;
      RECT 443.54 20.825 443.71 21.835 ;
      RECT 456.34 20.74 456.875 21.42 ;
      RECT 454.925 20.39 456.875 20.74 ;
      RECT 455.65 20.925 455.82 21.455 ;
      RECT 454.615 21.09 455.07 21.64 ;
      RECT 454.615 21.64 456.545 21.81 ;
      RECT 457.22 18.195 457.94 19.445 ;
      RECT 457.1 21.04 458.515 21.34 ;
      RECT 464.155 20.655 464.325 23.365 ;
      RECT 461.62 20.655 462.57 21.905 ;
      RECT 462.055 21.905 462.565 23.425 ;
      RECT 463.275 20.655 463.445 23.365 ;
      RECT 462.415 23.915 464.1 24.085 ;
      RECT 12.7 27.93 14.72 28.68 ;
      RECT 18.92 31.065 19.09 33.775 ;
      RECT 17.36 31.065 17.53 33.775 ;
      RECT 16.08 31.065 16.25 33.775 ;
      RECT 18.14 31.065 18.31 33.775 ;
      RECT 15.85 53.095 24.335 53.265 ;
      RECT 24.04 52.565 24.335 53.095 ;
      RECT 24.165 51.935 24.335 52.565 ;
      RECT 15.85 42.71 16.02 53.095 ;
      RECT 15.685 41.775 16.02 42.71 ;
      RECT 18.33 41.775 19.34 53.095 ;
      RECT 24.04 41.775 24.335 51.935 ;
      RECT 14.665 41.605 24.335 41.775 ;
      RECT 14.665 41.57 21.1 41.605 ;
      RECT 24.04 39.135 24.335 41.605 ;
      RECT 20.335 38.545 21.1 41.57 ;
      RECT 22.69 41.13 22.86 41.605 ;
      RECT 22.69 38.545 22.86 39.04 ;
      RECT 22.685 39.04 22.86 41.13 ;
      RECT 24.165 37.025 24.335 39.135 ;
      RECT 20.335 36.775 20.505 38.545 ;
      RECT 14.665 36.4 14.835 41.57 ;
      RECT 20.335 36.4 21.1 36.775 ;
      RECT 14.665 35.05 21.1 36.4 ;
      RECT 20.335 34.025 21.1 35.05 ;
      RECT 20.335 32.905 20.505 34.025 ;
      RECT 24.04 30.35 24.335 37.025 ;
      RECT 24.165 29.845 24.335 30.35 ;
      RECT 14.665 29.88 14.835 35.05 ;
      RECT 20.335 29.88 21.1 32.905 ;
      RECT 14.665 29.845 21.1 29.88 ;
      RECT 14.665 29.675 24.335 29.845 ;
      RECT 15.6 30.645 19.57 30.815 ;
      RECT 15.6 30.815 15.77 34.085 ;
      RECT 19.4 30.815 19.57 34.085 ;
      RECT 23.57 30.195 23.74 32.905 ;
      RECT 22.69 30.195 22.86 32.905 ;
      RECT 24.535 29.49 24.705 30.665 ;
      RECT 24.535 30.665 26.15 30.835 ;
      RECT 22.545 29.32 24.705 29.49 ;
      RECT 24.895 30.295 26.15 30.465 ;
      RECT 24.895 29.15 25.065 30.295 ;
      RECT 21.755 28.98 25.065 29.15 ;
      RECT 21.755 29.15 22.285 29.49 ;
      RECT 21.745 30.195 21.98 33.065 ;
      RECT 22.915 33.455 23.585 33.625 ;
      RECT 21.155 33.455 22.635 33.625 ;
      RECT 28.1 32.665 28.27 33.335 ;
      RECT 28.1 31.485 28.27 32.155 ;
      RECT 27.475 30.425 27.645 36.58 ;
      RECT 51.3 30.425 51.47 36.59 ;
      RECT 27.475 30.255 51.47 30.425 ;
      RECT 49.99 36.75 51.47 36.76 ;
      RECT 27.475 36.59 51.47 36.75 ;
      RECT 27.475 36.58 50.1 36.59 ;
      RECT 32.12 27.305 34.83 27.475 ;
      RECT 39.42 27.305 42.13 27.475 ;
      RECT 38.81 32.665 38.98 33.335 ;
      RECT 38.81 31.485 38.98 32.155 ;
      RECT 39.69 32.665 39.86 33.335 ;
      RECT 39.69 31.485 39.86 32.155 ;
      RECT 44.54 27.4 45.21 27.9 ;
      RECT 45.72 27.4 46.39 27.9 ;
      RECT 48.16 25.785 48.81 26.115 ;
      RECT 48.16 27.045 48.81 27.375 ;
      RECT 48.16 26.415 48.81 26.745 ;
      RECT 48.16 27.675 48.81 28.005 ;
      RECT 54.13 31.89 54.3 32.56 ;
      RECT 50.4 32.665 50.57 33.335 ;
      RECT 50.4 31.485 50.57 32.155 ;
      RECT 54.55 32.755 55.56 32.925 ;
      RECT 54.55 31.575 55.56 31.745 ;
      RECT 53.625 31.05 53.795 33.355 ;
      RECT 53.625 33.355 56.195 33.525 ;
      RECT 53.625 30.88 56.195 31.05 ;
      RECT 56.025 31.05 56.195 33.355 ;
      RECT 59.81 31.89 59.98 32.56 ;
      RECT 60.23 32.755 61.24 32.925 ;
      RECT 60.23 31.575 61.24 31.745 ;
      RECT 59.275 33.355 61.845 33.525 ;
      RECT 424.14 23.04 425.17 23.21 ;
      RECT 423.88 22.155 424.415 22.73 ;
      RECT 424.325 27.23 428.565 27.4 ;
      RECT 428.395 23.71 428.925 23.88 ;
      RECT 424.325 23.78 425.07 23.95 ;
      RECT 424.47 23.71 425 23.78 ;
      RECT 424.325 23.95 424.495 27.23 ;
      RECT 428.395 23.88 428.565 27.23 ;
      RECT 425.34 23.66 425.51 24.35 ;
      RECT 425.205 24.35 425.51 27.06 ;
      RECT 425.34 22.935 425.59 23.605 ;
      RECT 425.34 23.605 425.555 23.66 ;
      RECT 425.385 21.835 425.555 22.935 ;
      RECT 425.36 20.825 425.555 21.835 ;
      RECT 423.48 20.815 423.65 23.87 ;
      RECT 424.44 20.825 424.61 21.835 ;
      RECT 427.34 19.79 427.87 19.96 ;
      RECT 427.34 19.96 427.51 20.66 ;
      RECT 427.34 18.16 427.51 19.79 ;
      RECT 428.52 19.31 431.05 19.48 ;
      RECT 429.49 20.89 431.05 21.06 ;
      RECT 428.52 19.48 428.69 20.66 ;
      RECT 429.49 21.06 429.66 22.4 ;
      RECT 430.35 21.06 430.52 22.4 ;
      RECT 430.88 19.48 431.05 20.89 ;
      RECT 428.52 18.16 428.69 19.31 ;
      RECT 426.52 23.71 427.05 23.88 ;
      RECT 426.7 22.935 426.87 23.71 ;
      RECT 427.34 21.23 427.51 22.4 ;
      RECT 428.2 21.23 428.37 22.4 ;
      RECT 429.315 22.6 430.665 22.77 ;
      RECT 429.315 22.57 430.565 22.6 ;
      RECT 429.06 21.23 429.23 22.4 ;
      RECT 430.78 21.23 430.95 22.4 ;
      RECT 429.92 21.23 430.09 22.4 ;
      RECT 429.195 19.79 429.87 19.96 ;
      RECT 429.7 19.65 429.87 19.79 ;
      RECT 429.7 19.96 429.87 20.66 ;
      RECT 430.645 22.94 431.175 23.11 ;
      RECT 430.645 23.805 431.61 23.975 ;
      RECT 431.125 23.985 431.795 24.155 ;
      RECT 433 26.625 433.38 27.645 ;
      RECT 430.645 23.11 430.955 23.805 ;
      RECT 431.125 23.975 431.61 23.985 ;
      RECT 431.24 27.645 433.38 27.735 ;
      RECT 431.24 24.155 431.61 27.645 ;
      RECT 431.125 27.735 433.38 27.905 ;
      RECT 426.965 24.08 427.225 27.06 ;
      RECT 425.68 23.78 426.35 23.95 ;
      RECT 425.76 23.04 426.29 23.21 ;
      RECT 425.76 23.21 426.255 23.78 ;
      RECT 426.085 23.95 426.255 27.06 ;
      RECT 427.425 24.08 427.685 27.06 ;
      RECT 430.785 24.145 430.955 24.375 ;
      RECT 430.785 24.375 431.07 27.085 ;
      RECT 426.31 27.655 429.845 27.905 ;
      RECT 429.315 25.395 429.845 27.655 ;
      RECT 428.975 24.37 429.145 27.37 ;
      RECT 430.32 24.395 430.49 27.475 ;
      RECT 434.215 20.5 435.225 20.67 ;
      RECT 434.695 20.44 435.225 20.5 ;
      RECT 432.925 20.5 433.935 20.67 ;
      RECT 432.925 20.44 433.455 20.5 ;
      RECT 432.165 23.125 432.785 23.455 ;
      RECT 432.46 23.71 433.38 23.88 ;
      RECT 432.46 23.455 432.785 23.71 ;
      RECT 433.21 23.88 433.38 25.045 ;
      RECT 432.82 20.84 432.99 22.635 ;
      RECT 433.04 23.07 433.71 23.24 ;
      RECT 433.11 22.94 433.64 23.07 ;
      RECT 433.34 22.565 433.87 22.735 ;
      RECT 433.7 21.625 433.87 22.565 ;
      RECT 434.28 22.565 434.81 22.735 ;
      RECT 434.28 21.625 434.45 22.565 ;
      RECT 431.825 22.55 432.11 22.72 ;
      RECT 431.825 22.72 431.995 23.625 ;
      RECT 431.825 23.625 432.29 23.795 ;
      RECT 432.12 23.795 432.29 24.375 ;
      RECT 431.94 21.625 432.11 22.55 ;
      RECT 432.12 24.375 432.83 24.845 ;
      RECT 432.66 24.845 432.83 27.085 ;
      RECT 435.365 23.125 435.985 23.455 ;
      RECT 434.77 23.71 435.69 23.88 ;
      RECT 435.365 23.455 435.69 23.71 ;
      RECT 434.77 23.88 434.94 25.045 ;
      RECT 435.16 20.84 435.33 22.635 ;
      RECT 434.44 23.07 435.11 23.24 ;
      RECT 434.51 22.94 435.04 23.07 ;
      RECT 436.04 22.55 436.325 22.72 ;
      RECT 436.155 22.72 436.325 23.625 ;
      RECT 435.86 23.625 436.325 23.795 ;
      RECT 435.86 23.795 436.03 24.375 ;
      RECT 436.04 21.625 436.21 22.55 ;
      RECT 435.32 24.375 436.03 24.845 ;
      RECT 435.32 24.845 435.49 27.085 ;
      RECT 433.31 25.52 434.84 26.27 ;
      RECT 433.55 26.27 434.6 27.475 ;
      RECT 433.55 24.375 434.6 25.52 ;
      RECT 431.78 24.375 431.95 27.475 ;
      RECT 436.355 23.985 437.025 24.155 ;
      RECT 436.54 23.805 437.505 23.975 ;
      RECT 434.77 26.625 435.15 27.645 ;
      RECT 436.975 22.94 437.505 23.11 ;
      RECT 436.54 23.975 437.025 23.985 ;
      RECT 437.195 23.11 437.505 23.805 ;
      RECT 434.77 27.645 436.91 27.735 ;
      RECT 436.54 24.155 436.91 27.645 ;
      RECT 434.77 27.735 437.025 27.905 ;
      RECT 436.2 24.375 436.37 27.475 ;
      RECT 437.1 19.31 439.63 19.48 ;
      RECT 437.1 20.89 438.66 21.06 ;
      RECT 437.1 19.48 437.27 20.89 ;
      RECT 437.63 21.06 437.8 22.4 ;
      RECT 438.49 21.06 438.66 22.4 ;
      RECT 439.46 19.48 439.63 20.66 ;
      RECT 439.46 18.16 439.63 19.31 ;
      RECT 437.2 21.23 437.37 22.4 ;
      RECT 438.06 21.23 438.23 22.4 ;
      RECT 438.92 21.23 439.09 22.4 ;
      RECT 439.78 21.23 439.95 22.4 ;
      RECT 438.28 19.79 438.955 19.96 ;
      RECT 438.28 19.65 438.45 19.79 ;
      RECT 438.28 19.96 438.45 20.66 ;
      RECT 440.28 19.79 440.81 19.96 ;
      RECT 440.64 19.96 440.81 20.66 ;
      RECT 440.64 18.16 440.81 19.79 ;
      RECT 440.64 21.23 440.81 22.4 ;
      RECT 408.295 22.6 409.645 22.77 ;
      RECT 408.295 22.57 409.545 22.6 ;
      RECT 411.145 23.125 411.765 23.455 ;
      RECT 411.44 23.71 412.36 23.88 ;
      RECT 411.44 23.455 411.765 23.71 ;
      RECT 412.19 23.88 412.36 25.045 ;
      RECT 408.04 21.23 408.21 22.4 ;
      RECT 409.76 21.23 409.93 22.4 ;
      RECT 408.9 21.23 409.07 22.4 ;
      RECT 408.175 19.79 408.85 19.96 ;
      RECT 408.68 19.65 408.85 19.79 ;
      RECT 408.68 19.96 408.85 20.66 ;
      RECT 409.625 22.94 410.155 23.11 ;
      RECT 409.625 23.805 410.59 23.975 ;
      RECT 410.105 23.985 410.775 24.155 ;
      RECT 411.98 26.625 412.36 27.645 ;
      RECT 409.625 23.11 409.935 23.805 ;
      RECT 410.105 23.975 410.59 23.985 ;
      RECT 410.22 27.645 412.36 27.735 ;
      RECT 410.22 24.155 410.59 27.645 ;
      RECT 410.105 27.735 412.36 27.905 ;
      RECT 410.805 22.55 411.09 22.72 ;
      RECT 410.805 22.72 410.975 23.625 ;
      RECT 410.805 23.625 411.27 23.795 ;
      RECT 411.1 23.795 411.27 24.375 ;
      RECT 410.92 21.625 411.09 22.55 ;
      RECT 411.1 24.375 411.81 24.845 ;
      RECT 411.64 24.845 411.81 27.085 ;
      RECT 413.195 20.5 414.205 20.67 ;
      RECT 413.675 20.44 414.205 20.5 ;
      RECT 411.905 20.5 412.915 20.67 ;
      RECT 411.905 20.44 412.435 20.5 ;
      RECT 411.8 20.84 411.97 22.635 ;
      RECT 413.42 23.07 414.09 23.24 ;
      RECT 413.49 22.94 414.02 23.07 ;
      RECT 412.02 23.07 412.69 23.24 ;
      RECT 412.09 22.94 412.62 23.07 ;
      RECT 413.26 22.565 413.79 22.735 ;
      RECT 413.26 21.625 413.43 22.565 ;
      RECT 412.32 22.565 412.85 22.735 ;
      RECT 412.68 21.625 412.85 22.565 ;
      RECT 410.76 24.375 410.93 27.475 ;
      RECT 409.765 24.145 409.935 24.375 ;
      RECT 409.765 24.375 410.05 27.085 ;
      RECT 405.29 27.655 408.825 27.905 ;
      RECT 408.295 25.395 408.825 27.655 ;
      RECT 409.3 24.395 409.47 27.475 ;
      RECT 414.345 23.125 414.965 23.455 ;
      RECT 414.345 23.455 414.67 23.71 ;
      RECT 413.75 23.71 414.67 23.88 ;
      RECT 413.75 23.88 413.92 25.045 ;
      RECT 412.29 25.52 413.82 26.27 ;
      RECT 412.53 26.27 413.58 27.475 ;
      RECT 412.53 24.375 413.58 25.52 ;
      RECT 414.14 20.84 414.31 22.635 ;
      RECT 417.9 21.23 418.07 22.4 ;
      RECT 416.08 19.31 418.61 19.48 ;
      RECT 416.08 20.89 417.64 21.06 ;
      RECT 416.08 19.48 416.25 20.89 ;
      RECT 416.61 21.06 416.78 22.4 ;
      RECT 417.47 21.06 417.64 22.4 ;
      RECT 418.44 19.48 418.61 20.66 ;
      RECT 418.44 18.16 418.61 19.31 ;
      RECT 416.18 21.23 416.35 22.4 ;
      RECT 417.04 21.23 417.21 22.4 ;
      RECT 417.26 19.79 417.935 19.96 ;
      RECT 417.26 19.65 417.43 19.79 ;
      RECT 417.26 19.96 417.43 20.66 ;
      RECT 418.76 21.23 418.93 22.4 ;
      RECT 419.26 19.79 419.79 19.96 ;
      RECT 419.62 19.96 419.79 20.66 ;
      RECT 419.62 18.16 419.79 19.79 ;
      RECT 414.84 23.795 415.01 24.375 ;
      RECT 414.84 23.625 415.305 23.795 ;
      RECT 415.135 22.72 415.305 23.625 ;
      RECT 415.02 22.55 415.305 22.72 ;
      RECT 414.3 24.375 415.01 24.845 ;
      RECT 415.02 21.625 415.19 22.55 ;
      RECT 414.3 24.845 414.47 27.085 ;
      RECT 416.465 22.6 417.815 22.77 ;
      RECT 416.565 22.57 417.815 22.6 ;
      RECT 415.335 23.985 416.005 24.155 ;
      RECT 415.52 23.805 416.485 23.975 ;
      RECT 413.75 26.625 414.13 27.645 ;
      RECT 415.955 22.94 416.485 23.11 ;
      RECT 415.52 23.975 416.005 23.985 ;
      RECT 415.52 24.155 415.89 27.645 ;
      RECT 416.175 23.11 416.485 23.805 ;
      RECT 413.75 27.645 415.89 27.735 ;
      RECT 413.75 27.735 416.005 27.905 ;
      RECT 415.18 24.375 415.35 27.475 ;
      RECT 416.175 24.145 416.345 24.375 ;
      RECT 416.06 24.375 416.345 27.085 ;
      RECT 417.285 27.655 420.82 27.905 ;
      RECT 417.285 25.395 417.815 27.655 ;
      RECT 416.64 24.395 416.81 27.475 ;
      RECT 418.205 23.71 418.735 23.88 ;
      RECT 418.565 27.23 422.805 27.4 ;
      RECT 422.06 23.78 422.805 23.95 ;
      RECT 422.13 23.71 422.66 23.78 ;
      RECT 418.565 23.88 418.735 27.23 ;
      RECT 422.635 23.95 422.805 27.23 ;
      RECT 419.445 24.08 419.705 27.06 ;
      RECT 417.985 24.37 418.155 27.37 ;
      RECT 422.675 19.94 422.845 20.61 ;
      RECT 424.285 19.94 424.455 20.61 ;
      RECT 419.905 24.08 420.165 27.06 ;
      RECT 419.62 21.23 419.79 22.4 ;
      RECT 420.08 23.71 420.61 23.88 ;
      RECT 420.26 22.935 420.43 23.71 ;
      RECT 422.82 23.21 422.99 23.605 ;
      RECT 422.82 22.935 422.99 23.04 ;
      RECT 421.96 23.04 422.99 23.21 ;
      RECT 422.715 22.155 423.25 22.73 ;
      RECT 420.78 23.78 421.45 23.95 ;
      RECT 420.84 23.04 421.37 23.21 ;
      RECT 420.875 23.21 421.37 23.78 ;
      RECT 420.875 23.95 421.045 27.06 ;
      RECT 421.62 23.66 421.79 24.35 ;
      RECT 421.62 24.35 421.925 27.06 ;
      RECT 421.54 22.935 421.79 23.605 ;
      RECT 421.575 23.605 421.79 23.66 ;
      RECT 421.575 21.835 421.745 22.935 ;
      RECT 421.575 20.825 421.77 21.835 ;
      RECT 422.52 20.825 422.69 21.835 ;
      RECT 424.14 23.21 424.31 23.605 ;
      RECT 424.14 22.935 424.31 23.04 ;
      RECT 300.845 20.5 301.855 20.67 ;
      RECT 300.965 20.47 301.855 20.5 ;
      RECT 300.845 21.36 301.855 21.53 ;
      RECT 308.155 20.855 309.505 21.085 ;
      RECT 308.155 24.815 309.505 24.985 ;
      RECT 308.155 18.575 309.505 18.745 ;
      RECT 308.155 23.255 309.505 23.425 ;
      RECT 308.155 21.695 309.505 21.865 ;
      RECT 308.155 20.135 309.505 20.305 ;
      RECT 308.155 22.475 309.505 22.645 ;
      RECT 308.155 19.355 309.505 19.525 ;
      RECT 304.315 25.745 307.025 25.915 ;
      RECT 304.315 23.465 307.025 23.635 ;
      RECT 304.315 21.185 307.025 21.355 ;
      RECT 304.315 18.905 307.025 19.075 ;
      RECT 308.155 24.035 309.505 24.205 ;
      RECT 312.825 19.17 313.155 19.935 ;
      RECT 314.625 20.79 315.635 20.96 ;
      RECT 314.625 23.13 315.635 23.3 ;
      RECT 314.625 25.47 316.025 25.64 ;
      RECT 315.855 21.015 316.025 25.47 ;
      RECT 314.625 18.065 315.635 18.235 ;
      RECT 314.625 18.525 315.635 18.695 ;
      RECT 314.625 21.57 315.635 21.74 ;
      RECT 314.625 22.35 315.635 22.52 ;
      RECT 314.625 24.69 315.635 24.86 ;
      RECT 314.625 23.91 315.635 24.08 ;
      RECT 320.085 23.975 320.815 24.145 ;
      RECT 320.085 24.145 320.735 24.225 ;
      RECT 320.085 23.895 320.735 23.975 ;
      RECT 320.225 24.525 320.875 24.855 ;
      RECT 320.825 22.635 321.475 22.965 ;
      RECT 320.225 23.265 320.875 23.595 ;
      RECT 324.625 24.525 325.275 24.855 ;
      RECT 323.595 23.895 324.245 24.225 ;
      RECT 323.595 23.265 324.245 23.595 ;
      RECT 324.625 23.895 325.275 24.225 ;
      RECT 323.595 24.525 324.245 24.855 ;
      RECT 324.625 23.265 325.275 23.595 ;
      RECT 329.055 24.605 329.785 24.775 ;
      RECT 329.135 24.775 329.785 24.855 ;
      RECT 329.135 24.525 329.785 24.605 ;
      RECT 329.025 23.975 329.615 24.145 ;
      RECT 329.025 24.145 329.535 24.225 ;
      RECT 329.025 23.895 329.535 23.975 ;
      RECT 332.395 23.895 333.045 24.225 ;
      RECT 327.995 23.265 328.645 23.595 ;
      RECT 328.135 24.145 328.305 24.225 ;
      RECT 328.135 23.895 328.305 23.975 ;
      RECT 328.475 24.145 328.645 24.225 ;
      RECT 328.055 23.975 328.645 24.145 ;
      RECT 328.475 23.895 328.645 23.975 ;
      RECT 330.425 25.155 331.075 25.485 ;
      RECT 332.425 23.265 333.075 23.595 ;
      RECT 333.825 23.895 334.475 24.225 ;
      RECT 332.825 24.525 333.475 24.855 ;
      RECT 341.195 22.635 341.845 22.965 ;
      RECT 341.195 23.265 341.845 23.595 ;
      RECT 341.195 25.155 341.845 25.485 ;
      RECT 341.195 23.895 341.845 24.225 ;
      RECT 341.195 24.525 341.845 24.855 ;
      RECT 347.875 23.025 350.585 23.195 ;
      RECT 347.875 19.185 350.585 19.355 ;
      RECT 347.875 21.745 350.585 21.915 ;
      RECT 347.875 20.465 350.585 20.635 ;
      RECT 351.525 21.745 354.235 21.915 ;
      RECT 351.525 23.025 354.235 23.195 ;
      RECT 351.525 27.305 354.235 27.475 ;
      RECT 351.525 23.195 353.91 27.305 ;
      RECT 351.525 21.915 353.91 23.025 ;
      RECT 351.525 20.465 354.235 20.635 ;
      RECT 355.175 23.025 357.885 23.195 ;
      RECT 355.175 20.465 357.885 20.635 ;
      RECT 355.175 19.185 357.885 19.355 ;
      RECT 351.525 19.185 354.235 19.355 ;
      RECT 355.175 21.745 357.885 21.915 ;
      RECT 358.105 21.575 358.285 22.11 ;
      RECT 358.105 22.11 358.275 22.505 ;
      RECT 358.105 21.155 358.275 21.575 ;
      RECT 358.105 26.92 358.275 27.115 ;
      RECT 357.98 23.58 358.275 26.92 ;
      RECT 358.105 23.385 358.275 23.58 ;
      RECT 363.74 24.64 365.065 25.05 ;
      RECT 363.395 19.075 363.935 24.47 ;
      RECT 364.87 19.075 365.41 24.47 ;
      RECT 370.345 24.64 371.67 25.05 ;
      RECT 371.475 19.075 372.015 24.47 ;
      RECT 370 19.075 370.54 24.47 ;
      RECT 403.265 19.94 403.435 20.61 ;
      RECT 404.365 21.835 404.535 22.935 ;
      RECT 404.32 22.935 404.57 23.605 ;
      RECT 404.32 23.605 404.535 23.66 ;
      RECT 404.185 24.35 404.49 27.06 ;
      RECT 404.32 23.66 404.49 24.35 ;
      RECT 404.34 20.825 404.535 21.835 ;
      RECT 403.42 20.825 403.59 21.835 ;
      RECT 406.32 19.79 406.85 19.96 ;
      RECT 406.32 19.96 406.49 20.66 ;
      RECT 406.32 18.16 406.49 19.79 ;
      RECT 406.32 21.23 406.49 22.4 ;
      RECT 407.18 21.23 407.35 22.4 ;
      RECT 407.5 19.31 410.03 19.48 ;
      RECT 408.47 20.89 410.03 21.06 ;
      RECT 407.5 19.48 407.67 20.66 ;
      RECT 408.47 21.06 408.64 22.4 ;
      RECT 409.33 21.06 409.5 22.4 ;
      RECT 409.86 19.48 410.03 20.89 ;
      RECT 407.5 18.16 407.67 19.31 ;
      RECT 403.12 23.21 403.29 23.605 ;
      RECT 403.12 22.935 403.29 23.04 ;
      RECT 403.12 23.04 404.15 23.21 ;
      RECT 402.86 22.155 403.395 22.73 ;
      RECT 403.305 27.23 407.545 27.4 ;
      RECT 407.375 23.71 407.905 23.88 ;
      RECT 403.305 23.78 404.05 23.95 ;
      RECT 403.45 23.71 403.98 23.78 ;
      RECT 403.305 23.95 403.475 27.23 ;
      RECT 407.375 23.88 407.545 27.23 ;
      RECT 405.5 23.71 406.03 23.88 ;
      RECT 405.68 22.935 405.85 23.71 ;
      RECT 405.945 24.08 406.205 27.06 ;
      RECT 404.66 23.78 405.33 23.95 ;
      RECT 404.74 23.04 405.27 23.21 ;
      RECT 404.74 23.21 405.235 23.78 ;
      RECT 405.065 23.95 405.235 27.06 ;
      RECT 406.405 24.08 406.665 27.06 ;
      RECT 407.955 24.37 408.125 27.37 ;
      RECT 258.655 21.61 258.825 24.645 ;
      RECT 258.65 19.745 258.91 20.385 ;
      RECT 258.665 18.945 258.865 19.745 ;
      RECT 258.695 20.385 258.865 21.025 ;
      RECT 259.73 18.04 260.87 18.21 ;
      RECT 259.805 18.21 260.695 18.27 ;
      RECT 257.8 19.795 258.415 21.225 ;
      RECT 257.8 19.625 258.48 19.795 ;
      RECT 257.8 21.225 258.475 21.395 ;
      RECT 258.545 25.215 258.805 26.145 ;
      RECT 257.875 24.955 258.805 25.215 ;
      RECT 258.545 26.145 259.685 26.405 ;
      RECT 259.28 26.405 259.45 27.1 ;
      RECT 259.28 26.09 259.45 26.145 ;
      RECT 260.09 25.13 263.995 25.3 ;
      RECT 268.485 23.85 268.655 26.56 ;
      RECT 268.485 19.87 268.655 22.58 ;
      RECT 267.205 23.85 267.375 26.56 ;
      RECT 267.205 19.87 267.375 22.58 ;
      RECT 265.925 23.85 266.095 26.56 ;
      RECT 265.925 19.87 266.095 22.58 ;
      RECT 263.485 19.87 263.655 24.62 ;
      RECT 264.765 19.87 264.935 24.62 ;
      RECT 263.985 21.22 264.53 23.41 ;
      RECT 263.985 21.12 264.515 21.22 ;
      RECT 266.025 22.75 278.67 23.68 ;
      RECT 273.605 19.87 273.775 22.58 ;
      RECT 272.325 23.85 272.495 26.56 ;
      RECT 272.325 19.87 272.495 22.58 ;
      RECT 271.045 23.85 271.215 26.56 ;
      RECT 271.045 19.87 271.215 22.58 ;
      RECT 269.765 23.85 269.935 26.56 ;
      RECT 269.765 19.87 269.935 22.58 ;
      RECT 273.605 23.85 273.775 26.56 ;
      RECT 278.725 23.85 278.895 26.56 ;
      RECT 278.725 19.87 278.895 22.58 ;
      RECT 277.445 23.85 277.615 26.56 ;
      RECT 277.445 19.87 277.615 22.58 ;
      RECT 276.165 23.85 276.335 26.56 ;
      RECT 276.165 19.87 276.335 22.58 ;
      RECT 274.885 23.85 275.055 26.56 ;
      RECT 274.885 19.87 275.055 22.58 ;
      RECT 279.605 19.87 279.775 22.58 ;
      RECT 280.485 23.85 280.655 26.56 ;
      RECT 279.605 23.85 279.775 26.56 ;
      RECT 278.95 22.75 284.01 23.68 ;
      RECT 280.485 19.87 280.655 22.58 ;
      RECT 286.17 3.825 286.34 23.71 ;
      RECT 285.52 23.765 285.94 24.295 ;
      RECT 284.005 19.87 284.175 22.58 ;
      RECT 284.005 23.85 284.175 26.56 ;
      RECT 281.365 19.87 281.535 22.58 ;
      RECT 283.125 19.87 283.295 22.58 ;
      RECT 281.365 23.85 281.535 26.56 ;
      RECT 283.125 23.85 283.295 26.56 ;
      RECT 282.245 19.87 282.415 22.58 ;
      RECT 282.245 23.85 282.415 26.56 ;
      RECT 287.525 19.965 288.925 20.135 ;
      RECT 288.755 18.36 288.925 19.965 ;
      RECT 290.655 19.965 292.085 20.135 ;
      RECT 290.655 18.36 290.825 19.965 ;
      RECT 287.525 18.135 288.535 18.305 ;
      RECT 291.075 18.135 292.085 18.305 ;
      RECT 290.655 20.305 290.825 21.19 ;
      RECT 287.525 22.525 288.535 22.695 ;
      RECT 288.755 20.305 288.925 21.19 ;
      RECT 290.655 21.47 290.825 23.46 ;
      RECT 288.755 21.755 288.925 23.46 ;
      RECT 287.525 21.245 288.535 21.415 ;
      RECT 287.525 19.415 288.535 19.585 ;
      RECT 291.075 19.415 292.085 19.585 ;
      RECT 291.075 21.245 292.085 21.415 ;
      RECT 291.075 22.525 292.085 22.695 ;
      RECT 286.61 24.275 286.78 24.295 ;
      RECT 286.61 23.765 286.99 24.275 ;
      RECT 287.525 24.56 288.185 24.755 ;
      RECT 287.525 24.355 288.535 24.56 ;
      RECT 287.525 23.245 288.115 24.055 ;
      RECT 287.525 23.075 288.535 23.245 ;
      RECT 291.075 23.075 292.085 23.245 ;
      RECT 288.755 24.16 288.925 24.3 ;
      RECT 288.34 23.63 288.925 24.16 ;
      RECT 290.655 24.14 290.825 24.3 ;
      RECT 290.655 23.97 291.415 24.14 ;
      RECT 290.655 23.63 290.825 23.97 ;
      RECT 288.395 25.065 288.925 25.235 ;
      RECT 288.755 25.235 288.925 26.46 ;
      RECT 288.755 24.58 288.925 25.065 ;
      RECT 290.655 25.065 291.185 25.235 ;
      RECT 290.655 25.235 290.825 25.38 ;
      RECT 290.655 24.58 290.825 25.065 ;
      RECT 291.075 24.355 292.085 24.525 ;
      RECT 291.075 25.435 292.085 25.605 ;
      RECT 287.525 25.435 288.535 25.605 ;
      RECT 296.4 24.345 299.22 24.525 ;
      RECT 296.4 21.455 296.58 24.345 ;
      RECT 296.4 20.535 299.22 20.715 ;
      RECT 296.4 20.715 296.58 20.845 ;
      RECT 299.04 20.715 299.22 24.345 ;
      RECT 295.225 21.015 297.08 21.285 ;
      RECT 295.225 21.285 295.395 21.605 ;
      RECT 296.91 21.285 297.08 23.71 ;
      RECT 296.4 25.5 299.22 25.68 ;
      RECT 296.4 25.68 296.58 34.06 ;
      RECT 296.4 34.06 299.22 34.24 ;
      RECT 299.04 25.68 299.22 34.06 ;
      RECT 296.9 18 298.37 18.17 ;
      RECT 296.9 18.17 297.07 18.955 ;
      RECT 297.3 21.125 298.31 21.295 ;
      RECT 297.3 23.765 298.31 23.935 ;
      RECT 297.36 18.55 298.37 18.72 ;
      RECT 297.36 19.01 298.37 19.18 ;
      RECT 297.3 22.005 298.31 22.175 ;
      RECT 297.3 22.885 298.31 23.055 ;
      RECT 300.415 22.57 300.585 27.125 ;
      RECT 300.045 19.005 300.585 19.535 ;
      RECT 300.415 19.535 300.585 19.725 ;
      RECT 300.415 20.295 300.585 21.735 ;
      RECT 300.845 20.07 301.855 20.24 ;
      RECT 300.845 21.79 301.855 21.96 ;
      RECT 300.845 18.37 301.855 18.54 ;
      RECT 300.845 18.83 301.855 19 ;
      RECT 300.845 19.29 301.855 19.46 ;
      RECT 300.845 22.46 301.855 22.63 ;
      RECT 300.845 20.93 301.855 21.1 ;
      RECT 300.845 23.64 301.855 23.81 ;
      RECT 300.845 24.82 301.855 24.99 ;
      RECT 154.585 19.08 154.755 23.495 ;
      RECT 155.62 22.01 155.88 22.655 ;
      RECT 155.665 22.655 155.835 25.87 ;
      RECT 155.665 19.08 155.835 22.01 ;
      RECT 153.46 19.565 153.72 20.6 ;
      RECT 153.505 20.6 153.675 25.87 ;
      RECT 153.505 19.08 153.675 19.565 ;
      RECT 164.01 18.25 165.335 18.66 ;
      RECT 163.665 18.83 164.205 24.225 ;
      RECT 165.14 18.83 165.68 24.225 ;
      RECT 170.25 18.83 170.79 24.225 ;
      RECT 170.595 18.25 171.92 18.66 ;
      RECT 171.725 18.83 172.265 24.225 ;
      RECT 176.975 23.665 178.995 24.415 ;
      RECT 211.01 23.665 213.03 24.415 ;
      RECT 218.085 18.25 219.41 18.66 ;
      RECT 219.215 18.83 219.755 24.225 ;
      RECT 217.74 18.83 218.28 24.225 ;
      RECT 224.67 18.25 225.995 18.66 ;
      RECT 224.325 18.83 224.865 24.225 ;
      RECT 225.8 18.83 226.34 24.225 ;
      RECT 234.125 22.01 234.385 22.655 ;
      RECT 234.17 22.655 234.34 25.87 ;
      RECT 234.17 19.08 234.34 22.01 ;
      RECT 233.575 19.055 233.745 26.47 ;
      RECT 239.155 24.97 239.325 26.47 ;
      RECT 239.155 24.8 244.845 24.97 ;
      RECT 233.575 26.47 239.325 26.64 ;
      RECT 235.205 23.495 235.465 25 ;
      RECT 235.25 25 235.42 25.87 ;
      RECT 235.25 19.08 235.42 23.495 ;
      RECT 238.445 19.565 238.705 20.6 ;
      RECT 238.49 20.6 238.66 25.87 ;
      RECT 238.49 19.08 238.66 19.565 ;
      RECT 239.5 22.015 239.76 22.655 ;
      RECT 239.545 22.655 239.715 24.28 ;
      RECT 239.545 19.53 239.715 22.015 ;
      RECT 237.365 23.495 237.625 25 ;
      RECT 237.41 25 237.58 25.87 ;
      RECT 237.41 19.08 237.58 23.495 ;
      RECT 236.285 19.565 236.545 20.6 ;
      RECT 236.33 20.6 236.5 25.87 ;
      RECT 236.33 19.08 236.5 19.565 ;
      RECT 239.77 18.85 244.79 19.02 ;
      RECT 239.605 25.475 239.775 27.495 ;
      RECT 236.735 18.82 237.16 26.185 ;
      RECT 234.49 18.65 238.435 18.82 ;
      RECT 237.75 22.94 238.28 23.11 ;
      RECT 237.815 23.11 238.24 26.185 ;
      RECT 237.815 18.82 238.24 22.94 ;
      RECT 240.285 25.39 245.035 25.56 ;
      RECT 244.845 19.53 245.015 19.565 ;
      RECT 244.8 19.565 245.06 24.34 ;
      RECT 243.285 19.53 243.455 19.565 ;
      RECT 243.24 19.565 243.5 24.34 ;
      RECT 242.62 22.015 242.88 22.655 ;
      RECT 242.665 22.655 242.835 24.28 ;
      RECT 242.665 19.53 242.835 22.015 ;
      RECT 245.71 25.675 245.97 26.655 ;
      RECT 245.755 23.885 245.925 25.675 ;
      RECT 245.305 22.19 245.695 22.84 ;
      RECT 245.305 22.84 247.25 23.235 ;
      RECT 241.06 22.015 241.32 22.655 ;
      RECT 241.105 22.655 241.275 24.28 ;
      RECT 241.105 19.53 241.275 22.015 ;
      RECT 244.02 22.7 244.28 23.34 ;
      RECT 244.065 23.34 244.235 24.28 ;
      RECT 244.065 19.53 244.235 22.7 ;
      RECT 241.84 20.875 242.1 21.515 ;
      RECT 241.885 21.515 242.055 24.28 ;
      RECT 241.885 19.53 242.055 20.875 ;
      RECT 240.28 20.875 240.54 21.515 ;
      RECT 240.325 21.515 240.495 24.28 ;
      RECT 240.325 19.53 240.495 20.875 ;
      RECT 247.115 19.775 252.825 19.945 ;
      RECT 250.23 20.24 250.49 21.31 ;
      RECT 248.67 20.24 248.93 21.31 ;
      RECT 247.11 20.24 247.37 21.31 ;
      RECT 246.015 20.815 246.69 21.145 ;
      RECT 247.42 22.67 247.68 23.405 ;
      RECT 246.49 23.405 247.68 23.71 ;
      RECT 246.015 21.145 246.605 22.08 ;
      RECT 246.015 19.325 246.605 20.815 ;
      RECT 246.49 23.71 246.75 26.595 ;
      RECT 246.015 22.08 248.66 22.67 ;
      RECT 249.495 20.3 249.665 21.655 ;
      RECT 247.89 21.125 248.15 21.765 ;
      RECT 247.935 20.3 248.105 21.125 ;
      RECT 251.055 20.3 251.225 21.57 ;
      RECT 250.23 25.675 250.49 26.655 ;
      RECT 250.275 23.885 250.445 25.675 ;
      RECT 248.67 25.675 248.93 26.655 ;
      RECT 248.715 23.885 248.885 25.675 ;
      RECT 247.89 23.495 248.15 26.595 ;
      RECT 247.27 25.675 247.53 26.655 ;
      RECT 247.315 23.885 247.485 25.675 ;
      RECT 249.495 23.67 249.665 26.595 ;
      RECT 248.94 22.08 250.22 22.67 ;
      RECT 250.5 22.08 252.38 22.67 ;
      RECT 251.055 23.67 251.225 26.595 ;
      RECT 254.575 24.795 257.655 25.31 ;
      RECT 254.575 23.36 255.065 24.795 ;
      RECT 257.225 25.31 257.655 25.36 ;
      RECT 257.225 25.36 257.765 28.03 ;
      RECT 257.225 28.03 257.755 28.2 ;
      RECT 253.615 23.36 254.025 23.375 ;
      RECT 253.615 21.34 254.025 22.85 ;
      RECT 253.615 22.85 255.065 23.36 ;
      RECT 251.79 20.24 252.05 21.31 ;
      RECT 251.79 25.675 252.05 26.655 ;
      RECT 251.835 23.885 252.005 25.675 ;
      RECT 254.145 23.61 254.315 26.08 ;
      RECT 253.265 20.41 253.435 25.94 ;
      RECT 255.46 21.085 255.63 24.2 ;
      RECT 254.11 19.55 255.63 21.085 ;
      RECT 252.615 23.67 252.785 26.595 ;
      RECT 252.615 20.3 252.785 21.57 ;
      RECT 255.8 19.96 256.31 24.415 ;
      RECT 257.3 21.33 257.595 22.705 ;
      RECT 257.375 22.705 257.545 24.32 ;
      RECT 257.305 18.94 257.595 21.33 ;
      RECT 255.86 25.73 256.44 26.865 ;
      RECT 256.535 21.225 257.08 21.395 ;
      RECT 259.865 19.87 260.035 24.62 ;
      RECT 260.645 19.87 260.815 24.62 ;
      RECT 261.425 19.87 261.595 24.62 ;
      RECT 262.205 19.87 262.375 24.62 ;
      RECT 118.79 19.87 118.96 22.58 ;
      RECT 120.07 23.85 120.24 26.56 ;
      RECT 120.07 19.87 120.24 22.58 ;
      RECT 121.35 23.85 121.52 26.56 ;
      RECT 121.35 19.87 121.52 22.58 ;
      RECT 122.63 23.85 122.8 26.56 ;
      RECT 122.63 19.87 122.8 22.58 ;
      RECT 123.91 23.85 124.08 26.56 ;
      RECT 123.91 19.87 124.08 22.58 ;
      RECT 129.97 19.87 130.14 24.62 ;
      RECT 129.19 19.87 129.36 24.62 ;
      RECT 128.41 19.87 128.58 24.62 ;
      RECT 127.63 19.87 127.8 24.62 ;
      RECT 126.35 19.87 126.52 24.62 ;
      RECT 125.07 19.87 125.24 24.62 ;
      RECT 129.135 18.04 130.275 18.21 ;
      RECT 129.31 18.21 130.2 18.27 ;
      RECT 125.475 21.22 126.02 23.41 ;
      RECT 125.49 21.12 126.02 21.22 ;
      RECT 126.01 25.13 129.915 25.3 ;
      RECT 131.18 21.61 131.35 24.645 ;
      RECT 131.095 19.745 131.355 20.385 ;
      RECT 131.14 18.945 131.34 19.745 ;
      RECT 131.14 20.385 131.31 21.025 ;
      RECT 131.59 19.795 132.205 21.225 ;
      RECT 131.525 19.625 132.205 19.795 ;
      RECT 131.53 21.225 132.205 21.395 ;
      RECT 131.2 24.955 132.13 25.215 ;
      RECT 131.2 25.215 131.46 26.145 ;
      RECT 130.32 26.145 131.46 26.405 ;
      RECT 130.555 26.405 130.725 27.1 ;
      RECT 130.555 26.09 130.725 26.145 ;
      RECT 135.69 23.61 135.86 26.08 ;
      RECT 134.375 21.085 134.545 24.2 ;
      RECT 134.375 19.55 135.895 21.085 ;
      RECT 133.695 19.96 134.205 24.415 ;
      RECT 132.41 21.33 132.705 22.705 ;
      RECT 132.46 22.705 132.63 24.32 ;
      RECT 132.41 18.94 132.7 21.33 ;
      RECT 133.565 25.73 134.145 26.865 ;
      RECT 132.925 21.225 133.47 21.395 ;
      RECT 132.24 25.36 132.78 28.03 ;
      RECT 132.35 25.31 132.78 25.36 ;
      RECT 132.25 28.03 132.78 28.2 ;
      RECT 132.35 24.795 135.43 25.31 ;
      RECT 134.94 23.36 135.43 24.795 ;
      RECT 135.98 23.36 136.39 23.375 ;
      RECT 135.98 21.34 136.39 22.85 ;
      RECT 134.94 22.85 136.39 23.36 ;
      RECT 137.18 19.775 142.89 19.945 ;
      RECT 136.57 20.41 136.74 25.94 ;
      RECT 137.22 23.67 137.39 26.595 ;
      RECT 139.515 25.675 139.775 26.655 ;
      RECT 139.56 23.885 139.73 25.675 ;
      RECT 137.22 20.3 137.39 21.57 ;
      RECT 137.955 20.24 138.215 21.31 ;
      RECT 138.78 20.3 138.95 21.57 ;
      RECT 139.515 20.24 139.775 21.31 ;
      RECT 137.625 22.08 139.505 22.67 ;
      RECT 138.78 23.67 138.95 26.595 ;
      RECT 139.785 22.08 141.065 22.67 ;
      RECT 137.955 25.675 138.215 26.655 ;
      RECT 138 23.885 138.17 25.675 ;
      RECT 141.075 25.675 141.335 26.655 ;
      RECT 141.12 23.885 141.29 25.675 ;
      RECT 141.075 20.24 141.335 21.31 ;
      RECT 140.34 23.67 140.51 26.595 ;
      RECT 142.325 22.67 142.585 23.405 ;
      RECT 142.325 23.405 143.515 23.71 ;
      RECT 143.315 20.815 143.99 21.145 ;
      RECT 141.345 22.08 143.99 22.67 ;
      RECT 143.4 21.145 143.99 22.08 ;
      RECT 143.4 19.325 143.99 20.815 ;
      RECT 143.255 23.71 143.515 26.595 ;
      RECT 140.34 20.3 140.51 21.655 ;
      RECT 144.97 25.39 149.72 25.56 ;
      RECT 144.99 19.53 145.16 19.565 ;
      RECT 144.945 19.565 145.205 24.34 ;
      RECT 146.55 19.53 146.72 19.565 ;
      RECT 146.505 19.565 146.765 24.34 ;
      RECT 147.125 22.015 147.385 22.655 ;
      RECT 147.17 22.655 147.34 24.28 ;
      RECT 147.17 19.53 147.34 22.015 ;
      RECT 141.855 23.495 142.115 26.595 ;
      RECT 142.475 25.675 142.735 26.655 ;
      RECT 142.52 23.885 142.69 25.675 ;
      RECT 144.035 25.675 144.295 26.655 ;
      RECT 144.08 23.885 144.25 25.675 ;
      RECT 142.635 20.24 142.895 21.31 ;
      RECT 145.215 18.85 150.235 19.02 ;
      RECT 144.31 22.19 144.7 22.84 ;
      RECT 142.755 22.84 144.7 23.235 ;
      RECT 145.725 22.7 145.985 23.34 ;
      RECT 145.77 23.34 145.94 24.28 ;
      RECT 145.77 19.53 145.94 22.7 ;
      RECT 145.16 24.8 150.85 24.97 ;
      RECT 150.68 24.97 150.85 26.47 ;
      RECT 156.26 19.055 156.43 26.47 ;
      RECT 150.68 26.47 156.43 26.64 ;
      RECT 141.855 21.125 142.115 21.765 ;
      RECT 141.9 20.3 142.07 21.125 ;
      RECT 151.3 19.565 151.56 20.6 ;
      RECT 151.345 20.6 151.515 25.87 ;
      RECT 151.345 19.08 151.515 19.565 ;
      RECT 150.245 22.015 150.505 22.655 ;
      RECT 150.29 22.655 150.46 24.28 ;
      RECT 150.29 19.53 150.46 22.015 ;
      RECT 152.38 23.495 152.64 25 ;
      RECT 152.425 25 152.595 25.87 ;
      RECT 152.425 19.08 152.595 23.495 ;
      RECT 150.23 25.475 150.4 27.495 ;
      RECT 152.845 18.82 153.27 26.185 ;
      RECT 151.57 18.65 155.515 18.82 ;
      RECT 151.725 22.94 152.255 23.11 ;
      RECT 151.765 23.11 152.19 26.185 ;
      RECT 151.765 18.82 152.19 22.94 ;
      RECT 148.685 22.015 148.945 22.655 ;
      RECT 148.73 22.655 148.9 24.28 ;
      RECT 148.73 19.53 148.9 22.015 ;
      RECT 147.905 20.875 148.165 21.515 ;
      RECT 147.95 21.515 148.12 24.28 ;
      RECT 147.95 19.53 148.12 20.875 ;
      RECT 149.465 20.875 149.725 21.515 ;
      RECT 149.51 21.515 149.68 24.28 ;
      RECT 149.51 19.53 149.68 20.875 ;
      RECT 154.54 23.495 154.8 25 ;
      RECT 154.585 25 154.755 25.87 ;
      RECT 69.13 23.265 69.78 23.595 ;
      RECT 76.85 19.17 77.18 19.935 ;
      RECT 73.98 25.47 75.38 25.64 ;
      RECT 73.98 21.015 74.15 25.47 ;
      RECT 74.37 20.79 75.38 20.96 ;
      RECT 74.37 23.13 75.38 23.3 ;
      RECT 74.37 18.065 75.38 18.235 ;
      RECT 74.37 18.525 75.38 18.695 ;
      RECT 74.37 21.57 75.38 21.74 ;
      RECT 74.37 22.35 75.38 22.52 ;
      RECT 74.37 24.69 75.38 24.86 ;
      RECT 74.37 23.91 75.38 24.08 ;
      RECT 80.5 20.855 81.85 21.085 ;
      RECT 80.5 20.135 81.85 20.305 ;
      RECT 80.5 24.815 81.85 24.985 ;
      RECT 80.5 18.575 81.85 18.745 ;
      RECT 80.5 23.255 81.85 23.425 ;
      RECT 80.5 21.695 81.85 21.865 ;
      RECT 80.5 22.475 81.85 22.645 ;
      RECT 80.5 19.355 81.85 19.525 ;
      RECT 82.98 25.745 85.69 25.915 ;
      RECT 82.98 23.465 85.69 23.635 ;
      RECT 82.98 21.185 85.69 21.355 ;
      RECT 82.98 18.905 85.69 19.075 ;
      RECT 80.5 24.035 81.85 24.205 ;
      RECT 89.42 22.57 89.59 27.125 ;
      RECT 89.42 19.005 89.96 19.535 ;
      RECT 89.42 19.535 89.59 19.725 ;
      RECT 89.42 20.295 89.59 21.735 ;
      RECT 88.15 20.07 89.16 20.24 ;
      RECT 88.15 21.79 89.16 21.96 ;
      RECT 88.15 18.37 89.16 18.54 ;
      RECT 88.15 18.83 89.16 19 ;
      RECT 88.15 19.29 89.16 19.46 ;
      RECT 88.15 22.46 89.16 22.63 ;
      RECT 88.15 20.93 89.16 21.1 ;
      RECT 88.15 23.64 89.16 23.81 ;
      RECT 88.15 24.82 89.16 24.99 ;
      RECT 88.15 20.5 89.16 20.67 ;
      RECT 88.15 20.47 89.04 20.5 ;
      RECT 88.15 21.36 89.16 21.53 ;
      RECT 90.785 24.345 93.605 24.525 ;
      RECT 93.425 21.455 93.605 24.345 ;
      RECT 90.785 20.535 93.605 20.715 ;
      RECT 93.425 20.715 93.605 20.845 ;
      RECT 90.785 20.715 90.965 24.345 ;
      RECT 92.925 21.015 94.78 21.285 ;
      RECT 94.61 21.285 94.78 21.605 ;
      RECT 92.925 21.285 93.095 23.71 ;
      RECT 90.785 25.5 93.605 25.68 ;
      RECT 93.425 25.68 93.605 34.06 ;
      RECT 90.785 34.06 93.605 34.24 ;
      RECT 90.785 25.68 90.965 34.06 ;
      RECT 91.635 18 93.105 18.17 ;
      RECT 92.935 18.17 93.105 18.955 ;
      RECT 91.695 21.125 92.705 21.295 ;
      RECT 91.695 23.765 92.705 23.935 ;
      RECT 91.635 18.55 92.645 18.72 ;
      RECT 91.635 19.01 92.645 19.18 ;
      RECT 91.695 22.005 92.705 22.175 ;
      RECT 91.695 22.885 92.705 23.055 ;
      RECT 97.92 23.075 98.93 23.245 ;
      RECT 99.18 24.14 99.35 24.3 ;
      RECT 98.59 23.97 99.35 24.14 ;
      RECT 99.18 23.63 99.35 23.97 ;
      RECT 99.18 20.305 99.35 21.19 ;
      RECT 99.18 21.47 99.35 23.46 ;
      RECT 97.92 19.965 99.35 20.135 ;
      RECT 99.18 18.36 99.35 19.965 ;
      RECT 98.82 25.065 99.35 25.235 ;
      RECT 99.18 25.235 99.35 25.38 ;
      RECT 99.18 24.58 99.35 25.065 ;
      RECT 97.92 18.135 98.93 18.305 ;
      RECT 97.92 24.355 98.93 24.525 ;
      RECT 97.92 19.415 98.93 19.585 ;
      RECT 97.92 21.245 98.93 21.415 ;
      RECT 97.92 22.525 98.93 22.695 ;
      RECT 97.92 25.435 98.93 25.605 ;
      RECT 101.08 20.305 101.25 21.19 ;
      RECT 101.08 19.965 102.48 20.135 ;
      RECT 101.08 18.36 101.25 19.965 ;
      RECT 101.47 18.135 102.48 18.305 ;
      RECT 101.47 19.415 102.48 19.585 ;
      RECT 105.83 19.87 106 22.58 ;
      RECT 106.71 19.87 106.88 22.58 ;
      RECT 101.89 23.245 102.48 24.055 ;
      RECT 101.47 23.075 102.48 23.245 ;
      RECT 101.08 24.16 101.25 24.3 ;
      RECT 101.08 23.63 101.665 24.16 ;
      RECT 101.47 24.355 102.48 24.56 ;
      RECT 101.82 24.56 102.48 24.755 ;
      RECT 101.47 22.525 102.48 22.695 ;
      RECT 101.08 21.755 101.25 23.46 ;
      RECT 101.08 25.065 101.61 25.235 ;
      RECT 101.08 25.235 101.25 26.46 ;
      RECT 101.08 24.58 101.25 25.065 ;
      RECT 101.47 21.245 102.48 21.415 ;
      RECT 103.225 24.275 103.395 24.295 ;
      RECT 103.015 23.765 103.395 24.275 ;
      RECT 101.47 25.435 102.48 25.605 ;
      RECT 103.665 3.825 103.835 23.71 ;
      RECT 104.065 23.765 104.485 24.295 ;
      RECT 105.83 23.85 106 26.56 ;
      RECT 105.995 22.75 111.055 23.68 ;
      RECT 106.71 23.85 106.88 26.56 ;
      RECT 111.11 23.85 111.28 26.56 ;
      RECT 111.11 19.87 111.28 22.58 ;
      RECT 112.39 23.85 112.56 26.56 ;
      RECT 112.39 19.87 112.56 22.58 ;
      RECT 110.23 19.87 110.4 22.58 ;
      RECT 108.47 19.87 108.64 22.58 ;
      RECT 109.35 23.85 109.52 26.56 ;
      RECT 110.23 23.85 110.4 26.56 ;
      RECT 108.47 23.85 108.64 26.56 ;
      RECT 107.59 19.87 107.76 22.58 ;
      RECT 109.35 19.87 109.52 22.58 ;
      RECT 107.59 23.85 107.76 26.56 ;
      RECT 117.51 23.85 117.68 26.56 ;
      RECT 117.51 19.87 117.68 22.58 ;
      RECT 113.67 23.85 113.84 26.56 ;
      RECT 113.67 19.87 113.84 22.58 ;
      RECT 114.95 23.85 115.12 26.56 ;
      RECT 114.95 19.87 115.12 22.58 ;
      RECT 116.23 23.85 116.4 26.56 ;
      RECT 116.23 19.87 116.4 22.58 ;
      RECT 111.335 22.75 123.98 23.68 ;
      RECT 118.79 23.85 118.96 26.56 ;
      RECT 442.16 17.155 442.33 18.735 ;
      RECT 441.68 20.825 442.33 21.835 ;
      RECT 439.19 22.765 440.54 22.77 ;
      RECT 442.16 18.905 442.33 20.825 ;
      RECT 441.82 16.775 441.99 17.385 ;
      RECT 444.5 16.775 444.67 17.385 ;
      RECT 441.82 16.605 444.67 16.775 ;
      RECT 438.78 18.225 439.11 19.075 ;
      RECT 438.86 17.615 439.03 18.225 ;
      RECT 439.46 16.86 440.33 17.87 ;
      RECT 439.8 17.87 440.33 18.905 ;
      RECT 442.5 20.07 443.03 20.24 ;
      RECT 442.62 17.155 442.79 20.07 ;
      RECT 440.98 21.975 441.51 22.145 ;
      RECT 441.34 16.85 441.51 21.975 ;
      RECT 448.085 15.745 448.615 15.915 ;
      RECT 448.285 15.915 448.615 15.985 ;
      RECT 448.285 15.505 448.615 15.745 ;
      RECT 448.275 14.04 448.605 15.335 ;
      RECT 448.15 13.335 451.05 13.585 ;
      RECT 450.085 14.04 450.415 15.335 ;
      RECT 448.16 13.585 451.04 14.04 ;
      RECT 448.295 16.155 448.545 17.2 ;
      RECT 448.15 17.37 451.04 17.925 ;
      RECT 449.155 16.155 449.485 17.2 ;
      RECT 448.15 17.925 451.22 18.175 ;
      RECT 450.085 16.155 450.415 17.2 ;
      RECT 448.16 17.2 451.04 17.37 ;
      RECT 443.675 18.735 444.205 18.905 ;
      RECT 443.45 16.965 444.205 17.135 ;
      RECT 444.035 17.135 444.205 18.735 ;
      RECT 444.035 18.905 444.205 20.825 ;
      RECT 444 20.825 444.205 21.835 ;
      RECT 442.96 17.155 443.25 19.575 ;
      RECT 443.2 19.865 443.5 20.5 ;
      RECT 442.96 19.575 443.5 19.865 ;
      RECT 442.96 20.5 443.5 20.655 ;
      RECT 442.96 22.67 443.49 22.84 ;
      RECT 442.96 20.655 443.37 22.67 ;
      RECT 448.725 16.155 448.975 16.935 ;
      RECT 448.805 15.335 448.975 16.155 ;
      RECT 448.805 14.395 449.895 15.335 ;
      RECT 449.145 14.305 449.895 14.395 ;
      RECT 449.655 15.335 449.895 15.505 ;
      RECT 449.655 15.505 450.415 15.985 ;
      RECT 449.145 15.505 449.475 15.985 ;
      RECT 454.075 12.275 454.585 15.045 ;
      RECT 450.585 14.305 450.915 16.935 ;
      RECT 459.25 16.735 459.42 19.445 ;
      RECT 460.13 18.195 460.85 19.445 ;
      RECT 460.13 16.675 460.64 18.195 ;
      RECT 457.935 12.275 459.255 15.045 ;
      RECT 455.295 12.275 455.465 14.985 ;
      RECT 456.175 12.275 456.345 14.985 ;
      RECT 459.19 15.535 460.79 15.705 ;
      RECT 459.965 12.275 460.135 14.985 ;
      RECT 454.64 15.535 457.88 15.705 ;
      RECT 456.34 16.735 456.51 19.445 ;
      RECT 457.055 12.275 457.225 14.985 ;
      RECT 464.16 16.735 464.33 19.445 ;
      RECT 464.325 12.275 464.495 14.985 ;
      RECT 462.73 18.195 463.45 19.445 ;
      RECT 462.94 16.675 463.45 18.195 ;
      RECT 461.655 15.045 461.905 15.165 ;
      RECT 460.845 12.275 462.735 15.045 ;
      RECT 462.55 15.535 464.27 15.705 ;
      RECT 463.445 12.275 463.615 14.985 ;
      RECT 18.335 24.64 19.66 25.05 ;
      RECT 17.99 19.075 18.53 24.47 ;
      RECT 19.465 19.075 20.005 24.47 ;
      RECT 24.94 24.64 26.265 25.05 ;
      RECT 24.595 19.075 25.135 24.47 ;
      RECT 26.07 19.075 26.61 24.47 ;
      RECT 31.72 21.575 31.9 22.11 ;
      RECT 31.73 22.11 31.9 22.505 ;
      RECT 31.73 21.155 31.9 21.575 ;
      RECT 35.77 21.745 38.48 21.915 ;
      RECT 35.77 23.025 38.48 23.195 ;
      RECT 35.77 27.305 38.48 27.475 ;
      RECT 36.095 23.195 38.48 27.305 ;
      RECT 36.095 21.915 38.48 23.025 ;
      RECT 31.73 26.92 31.9 27.115 ;
      RECT 31.73 23.58 32.025 26.92 ;
      RECT 31.73 23.385 31.9 23.58 ;
      RECT 35.77 20.465 38.48 20.635 ;
      RECT 32.12 23.025 34.83 23.195 ;
      RECT 32.12 20.465 34.83 20.635 ;
      RECT 32.12 19.185 34.83 19.355 ;
      RECT 35.77 19.185 38.48 19.355 ;
      RECT 32.12 21.745 34.83 21.915 ;
      RECT 39.42 23.025 42.13 23.195 ;
      RECT 39.42 19.185 42.13 19.355 ;
      RECT 39.42 21.745 42.13 21.915 ;
      RECT 39.42 20.465 42.13 20.635 ;
      RECT 48.16 22.635 48.81 22.965 ;
      RECT 48.16 23.265 48.81 23.595 ;
      RECT 48.16 25.155 48.81 25.485 ;
      RECT 48.16 23.895 48.81 24.225 ;
      RECT 48.16 24.525 48.81 24.855 ;
      RECT 60.39 23.975 60.98 24.145 ;
      RECT 60.47 24.145 60.98 24.225 ;
      RECT 60.47 23.895 60.98 23.975 ;
      RECT 60.22 24.605 60.95 24.775 ;
      RECT 60.22 24.775 60.87 24.855 ;
      RECT 60.22 24.525 60.87 24.605 ;
      RECT 56.96 23.895 57.61 24.225 ;
      RECT 56.93 23.265 57.58 23.595 ;
      RECT 58.93 25.155 59.58 25.485 ;
      RECT 55.53 23.895 56.18 24.225 ;
      RECT 56.53 24.525 57.18 24.855 ;
      RECT 64.73 24.525 65.38 24.855 ;
      RECT 65.76 23.895 66.41 24.225 ;
      RECT 65.76 23.265 66.41 23.595 ;
      RECT 64.73 23.895 65.38 24.225 ;
      RECT 65.76 24.525 66.41 24.855 ;
      RECT 64.73 23.265 65.38 23.595 ;
      RECT 61.36 23.265 62.01 23.595 ;
      RECT 61.7 24.145 61.87 24.225 ;
      RECT 61.7 23.895 61.87 23.975 ;
      RECT 61.36 24.145 61.53 24.225 ;
      RECT 61.36 23.975 61.95 24.145 ;
      RECT 61.36 23.895 61.53 23.975 ;
      RECT 69.19 23.975 69.92 24.145 ;
      RECT 69.27 24.145 69.92 24.225 ;
      RECT 69.27 23.895 69.92 23.975 ;
      RECT 69.13 24.525 69.78 24.855 ;
      RECT 68.53 22.635 69.18 22.965 ;
      RECT 417.67 13.54 417.84 14.59 ;
      RECT 415.91 13.54 416.08 14.59 ;
      RECT 417.76 18.225 418.09 19.075 ;
      RECT 417.84 17.615 418.01 18.225 ;
      RECT 419.43 13.54 419.6 14.59 ;
      RECT 418.44 16.86 419.31 17.87 ;
      RECT 418.78 17.87 419.31 18.905 ;
      RECT 422.95 12.03 423.12 12.56 ;
      RECT 421.19 12.03 421.36 12.36 ;
      RECT 424.71 12.03 424.88 12.56 ;
      RECT 419.96 21.975 420.49 22.145 ;
      RECT 420.32 16.85 420.49 21.975 ;
      RECT 422.655 18.735 423.185 18.905 ;
      RECT 422.43 16.965 423.185 17.135 ;
      RECT 423.015 17.135 423.185 18.735 ;
      RECT 423.015 18.905 423.185 20.825 ;
      RECT 422.98 20.825 423.185 21.835 ;
      RECT 422.95 13.54 423.12 14.59 ;
      RECT 422.95 12.98 423.12 13.31 ;
      RECT 421.19 12.98 421.36 13.31 ;
      RECT 420.78 18.735 421.31 18.905 ;
      RECT 420.66 21.835 420.83 22.595 ;
      RECT 418.17 22.595 420.83 22.765 ;
      RECT 421.14 17.155 421.31 18.735 ;
      RECT 420.66 20.825 421.31 21.835 ;
      RECT 418.17 22.765 419.52 22.77 ;
      RECT 421.14 18.905 421.31 20.825 ;
      RECT 421.94 17.155 422.23 19.575 ;
      RECT 422.18 19.865 422.48 20.5 ;
      RECT 421.94 19.575 422.48 19.865 ;
      RECT 421.94 20.5 422.48 20.655 ;
      RECT 421.94 22.67 422.47 22.84 ;
      RECT 421.94 20.655 422.35 22.67 ;
      RECT 420.8 16.775 420.97 17.385 ;
      RECT 423.48 16.775 423.65 17.385 ;
      RECT 426.16 16.775 426.33 17.385 ;
      RECT 420.8 16.605 426.33 16.775 ;
      RECT 421.19 13.54 421.36 14.59 ;
      RECT 421.48 20.07 422.01 20.24 ;
      RECT 421.6 17.155 421.77 20.07 ;
      RECT 424.71 13.54 424.88 14.59 ;
      RECT 423.945 18.735 424.475 18.905 ;
      RECT 423.945 16.965 424.7 17.135 ;
      RECT 423.945 17.135 424.115 18.735 ;
      RECT 423.945 18.905 424.115 20.825 ;
      RECT 423.945 20.825 424.15 21.835 ;
      RECT 424.71 12.78 424.88 13.31 ;
      RECT 424.9 17.155 425.19 19.575 ;
      RECT 424.65 19.865 424.95 20.5 ;
      RECT 424.65 19.575 425.19 19.865 ;
      RECT 424.65 20.5 425.19 20.655 ;
      RECT 424.66 22.67 425.19 22.84 ;
      RECT 424.78 20.655 425.19 22.67 ;
      RECT 425.12 20.07 425.65 20.24 ;
      RECT 425.36 17.155 425.53 20.07 ;
      RECT 429.83 11.45 431.86 11.62 ;
      RECT 425.82 18.735 426.35 18.905 ;
      RECT 426.3 21.835 426.47 22.595 ;
      RECT 426.3 22.595 428.96 22.765 ;
      RECT 425.82 17.155 425.99 18.735 ;
      RECT 425.82 20.825 426.47 21.835 ;
      RECT 427.61 22.765 428.96 22.77 ;
      RECT 425.82 18.905 425.99 20.825 ;
      RECT 430.77 12.02 430.94 14.73 ;
      RECT 426.98 17.87 427.17 20.89 ;
      RECT 426.98 16.52 429.87 16.69 ;
      RECT 426.98 20.89 428.8 21.06 ;
      RECT 427.77 21.06 427.94 22.4 ;
      RECT 428.63 21.06 428.8 22.4 ;
      RECT 426.98 16.69 427.51 17.87 ;
      RECT 429.7 16.69 429.87 19.14 ;
      RECT 430.52 18.735 431.05 18.905 ;
      RECT 430.88 18.905 431.05 19.14 ;
      RECT 430.88 16.86 431.05 18.735 ;
      RECT 429.04 18.225 429.37 19.075 ;
      RECT 429.12 17.615 429.29 18.225 ;
      RECT 427.82 16.86 428.69 17.87 ;
      RECT 427.82 17.87 428.35 18.905 ;
      RECT 426.64 21.975 427.17 22.145 ;
      RECT 426.64 16.85 426.81 21.975 ;
      RECT 433.3 11.45 434.99 11.62 ;
      RECT 433.88 12.02 434.05 14.73 ;
      RECT 431.185 15.285 431.855 15.455 ;
      RECT 431.245 14.76 431.775 15.285 ;
      RECT 432.945 15.28 433.615 15.45 ;
      RECT 433.005 15.13 433.535 15.28 ;
      RECT 434.77 20.04 435.315 20.21 ;
      RECT 434.77 20.21 434.94 20.24 ;
      RECT 434.77 17.24 434.94 20.04 ;
      RECT 433.99 17.24 434.16 19.95 ;
      RECT 435.55 17.24 435.72 19.95 ;
      RECT 432.835 20.04 433.38 20.21 ;
      RECT 433.21 20.21 433.38 20.24 ;
      RECT 433.21 17.24 433.38 20.04 ;
      RECT 432.43 17.24 432.6 19.95 ;
      RECT 432.55 16.89 435.6 17.025 ;
      RECT 432.39 16.72 435.76 16.89 ;
      RECT 436.38 21.96 436.91 22.13 ;
      RECT 436.495 23.31 437.025 23.48 ;
      RECT 436.495 22.13 436.805 23.31 ;
      RECT 436.52 16.85 436.69 21.96 ;
      RECT 431.24 21.96 431.77 22.13 ;
      RECT 431.125 23.31 431.655 23.48 ;
      RECT 431.345 22.13 431.655 23.31 ;
      RECT 431.46 16.85 431.63 21.96 ;
      RECT 441.06 10.73 441.23 11.06 ;
      RECT 439.09 11.56 439.26 12.75 ;
      RECT 439.09 11.23 439.81 11.56 ;
      RECT 443.03 11.56 443.2 12.75 ;
      RECT 442.48 11.23 443.2 11.56 ;
      RECT 441.06 11.23 441.23 11.56 ;
      RECT 439.64 11.73 439.81 12.74 ;
      RECT 441.06 11.73 441.23 12.74 ;
      RECT 442.48 11.73 442.65 12.74 ;
      RECT 440.98 17.87 441.17 20.89 ;
      RECT 438.28 16.52 441.17 16.69 ;
      RECT 439.35 20.89 441.17 21.06 ;
      RECT 439.35 21.06 439.52 22.4 ;
      RECT 440.21 21.06 440.38 22.4 ;
      RECT 440.64 16.69 441.17 17.87 ;
      RECT 438.28 16.69 438.45 19.14 ;
      RECT 437.1 18.735 437.63 18.905 ;
      RECT 437.1 18.905 437.27 19.14 ;
      RECT 437.1 16.86 437.27 18.735 ;
      RECT 441.8 18.735 442.33 18.905 ;
      RECT 441.68 21.835 441.85 22.595 ;
      RECT 439.19 22.595 441.85 22.765 ;
      RECT 351.525 15.345 354.235 15.515 ;
      RECT 351.525 14.065 354.235 14.235 ;
      RECT 355.175 11.505 357.885 11.675 ;
      RECT 358.105 13.165 358.275 20.525 ;
      RECT 358.105 10.605 358.275 12.565 ;
      RECT 362.22 17.505 366.595 18.205 ;
      RECT 362.22 18.205 362.92 25.335 ;
      RECT 365.895 18.205 366.595 25.335 ;
      RECT 362.22 25.335 366.595 26.045 ;
      RECT 368.815 17.505 373.19 18.205 ;
      RECT 368.815 18.205 369.515 25.335 ;
      RECT 372.49 18.205 373.19 25.335 ;
      RECT 368.815 25.335 373.19 26.045 ;
      RECT 375.285 17.35 377.305 18.1 ;
      RECT 405.96 16.52 408.85 16.69 ;
      RECT 405.96 17.87 406.15 20.89 ;
      RECT 405.96 20.89 407.78 21.06 ;
      RECT 406.75 21.06 406.92 22.4 ;
      RECT 407.61 21.06 407.78 22.4 ;
      RECT 405.96 16.69 406.49 17.87 ;
      RECT 408.68 16.69 408.85 19.14 ;
      RECT 405.62 21.975 406.15 22.145 ;
      RECT 405.62 16.85 405.79 21.975 ;
      RECT 403.92 12.03 404.09 12.56 ;
      RECT 407.11 12.03 407.28 12.56 ;
      RECT 402.925 18.735 403.455 18.905 ;
      RECT 402.925 16.965 403.68 17.135 ;
      RECT 402.925 17.135 403.095 18.735 ;
      RECT 402.925 18.905 403.095 20.825 ;
      RECT 402.925 20.825 403.13 21.835 ;
      RECT 402.46 16.775 402.63 17.385 ;
      RECT 402.46 16.605 405.31 16.775 ;
      RECT 405.14 16.775 405.31 17.385 ;
      RECT 405.68 12.77 405.85 14.59 ;
      RECT 403.92 13.525 404.09 14.59 ;
      RECT 403.92 12.78 404.09 13.355 ;
      RECT 404.8 18.735 405.33 18.905 ;
      RECT 405.28 21.835 405.45 22.595 ;
      RECT 405.28 22.595 407.94 22.765 ;
      RECT 404.8 17.155 404.97 18.735 ;
      RECT 404.8 20.825 405.45 21.835 ;
      RECT 406.59 22.765 407.94 22.77 ;
      RECT 404.8 18.905 404.97 20.825 ;
      RECT 403.88 17.155 404.17 19.575 ;
      RECT 403.63 19.865 403.93 20.5 ;
      RECT 403.63 19.575 404.17 19.865 ;
      RECT 403.63 20.5 404.17 20.655 ;
      RECT 403.64 22.67 404.17 22.84 ;
      RECT 403.76 20.655 404.17 22.67 ;
      RECT 404.1 20.07 404.63 20.24 ;
      RECT 404.34 17.155 404.51 20.07 ;
      RECT 407.11 13.54 407.28 14.59 ;
      RECT 407.11 12.78 407.28 13.31 ;
      RECT 406.8 16.86 407.67 17.87 ;
      RECT 406.8 17.87 407.33 18.905 ;
      RECT 441.095 30.475 441.625 30.645 ;
      RECT 413.485 30.475 414.02 30.645 ;
      RECT 413.485 30.645 413.665 30.735 ;
      RECT 413.485 28.325 413.665 30.475 ;
      RECT 432.35 30.475 432.885 30.645 ;
      RECT 432.705 30.645 432.885 30.735 ;
      RECT 435.535 30.475 436.07 30.645 ;
      RECT 435.535 30.645 435.715 30.79 ;
      RECT 435.535 28.69 435.715 30.475 ;
      RECT 441.445 30.645 441.625 30.79 ;
      RECT 441.445 28.69 441.625 30.475 ;
      RECT 444.5 20.815 444.67 22.835 ;
      RECT 413.485 28.15 444.675 28.155 ;
      RECT 413.91 28.325 444.675 28.33 ;
      RECT 432.705 28.335 432.885 30.475 ;
      RECT 402.46 28.155 444.675 28.325 ;
      RECT 432.705 28.33 444.675 28.335 ;
      RECT 402.46 17.555 402.63 28.155 ;
      RECT 435.535 28.335 441.625 28.69 ;
      RECT 444.495 22.835 444.675 28.15 ;
      RECT 408.87 12.03 409.04 12.56 ;
      RECT 408.87 12.98 409.04 13.31 ;
      RECT 408.02 18.225 408.35 19.075 ;
      RECT 408.1 17.615 408.27 18.225 ;
      RECT 408.87 13.54 409.04 14.59 ;
      RECT 409.5 18.735 410.03 18.905 ;
      RECT 409.86 18.905 410.03 19.14 ;
      RECT 409.86 16.86 410.03 18.735 ;
      RECT 410.63 13.54 410.8 14.59 ;
      RECT 410.63 12.03 410.8 12.56 ;
      RECT 410.63 12.78 410.8 13.31 ;
      RECT 411.41 17.24 411.58 19.95 ;
      RECT 411.53 16.89 414.58 17.025 ;
      RECT 411.37 16.72 414.74 16.89 ;
      RECT 410.22 21.96 410.75 22.13 ;
      RECT 410.105 23.31 410.635 23.48 ;
      RECT 410.325 22.13 410.635 23.31 ;
      RECT 410.44 16.85 410.61 21.96 ;
      RECT 412.39 12.03 412.56 12.56 ;
      RECT 412.39 12.98 412.56 13.31 ;
      RECT 413.75 20.04 414.295 20.21 ;
      RECT 413.75 20.21 413.92 20.24 ;
      RECT 413.75 17.24 413.92 20.04 ;
      RECT 412.97 17.24 413.14 19.95 ;
      RECT 411.815 20.04 412.36 20.21 ;
      RECT 412.19 20.21 412.36 20.24 ;
      RECT 412.19 17.24 412.36 20.04 ;
      RECT 412.39 13.54 412.56 14.59 ;
      RECT 417.26 16.52 420.15 16.69 ;
      RECT 419.96 17.87 420.15 20.89 ;
      RECT 418.33 20.89 420.15 21.06 ;
      RECT 418.33 21.06 418.5 22.4 ;
      RECT 419.19 21.06 419.36 22.4 ;
      RECT 417.26 16.69 417.43 19.14 ;
      RECT 419.62 16.69 420.15 17.87 ;
      RECT 414.15 12.03 414.32 12.56 ;
      RECT 414.15 12.98 414.32 13.31 ;
      RECT 417.67 12.03 417.84 12.56 ;
      RECT 415.91 12.03 416.08 12.56 ;
      RECT 415.91 12.98 416.08 13.31 ;
      RECT 417.67 12.98 417.84 13.31 ;
      RECT 419.43 12.03 419.6 12.56 ;
      RECT 419.43 12.98 419.6 13.31 ;
      RECT 414.53 17.24 414.7 19.95 ;
      RECT 414.15 13.54 414.32 14.59 ;
      RECT 415.36 21.96 415.89 22.13 ;
      RECT 415.475 23.31 416.005 23.48 ;
      RECT 415.475 22.13 415.785 23.31 ;
      RECT 415.5 16.85 415.67 21.96 ;
      RECT 416.08 18.735 416.61 18.905 ;
      RECT 416.08 18.905 416.25 19.14 ;
      RECT 416.08 16.86 416.25 18.735 ;
      RECT 297.36 15.69 298.37 15.78 ;
      RECT 296.97 14.105 297.14 15.52 ;
      RECT 296.83 16.385 297 17.3 ;
      RECT 296.4 17.485 296.57 17.83 ;
      RECT 296.4 17.3 297 17.485 ;
      RECT 297.3 11.935 298.31 12.105 ;
      RECT 297.36 14.83 298.37 15 ;
      RECT 297.36 17.54 298.37 17.71 ;
      RECT 297.36 16.16 298.37 16.33 ;
      RECT 297.3 10.175 298.31 10.345 ;
      RECT 297.3 11.055 298.31 11.225 ;
      RECT 297.36 17.08 298.37 17.25 ;
      RECT 297.36 16.62 298.37 16.79 ;
      RECT 300.415 13.325 300.585 15.785 ;
      RECT 298.62 16.42 298.79 18.435 ;
      RECT 300.415 10.84 300.585 12.28 ;
      RECT 300.845 11.905 301.855 12.105 ;
      RECT 302.085 15.655 302.255 16.755 ;
      RECT 302.085 14.275 302.255 15.375 ;
      RECT 300.415 16.42 300.585 18.255 ;
      RECT 300.845 17.82 302.255 17.99 ;
      RECT 302.085 17.99 302.255 18.775 ;
      RECT 300.845 10.615 301.855 10.785 ;
      RECT 300.845 12.335 301.855 12.505 ;
      RECT 300.845 17.36 301.855 17.53 ;
      RECT 300.845 14.05 301.855 14.22 ;
      RECT 300.845 13.59 301.855 13.76 ;
      RECT 300.845 15.43 301.855 15.6 ;
      RECT 300.845 16.81 301.855 16.98 ;
      RECT 300.845 11.475 301.855 11.645 ;
      RECT 300.845 14.51 301.855 14.68 ;
      RECT 300.845 14.97 301.855 15.14 ;
      RECT 300.845 16.35 301.855 16.52 ;
      RECT 300.845 15.89 301.855 16.06 ;
      RECT 300.845 11.045 301.855 11.215 ;
      RECT 307.575 16.265 307.745 27.99 ;
      RECT 308.155 14.675 309.505 14.845 ;
      RECT 308.155 17.795 309.505 17.965 ;
      RECT 308.155 16.235 309.505 16.405 ;
      RECT 308.155 13.115 309.505 13.285 ;
      RECT 308.155 11.555 309.505 11.725 ;
      RECT 304.315 16.625 307.025 16.795 ;
      RECT 304.315 14.345 307.025 14.515 ;
      RECT 304.315 12.065 307.025 12.235 ;
      RECT 308.155 13.895 309.505 14.065 ;
      RECT 308.155 12.335 309.505 12.505 ;
      RECT 308.155 10.775 309.505 10.945 ;
      RECT 308.155 17.015 309.505 17.185 ;
      RECT 314.055 14.95 314.225 18.47 ;
      RECT 312.825 13.23 313.155 14.25 ;
      RECT 314.625 17.085 315.635 17.255 ;
      RECT 314.415 12.625 315.545 12.795 ;
      RECT 314.415 12.795 314.585 13.65 ;
      RECT 309.725 15.52 310.375 16.125 ;
      RECT 314.625 10.065 315.635 10.235 ;
      RECT 314.625 15.185 315.635 15.355 ;
      RECT 314.625 14.725 315.635 14.895 ;
      RECT 314.625 16.165 315.635 16.335 ;
      RECT 314.875 13.705 315.545 13.875 ;
      RECT 314.625 15.705 315.635 15.875 ;
      RECT 314.625 17.545 315.635 17.715 ;
      RECT 319.885 13.665 321.02 14.335 ;
      RECT 319.885 15.02 320.475 15.19 ;
      RECT 319.885 15.19 320.055 15.515 ;
      RECT 319.885 14.845 320.055 15.02 ;
      RECT 319.885 18.085 320.475 18.255 ;
      RECT 319.885 18.255 320.055 18.53 ;
      RECT 319.885 17.86 320.055 18.085 ;
      RECT 319.885 16.71 320.475 16.88 ;
      RECT 319.885 16.88 320.055 17.35 ;
      RECT 319.885 16.68 320.055 16.71 ;
      RECT 330.005 16.71 330.705 16.88 ;
      RECT 330.535 16.655 330.705 16.71 ;
      RECT 330.535 18.445 330.705 18.505 ;
      RECT 330.005 18.275 330.705 18.445 ;
      RECT 330.535 16.88 330.705 18.275 ;
      RECT 331.075 16.72 331.775 16.89 ;
      RECT 331.075 16.655 331.245 16.72 ;
      RECT 331.075 18.29 331.245 18.505 ;
      RECT 331.075 18.12 331.775 18.29 ;
      RECT 331.075 16.89 331.245 18.12 ;
      RECT 330.005 14.915 330.705 15.085 ;
      RECT 330.535 15.085 330.705 15.515 ;
      RECT 330.005 13.725 330.705 13.895 ;
      RECT 330.535 13.665 330.705 13.725 ;
      RECT 330.535 13.895 330.705 14.915 ;
      RECT 331.075 15.285 331.775 15.455 ;
      RECT 331.075 15.455 331.245 15.515 ;
      RECT 331.075 13.705 331.775 13.875 ;
      RECT 331.075 13.665 331.245 13.705 ;
      RECT 331.075 13.875 331.245 15.285 ;
      RECT 341.42 16.89 341.895 17.325 ;
      RECT 340.89 16.72 341.895 16.89 ;
      RECT 341.42 16.655 341.895 16.72 ;
      RECT 341.305 13.705 341.895 13.875 ;
      RECT 341.725 13.875 341.895 14.335 ;
      RECT 341.725 13.665 341.895 13.705 ;
      RECT 341.195 18.12 341.895 18.29 ;
      RECT 341.725 18.29 341.895 18.505 ;
      RECT 341.725 17.835 341.895 18.12 ;
      RECT 341.195 15.095 341.895 15.265 ;
      RECT 341.725 15.265 341.895 15.515 ;
      RECT 341.725 14.845 341.895 15.095 ;
      RECT 347.875 10.225 350.585 10.395 ;
      RECT 347.875 11.505 350.585 11.675 ;
      RECT 347.875 14.065 350.585 14.235 ;
      RECT 347.875 16.625 350.585 16.795 ;
      RECT 347.875 17.905 350.585 18.075 ;
      RECT 347.875 15.345 350.585 15.515 ;
      RECT 347.875 12.785 350.585 12.955 ;
      RECT 355.175 10.225 357.885 10.395 ;
      RECT 355.175 17.905 357.885 18.075 ;
      RECT 355.175 15.345 357.885 15.515 ;
      RECT 355.175 12.785 357.885 12.955 ;
      RECT 354.035 17.515 354.625 17.685 ;
      RECT 354.035 14.955 354.625 15.125 ;
      RECT 354.455 13.175 354.625 14.955 ;
      RECT 354.035 15.735 354.625 15.905 ;
      RECT 354.455 15.125 354.625 15.735 ;
      RECT 354.035 18.295 354.625 18.465 ;
      RECT 354.455 15.905 354.625 17.515 ;
      RECT 354.455 17.685 354.625 18.295 ;
      RECT 354.455 18.465 354.625 27.115 ;
      RECT 355.175 16.625 357.885 16.795 ;
      RECT 355.175 14.065 357.885 14.235 ;
      RECT 351.525 17.905 354.235 18.075 ;
      RECT 351.525 16.625 354.235 16.795 ;
      RECT 268.3 11.1 268.81 11.43 ;
      RECT 268.29 17.7 268.82 17.87 ;
      RECT 268.3 17.51 268.81 17.7 ;
      RECT 264.23 11.1 264.74 11.43 ;
      RECT 264.23 17.51 264.74 17.84 ;
      RECT 264.3 13.85 264.67 17.51 ;
      RECT 264.3 11.43 264.67 13.59 ;
      RECT 263.41 13.59 264.67 13.85 ;
      RECT 263.41 13.85 263.58 17.345 ;
      RECT 263.41 11.6 263.58 13.59 ;
      RECT 266.6 11.6 266.77 17.345 ;
      RECT 266.72 11.26 267.25 11.43 ;
      RECT 267.08 11.43 267.25 11.6 ;
      RECT 267.15 12.61 267.32 17.345 ;
      RECT 267.08 11.6 267.32 12.61 ;
      RECT 266.06 11.43 266.43 17.51 ;
      RECT 265.99 11.1 266.5 11.43 ;
      RECT 265.99 17.51 266.5 17.84 ;
      RECT 267.49 11.43 267.86 17.51 ;
      RECT 267.42 11.1 267.93 11.43 ;
      RECT 267.42 17.51 267.93 17.84 ;
      RECT 263.53 11.26 264.06 11.43 ;
      RECT 263.89 11.43 264.06 11.6 ;
      RECT 263.89 11.6 264.13 13.42 ;
      RECT 265.72 11.6 265.89 13.21 ;
      RECT 265.61 10.39 266.14 10.56 ;
      RECT 265.63 10.56 266.14 10.59 ;
      RECT 265.63 10.26 266.14 10.39 ;
      RECT 267.39 10.39 268 10.56 ;
      RECT 267.39 10.56 267.9 10.59 ;
      RECT 267.39 10.26 267.9 10.39 ;
      RECT 268.03 11.6 268.2 13.21 ;
      RECT 263.96 14.33 264.13 17.04 ;
      RECT 265.72 14.33 265.89 17.04 ;
      RECT 265.72 13.83 265.89 14.16 ;
      RECT 268.03 14.33 268.2 17.04 ;
      RECT 268.03 13.83 268.2 14.16 ;
      RECT 269.25 11.43 269.62 17.51 ;
      RECT 269.18 11.1 269.69 11.43 ;
      RECT 269.17 17.7 269.7 17.87 ;
      RECT 269.18 17.51 269.69 17.7 ;
      RECT 261.72 18.04 275.225 18.21 ;
      RECT 262.795 18.21 267.285 18.265 ;
      RECT 271.255 17.27 275.225 18.04 ;
      RECT 271.255 13.9 271.425 17.27 ;
      RECT 275.055 13.9 275.225 17.27 ;
      RECT 269.79 11.6 269.96 13.42 ;
      RECT 270.955 12.9 272.885 13.18 ;
      RECT 272.08 13.18 272.36 13.76 ;
      RECT 272.08 13.76 272.885 14.04 ;
      RECT 272.715 11.72 272.885 12.9 ;
      RECT 272.355 14.04 272.885 14.16 ;
      RECT 270.955 11.72 271.125 12.9 ;
      RECT 272.715 14.16 272.885 16.92 ;
      RECT 271.835 11.72 272.005 12.73 ;
      RECT 274.475 12.725 274.94 13.005 ;
      RECT 273.26 13.52 273.54 13.72 ;
      RECT 274.475 14.21 274.645 16.92 ;
      RECT 272.53 13.35 273.54 13.52 ;
      RECT 274.475 11.72 274.645 12.725 ;
      RECT 274.66 13.005 274.94 13.72 ;
      RECT 273.26 13.72 274.94 13.77 ;
      RECT 274.475 14 274.885 14.21 ;
      RECT 273.26 13.77 274.885 14 ;
      RECT 269.79 14.33 269.96 17.04 ;
      RECT 271.835 14.21 272.005 16.92 ;
      RECT 273.82 13.35 274.49 13.52 ;
      RECT 273.595 14.21 273.765 16.92 ;
      RECT 275.355 11.72 275.525 12.73 ;
      RECT 279.37 12.9 279.9 12.95 ;
      RECT 279.38 13.07 281.675 13.12 ;
      RECT 279.37 12.95 281.675 13.07 ;
      RECT 275.635 14.17 275.805 18.92 ;
      RECT 276.12 12.95 276.79 13.12 ;
      RECT 276.26 12.91 276.79 12.95 ;
      RECT 277.07 12.95 277.74 13.12 ;
      RECT 277.26 13.12 277.79 13.32 ;
      RECT 278.07 12.95 279.1 13.15 ;
      RECT 278.07 13.15 278.6 13.32 ;
      RECT 278.535 13.66 280.865 13.74 ;
      RECT 275.985 13.49 280.735 13.57 ;
      RECT 275.985 13.57 280.865 13.66 ;
      RECT 278.275 14.17 278.445 18.92 ;
      RECT 280.035 14.17 280.205 18.92 ;
      RECT 276.515 14.17 276.685 18.92 ;
      RECT 277.395 14.17 277.565 18.92 ;
      RECT 279.155 14.17 279.325 18.92 ;
      RECT 281.465 14.17 281.635 18.92 ;
      RECT 283.225 14.17 283.395 18.92 ;
      RECT 280.915 14.17 281.085 18.92 ;
      RECT 281.505 13.49 282.175 13.66 ;
      RECT 283.805 13.9 283.975 18.9 ;
      RECT 290.655 16.855 292.085 17.025 ;
      RECT 290.655 15.25 290.825 16.855 ;
      RECT 290.655 14.445 291.395 14.615 ;
      RECT 290.655 14.615 290.825 14.97 ;
      RECT 290.655 13.97 290.825 14.445 ;
      RECT 290.655 17.195 290.825 18.08 ;
      RECT 291.055 13.665 292.085 13.915 ;
      RECT 290.245 13.265 292.505 13.435 ;
      RECT 290.245 25.915 292.505 26.085 ;
      RECT 292.335 13.435 292.505 25.915 ;
      RECT 290.245 13.435 290.415 25.915 ;
      RECT 291.055 16.305 292.085 16.475 ;
      RECT 288.755 13.97 288.925 14.97 ;
      RECT 287.525 16.855 288.925 17.025 ;
      RECT 288.755 15.25 288.925 16.855 ;
      RECT 288.755 17.195 288.925 18.08 ;
      RECT 291.075 15.025 292.15 15.195 ;
      RECT 287.525 13.745 288.535 13.915 ;
      RECT 287.525 15.025 288.535 15.195 ;
      RECT 287.525 16.305 288.535 16.475 ;
      RECT 287.525 10.125 288.535 10.295 ;
      RECT 291.075 10.105 292.085 10.275 ;
      RECT 296.4 13.46 299.22 13.52 ;
      RECT 296.32 13.52 299.22 13.64 ;
      RECT 296.32 16 296.58 16.9 ;
      RECT 296.4 16.9 296.58 17.085 ;
      RECT 299.04 13.64 299.22 19.485 ;
      RECT 296.4 18.055 296.58 19.485 ;
      RECT 296.4 14.585 296.58 16 ;
      RECT 296.32 13.64 296.58 14.585 ;
      RECT 296.4 19.485 299.22 19.77 ;
      RECT 297.36 14.14 298.79 14.31 ;
      RECT 297.36 14.05 298.37 14.14 ;
      RECT 298.62 14.31 298.79 15.725 ;
      RECT 296.97 15.52 298.37 15.69 ;
      RECT 247.195 19.135 253.325 19.5 ;
      RECT 246.66 18.04 249.86 18.855 ;
      RECT 245.23 18.855 249.86 18.88 ;
      RECT 250.73 18.21 255.935 18.88 ;
      RECT 245.23 19.03 253.325 19.135 ;
      RECT 245.23 18.88 255.935 18.92 ;
      RECT 245.23 18.92 255.82 19.03 ;
      RECT 243.39 14.33 243.56 17.04 ;
      RECT 243.39 13.83 243.56 14.16 ;
      RECT 245.7 14.33 245.87 17.04 ;
      RECT 245.15 14.33 245.32 17.04 ;
      RECT 250.65 11.725 250.82 17.345 ;
      RECT 246.58 11.725 246.75 17.345 ;
      RECT 250.11 11.43 250.48 17.51 ;
      RECT 250.04 11.1 250.55 11.43 ;
      RECT 250.03 17.51 250.56 18.67 ;
      RECT 246.92 11.43 247.29 17.51 ;
      RECT 246.85 11.1 247.36 11.43 ;
      RECT 246.85 17.51 247.36 17.84 ;
      RECT 250.99 11.43 251.36 17.51 ;
      RECT 250.91 11.26 251.44 11.43 ;
      RECT 250.92 17.51 251.43 17.84 ;
      RECT 250.92 11.1 251.43 11.26 ;
      RECT 246.04 11.43 246.41 17.51 ;
      RECT 245.97 11.1 246.48 11.43 ;
      RECT 245.96 17.51 246.49 18.67 ;
      RECT 248.46 11.26 248.99 11.43 ;
      RECT 248.82 11.6 249.06 17.345 ;
      RECT 248.82 11.43 248.99 11.6 ;
      RECT 248.34 11.6 248.51 17.345 ;
      RECT 249.23 11.43 249.6 17.51 ;
      RECT 249.16 11.1 249.67 11.43 ;
      RECT 249.16 17.51 249.67 17.84 ;
      RECT 247.8 11.43 248.17 17.51 ;
      RECT 247.73 11.1 248.24 11.43 ;
      RECT 247.73 17.51 248.24 17.84 ;
      RECT 249.77 11.6 249.94 13.21 ;
      RECT 247.46 11.6 247.63 13.21 ;
      RECT 249.77 13.83 249.94 14.16 ;
      RECT 247.46 13.83 247.63 14.16 ;
      RECT 249.15 10.39 249.68 10.56 ;
      RECT 249.17 10.56 249.68 10.59 ;
      RECT 249.17 10.26 249.68 10.39 ;
      RECT 251.53 11.6 251.7 13.42 ;
      RECT 249.77 14.33 249.94 17.04 ;
      RECT 247.46 14.33 247.63 17.04 ;
      RECT 251.53 14.33 251.7 17.04 ;
      RECT 256.15 11.725 256.32 17.345 ;
      RECT 252.96 11.725 253.13 17.345 ;
      RECT 257.37 11.43 257.74 17.51 ;
      RECT 257.3 11.1 257.81 11.43 ;
      RECT 257.3 17.51 257.81 17.84 ;
      RECT 256.49 11.43 256.86 17.51 ;
      RECT 256.42 11.1 256.93 11.43 ;
      RECT 256.41 17.7 256.94 17.87 ;
      RECT 256.42 17.51 256.93 17.7 ;
      RECT 253.3 11.43 253.67 17.51 ;
      RECT 253.23 11.1 253.74 11.43 ;
      RECT 253.22 17.7 253.75 17.87 ;
      RECT 253.23 17.51 253.74 17.7 ;
      RECT 255.54 11.1 256.05 11.43 ;
      RECT 255.54 17.51 256.05 17.84 ;
      RECT 255.61 13.85 255.98 17.51 ;
      RECT 255.61 11.43 255.98 13.59 ;
      RECT 254.72 13.59 255.98 13.85 ;
      RECT 254.72 13.85 254.89 17.345 ;
      RECT 254.72 11.6 254.89 13.59 ;
      RECT 252.42 11.43 252.79 17.51 ;
      RECT 252.35 11.1 252.86 11.43 ;
      RECT 252.34 17.7 252.87 17.87 ;
      RECT 252.35 17.51 252.86 17.7 ;
      RECT 254.18 11.43 254.55 17.51 ;
      RECT 254.11 11.1 254.62 11.43 ;
      RECT 254.11 17.51 254.62 17.84 ;
      RECT 252.08 11.6 252.25 13.42 ;
      RECT 253.84 11.6 254.01 13.21 ;
      RECT 255.27 11.6 255.44 13.42 ;
      RECT 257.03 11.6 257.2 13.21 ;
      RECT 252.08 14.33 252.25 17.04 ;
      RECT 255.27 14.33 255.44 17.04 ;
      RECT 253.84 14.33 254.01 17.04 ;
      RECT 253.84 13.83 254.01 14.16 ;
      RECT 257.03 14.33 257.2 17.04 ;
      RECT 257.03 13.83 257.2 14.16 ;
      RECT 257.91 11.725 258.08 17.345 ;
      RECT 261.65 11.725 261.82 17.345 ;
      RECT 261.99 11.43 262.36 17.51 ;
      RECT 261.92 11.1 262.43 11.43 ;
      RECT 261.91 17.7 262.44 17.87 ;
      RECT 261.92 17.51 262.43 17.7 ;
      RECT 258.25 11.43 258.62 17.51 ;
      RECT 258.18 11.1 258.69 11.43 ;
      RECT 259.035 18.875 259.565 19.045 ;
      RECT 258.18 17.515 259.44 17.84 ;
      RECT 258.18 17.51 258.69 17.515 ;
      RECT 259.035 17.84 259.44 18.875 ;
      RECT 261.11 11.43 261.48 17.51 ;
      RECT 261.04 11.1 261.55 11.43 ;
      RECT 261.04 18.465 261.575 18.635 ;
      RECT 261.04 17.51 261.55 18.465 ;
      RECT 259.34 11.6 259.51 17.345 ;
      RECT 259.68 11.43 260.05 17.51 ;
      RECT 259.61 11.1 260.12 11.43 ;
      RECT 259.61 17.51 260.12 17.84 ;
      RECT 262.87 11.43 263.24 17.51 ;
      RECT 262.8 11.1 263.31 11.43 ;
      RECT 262.8 17.51 263.31 17.84 ;
      RECT 259.15 10.39 259.68 10.56 ;
      RECT 259.16 10.56 259.67 10.59 ;
      RECT 259.16 10.26 259.67 10.39 ;
      RECT 258.79 14.33 258.96 17.04 ;
      RECT 258.79 11.6 258.96 13.42 ;
      RECT 260.22 11.6 260.39 13.21 ;
      RECT 260.22 14.33 260.39 17.04 ;
      RECT 260.22 13.83 260.39 14.16 ;
      RECT 260.77 14.33 260.94 17.04 ;
      RECT 262.53 14.33 262.7 17.04 ;
      RECT 262.53 11.6 262.7 13.21 ;
      RECT 260.77 11.6 260.94 13.42 ;
      RECT 262.53 13.83 262.7 14.16 ;
      RECT 264.84 11.725 265.01 17.345 ;
      RECT 268.91 11.725 269.08 17.345 ;
      RECT 265.18 11.43 265.55 17.51 ;
      RECT 265.1 11.26 265.63 11.43 ;
      RECT 265.11 17.51 265.62 17.84 ;
      RECT 265.11 11.1 265.62 11.26 ;
      RECT 268.37 11.43 268.74 17.51 ;
      RECT 144.865 17.295 145.395 17.465 ;
      RECT 145.025 11.43 145.395 17.295 ;
      RECT 144.955 17.465 145.395 17.51 ;
      RECT 142.715 11.43 143.085 17.51 ;
      RECT 142.645 11.1 143.155 11.43 ;
      RECT 142.645 17.51 143.155 17.84 ;
      RECT 145.905 11.43 146.275 17.51 ;
      RECT 145.825 11.26 146.355 11.43 ;
      RECT 145.835 17.51 146.345 17.84 ;
      RECT 145.835 11.1 146.345 11.26 ;
      RECT 147.325 11.6 147.495 17.345 ;
      RECT 146.785 11.43 147.155 17.51 ;
      RECT 146.715 11.1 147.225 11.43 ;
      RECT 146.705 17.51 147.235 18.27 ;
      RECT 141.835 11.43 142.205 17.51 ;
      RECT 141.765 11.1 142.275 11.43 ;
      RECT 141.765 17.51 142.275 17.84 ;
      RECT 142.375 11.6 142.545 13.21 ;
      RECT 142.375 13.83 142.545 14.16 ;
      RECT 146.445 11.6 146.615 13.21 ;
      RECT 144.135 11.6 144.305 13.42 ;
      RECT 144.685 11.6 144.855 13.42 ;
      RECT 146.445 13.83 146.615 14.16 ;
      RECT 142.375 14.33 142.545 17.04 ;
      RECT 144.685 14.33 144.855 17.04 ;
      RECT 146.445 14.33 146.615 17.04 ;
      RECT 144.135 14.33 144.305 17.04 ;
      RECT 148.875 15.14 149.545 15.31 ;
      RECT 151.23 11.36 151.76 11.53 ;
      RECT 151.23 11.53 151.4 13.505 ;
      RECT 151.23 10.795 151.4 11.36 ;
      RECT 152.81 15.225 157.66 15.395 ;
      RECT 148.02 11.6 148.19 13.41 ;
      RECT 150.65 14.185 154.32 14.355 ;
      RECT 150.47 10.86 151 11.03 ;
      RECT 153.91 10.86 154.44 11.03 ;
      RECT 150.65 11.03 150.82 14.185 ;
      RECT 150.65 10.855 150.82 10.86 ;
      RECT 154.15 11.03 154.32 14.185 ;
      RECT 154.15 10.855 154.32 10.86 ;
      RECT 152.01 10.795 152.18 14.185 ;
      RECT 153.57 10.795 153.74 14.185 ;
      RECT 148.755 17.235 149.645 17.615 ;
      RECT 152.91 16.505 157.66 16.675 ;
      RECT 150.06 14.655 155.27 14.825 ;
      RECT 144.215 18.44 148.19 18.66 ;
      RECT 131.405 18.04 139.275 18.21 ;
      RECT 148.02 13.83 148.19 18.04 ;
      RECT 147.405 18.04 148.19 18.44 ;
      RECT 144.215 18.04 146.535 18.44 ;
      RECT 144.395 19.135 144.775 21.15 ;
      RECT 144.395 18.66 144.775 18.855 ;
      RECT 131.995 18.21 132.885 18.3 ;
      RECT 136.68 19.135 142.81 19.5 ;
      RECT 140.145 18.04 143.345 18.855 ;
      RECT 140.145 18.855 144.775 18.88 ;
      RECT 134.07 18.21 139.275 18.88 ;
      RECT 136.68 19.03 144.775 19.135 ;
      RECT 134.07 18.88 144.775 18.92 ;
      RECT 134.185 18.92 144.775 19.03 ;
      RECT 149.87 15.35 152.43 18.455 ;
      RECT 158.075 14.42 160.095 15.17 ;
      RECT 164.01 13.63 165.335 14.04 ;
      RECT 162.48 17.255 166.855 17.965 ;
      RECT 162.48 17.965 163.18 25.095 ;
      RECT 166.155 17.965 166.855 25.095 ;
      RECT 162.48 25.095 166.855 25.795 ;
      RECT 169.075 17.255 173.45 17.965 ;
      RECT 169.075 17.965 169.775 25.095 ;
      RECT 172.75 17.965 173.45 25.095 ;
      RECT 169.075 25.095 173.45 25.795 ;
      RECT 170.595 13.63 171.92 14.04 ;
      RECT 216.555 17.255 220.93 17.965 ;
      RECT 216.555 17.965 217.255 25.095 ;
      RECT 220.23 17.965 220.93 25.095 ;
      RECT 216.555 25.095 220.93 25.795 ;
      RECT 218.085 13.63 219.41 14.04 ;
      RECT 224.67 13.63 225.995 14.04 ;
      RECT 223.15 17.255 227.525 17.965 ;
      RECT 223.15 17.965 223.85 25.095 ;
      RECT 226.825 17.965 227.525 25.095 ;
      RECT 223.15 25.095 227.525 25.795 ;
      RECT 232.345 15.225 237.195 15.395 ;
      RECT 229.91 14.42 231.93 15.17 ;
      RECT 232.345 16.505 237.095 16.675 ;
      RECT 238.245 11.36 238.775 11.53 ;
      RECT 238.605 11.53 238.775 13.505 ;
      RECT 238.605 10.795 238.775 11.36 ;
      RECT 235.685 14.185 239.355 14.355 ;
      RECT 235.565 10.86 236.095 11.03 ;
      RECT 239.005 10.86 239.535 11.03 ;
      RECT 235.685 11.03 235.855 14.185 ;
      RECT 235.685 10.855 235.855 10.86 ;
      RECT 239.185 11.03 239.355 14.185 ;
      RECT 239.185 10.855 239.355 10.86 ;
      RECT 236.265 10.795 236.435 14.185 ;
      RECT 237.825 10.795 237.995 14.185 ;
      RECT 234.735 14.655 239.945 14.825 ;
      RECT 237.575 15.35 240.135 18.455 ;
      RECT 244.27 11.725 244.44 17.345 ;
      RECT 243.73 11.43 244.1 17.51 ;
      RECT 243.65 11.26 244.18 11.43 ;
      RECT 243.66 17.51 244.17 17.84 ;
      RECT 243.66 11.1 244.17 11.26 ;
      RECT 244.54 11.1 245.05 11.43 ;
      RECT 244.54 17.51 245.05 17.84 ;
      RECT 244.61 17.295 245.14 17.465 ;
      RECT 244.61 11.43 244.98 17.295 ;
      RECT 244.61 17.465 245.05 17.51 ;
      RECT 242.51 11.6 242.68 17.345 ;
      RECT 242.85 11.43 243.22 17.51 ;
      RECT 242.78 11.1 243.29 11.43 ;
      RECT 242.77 17.51 243.3 18.27 ;
      RECT 241.815 11.6 241.985 13.41 ;
      RECT 243.39 11.6 243.56 13.21 ;
      RECT 245.7 11.6 245.87 13.42 ;
      RECT 245.15 11.6 245.32 13.42 ;
      RECT 240.46 15.14 241.13 15.31 ;
      RECT 240.36 17.235 241.25 17.615 ;
      RECT 241.815 18.44 245.79 18.66 ;
      RECT 250.73 18.04 258.6 18.21 ;
      RECT 241.815 13.83 241.985 18.04 ;
      RECT 241.815 18.04 242.6 18.44 ;
      RECT 243.47 18.04 245.79 18.44 ;
      RECT 245.23 19.135 245.61 21.15 ;
      RECT 245.23 18.66 245.61 18.855 ;
      RECT 257.12 18.21 258.01 18.3 ;
      RECT 123.865 10.39 124.395 10.56 ;
      RECT 123.865 10.56 124.375 10.59 ;
      RECT 123.865 10.26 124.375 10.39 ;
      RECT 120.045 14.33 120.215 17.04 ;
      RECT 121.805 14.33 121.975 17.04 ;
      RECT 121.805 13.83 121.975 14.16 ;
      RECT 124.115 14.33 124.285 17.04 ;
      RECT 124.115 13.83 124.285 14.16 ;
      RECT 124.995 11.725 125.165 17.345 ;
      RECT 128.185 11.725 128.355 17.345 ;
      RECT 125.265 11.1 125.775 11.43 ;
      RECT 125.265 17.51 125.775 17.84 ;
      RECT 125.335 13.85 125.705 17.51 ;
      RECT 125.335 11.43 125.705 13.59 ;
      RECT 125.335 13.59 126.595 13.85 ;
      RECT 126.425 13.85 126.595 17.345 ;
      RECT 126.425 11.6 126.595 13.59 ;
      RECT 128.525 11.43 128.895 17.51 ;
      RECT 128.455 11.1 128.965 11.43 ;
      RECT 128.43 18.465 128.965 18.635 ;
      RECT 128.455 17.51 128.965 18.465 ;
      RECT 124.455 11.43 124.825 17.51 ;
      RECT 124.375 11.26 124.905 11.43 ;
      RECT 124.385 17.51 124.895 17.84 ;
      RECT 124.385 11.1 124.895 11.26 ;
      RECT 127.645 11.43 128.015 17.51 ;
      RECT 127.575 11.1 128.085 11.43 ;
      RECT 127.565 17.7 128.095 17.87 ;
      RECT 127.575 17.51 128.085 17.7 ;
      RECT 129.955 11.43 130.325 17.51 ;
      RECT 129.885 11.1 130.395 11.43 ;
      RECT 129.885 17.51 130.395 17.84 ;
      RECT 126.765 11.43 127.135 17.51 ;
      RECT 126.695 11.1 127.205 11.43 ;
      RECT 126.695 17.51 127.205 17.84 ;
      RECT 127.305 11.6 127.475 13.21 ;
      RECT 125.945 11.26 126.475 11.43 ;
      RECT 125.945 11.43 126.115 11.6 ;
      RECT 125.875 11.6 126.115 13.42 ;
      RECT 127.305 13.83 127.475 14.16 ;
      RECT 129.065 11.6 129.235 13.42 ;
      RECT 129.615 11.6 129.785 13.21 ;
      RECT 129.615 13.83 129.785 14.16 ;
      RECT 127.305 14.33 127.475 17.04 ;
      RECT 125.875 14.33 126.045 17.04 ;
      RECT 129.065 14.33 129.235 17.04 ;
      RECT 129.615 14.33 129.785 17.04 ;
      RECT 130.325 10.39 130.855 10.56 ;
      RECT 130.335 10.56 130.845 10.59 ;
      RECT 130.335 10.26 130.845 10.39 ;
      RECT 131.925 11.725 132.095 17.345 ;
      RECT 131.385 11.43 131.755 17.51 ;
      RECT 131.315 11.1 131.825 11.43 ;
      RECT 130.44 18.875 130.97 19.045 ;
      RECT 130.565 17.515 131.825 17.84 ;
      RECT 131.315 17.51 131.825 17.515 ;
      RECT 130.565 17.84 130.97 18.875 ;
      RECT 132.265 11.43 132.635 17.51 ;
      RECT 132.195 11.1 132.705 11.43 ;
      RECT 132.195 17.51 132.705 17.84 ;
      RECT 133.145 11.43 133.515 17.51 ;
      RECT 133.075 11.1 133.585 11.43 ;
      RECT 133.065 17.7 133.595 17.87 ;
      RECT 133.075 17.51 133.585 17.7 ;
      RECT 130.495 11.6 130.665 17.345 ;
      RECT 132.805 14.33 132.975 17.04 ;
      RECT 131.045 14.33 131.215 17.04 ;
      RECT 132.805 11.6 132.975 13.21 ;
      RECT 131.045 11.6 131.215 13.42 ;
      RECT 132.805 13.83 132.975 14.16 ;
      RECT 134.565 14.33 134.735 17.04 ;
      RECT 134.565 11.6 134.735 13.42 ;
      RECT 133.685 11.725 133.855 17.345 ;
      RECT 133.955 17.51 134.465 17.84 ;
      RECT 133.955 11.1 134.465 11.43 ;
      RECT 134.025 13.85 134.395 17.51 ;
      RECT 134.025 11.43 134.395 13.59 ;
      RECT 134.025 13.59 135.285 13.85 ;
      RECT 135.115 13.85 135.285 17.345 ;
      RECT 135.115 11.6 135.285 13.59 ;
      RECT 135.385 17.51 135.895 17.84 ;
      RECT 135.455 11.43 135.825 17.51 ;
      RECT 135.385 11.1 135.895 11.43 ;
      RECT 139.185 11.725 139.355 17.345 ;
      RECT 136.875 11.725 137.045 17.345 ;
      RECT 138.645 11.43 139.015 17.51 ;
      RECT 138.565 11.26 139.095 11.43 ;
      RECT 138.575 17.51 139.085 17.84 ;
      RECT 138.575 11.1 139.085 11.26 ;
      RECT 137.215 11.43 137.585 17.51 ;
      RECT 137.145 11.1 137.655 11.43 ;
      RECT 137.135 17.7 137.665 17.87 ;
      RECT 137.145 17.51 137.655 17.7 ;
      RECT 139.525 11.43 139.895 17.51 ;
      RECT 139.455 11.1 139.965 11.43 ;
      RECT 139.445 17.51 139.975 18.67 ;
      RECT 136.335 11.43 136.705 17.51 ;
      RECT 136.265 11.1 136.775 11.43 ;
      RECT 136.255 17.7 136.785 17.87 ;
      RECT 136.265 17.51 136.775 17.7 ;
      RECT 141.015 11.26 141.545 11.43 ;
      RECT 140.945 11.6 141.185 17.345 ;
      RECT 141.015 11.43 141.185 11.6 ;
      RECT 141.495 11.6 141.665 17.345 ;
      RECT 140.405 11.43 140.775 17.51 ;
      RECT 140.335 11.1 140.845 11.43 ;
      RECT 140.335 17.51 140.845 17.84 ;
      RECT 135.995 11.6 136.165 13.21 ;
      RECT 135.995 13.83 136.165 14.16 ;
      RECT 137.755 11.6 137.925 13.42 ;
      RECT 138.305 11.6 138.475 13.42 ;
      RECT 140.065 11.6 140.235 13.21 ;
      RECT 140.065 13.83 140.235 14.16 ;
      RECT 140.325 10.39 140.855 10.56 ;
      RECT 140.325 10.56 140.835 10.59 ;
      RECT 140.325 10.26 140.835 10.39 ;
      RECT 135.995 14.33 136.165 17.04 ;
      RECT 137.755 14.33 137.925 17.04 ;
      RECT 138.305 14.33 138.475 17.04 ;
      RECT 140.065 14.33 140.235 17.04 ;
      RECT 143.255 11.725 143.425 17.345 ;
      RECT 145.565 11.725 145.735 17.345 ;
      RECT 143.595 11.43 143.965 17.51 ;
      RECT 143.525 11.1 144.035 11.43 ;
      RECT 143.515 17.51 144.045 18.67 ;
      RECT 144.955 11.1 145.465 11.43 ;
      RECT 144.955 17.51 145.465 17.84 ;
      RECT 88.15 16.35 89.16 16.52 ;
      RECT 88.15 15.89 89.16 16.06 ;
      RECT 88.15 11.045 89.16 11.215 ;
      RECT 90.785 13.64 90.965 19.485 ;
      RECT 90.785 13.46 93.605 13.52 ;
      RECT 90.785 13.52 93.685 13.64 ;
      RECT 93.425 16 93.685 16.9 ;
      RECT 93.425 16.9 93.605 17.085 ;
      RECT 93.425 18.055 93.605 19.485 ;
      RECT 93.425 14.585 93.605 16 ;
      RECT 93.425 13.64 93.685 14.585 ;
      RECT 90.785 19.485 93.605 19.77 ;
      RECT 91.215 16.42 91.385 18.435 ;
      RECT 91.215 14.14 92.645 14.31 ;
      RECT 91.635 14.05 92.645 14.14 ;
      RECT 91.215 14.31 91.385 15.725 ;
      RECT 91.635 15.52 93.035 15.69 ;
      RECT 91.635 15.69 92.645 15.78 ;
      RECT 92.865 14.105 93.035 15.52 ;
      RECT 93.005 16.385 93.175 17.3 ;
      RECT 93.435 17.485 93.605 17.83 ;
      RECT 93.005 17.3 93.605 17.485 ;
      RECT 91.695 11.935 92.705 12.105 ;
      RECT 91.635 14.83 92.645 15 ;
      RECT 91.635 17.54 92.645 17.71 ;
      RECT 91.635 16.16 92.645 16.33 ;
      RECT 91.695 10.175 92.705 10.345 ;
      RECT 91.695 11.055 92.705 11.225 ;
      RECT 91.635 17.08 92.645 17.25 ;
      RECT 91.635 16.62 92.645 16.79 ;
      RECT 97.92 16.855 99.35 17.025 ;
      RECT 99.18 15.25 99.35 16.855 ;
      RECT 98.61 14.445 99.35 14.615 ;
      RECT 99.18 14.615 99.35 14.97 ;
      RECT 99.18 13.97 99.35 14.445 ;
      RECT 99.18 17.195 99.35 18.08 ;
      RECT 97.92 13.665 98.95 13.915 ;
      RECT 97.5 13.265 99.76 13.435 ;
      RECT 97.5 25.915 99.76 26.085 ;
      RECT 97.5 13.435 97.67 25.915 ;
      RECT 99.59 13.435 99.76 25.915 ;
      RECT 97.855 15.025 98.93 15.195 ;
      RECT 97.92 16.305 98.95 16.475 ;
      RECT 97.92 10.105 98.93 10.275 ;
      RECT 101.08 13.97 101.25 14.97 ;
      RECT 101.08 16.855 102.48 17.025 ;
      RECT 101.08 15.25 101.25 16.855 ;
      RECT 101.08 17.195 101.25 18.08 ;
      RECT 101.47 13.745 102.48 13.915 ;
      RECT 101.47 15.025 102.48 15.195 ;
      RECT 101.47 16.305 102.48 16.475 ;
      RECT 106.61 14.17 106.78 18.92 ;
      RECT 101.47 10.125 102.48 10.295 ;
      RECT 106.03 13.9 106.2 18.9 ;
      RECT 110.105 12.9 110.635 12.95 ;
      RECT 108.33 13.07 110.625 13.12 ;
      RECT 108.33 12.95 110.635 13.07 ;
      RECT 108.92 14.17 109.09 18.92 ;
      RECT 108.37 14.17 108.54 18.92 ;
      RECT 112.265 12.95 112.935 13.12 ;
      RECT 112.215 13.12 112.745 13.32 ;
      RECT 110.905 12.95 111.935 13.15 ;
      RECT 111.405 13.15 111.935 13.32 ;
      RECT 107.83 13.49 108.5 13.66 ;
      RECT 109.14 13.66 111.47 13.74 ;
      RECT 109.27 13.49 114.02 13.57 ;
      RECT 109.14 13.57 114.02 13.66 ;
      RECT 111.56 14.17 111.73 18.92 ;
      RECT 109.8 14.17 109.97 18.92 ;
      RECT 112.44 14.17 112.61 18.92 ;
      RECT 110.68 14.17 110.85 18.92 ;
      RECT 114.78 18.04 128.285 18.21 ;
      RECT 122.72 18.21 127.21 18.265 ;
      RECT 114.78 17.27 118.75 18.04 ;
      RECT 118.58 13.9 118.75 17.27 ;
      RECT 114.78 13.9 114.95 17.27 ;
      RECT 114.48 11.72 114.65 12.73 ;
      RECT 115.065 12.725 115.53 13.005 ;
      RECT 116.465 13.52 116.745 13.72 ;
      RECT 115.36 14.21 115.53 16.92 ;
      RECT 116.465 13.35 117.475 13.52 ;
      RECT 115.36 11.72 115.53 12.725 ;
      RECT 115.065 13.005 115.345 13.72 ;
      RECT 115.065 13.72 116.745 13.77 ;
      RECT 115.12 14 115.53 14.21 ;
      RECT 115.12 13.77 116.745 14 ;
      RECT 114.2 14.17 114.37 18.92 ;
      RECT 113.215 12.95 113.885 13.12 ;
      RECT 113.215 12.91 113.745 12.95 ;
      RECT 115.515 13.35 116.185 13.52 ;
      RECT 116.24 14.21 116.41 16.92 ;
      RECT 113.32 14.17 113.49 18.92 ;
      RECT 118 14.21 118.17 16.92 ;
      RECT 117.12 13.76 117.925 14.04 ;
      RECT 117.645 13.18 117.925 13.76 ;
      RECT 117.12 12.9 119.05 13.18 ;
      RECT 117.12 14.04 117.65 14.16 ;
      RECT 117.12 11.72 117.29 12.9 ;
      RECT 117.12 14.16 117.29 16.92 ;
      RECT 118.88 11.72 119.05 12.9 ;
      RECT 118 11.72 118.17 12.73 ;
      RECT 120.925 11.725 121.095 17.345 ;
      RECT 120.385 11.43 120.755 17.51 ;
      RECT 120.315 11.1 120.825 11.43 ;
      RECT 120.305 17.7 120.835 17.87 ;
      RECT 120.315 17.51 120.825 17.7 ;
      RECT 121.265 11.43 121.635 17.51 ;
      RECT 121.195 11.1 121.705 11.43 ;
      RECT 121.185 17.7 121.715 17.87 ;
      RECT 121.195 17.51 121.705 17.7 ;
      RECT 123.235 11.6 123.405 17.345 ;
      RECT 122.755 11.26 123.285 11.43 ;
      RECT 122.755 11.43 122.925 11.6 ;
      RECT 122.685 12.61 122.855 17.345 ;
      RECT 122.685 11.6 122.925 12.61 ;
      RECT 123.575 11.43 123.945 17.51 ;
      RECT 123.505 11.1 124.015 11.43 ;
      RECT 123.505 17.51 124.015 17.84 ;
      RECT 122.145 11.43 122.515 17.51 ;
      RECT 122.075 11.1 122.585 11.43 ;
      RECT 122.075 17.51 122.585 17.84 ;
      RECT 120.045 11.6 120.215 13.42 ;
      RECT 121.805 11.6 121.975 13.21 ;
      RECT 122.005 10.39 122.615 10.56 ;
      RECT 122.105 10.56 122.615 10.59 ;
      RECT 122.105 10.26 122.615 10.39 ;
      RECT 124.115 11.6 124.285 13.21 ;
      RECT 441.77 9.05 441.94 13.24 ;
      RECT 442.14 9.05 442.31 13.24 ;
      RECT 442.48 9.55 442.65 10.56 ;
      RECT 12.7 17.35 14.72 18.1 ;
      RECT 16.815 17.505 21.19 18.205 ;
      RECT 16.815 18.205 17.515 25.335 ;
      RECT 20.49 18.205 21.19 25.335 ;
      RECT 16.815 25.335 21.19 26.045 ;
      RECT 23.41 17.505 27.785 18.205 ;
      RECT 23.41 18.205 24.11 25.335 ;
      RECT 27.085 18.205 27.785 25.335 ;
      RECT 23.41 25.335 27.785 26.045 ;
      RECT 31.73 13.165 31.9 20.525 ;
      RECT 31.73 10.605 31.9 12.565 ;
      RECT 32.12 10.225 34.83 10.395 ;
      RECT 32.12 17.905 34.83 18.075 ;
      RECT 32.12 15.345 34.83 15.515 ;
      RECT 32.12 12.785 34.83 12.955 ;
      RECT 35.38 17.515 35.97 17.685 ;
      RECT 35.38 14.955 35.97 15.125 ;
      RECT 35.38 13.175 35.55 14.955 ;
      RECT 35.38 15.735 35.97 15.905 ;
      RECT 35.38 15.125 35.55 15.735 ;
      RECT 35.38 18.295 35.97 18.465 ;
      RECT 35.38 15.905 35.55 17.515 ;
      RECT 35.38 17.685 35.55 18.295 ;
      RECT 35.38 18.465 35.55 27.115 ;
      RECT 32.12 16.625 34.83 16.795 ;
      RECT 32.12 14.065 34.83 14.235 ;
      RECT 35.77 17.905 38.48 18.075 ;
      RECT 35.77 16.625 38.48 16.795 ;
      RECT 35.77 15.345 38.48 15.515 ;
      RECT 35.77 14.065 38.48 14.235 ;
      RECT 32.12 11.505 34.83 11.675 ;
      RECT 39.42 10.225 42.13 10.395 ;
      RECT 39.42 11.505 42.13 11.675 ;
      RECT 39.42 14.065 42.13 14.235 ;
      RECT 39.42 16.625 42.13 16.795 ;
      RECT 39.42 17.905 42.13 18.075 ;
      RECT 39.42 15.345 42.13 15.515 ;
      RECT 39.42 12.785 42.13 12.955 ;
      RECT 48.11 16.89 48.585 17.325 ;
      RECT 48.11 16.72 49.115 16.89 ;
      RECT 48.11 16.655 48.585 16.72 ;
      RECT 48.11 13.705 48.7 13.875 ;
      RECT 48.11 13.875 48.28 14.335 ;
      RECT 48.11 13.665 48.28 13.705 ;
      RECT 48.11 18.12 48.81 18.29 ;
      RECT 48.11 18.29 48.28 18.505 ;
      RECT 48.11 17.835 48.28 18.12 ;
      RECT 48.11 15.095 48.81 15.265 ;
      RECT 48.11 15.265 48.28 15.515 ;
      RECT 48.11 14.845 48.28 15.095 ;
      RECT 59.3 18.275 60 18.445 ;
      RECT 59.3 18.445 59.47 18.505 ;
      RECT 59.3 16.71 60 16.88 ;
      RECT 59.3 16.655 59.47 16.71 ;
      RECT 59.3 16.88 59.47 18.275 ;
      RECT 58.23 16.72 58.93 16.89 ;
      RECT 58.76 16.655 58.93 16.72 ;
      RECT 58.76 18.29 58.93 18.505 ;
      RECT 58.23 18.12 58.93 18.29 ;
      RECT 58.76 16.89 58.93 18.12 ;
      RECT 59.3 14.915 60 15.085 ;
      RECT 59.3 15.085 59.47 15.515 ;
      RECT 59.3 13.725 60 13.895 ;
      RECT 59.3 13.665 59.47 13.725 ;
      RECT 59.3 13.895 59.47 14.915 ;
      RECT 58.23 15.285 58.93 15.455 ;
      RECT 58.76 15.455 58.93 15.515 ;
      RECT 58.23 13.705 58.93 13.875 ;
      RECT 58.76 13.665 58.93 13.705 ;
      RECT 58.76 13.875 58.93 15.285 ;
      RECT 68.985 13.665 70.12 14.335 ;
      RECT 69.53 18.085 70.12 18.255 ;
      RECT 69.95 18.255 70.12 18.53 ;
      RECT 69.95 17.86 70.12 18.085 ;
      RECT 69.53 16.71 70.12 16.88 ;
      RECT 69.95 16.88 70.12 17.35 ;
      RECT 69.95 16.68 70.12 16.71 ;
      RECT 69.53 15.02 70.12 15.19 ;
      RECT 69.95 15.19 70.12 15.515 ;
      RECT 69.95 14.845 70.12 15.02 ;
      RECT 75.78 14.95 75.95 18.47 ;
      RECT 76.85 13.23 77.18 14.25 ;
      RECT 74.37 17.085 75.38 17.255 ;
      RECT 74.46 12.625 75.59 12.795 ;
      RECT 75.42 12.795 75.59 13.65 ;
      RECT 74.37 10.065 75.38 10.235 ;
      RECT 74.37 15.185 75.38 15.355 ;
      RECT 74.37 14.725 75.38 14.895 ;
      RECT 74.37 16.165 75.38 16.335 ;
      RECT 74.46 13.705 75.13 13.875 ;
      RECT 74.37 17.545 75.38 17.715 ;
      RECT 74.37 15.705 75.38 15.875 ;
      RECT 82.26 16.265 82.43 27.99 ;
      RECT 79.63 15.52 80.28 16.125 ;
      RECT 80.5 14.675 81.85 14.845 ;
      RECT 80.5 17.795 81.85 17.965 ;
      RECT 80.5 16.235 81.85 16.405 ;
      RECT 80.5 13.115 81.85 13.285 ;
      RECT 80.5 11.555 81.85 11.725 ;
      RECT 82.98 16.625 85.69 16.795 ;
      RECT 82.98 14.345 85.69 14.515 ;
      RECT 82.98 12.065 85.69 12.235 ;
      RECT 80.5 13.895 81.85 14.065 ;
      RECT 80.5 12.335 81.85 12.505 ;
      RECT 80.5 10.775 81.85 10.945 ;
      RECT 80.5 17.015 81.85 17.185 ;
      RECT 89.42 13.325 89.59 15.785 ;
      RECT 89.42 10.84 89.59 12.28 ;
      RECT 88.15 11.905 89.16 12.105 ;
      RECT 87.75 15.655 87.92 16.755 ;
      RECT 87.75 14.275 87.92 15.375 ;
      RECT 89.42 16.42 89.59 18.255 ;
      RECT 87.75 17.82 89.16 17.99 ;
      RECT 87.75 17.99 87.92 18.775 ;
      RECT 88.15 10.615 89.16 10.785 ;
      RECT 88.15 12.335 89.16 12.505 ;
      RECT 88.15 17.36 89.16 17.53 ;
      RECT 88.15 14.05 89.16 14.22 ;
      RECT 88.15 13.59 89.16 13.76 ;
      RECT 88.15 15.43 89.16 15.6 ;
      RECT 88.15 16.81 89.16 16.98 ;
      RECT 88.15 11.475 89.16 11.645 ;
      RECT 88.15 14.51 89.16 14.68 ;
      RECT 88.15 14.97 89.16 15.14 ;
      RECT 410.97 8.68 411.34 14.76 ;
      RECT 410.9 14.76 411.41 15.09 ;
      RECT 410.02 8.35 410.53 8.68 ;
      RECT 410.02 14.76 410.53 15.09 ;
      RECT 410.09 8.68 410.46 14.76 ;
      RECT 408.26 8.35 409.65 8.68 ;
      RECT 408.26 14.76 409.65 15.09 ;
      RECT 409.21 8.68 409.58 14.76 ;
      RECT 408.33 8.68 408.7 14.76 ;
      RECT 413.27 8.85 413.44 14.59 ;
      RECT 411.51 8.85 411.68 14.59 ;
      RECT 409.75 8.83 409.92 14.59 ;
      RECT 410.63 9.15 410.8 11.86 ;
      RECT 408.87 9.15 409.04 11.86 ;
      RECT 412.39 9.15 412.56 11.86 ;
      RECT 417.06 8.35 417.57 8.68 ;
      RECT 417.13 8.68 417.5 14.76 ;
      RECT 417.06 14.76 417.57 15.09 ;
      RECT 416.25 8.68 416.62 14.76 ;
      RECT 415.37 8.68 415.74 14.76 ;
      RECT 416.18 8.65 416.69 8.68 ;
      RECT 415.295 8.35 416.69 8.65 ;
      RECT 415.295 8.65 415.805 8.68 ;
      RECT 416.18 14.76 416.69 14.79 ;
      RECT 415.3 14.79 416.69 15.09 ;
      RECT 415.3 14.76 415.81 14.79 ;
      RECT 418.89 8.68 419.26 14.76 ;
      RECT 419.77 8.68 420.14 14.76 ;
      RECT 418.82 8.65 419.33 8.68 ;
      RECT 418.82 14.76 419.33 14.79 ;
      RECT 418.82 8.35 420.21 8.65 ;
      RECT 419.7 8.65 420.21 8.68 ;
      RECT 418.82 14.79 420.21 15.09 ;
      RECT 419.7 14.76 420.21 14.79 ;
      RECT 417.94 8.35 418.45 8.68 ;
      RECT 418.01 8.68 418.38 14.76 ;
      RECT 417.94 14.76 418.45 15.09 ;
      RECT 416.79 8.85 416.96 14.59 ;
      RECT 418.55 8.85 418.72 14.59 ;
      RECT 415.03 8.85 415.2 14.59 ;
      RECT 417.67 9.15 417.84 11.86 ;
      RECT 415.91 9.15 416.08 11.86 ;
      RECT 414.15 9.15 414.32 11.86 ;
      RECT 419.43 9.15 419.6 11.86 ;
      RECT 424.1 8.35 424.61 8.68 ;
      RECT 424.17 8.68 424.54 14.76 ;
      RECT 424.1 14.76 424.61 15.09 ;
      RECT 423.29 8.68 423.66 14.76 ;
      RECT 422.41 8.68 422.78 14.76 ;
      RECT 423.22 8.65 423.73 8.68 ;
      RECT 423.22 14.76 423.73 14.79 ;
      RECT 422.335 8.35 423.73 8.65 ;
      RECT 422.335 8.65 422.845 8.68 ;
      RECT 422.34 14.79 423.73 15.09 ;
      RECT 422.34 14.76 422.85 14.79 ;
      RECT 420.65 8.68 421.02 14.76 ;
      RECT 421.53 8.68 421.9 14.76 ;
      RECT 420.58 8.65 421.09 8.68 ;
      RECT 420.58 14.76 421.09 14.79 ;
      RECT 420.58 8.35 421.97 8.65 ;
      RECT 421.46 8.65 421.97 8.68 ;
      RECT 420.58 14.79 421.97 15.09 ;
      RECT 421.46 14.76 421.97 14.79 ;
      RECT 423.83 8.85 424 14.59 ;
      RECT 420.31 8.85 420.48 14.59 ;
      RECT 422.07 8.85 422.24 14.59 ;
      RECT 424.71 9.15 424.88 11.86 ;
      RECT 422.95 9.15 423.12 11.86 ;
      RECT 421.19 9.15 421.36 11.86 ;
      RECT 430.77 9.96 430.94 11.015 ;
      RECT 428.21 9.96 428.38 11.015 ;
      RECT 402.46 15.87 402.63 16.435 ;
      RECT 402.46 15.7 438.335 15.87 ;
      RECT 402.85 15.685 442.22 15.7 ;
      RECT 434.46 15.625 442.22 15.685 ;
      RECT 425.405 14.6 430.36 15.685 ;
      RECT 434.46 13.565 443.2 15.625 ;
      RECT 426.97 13.54 430.36 14.6 ;
      RECT 434.46 13.34 438.335 13.565 ;
      RECT 429.83 13.14 430.36 13.54 ;
      RECT 435.74 13.28 438.335 13.34 ;
      RECT 434.46 13.14 434.99 13.34 ;
      RECT 435.74 13.14 438.355 13.28 ;
      RECT 426.97 13.125 429.1 13.54 ;
      RECT 437.465 13.11 438.355 13.14 ;
      RECT 425.405 13.08 426.34 14.6 ;
      RECT 402.46 12.78 402.63 15.7 ;
      RECT 437.485 12.165 438.335 13.11 ;
      RECT 426.97 12.09 428.38 13.125 ;
      RECT 436.44 12.09 436.61 13.14 ;
      RECT 437.465 11.275 438.355 12.165 ;
      RECT 437.485 9.31 438.335 11.275 ;
      RECT 437.465 8.93 438.355 9.31 ;
      RECT 426.97 8.93 427.5 12.09 ;
      RECT 426.97 8.42 438.355 8.93 ;
      RECT 428.09 9.49 436.73 9.71 ;
      RECT 428.255 9.18 436.705 9.49 ;
      RECT 429.49 9.96 429.66 13.1 ;
      RECT 432.42 11.45 432.95 11.62 ;
      RECT 432.6 11.62 432.77 14.73 ;
      RECT 432.6 9.96 432.77 11.45 ;
      RECT 433.88 9.96 434.05 11.015 ;
      RECT 431.9 11.82 432.43 11.99 ;
      RECT 432.05 9.96 432.22 11.82 ;
      RECT 432.05 11.99 432.22 14.73 ;
      RECT 436.44 9.96 436.61 11.015 ;
      RECT 435.16 12.54 435.74 12.71 ;
      RECT 435.16 12.71 435.33 13.1 ;
      RECT 435.16 9.96 435.33 12.54 ;
      RECT 439.09 8.01 443.2 8.88 ;
      RECT 438.73 9.54 439.26 9.71 ;
      RECT 443.03 8.88 443.2 9.54 ;
      RECT 442.82 9.54 443.35 9.71 ;
      RECT 439.09 8.88 439.26 9.54 ;
      RECT 439.09 10.56 439.38 10.73 ;
      RECT 439.09 9.71 439.26 10.56 ;
      RECT 439.09 10.73 439.81 11.06 ;
      RECT 442.48 10.73 443.2 11.06 ;
      RECT 443.03 9.71 443.2 10.73 ;
      RECT 439.64 9.55 439.81 10.56 ;
      RECT 439.98 9.05 440.15 13.24 ;
      RECT 440.35 9.05 440.52 13.24 ;
      RECT 441.06 9.55 441.23 10.56 ;
      RECT 440.72 9.38 440.89 12.91 ;
      RECT 440.72 9.05 441.57 9.38 ;
      RECT 440.72 12.91 441.57 13.24 ;
      RECT 441.4 9.38 441.57 12.91 ;
      RECT 368.815 5.135 369.515 12.265 ;
      RECT 368.815 4.425 373.19 5.135 ;
      RECT 368.815 12.265 373.19 12.965 ;
      RECT 372.49 5.135 373.19 12.265 ;
      RECT 371.475 6 372.015 11.395 ;
      RECT 370 6 370.54 11.395 ;
      RECT 375.665 3.905 378.175 4.075 ;
      RECT 375.665 4.075 375.835 15.315 ;
      RECT 375.665 15.315 378.175 15.485 ;
      RECT 378.005 4.075 378.175 15.315 ;
      RECT 376.47 4.315 377.37 4.485 ;
      RECT 376.585 4.485 377.255 14.905 ;
      RECT 376.06 14.905 377.37 15.075 ;
      RECT 388.74 6.62 388.91 7.63 ;
      RECT 388.74 4.95 388.91 5.96 ;
      RECT 386.27 9.66 386.6 10.31 ;
      RECT 386.9 9.66 387.23 10.31 ;
      RECT 389.42 9.66 389.75 10.31 ;
      RECT 390.05 9.66 390.38 10.31 ;
      RECT 388.79 9.66 389.12 10.31 ;
      RECT 388.16 9.66 388.49 10.31 ;
      RECT 387.53 9.66 387.86 10.31 ;
      RECT 388.15 4.65 388.33 8.125 ;
      RECT 392.84 4.65 393.02 5.79 ;
      RECT 401.145 8.305 401.325 12.285 ;
      RECT 402.46 5.97 402.64 8.01 ;
      RECT 392.84 5.79 402.64 5.97 ;
      RECT 401.145 8.01 425.58 8.125 ;
      RECT 402.46 8.18 402.63 12.17 ;
      RECT 425.405 8.18 425.575 12.56 ;
      RECT 388.15 4.47 393.02 4.65 ;
      RECT 388.15 8.18 401.325 8.305 ;
      RECT 388.15 8.125 425.58 8.18 ;
      RECT 390.5 6.62 390.67 7.63 ;
      RECT 389.62 6.62 389.79 7.63 ;
      RECT 390.5 4.95 390.67 5.96 ;
      RECT 389.62 4.95 389.79 5.96 ;
      RECT 395.77 3.17 395.94 4.195 ;
      RECT 395.18 4.845 401.93 5.025 ;
      RECT 395.18 2.64 401.93 2.82 ;
      RECT 401.75 2.82 401.93 4.845 ;
      RECT 395.18 2.82 395.36 4.845 ;
      RECT 391.38 6.62 391.55 7.63 ;
      RECT 391.38 4.95 391.55 5.96 ;
      RECT 396.18 6.62 396.35 7.63 ;
      RECT 394.9 6.62 395.07 7.63 ;
      RECT 394.02 6.62 394.19 7.63 ;
      RECT 392.26 4.95 392.43 5.96 ;
      RECT 395.125 6.22 396.655 6.39 ;
      RECT 388.965 6.22 394.955 6.39 ;
      RECT 395.865 4.425 396.545 4.595 ;
      RECT 393.14 6.62 393.31 7.63 ;
      RECT 392.26 6.62 392.43 7.63 ;
      RECT 390.68 9.66 391.01 10.31 ;
      RECT 391.31 9.66 391.64 10.31 ;
      RECT 393.2 9.66 393.53 10.31 ;
      RECT 393.83 9.66 394.16 10.31 ;
      RECT 391.94 9.66 392.27 10.31 ;
      RECT 392.57 9.66 392.9 10.31 ;
      RECT 396.35 9.66 396.68 10.68 ;
      RECT 395.72 9.66 396.05 10.68 ;
      RECT 395.09 9.66 395.42 10.68 ;
      RECT 394.46 9.66 394.79 10.68 ;
      RECT 396.85 3.17 397.02 4.18 ;
      RECT 396.715 4.425 398.955 4.595 ;
      RECT 397.93 3.17 398.1 4.195 ;
      RECT 399.01 3.17 399.18 4.18 ;
      RECT 401.17 3.17 401.34 4.18 ;
      RECT 400.6 3.605 400.83 4.425 ;
      RECT 399.235 4.425 401.115 4.595 ;
      RECT 400.09 3.17 400.26 4.195 ;
      RECT 396.73 6.62 396.9 7.63 ;
      RECT 398.24 9.66 398.57 10.28 ;
      RECT 397.61 9.66 397.94 10.28 ;
      RECT 396.98 9.66 397.31 10.28 ;
      RECT 397.07 6.39 398.84 6.76 ;
      RECT 396.955 6.22 398.955 6.39 ;
      RECT 399.01 6.62 399.18 7.63 ;
      RECT 401.29 6.62 401.46 7.63 ;
      RECT 399.5 9.66 399.83 10.31 ;
      RECT 398.87 9.66 399.2 10.31 ;
      RECT 399.235 6.22 401.235 6.39 ;
      RECT 404.19 8.35 404.7 8.68 ;
      RECT 404.26 8.68 404.63 14.76 ;
      RECT 404.19 14.76 404.7 15.09 ;
      RECT 405.07 8.35 405.58 8.68 ;
      RECT 405.14 8.68 405.51 14.76 ;
      RECT 405.01 14.76 405.58 15.09 ;
      RECT 407.38 8.35 407.89 8.68 ;
      RECT 407.38 14.76 407.91 14.93 ;
      RECT 407.38 14.93 407.89 15.09 ;
      RECT 407.45 8.68 407.82 14.76 ;
      RECT 406.5 8.35 407.01 8.68 ;
      RECT 406.57 8.68 406.94 14.76 ;
      RECT 406.5 14.76 407.03 15.3 ;
      RECT 403.31 8.35 403.82 8.68 ;
      RECT 403.38 8.68 403.75 14.76 ;
      RECT 403.31 14.84 403.84 15.01 ;
      RECT 403.31 15.01 403.82 15.09 ;
      RECT 403.31 14.76 403.82 14.84 ;
      RECT 407.99 8.845 408.16 14.59 ;
      RECT 407.11 9.15 407.28 11.86 ;
      RECT 405.8 14.76 406.33 14.93 ;
      RECT 406.23 8.845 406.4 14.445 ;
      RECT 406.02 14.615 406.33 14.76 ;
      RECT 406.02 14.445 406.4 14.615 ;
      RECT 403.04 8.83 403.21 14.59 ;
      RECT 405.68 9.15 405.85 11.86 ;
      RECT 403.92 9.15 404.09 11.86 ;
      RECT 404.8 8.83 404.97 14.465 ;
      RECT 413.61 8.68 413.98 14.76 ;
      RECT 414.49 8.68 414.86 14.76 ;
      RECT 413.54 8.65 414.05 8.68 ;
      RECT 413.54 14.76 414.05 14.79 ;
      RECT 413.54 8.35 414.93 8.65 ;
      RECT 414.42 8.65 414.93 8.68 ;
      RECT 413.54 14.79 414.93 15.09 ;
      RECT 414.42 14.76 414.93 14.79 ;
      RECT 412.73 8.68 413.1 14.76 ;
      RECT 411.85 8.68 412.22 14.76 ;
      RECT 412.66 8.65 413.17 8.68 ;
      RECT 411.78 8.35 413.17 8.65 ;
      RECT 411.78 8.65 412.29 8.68 ;
      RECT 412.66 14.76 413.17 14.79 ;
      RECT 411.78 14.79 413.17 15.09 ;
      RECT 411.78 14.76 412.29 14.79 ;
      RECT 410.9 8.35 411.41 8.68 ;
      RECT 342.49 5.415 342.67 10.48 ;
      RECT 341.725 11.865 342.67 12.535 ;
      RECT 319.325 21.685 319.505 28.375 ;
      RECT 319.325 20.305 319.505 21.175 ;
      RECT 342.49 10.99 342.67 11.865 ;
      RECT 342.49 12.535 342.67 19.635 ;
      RECT 319.325 21.175 342.67 21.685 ;
      RECT 342.49 20.305 342.67 21.175 ;
      RECT 342.49 4.19 342.67 5.235 ;
      RECT 342.49 21.685 342.67 28.375 ;
      RECT 358.525 5.415 358.705 15.485 ;
      RECT 341.725 19.635 342.67 20.305 ;
      RECT 319.325 10.48 342.67 10.99 ;
      RECT 320.085 8.48 320.815 8.65 ;
      RECT 320.085 8.65 320.735 8.73 ;
      RECT 320.085 8.4 320.735 8.48 ;
      RECT 320.225 7.77 320.875 8.1 ;
      RECT 320.825 9.66 321.475 9.99 ;
      RECT 320.225 9.03 320.875 9.36 ;
      RECT 320.025 6.51 320.675 6.84 ;
      RECT 320.025 5.25 320.675 5.58 ;
      RECT 320.025 4.62 320.705 4.95 ;
      RECT 320.025 5.88 320.675 6.21 ;
      RECT 324.625 7.77 325.275 8.1 ;
      RECT 323.595 8.4 324.245 8.73 ;
      RECT 323.595 9.03 324.245 9.36 ;
      RECT 324.625 8.4 325.275 8.73 ;
      RECT 323.595 7.77 324.245 8.1 ;
      RECT 324.625 9.03 325.275 9.36 ;
      RECT 329.055 7.85 329.785 8.02 ;
      RECT 329.135 8.02 329.785 8.1 ;
      RECT 329.135 7.77 329.785 7.85 ;
      RECT 329.025 8.48 329.615 8.65 ;
      RECT 329.025 8.65 329.535 8.73 ;
      RECT 329.025 8.4 329.535 8.48 ;
      RECT 332.395 8.4 333.045 8.73 ;
      RECT 327.995 9.03 328.645 9.36 ;
      RECT 328.135 8.65 328.305 8.73 ;
      RECT 328.135 8.4 328.305 8.48 ;
      RECT 328.475 8.65 328.645 8.73 ;
      RECT 328.055 8.48 328.645 8.65 ;
      RECT 328.475 8.4 328.645 8.48 ;
      RECT 328.425 6.51 329.075 6.84 ;
      RECT 330.425 7.14 331.075 7.47 ;
      RECT 327.395 6.51 328.045 6.84 ;
      RECT 332.425 9.03 333.075 9.36 ;
      RECT 336.69 2.755 337.22 2.925 ;
      RECT 336.69 2.235 337.2 2.755 ;
      RECT 333.825 8.4 334.475 8.73 ;
      RECT 332.825 7.77 333.475 8.1 ;
      RECT 343.27 6.34 343.44 16.19 ;
      RECT 343.405 3.925 343.95 4.595 ;
      RECT 343.615 5.815 344.285 5.985 ;
      RECT 341.195 9.66 341.845 9.99 ;
      RECT 341.195 9.03 341.845 9.36 ;
      RECT 341.195 6.51 341.845 6.84 ;
      RECT 341.195 7.14 341.845 7.47 ;
      RECT 341.195 8.4 341.845 8.73 ;
      RECT 341.195 5.88 341.845 6.21 ;
      RECT 341.195 5.25 341.845 5.58 ;
      RECT 341.195 4.62 341.845 4.95 ;
      RECT 341.195 7.77 341.845 8.1 ;
      RECT 344.45 6.34 344.62 16.19 ;
      RECT 345.63 6.34 345.8 16.19 ;
      RECT 349.375 3.925 350.15 4.595 ;
      RECT 347.335 3.925 348.02 4.595 ;
      RECT 345.48 3.925 346.135 4.595 ;
      RECT 349.1 2.335 349.63 2.505 ;
      RECT 349.11 2.505 349.62 2.905 ;
      RECT 349.11 2.235 349.62 2.335 ;
      RECT 347.155 6.5 347.44 9.84 ;
      RECT 347.155 6.305 347.325 6.5 ;
      RECT 347.155 23.58 347.44 26.92 ;
      RECT 347.155 26.92 347.325 27.115 ;
      RECT 347.155 9.84 347.325 23.58 ;
      RECT 347.875 5.945 350.585 6.115 ;
      RECT 344.795 5.82 345.465 5.99 ;
      RECT 353.17 3.925 356.475 4.595 ;
      RECT 351.13 3.925 351.825 4.595 ;
      RECT 351.525 5.945 354.235 6.115 ;
      RECT 351.525 11.505 354.235 11.675 ;
      RECT 351.525 12.785 354.235 12.955 ;
      RECT 351.525 10.225 354.235 10.395 ;
      RECT 351.525 5.93 353.97 5.945 ;
      RECT 351.525 11.675 353.97 12.785 ;
      RECT 351.525 10.395 353.97 11.505 ;
      RECT 351.525 6.115 353.97 10.225 ;
      RECT 350.385 15.735 350.975 15.905 ;
      RECT 350.805 15.125 350.975 15.735 ;
      RECT 350.385 14.955 350.975 15.125 ;
      RECT 350.385 17.515 350.975 17.685 ;
      RECT 350.805 15.905 350.975 17.515 ;
      RECT 350.385 18.295 350.975 18.465 ;
      RECT 350.805 17.685 350.975 18.295 ;
      RECT 350.805 6.305 350.975 14.955 ;
      RECT 350.805 18.465 350.975 27.115 ;
      RECT 354.455 6.305 354.625 10.035 ;
      RECT 355.175 5.945 357.885 6.115 ;
      RECT 358.025 2.235 358.535 2.905 ;
      RECT 358.005 3.925 358.515 4.595 ;
      RECT 357.98 6.5 358.275 9.84 ;
      RECT 358.105 9.915 358.275 10.035 ;
      RECT 358.005 9.84 358.275 9.915 ;
      RECT 358.005 6.305 358.275 6.5 ;
      RECT 363.74 5.42 365.065 5.83 ;
      RECT 367.355 3.665 368.055 13.725 ;
      RECT 360.76 3.665 361.46 13.725 ;
      RECT 378.935 3.135 379.105 16.245 ;
      RECT 367.355 16.745 368.055 26.805 ;
      RECT 373.95 16.745 374.65 26.805 ;
      RECT 360.76 16.745 361.46 26.805 ;
      RECT 360.76 26.805 374.65 27.505 ;
      RECT 373.95 3.665 374.905 13.725 ;
      RECT 360.76 2.965 379.105 3.135 ;
      RECT 360.76 16.045 374.905 16.245 ;
      RECT 360.76 16.415 374.65 16.745 ;
      RECT 360.76 16.245 379.105 16.415 ;
      RECT 360.76 3.135 374.905 3.665 ;
      RECT 374.735 14.425 374.905 16.045 ;
      RECT 360.76 13.725 374.905 14.425 ;
      RECT 365.895 5.135 366.595 12.265 ;
      RECT 362.22 4.425 366.595 5.135 ;
      RECT 362.22 12.265 366.595 12.965 ;
      RECT 362.22 5.135 362.92 12.265 ;
      RECT 363.395 6 363.935 11.395 ;
      RECT 364.87 6 365.41 11.395 ;
      RECT 370.345 5.42 371.67 5.83 ;
      RECT 288.755 6.915 290.825 7.085 ;
      RECT 290.655 7.085 290.825 7.38 ;
      RECT 290.655 6.28 290.825 6.915 ;
      RECT 287.525 6.055 288.535 6.225 ;
      RECT 287.525 4.675 288.535 4.845 ;
      RECT 287.525 5.135 288.535 5.305 ;
      RECT 287.525 5.595 288.535 5.765 ;
      RECT 291.075 6.055 292.085 6.225 ;
      RECT 291.075 5.595 292.085 5.765 ;
      RECT 291.075 5.135 292.085 5.305 ;
      RECT 291.075 4.675 292.085 4.845 ;
      RECT 287.525 7.345 288.535 7.605 ;
      RECT 288.755 8.08 288.925 8.66 ;
      RECT 288.755 7.91 290.825 8.08 ;
      RECT 290.655 8.08 290.825 8.99 ;
      RECT 287.525 8.485 288.535 8.685 ;
      RECT 287.525 7.985 288.535 8.155 ;
      RECT 289.165 8.815 289.71 8.985 ;
      RECT 289.165 8.985 289.335 8.995 ;
      RECT 289.165 8.25 289.335 8.815 ;
      RECT 289.165 7.255 289.335 7.74 ;
      RECT 287.525 6.975 288.535 7.145 ;
      RECT 287.525 6.515 288.535 6.685 ;
      RECT 291.075 7.985 292.085 8.18 ;
      RECT 290.26 8.995 290.43 9.055 ;
      RECT 290.245 8.25 290.415 8.885 ;
      RECT 290.245 8.885 290.43 8.995 ;
      RECT 290.245 7.255 290.415 7.74 ;
      RECT 291.075 8.485 292.085 8.685 ;
      RECT 291.075 7.435 292.085 7.605 ;
      RECT 291.125 7.345 292.085 7.435 ;
      RECT 291.075 6.975 292.085 7.145 ;
      RECT 291.075 6.515 292.085 6.685 ;
      RECT 287.525 9.595 288.535 9.765 ;
      RECT 287.97 9.765 288.5 9.77 ;
      RECT 288.755 9.82 288.925 10.57 ;
      RECT 288.755 9.225 290.905 9.45 ;
      RECT 288.755 9.45 288.925 9.54 ;
      RECT 288.755 8.87 288.925 9.225 ;
      RECT 287.55 10.83 289.335 10.875 ;
      RECT 287.545 10.875 289.335 12.745 ;
      RECT 289.165 9.7 289.335 10.83 ;
      RECT 287.525 9.065 288.535 9.235 ;
      RECT 290.29 10.245 290.825 10.415 ;
      RECT 290.655 9.745 290.825 10.245 ;
      RECT 291.075 9.575 292.085 9.745 ;
      RECT 291.075 9.045 292.085 9.215 ;
      RECT 296.4 4.815 296.58 12.515 ;
      RECT 296.4 4.635 299.22 4.815 ;
      RECT 296.4 12.515 299.22 12.695 ;
      RECT 299.04 7.175 299.63 7.345 ;
      RECT 299.04 7.345 299.22 12.515 ;
      RECT 299.04 4.815 299.22 7.175 ;
      RECT 296.9 5.45 297.07 8.69 ;
      RECT 296.9 9.52 297.07 11.985 ;
      RECT 297.3 5.225 298.31 5.395 ;
      RECT 297.3 8.745 298.31 8.915 ;
      RECT 297.3 9.295 298.31 9.465 ;
      RECT 297.3 6.105 298.31 6.275 ;
      RECT 297.3 6.985 298.31 7.155 ;
      RECT 297.3 7.865 298.31 8.035 ;
      RECT 299.985 4.815 300.165 18.835 ;
      RECT 299.985 4.635 302.73 4.815 ;
      RECT 299.985 34.06 302.73 34.24 ;
      RECT 299.985 19.705 300.165 34.06 ;
      RECT 302.55 4.815 302.73 34.06 ;
      RECT 300.845 7.585 301.92 7.755 ;
      RECT 300.415 5.45 300.585 9.89 ;
      RECT 300.845 5.225 301.855 5.395 ;
      RECT 300.845 9.945 301.855 10.115 ;
      RECT 300.845 6.405 301.855 6.575 ;
      RECT 300.845 8.765 301.855 8.935 ;
      RECT 307.575 5.43 307.745 15.68 ;
      RECT 303.495 28.605 310.725 28.785 ;
      RECT 303.495 4.635 310.725 4.815 ;
      RECT 303.495 4.815 303.675 28.605 ;
      RECT 309.725 7.825 310.725 8.295 ;
      RECT 308.155 15.145 310.725 15.315 ;
      RECT 310.545 8.295 310.725 14.985 ;
      RECT 309.725 14.985 310.725 15.145 ;
      RECT 309.725 25.125 310.725 25.595 ;
      RECT 308.155 7.655 310.725 7.825 ;
      RECT 310.545 25.765 310.725 28.605 ;
      RECT 308.155 25.595 310.725 25.765 ;
      RECT 309.725 18.105 310.725 18.435 ;
      RECT 310.545 18.435 310.725 25.125 ;
      RECT 310.545 15.315 310.725 18.105 ;
      RECT 310.545 4.815 310.725 7.655 ;
      RECT 308.155 15.315 309.505 15.625 ;
      RECT 303.915 5.37 304.095 28.05 ;
      RECT 308.155 8.435 309.505 8.605 ;
      RECT 308.155 9.995 309.505 10.165 ;
      RECT 308.155 5.375 309.505 5.545 ;
      RECT 304.315 5.225 307.025 5.395 ;
      RECT 308.155 9.215 309.505 9.385 ;
      RECT 304.315 9.785 307.025 9.955 ;
      RECT 304.315 7.505 307.025 7.675 ;
      RECT 315.015 29.87 316.155 30.38 ;
      RECT 313.635 12.67 313.805 20.495 ;
      RECT 311.495 12.67 312.345 20.495 ;
      RECT 311.495 28.535 316.655 28.705 ;
      RECT 311.495 28.705 316.155 29.87 ;
      RECT 316.485 4.885 316.655 28.535 ;
      RECT 311.495 4.67 316.655 4.885 ;
      RECT 311.495 4.885 313.805 12.67 ;
      RECT 311.495 20.495 313.805 28.535 ;
      RECT 314.625 7.725 315.635 7.895 ;
      RECT 314.625 5.385 315.635 5.555 ;
      RECT 314.625 9.285 315.635 9.455 ;
      RECT 314.625 8.505 315.635 8.675 ;
      RECT 314.625 6.165 315.635 6.335 ;
      RECT 314.625 6.945 315.635 7.115 ;
      RECT 315.855 5.61 316.025 10.01 ;
      RECT 319.325 4.01 342.67 4.19 ;
      RECT 319.325 28.375 358.705 28.555 ;
      RECT 346.635 5.415 346.805 28.375 ;
      RECT 319.325 11.865 320.055 12.535 ;
      RECT 319.325 19.635 320.055 20.305 ;
      RECT 319.36 28.555 342.39 28.565 ;
      RECT 358.505 15.485 358.705 16.91 ;
      RECT 358.525 16.91 358.705 28.375 ;
      RECT 320.4 21.685 342.2 21.695 ;
      RECT 320.4 21.165 342.2 21.175 ;
      RECT 342.49 5.235 358.705 5.415 ;
      RECT 319.325 12.535 319.505 19.635 ;
      RECT 319.325 10.99 319.505 11.865 ;
      RECT 319.325 4.19 319.505 10.48 ;
      RECT 274 3.275 274.53 3.295 ;
      RECT 274.05 3.445 279.14 3.465 ;
      RECT 274 3.295 279.14 3.445 ;
      RECT 274 4.74 279.14 4.91 ;
      RECT 254.955 2.68 279.03 2.85 ;
      RECT 269.325 7.38 269.855 7.55 ;
      RECT 269.505 7.55 269.675 8.16 ;
      RECT 269.505 5.02 269.675 7.38 ;
      RECT 270.785 5.02 270.955 6.28 ;
      RECT 271.245 6.81 273.255 6.98 ;
      RECT 273.085 6.98 273.255 8.16 ;
      RECT 271.245 6.98 271.415 8.16 ;
      RECT 272.165 6.98 272.335 8.16 ;
      RECT 273.625 4.44 273.795 4.505 ;
      RECT 273.66 4.97 273.83 5.175 ;
      RECT 273.625 4.505 273.83 4.97 ;
      RECT 273.945 7.18 274.615 7.26 ;
      RECT 276.855 7.43 277.385 7.55 ;
      RECT 275.92 7.07 277.375 7.26 ;
      RECT 273.945 7.26 277.375 7.38 ;
      RECT 275.92 5.66 276.09 7.07 ;
      RECT 273.945 7.38 277.385 7.43 ;
      RECT 278.805 5.39 278.975 6.7 ;
      RECT 277.195 5.39 277.365 6.7 ;
      RECT 274.64 5.39 274.81 6.67 ;
      RECT 274.05 5.2 278.975 5.39 ;
      RECT 273.72 5.66 273.89 6.67 ;
      RECT 274.05 4.28 278.8 4.45 ;
      RECT 274.115 4.45 278.605 4.455 ;
      RECT 273.605 6.84 274.35 7.01 ;
      RECT 274.175 6.67 274.35 6.84 ;
      RECT 274.18 5.66 274.35 6.67 ;
      RECT 273.605 7.01 273.775 8.76 ;
      RECT 274.29 9.01 275.005 9.18 ;
      RECT 274.475 9.18 275.005 9.475 ;
      RECT 274.065 7.75 274.235 8.76 ;
      RECT 279.31 2.995 279.48 4.16 ;
      RECT 279.68 3.295 280.69 3.465 ;
      RECT 279.68 4.215 280.69 4.385 ;
      RECT 279.68 3.755 280.69 3.925 ;
      RECT 276.665 11.32 277.195 11.49 ;
      RECT 276.845 11.49 277.015 12.47 ;
      RECT 276.845 7.72 277.015 11.32 ;
      RECT 275.965 7.72 276.135 12.47 ;
      RECT 275.015 6.92 275.685 7.09 ;
      RECT 275.255 7.72 275.785 9.07 ;
      RECT 276.495 6.51 277.025 6.68 ;
      RECT 276.715 5.68 276.885 6.51 ;
      RECT 283.775 7.72 284.005 8.95 ;
      RECT 283.775 11.7 284.005 12.71 ;
      RECT 283.805 7.37 283.975 7.72 ;
      RECT 283.805 12.71 283.975 12.74 ;
      RECT 283.805 8.95 283.975 11.7 ;
      RECT 280.035 7.37 280.205 12.65 ;
      RECT 280.035 7.2 283.975 7.37 ;
      RECT 281.795 7.37 281.965 12.65 ;
      RECT 278.975 11.32 279.505 11.49 ;
      RECT 279.155 11.49 279.325 12.47 ;
      RECT 279.155 7.72 279.325 11.32 ;
      RECT 279.31 4.5 279.48 5.17 ;
      RECT 278.615 7.04 279.285 7.21 ;
      RECT 278.615 7.01 279.145 7.04 ;
      RECT 278.095 7.38 278.625 7.55 ;
      RECT 278.275 7.55 278.445 12.47 ;
      RECT 278.275 5.69 278.445 7.38 ;
      RECT 277.545 7.01 278.075 7.18 ;
      RECT 277.545 8.9 278.075 9.07 ;
      RECT 277.725 9.07 277.895 12.47 ;
      RECT 277.725 7.18 277.895 8.9 ;
      RECT 277.725 5.69 277.895 7.01 ;
      RECT 279.26 6.51 279.79 6.68 ;
      RECT 279.285 5.68 279.455 6.51 ;
      RECT 281.09 3.515 281.26 5.885 ;
      RECT 265.33 26.92 284.775 27.09 ;
      RECT 289.165 2.885 289.335 6.745 ;
      RECT 259.285 19.52 259.455 20.525 ;
      RECT 287.005 36.235 289.335 36.405 ;
      RECT 289.165 13.335 289.335 36.235 ;
      RECT 287.545 13.165 289.335 13.335 ;
      RECT 281.47 2.715 289.335 2.885 ;
      RECT 265.33 25.74 265.515 26.92 ;
      RECT 287.005 24.905 287.175 36.235 ;
      RECT 264.76 25.74 265.14 25.815 ;
      RECT 259.285 25.74 263.93 25.815 ;
      RECT 259.25 25.13 259.455 25.57 ;
      RECT 259.285 24.09 259.455 25.13 ;
      RECT 284.59 24.905 285.17 25.75 ;
      RECT 284.59 25.75 284.775 26.92 ;
      RECT 265.345 23.56 265.515 25.57 ;
      RECT 284.59 24.735 287.175 24.905 ;
      RECT 259.25 25.57 265.515 25.74 ;
      RECT 284.59 19.52 285.17 24.735 ;
      RECT 259.285 19.35 285.17 19.52 ;
      RECT 284.76 2.885 285.17 19.35 ;
      RECT 285.52 3.395 286.99 3.655 ;
      RECT 282.345 9.73 282.99 9.9 ;
      RECT 282.345 7.72 282.515 9.73 ;
      RECT 282.345 9.9 282.515 18.92 ;
      RECT 282.865 11.32 283.395 11.49 ;
      RECT 283.225 11.49 283.395 12.47 ;
      RECT 283.225 7.72 283.395 11.32 ;
      RECT 281.45 5.935 284.16 6.105 ;
      RECT 284.33 3.465 284.5 5.055 ;
      RECT 281.45 3.295 284.5 3.465 ;
      RECT 281.45 5.055 284.5 5.225 ;
      RECT 281.45 4.175 284.16 4.345 ;
      RECT 280.915 11.32 281.445 11.49 ;
      RECT 280.915 11.49 281.085 12.47 ;
      RECT 280.915 7.72 281.085 11.32 ;
      RECT 290.245 2.985 290.415 6.745 ;
      RECT 290.245 2.815 292.765 2.985 ;
      RECT 289.81 10.05 290.12 10.585 ;
      RECT 292.335 8.025 292.765 10.585 ;
      RECT 289.81 9.64 290.415 10.05 ;
      RECT 292.335 7.485 292.505 8.025 ;
      RECT 292.335 2.985 292.765 7.485 ;
      RECT 289.81 10.585 292.765 10.895 ;
      RECT 288.755 3.52 288.925 6 ;
      RECT 290.655 3.52 290.825 6 ;
      RECT 287.525 3.295 288.535 3.465 ;
      RECT 287.525 3.755 288.535 3.925 ;
      RECT 287.525 4.215 288.535 4.385 ;
      RECT 291.075 3.295 292.085 3.465 ;
      RECT 291.075 4.215 292.085 4.385 ;
      RECT 291.075 3.755 292.085 3.925 ;
      RECT 288.755 7.085 288.925 7.38 ;
      RECT 288.755 6.28 288.925 6.915 ;
      RECT 236.465 10.015 237.215 10.185 ;
      RECT 237.045 11.36 237.575 11.53 ;
      RECT 237.045 11.53 237.215 13.505 ;
      RECT 236.465 9.22 237 9.39 ;
      RECT 236.465 5.035 236.635 9.22 ;
      RECT 237.045 10.185 237.215 11.36 ;
      RECT 236.465 9.39 236.635 10.015 ;
      RECT 239.695 9.96 240.225 10.13 ;
      RECT 239.705 10.13 240.225 10.965 ;
      RECT 237.665 9.22 238.195 9.39 ;
      RECT 238.025 9.39 238.195 9.785 ;
      RECT 238.025 5.035 238.195 9.22 ;
      RECT 237.245 8.85 237.775 9.02 ;
      RECT 237.245 9.02 237.415 9.785 ;
      RECT 237.245 5.035 237.415 8.85 ;
      RECT 235.105 4.685 235.275 10.055 ;
      RECT 235.105 4.515 243.425 4.685 ;
      RECT 240.135 4.685 240.305 9.785 ;
      RECT 241.695 4.685 241.865 9.785 ;
      RECT 243.255 4.685 243.425 9.785 ;
      RECT 242.815 8.83 243.085 10.295 ;
      RECT 240.415 10.295 243.125 10.465 ;
      RECT 242.115 8.85 242.645 9.02 ;
      RECT 242.475 9.02 242.645 9.785 ;
      RECT 242.475 5.035 242.645 8.85 ;
      RECT 240.915 8.85 241.445 9.02 ;
      RECT 240.915 9.02 241.085 9.785 ;
      RECT 240.915 5.035 241.085 8.85 ;
      RECT 273.595 11.37 273.765 12.73 ;
      RECT 270.915 10.93 275.555 11.37 ;
      RECT 243.97 10.76 252.915 10.93 ;
      RECT 256.03 10.76 261.145 10.93 ;
      RECT 264.26 10.76 275.555 10.93 ;
      RECT 275.385 9.38 275.555 9.645 ;
      RECT 269.205 9.645 275.555 10.76 ;
      RECT 269.205 9.27 273.795 9.645 ;
      RECT 252.745 9.01 252.915 10.76 ;
      RECT 256.03 9.01 256.2 10.76 ;
      RECT 260.975 9.01 261.145 10.76 ;
      RECT 264.26 9.01 264.43 10.76 ;
      RECT 243.97 8.84 247.97 10.76 ;
      RECT 252.745 8.84 256.2 9.01 ;
      RECT 260.975 8.84 264.43 9.01 ;
      RECT 269.205 8.84 273.255 9.27 ;
      RECT 243.97 4.515 245.365 8.84 ;
      RECT 246.095 7.15 246.265 8.84 ;
      RECT 254.325 7.15 254.495 8.84 ;
      RECT 262.555 7.15 262.725 8.84 ;
      RECT 270.785 7.15 270.955 8.84 ;
      RECT 271.705 7.15 271.875 8.84 ;
      RECT 272.625 7.15 272.795 8.84 ;
      RECT 250.845 6.51 252.875 6.68 ;
      RECT 247.715 6.51 249.405 6.68 ;
      RECT 250.305 6.88 250.835 7.05 ;
      RECT 250.485 5.02 250.655 6.88 ;
      RECT 250.485 7.05 250.655 9.79 ;
      RECT 249.755 6.51 250.285 6.68 ;
      RECT 249.935 6.68 250.105 9.79 ;
      RECT 249.935 5.02 250.105 6.51 ;
      RECT 248.655 7.08 248.825 9.79 ;
      RECT 247.375 4.97 247.905 5.14 ;
      RECT 247.375 5.14 247.545 8.16 ;
      RECT 246.095 5.02 246.265 6.28 ;
      RECT 248.655 5.02 248.825 6.28 ;
      RECT 271.265 4.77 271.435 6.04 ;
      RECT 246.015 4.6 271.435 4.77 ;
      RECT 250.91 9.99 251.44 10.59 ;
      RECT 259.855 3.37 260.025 4.12 ;
      RECT 254.935 4.12 260.025 4.29 ;
      RECT 254.935 3.2 260.025 3.37 ;
      RECT 254.935 3.66 259.685 3.83 ;
      RECT 251.765 5.02 251.935 6.28 ;
      RECT 254.325 5.02 254.495 6.28 ;
      RECT 255.425 4.99 255.955 5.16 ;
      RECT 255.605 5.16 255.775 8.16 ;
      RECT 253.045 5.02 253.215 8.16 ;
      RECT 253.385 4.97 253.915 6.68 ;
      RECT 255.945 6.51 257.635 6.68 ;
      RECT 256.885 5.02 257.055 6.28 ;
      RECT 251.765 7.08 251.935 9.79 ;
      RECT 256.885 7.08 257.055 9.79 ;
      RECT 257.38 9.215 257.91 10.59 ;
      RECT 260.535 3.37 260.705 4.12 ;
      RECT 260.535 3.2 265.625 3.37 ;
      RECT 260.535 4.12 265.625 4.29 ;
      RECT 260.875 3.66 266.075 3.83 ;
      RECT 265.905 3.83 266.075 4.12 ;
      RECT 265.905 3.37 266.075 3.66 ;
      RECT 265.905 4.12 271.095 4.29 ;
      RECT 265.905 3.2 271.095 3.37 ;
      RECT 259.075 6.51 261.105 6.68 ;
      RECT 257.985 6.51 258.515 6.68 ;
      RECT 258.165 6.68 258.335 9.79 ;
      RECT 258.165 5.02 258.335 6.51 ;
      RECT 259.995 5.02 260.165 6.28 ;
      RECT 258.535 6.88 259.065 7.05 ;
      RECT 258.715 5.02 258.885 6.88 ;
      RECT 258.715 7.05 258.885 9.79 ;
      RECT 260.195 3.43 260.365 4.43 ;
      RECT 262.555 5.02 262.725 6.28 ;
      RECT 261.275 5.02 261.445 8.16 ;
      RECT 259.995 7.08 260.165 9.79 ;
      RECT 267.305 6.51 269.335 6.68 ;
      RECT 264.175 6.51 265.865 6.68 ;
      RECT 266.765 6.88 267.295 7.05 ;
      RECT 266.945 5.02 267.115 6.88 ;
      RECT 266.945 7.05 267.115 9.79 ;
      RECT 268.225 7.08 268.395 9.79 ;
      RECT 266.215 6.51 266.745 6.68 ;
      RECT 266.395 6.68 266.565 9.79 ;
      RECT 266.395 5.02 266.565 6.51 ;
      RECT 265.115 7.08 265.285 9.79 ;
      RECT 263.655 7.365 264.185 7.535 ;
      RECT 263.835 7.535 264.005 8.16 ;
      RECT 263.835 5.02 264.005 7.365 ;
      RECT 265.115 5.02 265.285 6.28 ;
      RECT 268.225 5.02 268.395 6.28 ;
      RECT 266.245 3.66 271.095 3.83 ;
      RECT 272.645 3.04 273.315 3.21 ;
      RECT 272.76 3.21 273.03 5.115 ;
      RECT 271.315 3.41 272.59 4.08 ;
      RECT 271.05 6.47 272.59 6.64 ;
      RECT 272.01 4.08 272.59 6.47 ;
      RECT 273.2 3.76 273.37 6.47 ;
      RECT 274.05 3.755 278.8 3.925 ;
      RECT 274.31 3.675 278.8 3.755 ;
      RECT 278.97 3.465 279.14 4.74 ;
      RECT 129.3 3.37 129.47 4.12 ;
      RECT 124.38 3.2 129.47 3.37 ;
      RECT 124.38 4.12 129.47 4.29 ;
      RECT 124.72 5.02 124.89 6.28 ;
      RECT 125.82 7.365 126.35 7.535 ;
      RECT 126 7.535 126.17 8.16 ;
      RECT 126 5.02 126.17 7.365 ;
      RECT 128.9 6.51 130.93 6.68 ;
      RECT 127.28 5.02 127.45 6.28 ;
      RECT 129.84 5.02 130.01 6.28 ;
      RECT 129.64 3.43 129.81 4.43 ;
      RECT 128.56 5.02 128.73 8.16 ;
      RECT 129.98 3.37 130.15 4.12 ;
      RECT 129.98 4.12 135.07 4.29 ;
      RECT 129.98 3.2 135.07 3.37 ;
      RECT 124.72 7.08 124.89 9.79 ;
      RECT 129.84 7.08 130.01 9.79 ;
      RECT 132.37 6.51 134.06 6.68 ;
      RECT 130.94 6.88 131.47 7.05 ;
      RECT 131.12 5.02 131.29 6.88 ;
      RECT 131.12 7.05 131.29 9.79 ;
      RECT 131.49 6.51 132.02 6.68 ;
      RECT 131.67 6.68 131.84 9.79 ;
      RECT 131.67 5.02 131.84 6.51 ;
      RECT 132.95 7.08 133.12 9.79 ;
      RECT 134.05 4.99 134.58 5.16 ;
      RECT 134.23 5.16 134.4 8.16 ;
      RECT 135.51 5.02 135.68 6.28 ;
      RECT 132.95 5.02 133.12 6.28 ;
      RECT 132.095 9.215 132.625 10.59 ;
      RECT 130.32 3.66 135.07 3.83 ;
      RECT 137.13 6.51 139.16 6.68 ;
      RECT 140.6 6.51 142.29 6.68 ;
      RECT 139.17 6.88 139.7 7.05 ;
      RECT 139.35 5.02 139.52 6.88 ;
      RECT 139.35 7.05 139.52 9.79 ;
      RECT 138.07 7.08 138.24 9.79 ;
      RECT 139.72 6.51 140.25 6.68 ;
      RECT 139.9 6.68 140.07 9.79 ;
      RECT 139.9 5.02 140.07 6.51 ;
      RECT 141.18 7.08 141.35 9.79 ;
      RECT 136.79 5.02 136.96 8.16 ;
      RECT 141.18 5.02 141.35 6.28 ;
      RECT 138.07 5.02 138.24 6.28 ;
      RECT 136.09 4.97 136.62 6.68 ;
      RECT 138.565 9.99 139.095 10.59 ;
      RECT 146.58 4.515 154.9 4.685 ;
      RECT 154.73 4.685 154.9 10.055 ;
      RECT 146.58 4.685 146.75 9.785 ;
      RECT 149.7 4.685 149.87 9.785 ;
      RECT 148.14 4.685 148.31 9.785 ;
      RECT 142.1 4.97 142.63 5.14 ;
      RECT 142.46 5.14 142.63 8.16 ;
      RECT 143.74 5.02 143.91 6.28 ;
      RECT 146.92 8.83 147.19 10.295 ;
      RECT 146.88 10.295 149.59 10.465 ;
      RECT 147.36 8.85 147.89 9.02 ;
      RECT 147.36 9.02 147.53 9.785 ;
      RECT 147.36 5.035 147.53 8.85 ;
      RECT 151.03 8.85 151.56 9.02 ;
      RECT 151.03 9.02 151.2 9.785 ;
      RECT 151.03 5.035 151.2 8.85 ;
      RECT 152.15 9.59 152.42 10.295 ;
      RECT 150.48 10.295 152.5 10.465 ;
      RECT 150.48 5.035 150.65 10.295 ;
      RECT 152.79 10.015 153.54 10.185 ;
      RECT 152.43 11.36 152.96 11.53 ;
      RECT 152.79 11.53 152.96 13.505 ;
      RECT 153.005 9.22 153.54 9.39 ;
      RECT 153.37 5.035 153.54 9.22 ;
      RECT 152.79 10.185 152.96 11.36 ;
      RECT 153.37 9.39 153.54 10.015 ;
      RECT 149.78 9.96 150.31 10.13 ;
      RECT 149.78 10.13 150.3 10.965 ;
      RECT 151.81 9.22 152.34 9.39 ;
      RECT 151.81 9.39 151.98 9.785 ;
      RECT 151.81 5.035 151.98 9.22 ;
      RECT 152.23 8.85 152.76 9.02 ;
      RECT 152.59 9.02 152.76 9.785 ;
      RECT 152.59 5.035 152.76 8.85 ;
      RECT 148.56 8.85 149.09 9.02 ;
      RECT 148.92 9.02 149.09 9.785 ;
      RECT 148.92 5.035 149.09 8.85 ;
      RECT 153.79 8.85 154.32 9.02 ;
      RECT 154.15 9.02 154.32 9.785 ;
      RECT 154.15 5.035 154.32 8.85 ;
      RECT 158.075 3.84 160.095 4.59 ;
      RECT 163.29 3.5 166 3.67 ;
      RECT 163.24 2.22 166 2.39 ;
      RECT 162.48 7.195 163.18 14.325 ;
      RECT 162.48 6.495 166.855 7.195 ;
      RECT 162.48 14.325 166.855 15.035 ;
      RECT 166.155 7.195 166.855 14.325 ;
      RECT 163.665 8.065 164.205 13.46 ;
      RECT 166.52 2.435 166.69 3.445 ;
      RECT 169.075 7.195 169.775 14.325 ;
      RECT 169.075 6.495 173.45 7.195 ;
      RECT 169.075 14.325 173.45 15.035 ;
      RECT 172.75 7.195 173.45 14.325 ;
      RECT 165.14 8.065 165.68 13.46 ;
      RECT 170.25 8.065 170.79 13.46 ;
      RECT 171.725 8.065 172.265 13.46 ;
      RECT 216.555 7.195 217.255 14.325 ;
      RECT 216.555 6.495 220.93 7.195 ;
      RECT 216.555 14.325 220.93 15.035 ;
      RECT 220.23 7.195 220.93 14.325 ;
      RECT 219.215 8.065 219.755 13.46 ;
      RECT 217.74 8.065 218.28 13.46 ;
      RECT 223.315 2.435 223.485 3.445 ;
      RECT 224.005 3.5 226.715 3.67 ;
      RECT 224.005 2.22 226.765 2.39 ;
      RECT 226.825 7.195 227.525 14.325 ;
      RECT 223.15 6.495 227.525 7.195 ;
      RECT 223.15 14.325 227.525 15.035 ;
      RECT 223.15 7.195 223.85 14.325 ;
      RECT 224.325 8.065 224.865 13.46 ;
      RECT 225.8 8.065 226.34 13.46 ;
      RECT 229.91 3.84 231.93 4.59 ;
      RECT 235.685 8.85 236.215 9.02 ;
      RECT 235.685 9.02 235.855 9.785 ;
      RECT 235.685 5.035 235.855 8.85 ;
      RECT 238.445 8.85 238.975 9.02 ;
      RECT 238.805 9.02 238.975 9.785 ;
      RECT 238.805 5.035 238.975 8.85 ;
      RECT 237.585 9.59 237.855 10.295 ;
      RECT 237.505 10.295 239.525 10.465 ;
      RECT 239.355 5.035 239.525 10.295 ;
      RECT 101.47 9.065 102.48 9.235 ;
      RECT 101.47 6.975 102.48 7.145 ;
      RECT 101.47 6.515 102.48 6.685 ;
      RECT 101.47 9.595 102.48 9.765 ;
      RECT 101.505 9.765 102.035 9.77 ;
      RECT 101.08 9.82 101.25 10.57 ;
      RECT 108.745 3.515 108.915 5.885 ;
      RECT 109.315 3.295 110.325 3.465 ;
      RECT 109.315 4.215 110.325 4.385 ;
      RECT 109.315 3.755 110.325 3.925 ;
      RECT 110.525 4.5 110.695 5.17 ;
      RECT 110.525 2.995 110.695 4.16 ;
      RECT 111.205 3.755 115.955 3.925 ;
      RECT 111.205 3.675 115.695 3.755 ;
      RECT 110.865 3.465 111.035 4.74 ;
      RECT 115.475 3.275 116.005 3.295 ;
      RECT 110.865 3.295 116.005 3.445 ;
      RECT 110.865 3.445 115.955 3.465 ;
      RECT 110.865 4.74 116.005 4.91 ;
      RECT 111.205 4.28 115.955 4.45 ;
      RECT 111.4 4.45 115.89 4.455 ;
      RECT 110.975 2.68 135.05 2.85 ;
      RECT 107.015 9.73 107.66 9.9 ;
      RECT 107.49 7.72 107.66 9.73 ;
      RECT 107.49 9.9 107.66 18.92 ;
      RECT 108.56 11.32 109.09 11.49 ;
      RECT 108.92 11.49 109.09 12.47 ;
      RECT 108.92 7.72 109.09 11.32 ;
      RECT 110.5 11.32 111.03 11.49 ;
      RECT 110.68 11.49 110.85 12.47 ;
      RECT 110.68 7.72 110.85 11.32 ;
      RECT 110.72 7.04 111.39 7.21 ;
      RECT 110.86 7.01 111.39 7.04 ;
      RECT 111.38 7.38 111.91 7.55 ;
      RECT 111.56 7.55 111.73 12.47 ;
      RECT 111.56 5.69 111.73 7.38 ;
      RECT 111.03 5.39 111.2 6.7 ;
      RECT 112.64 5.39 112.81 6.7 ;
      RECT 115.195 5.39 115.365 6.67 ;
      RECT 111.03 5.2 115.955 5.39 ;
      RECT 111.93 7.01 112.46 7.18 ;
      RECT 111.93 8.9 112.46 9.07 ;
      RECT 112.11 9.07 112.28 12.47 ;
      RECT 112.11 7.18 112.28 8.9 ;
      RECT 112.11 5.69 112.28 7.01 ;
      RECT 110.215 6.51 110.745 6.68 ;
      RECT 110.55 5.68 110.72 6.51 ;
      RECT 112.62 7.43 113.15 7.55 ;
      RECT 112.63 7.07 114.085 7.26 ;
      RECT 115.39 7.18 116.06 7.26 ;
      RECT 112.63 7.26 116.06 7.38 ;
      RECT 113.915 5.66 114.085 7.07 ;
      RECT 112.62 7.38 116.06 7.43 ;
      RECT 116.24 11.37 116.41 12.73 ;
      RECT 114.45 10.93 119.09 11.37 ;
      RECT 114.45 10.76 125.745 10.93 ;
      RECT 128.86 10.76 133.975 10.93 ;
      RECT 137.09 10.76 146.035 10.93 ;
      RECT 114.45 9.38 114.62 9.645 ;
      RECT 116.21 9.27 120.8 9.645 ;
      RECT 114.45 9.645 120.8 10.76 ;
      RECT 125.575 9.01 125.745 10.76 ;
      RECT 128.86 9.01 129.03 10.76 ;
      RECT 133.805 9.01 133.975 10.76 ;
      RECT 137.09 9.01 137.26 10.76 ;
      RECT 116.75 8.84 120.8 9.27 ;
      RECT 125.575 8.84 129.03 9.01 ;
      RECT 133.805 8.84 137.26 9.01 ;
      RECT 142.035 8.84 146.035 10.76 ;
      RECT 144.64 4.515 146.035 8.84 ;
      RECT 118.13 7.15 118.3 8.84 ;
      RECT 117.21 7.15 117.38 8.84 ;
      RECT 119.05 7.15 119.22 8.84 ;
      RECT 127.28 7.15 127.45 8.84 ;
      RECT 135.51 7.15 135.68 8.84 ;
      RECT 143.74 7.15 143.91 8.84 ;
      RECT 112.98 6.51 113.51 6.68 ;
      RECT 113.12 5.68 113.29 6.51 ;
      RECT 114.32 6.92 114.99 7.09 ;
      RECT 115.655 6.84 116.4 7.01 ;
      RECT 115.655 6.67 115.83 6.84 ;
      RECT 115.655 5.66 115.825 6.67 ;
      RECT 116.23 7.01 116.4 8.76 ;
      RECT 117.415 6.47 118.955 6.64 ;
      RECT 117.415 3.41 118.69 4.08 ;
      RECT 117.415 4.08 117.995 6.47 ;
      RECT 116.21 4.44 116.38 4.505 ;
      RECT 116.175 4.97 116.345 5.175 ;
      RECT 116.175 4.505 116.38 4.97 ;
      RECT 116.69 3.04 117.36 3.21 ;
      RECT 116.975 3.21 117.245 5.115 ;
      RECT 116.115 5.66 116.285 6.67 ;
      RECT 116.635 3.76 116.805 6.47 ;
      RECT 116.75 6.81 118.76 6.98 ;
      RECT 116.75 6.98 116.92 8.16 ;
      RECT 117.67 6.98 117.84 8.16 ;
      RECT 118.59 6.98 118.76 8.16 ;
      RECT 112.81 11.32 113.34 11.49 ;
      RECT 112.99 11.49 113.16 12.47 ;
      RECT 112.99 7.72 113.16 11.32 ;
      RECT 113.87 7.72 114.04 12.47 ;
      RECT 115 9.01 115.715 9.18 ;
      RECT 115 9.18 115.53 9.475 ;
      RECT 114.22 7.72 114.75 9.07 ;
      RECT 115.77 7.75 115.94 8.76 ;
      RECT 118.91 3.2 124.1 3.37 ;
      RECT 123.93 3.83 124.1 4.12 ;
      RECT 123.93 3.37 124.1 3.66 ;
      RECT 118.91 4.12 124.1 4.29 ;
      RECT 123.93 3.66 129.13 3.83 ;
      RECT 118.91 3.66 123.76 3.83 ;
      RECT 121.61 5.02 121.78 6.28 ;
      RECT 119.05 5.02 119.22 6.28 ;
      RECT 120.15 7.38 120.68 7.55 ;
      RECT 120.33 7.55 120.5 8.16 ;
      RECT 120.33 5.02 120.5 7.38 ;
      RECT 118.57 4.77 118.74 6.04 ;
      RECT 118.57 4.6 143.99 4.77 ;
      RECT 122.71 6.88 123.24 7.05 ;
      RECT 122.89 5.02 123.06 6.88 ;
      RECT 122.89 7.05 123.06 9.79 ;
      RECT 123.26 6.51 123.79 6.68 ;
      RECT 123.44 6.68 123.61 9.79 ;
      RECT 123.44 5.02 123.61 6.51 ;
      RECT 120.67 6.51 122.7 6.68 ;
      RECT 121.61 7.08 121.78 9.79 ;
      RECT 124.14 6.51 125.83 6.68 ;
      RECT 82.98 5.225 85.69 5.395 ;
      RECT 80.5 9.215 81.85 9.385 ;
      RECT 82.98 9.785 85.69 9.955 ;
      RECT 82.98 7.505 85.69 7.675 ;
      RECT 87.275 4.635 90.02 4.815 ;
      RECT 89.84 4.815 90.02 18.835 ;
      RECT 87.275 34.06 90.02 34.24 ;
      RECT 89.84 19.705 90.02 34.06 ;
      RECT 87.275 4.815 87.455 34.06 ;
      RECT 88.085 7.585 89.16 7.755 ;
      RECT 89.42 5.45 89.59 9.89 ;
      RECT 85.91 5.37 86.09 28.05 ;
      RECT 88.15 5.225 89.16 5.395 ;
      RECT 88.15 9.945 89.16 10.115 ;
      RECT 88.15 6.405 89.16 6.575 ;
      RECT 88.15 8.765 89.16 8.935 ;
      RECT 90.785 12.515 93.605 12.695 ;
      RECT 90.785 4.635 93.605 4.815 ;
      RECT 93.425 4.815 93.605 12.515 ;
      RECT 90.375 7.175 90.965 7.345 ;
      RECT 90.785 7.345 90.965 12.515 ;
      RECT 90.785 4.815 90.965 7.175 ;
      RECT 92.935 5.45 93.105 8.69 ;
      RECT 92.935 9.52 93.105 11.985 ;
      RECT 91.695 5.225 92.705 5.395 ;
      RECT 91.695 8.745 92.705 8.915 ;
      RECT 91.695 9.295 92.705 9.465 ;
      RECT 91.695 6.105 92.705 6.275 ;
      RECT 91.695 6.985 92.705 7.155 ;
      RECT 91.695 7.865 92.705 8.035 ;
      RECT 97.24 2.815 99.76 2.985 ;
      RECT 99.59 2.985 99.76 6.745 ;
      RECT 99.885 10.05 100.195 10.585 ;
      RECT 97.24 8.025 97.67 10.585 ;
      RECT 99.59 9.64 100.195 10.05 ;
      RECT 97.5 7.485 97.67 8.025 ;
      RECT 97.24 2.985 97.67 7.485 ;
      RECT 97.24 10.585 100.195 10.895 ;
      RECT 100.67 2.885 100.84 6.745 ;
      RECT 105.23 26.92 124.675 27.09 ;
      RECT 130.55 19.52 130.72 20.525 ;
      RECT 100.67 36.235 103 36.405 ;
      RECT 100.67 13.335 100.84 36.235 ;
      RECT 100.67 13.165 102.46 13.335 ;
      RECT 100.67 2.715 108.535 2.885 ;
      RECT 124.49 25.74 124.675 26.92 ;
      RECT 102.83 24.905 103 36.235 ;
      RECT 124.865 25.74 125.245 25.815 ;
      RECT 126.075 25.74 130.72 25.815 ;
      RECT 130.55 24.09 130.72 25.13 ;
      RECT 130.55 25.13 130.755 25.57 ;
      RECT 104.835 24.905 105.415 25.75 ;
      RECT 105.23 25.75 105.415 26.92 ;
      RECT 124.49 23.56 124.66 25.57 ;
      RECT 102.83 24.735 105.415 24.905 ;
      RECT 124.49 25.57 130.755 25.74 ;
      RECT 104.835 19.52 105.415 24.735 ;
      RECT 104.835 19.35 130.72 19.52 ;
      RECT 104.835 2.885 105.245 19.35 ;
      RECT 99.18 7.085 99.35 7.38 ;
      RECT 99.18 6.28 99.35 6.915 ;
      RECT 99.18 6.915 101.25 7.085 ;
      RECT 101.08 7.085 101.25 7.38 ;
      RECT 101.08 6.28 101.25 6.915 ;
      RECT 99.18 3.52 99.35 6 ;
      RECT 97.92 6.055 98.93 6.225 ;
      RECT 97.92 3.295 98.93 3.465 ;
      RECT 97.92 6.515 98.93 6.685 ;
      RECT 97.92 5.595 98.93 5.765 ;
      RECT 97.92 5.135 98.93 5.305 ;
      RECT 97.92 4.675 98.93 4.845 ;
      RECT 97.92 4.215 98.93 4.385 ;
      RECT 97.92 3.755 98.93 3.925 ;
      RECT 99.18 7.91 101.25 8.08 ;
      RECT 101.08 8.08 101.25 8.66 ;
      RECT 99.18 8.08 99.35 8.99 ;
      RECT 97.92 7.985 98.93 8.18 ;
      RECT 99.575 8.995 99.745 9.055 ;
      RECT 99.59 8.25 99.76 8.885 ;
      RECT 99.575 8.885 99.76 8.995 ;
      RECT 99.59 7.255 99.76 7.74 ;
      RECT 97.92 8.485 98.93 8.685 ;
      RECT 101.08 9.45 101.25 9.54 ;
      RECT 99.1 9.225 101.25 9.45 ;
      RECT 101.08 8.87 101.25 9.225 ;
      RECT 97.92 7.435 98.93 7.605 ;
      RECT 97.92 7.345 98.88 7.435 ;
      RECT 99.18 10.245 99.715 10.415 ;
      RECT 99.18 9.745 99.35 10.245 ;
      RECT 100.295 8.815 100.84 8.985 ;
      RECT 100.67 8.985 100.84 8.995 ;
      RECT 100.67 8.25 100.84 8.815 ;
      RECT 100.67 7.255 100.84 7.74 ;
      RECT 100.67 10.83 102.455 10.875 ;
      RECT 100.67 10.875 102.46 12.745 ;
      RECT 100.67 9.7 100.84 10.83 ;
      RECT 97.92 9.575 98.93 9.745 ;
      RECT 97.92 9.045 98.93 9.215 ;
      RECT 97.92 6.975 98.93 7.145 ;
      RECT 106.61 11.32 107.14 11.49 ;
      RECT 106.61 11.49 106.78 12.47 ;
      RECT 106.61 7.72 106.78 11.32 ;
      RECT 106 7.72 106.23 8.95 ;
      RECT 106 11.7 106.23 12.71 ;
      RECT 106.03 12.71 106.2 12.74 ;
      RECT 106.03 8.95 106.2 11.7 ;
      RECT 106.03 7.2 109.97 7.37 ;
      RECT 106.03 7.37 106.2 7.72 ;
      RECT 109.8 7.37 109.97 12.65 ;
      RECT 108.04 7.37 108.21 12.65 ;
      RECT 101.08 3.52 101.25 6 ;
      RECT 103.015 3.395 104.485 3.655 ;
      RECT 105.845 5.935 108.555 6.105 ;
      RECT 105.505 3.465 105.675 5.055 ;
      RECT 105.505 3.295 108.555 3.465 ;
      RECT 105.505 5.055 108.555 5.225 ;
      RECT 101.47 3.295 102.48 3.465 ;
      RECT 101.47 6.055 102.48 6.225 ;
      RECT 105.845 4.175 108.555 4.345 ;
      RECT 101.47 3.755 102.48 3.925 ;
      RECT 101.47 4.215 102.48 4.385 ;
      RECT 101.47 4.675 102.48 4.845 ;
      RECT 101.47 5.135 102.48 5.305 ;
      RECT 101.47 5.595 102.48 5.765 ;
      RECT 101.47 7.345 102.48 7.605 ;
      RECT 101.47 8.485 102.48 8.685 ;
      RECT 101.47 7.985 102.48 8.155 ;
      RECT 31.47 2.235 31.98 2.905 ;
      RECT 31.49 3.925 32 4.595 ;
      RECT 33.53 3.925 36.835 4.595 ;
      RECT 31.73 6.5 32.025 9.84 ;
      RECT 31.73 9.915 31.9 10.035 ;
      RECT 31.73 9.84 32 9.915 ;
      RECT 31.73 6.305 32 6.5 ;
      RECT 35.77 5.945 38.48 6.115 ;
      RECT 35.77 11.505 38.48 11.675 ;
      RECT 35.77 12.785 38.48 12.955 ;
      RECT 35.77 10.225 38.48 10.395 ;
      RECT 36.035 5.93 38.48 5.945 ;
      RECT 36.035 11.675 38.48 12.785 ;
      RECT 36.035 10.395 38.48 11.505 ;
      RECT 36.035 6.115 38.48 10.225 ;
      RECT 35.38 6.305 35.55 10.035 ;
      RECT 32.12 5.945 34.83 6.115 ;
      RECT 39.855 3.925 40.63 4.595 ;
      RECT 41.985 3.925 42.67 4.595 ;
      RECT 40.375 2.335 40.905 2.505 ;
      RECT 40.385 2.505 40.895 2.905 ;
      RECT 40.385 2.235 40.895 2.335 ;
      RECT 38.18 3.925 38.875 4.595 ;
      RECT 42.565 6.5 42.85 9.84 ;
      RECT 42.68 6.305 42.85 6.5 ;
      RECT 42.565 23.58 42.85 26.92 ;
      RECT 42.68 26.92 42.85 27.115 ;
      RECT 42.68 9.84 42.85 23.58 ;
      RECT 39.03 14.955 39.62 15.125 ;
      RECT 39.03 17.515 39.62 17.685 ;
      RECT 39.03 15.905 39.2 17.515 ;
      RECT 39.03 15.735 39.62 15.905 ;
      RECT 39.03 15.125 39.2 15.735 ;
      RECT 39.03 18.295 39.62 18.465 ;
      RECT 39.03 17.685 39.2 18.295 ;
      RECT 39.03 6.305 39.2 14.955 ;
      RECT 39.03 18.465 39.2 27.115 ;
      RECT 39.42 5.945 42.13 6.115 ;
      RECT 46.565 6.34 46.735 16.19 ;
      RECT 45.385 6.34 45.555 16.19 ;
      RECT 44.205 6.34 44.375 16.19 ;
      RECT 46.055 3.925 46.6 4.595 ;
      RECT 43.87 3.925 44.525 4.595 ;
      RECT 44.54 5.82 45.21 5.99 ;
      RECT 45.72 5.815 46.39 5.985 ;
      RECT 48.16 6.51 48.81 6.84 ;
      RECT 48.16 7.14 48.81 7.47 ;
      RECT 48.16 5.88 48.81 6.21 ;
      RECT 48.16 5.25 48.81 5.58 ;
      RECT 48.16 4.62 48.81 4.95 ;
      RECT 48.16 7.77 48.81 8.1 ;
      RECT 48.16 9.66 48.81 9.99 ;
      RECT 48.16 9.03 48.81 9.36 ;
      RECT 48.16 8.4 48.81 8.73 ;
      RECT 52.785 2.755 53.315 2.925 ;
      RECT 52.805 2.235 53.315 2.755 ;
      RECT 60.39 8.48 60.98 8.65 ;
      RECT 60.47 8.65 60.98 8.73 ;
      RECT 60.47 8.4 60.98 8.48 ;
      RECT 60.22 7.85 60.95 8.02 ;
      RECT 60.22 8.02 60.87 8.1 ;
      RECT 60.22 7.77 60.87 7.85 ;
      RECT 56.96 8.4 57.61 8.73 ;
      RECT 56.93 9.03 57.58 9.36 ;
      RECT 58.93 7.14 59.58 7.47 ;
      RECT 55.53 8.4 56.18 8.73 ;
      RECT 56.53 7.77 57.18 8.1 ;
      RECT 64.73 7.77 65.38 8.1 ;
      RECT 65.76 8.4 66.41 8.73 ;
      RECT 65.76 9.03 66.41 9.36 ;
      RECT 64.73 8.4 65.38 8.73 ;
      RECT 65.76 7.77 66.41 8.1 ;
      RECT 64.73 9.03 65.38 9.36 ;
      RECT 61.36 9.03 62.01 9.36 ;
      RECT 61.7 8.65 61.87 8.73 ;
      RECT 61.7 8.4 61.87 8.48 ;
      RECT 61.36 8.65 61.53 8.73 ;
      RECT 61.36 8.48 61.95 8.65 ;
      RECT 61.36 8.4 61.53 8.48 ;
      RECT 60.93 6.51 61.58 6.84 ;
      RECT 61.96 6.51 62.61 6.84 ;
      RECT 69.19 8.48 69.92 8.65 ;
      RECT 69.27 8.65 69.92 8.73 ;
      RECT 69.27 8.4 69.92 8.48 ;
      RECT 69.13 7.77 69.78 8.1 ;
      RECT 68.53 9.66 69.18 9.99 ;
      RECT 69.13 9.03 69.78 9.36 ;
      RECT 69.33 6.51 69.98 6.84 ;
      RECT 69.33 5.25 69.98 5.58 ;
      RECT 69.3 4.62 69.98 4.95 ;
      RECT 69.33 5.88 69.98 6.21 ;
      RECT 73.98 5.61 74.15 10.01 ;
      RECT 73.85 29.87 74.99 30.38 ;
      RECT 76.2 12.67 76.37 20.495 ;
      RECT 77.66 12.67 78.51 20.495 ;
      RECT 73.35 28.535 78.51 28.705 ;
      RECT 73.85 28.705 78.51 29.87 ;
      RECT 73.35 4.885 73.52 28.535 ;
      RECT 73.35 4.67 78.51 4.885 ;
      RECT 76.2 4.885 78.51 12.67 ;
      RECT 76.2 20.495 78.51 28.535 ;
      RECT 74.37 7.725 75.38 7.895 ;
      RECT 74.37 5.385 75.38 5.555 ;
      RECT 74.37 9.285 75.38 9.455 ;
      RECT 74.37 8.505 75.38 8.675 ;
      RECT 74.37 6.165 75.38 6.335 ;
      RECT 74.37 6.945 75.38 7.115 ;
      RECT 79.28 28.605 86.51 28.785 ;
      RECT 79.28 4.635 86.51 4.815 ;
      RECT 86.33 4.815 86.51 28.605 ;
      RECT 79.28 7.825 80.28 8.295 ;
      RECT 79.28 15.145 81.85 15.315 ;
      RECT 79.28 8.295 79.46 14.985 ;
      RECT 79.28 14.985 80.28 15.145 ;
      RECT 79.28 25.125 80.28 25.595 ;
      RECT 79.28 7.655 81.85 7.825 ;
      RECT 79.28 25.765 79.46 28.605 ;
      RECT 79.28 25.595 81.85 25.765 ;
      RECT 79.28 18.105 80.28 18.435 ;
      RECT 79.28 18.435 79.46 25.125 ;
      RECT 79.28 15.315 79.46 18.105 ;
      RECT 79.28 4.815 79.46 7.655 ;
      RECT 80.5 15.315 81.85 15.625 ;
      RECT 82.26 5.43 82.43 15.68 ;
      RECT 80.5 9.995 81.85 10.165 ;
      RECT 80.5 8.435 81.85 8.605 ;
      RECT 80.5 5.375 81.85 5.545 ;
      RECT 26.44 28.365 26.62 37.515 ;
      RECT 51.8 34.29 71.625 34.47 ;
      RECT 26.44 37.515 51.98 37.695 ;
      RECT 52.58 29.49 52.75 34.29 ;
      RECT 57.595 29.49 57.765 34.29 ;
      RECT 62.645 29.49 62.815 34.29 ;
      RECT 66.945 29.49 67.115 34.29 ;
      RECT 51.8 34.47 51.98 37.515 ;
      RECT 71.445 25.605 72.025 26 ;
      RECT 71.445 0.93 71.625 25.605 ;
      RECT 71.445 29.49 71.625 34.29 ;
      RECT 30.865 29.32 71.625 29.49 ;
      RECT 71.445 26 71.625 29.32 ;
      RECT 29.945 0.93 30.125 28.185 ;
      RECT 61.715 1.885 62.525 2.985 ;
      RECT 162.77 1.81 162.94 4.08 ;
      RECT 162.77 1.64 167.1 1.81 ;
      RECT 162.77 4.08 167.1 4.25 ;
      RECT 166.93 1.81 167.1 4.08 ;
      RECT 161.84 0.88 162.01 5.035 ;
      RECT 161.84 0.71 168.03 0.88 ;
      RECT 161.02 5.735 161.72 15.795 ;
      RECT 167.615 5.735 168.315 15.795 ;
      RECT 174.21 5.735 174.91 15.795 ;
      RECT 167.615 16.495 168.315 26.555 ;
      RECT 161.02 16.495 161.72 26.555 ;
      RECT 174.21 16.495 174.91 26.555 ;
      RECT 167.86 0.88 168.03 5.035 ;
      RECT 161.02 5.035 174.91 5.735 ;
      RECT 161.02 15.795 174.91 16.495 ;
      RECT 161.02 26.555 174.91 27.255 ;
      RECT 221.975 0.71 228.165 0.88 ;
      RECT 227.995 0.88 228.165 5.035 ;
      RECT 215.095 5.735 215.795 15.795 ;
      RECT 221.69 5.735 222.39 15.795 ;
      RECT 228.285 5.735 228.985 15.795 ;
      RECT 215.095 16.495 215.795 26.555 ;
      RECT 221.69 16.495 222.39 26.555 ;
      RECT 228.285 16.495 228.985 26.555 ;
      RECT 221.975 0.88 222.145 5.035 ;
      RECT 215.095 5.035 228.985 5.735 ;
      RECT 215.095 15.795 228.985 16.495 ;
      RECT 215.095 26.555 228.985 27.255 ;
      RECT 227.065 1.81 227.235 4.08 ;
      RECT 222.905 1.64 227.235 1.81 ;
      RECT 222.905 4.08 227.235 4.25 ;
      RECT 222.905 1.81 223.075 4.08 ;
      RECT 327.48 1.885 328.29 2.985 ;
      RECT 318.38 0.75 360.06 0.93 ;
      RECT 359.88 28.185 363.565 28.365 ;
      RECT 318.38 34.29 338.205 34.47 ;
      RECT 363.385 28.365 363.565 37.515 ;
      RECT 322.89 29.49 323.06 34.29 ;
      RECT 327.19 29.49 327.36 34.29 ;
      RECT 332.24 29.49 332.41 34.29 ;
      RECT 337.255 29.49 337.425 34.29 ;
      RECT 338.025 34.47 338.205 37.515 ;
      RECT 338.025 37.515 363.565 37.695 ;
      RECT 317.98 25.605 318.56 26 ;
      RECT 318.38 0.93 318.56 25.605 ;
      RECT 318.38 29.49 318.56 34.29 ;
      RECT 318.38 29.32 359.14 29.49 ;
      RECT 318.38 26 318.56 29.32 ;
      RECT 359.88 0.93 360.06 28.185 ;
      RECT 10.9 3.135 11.07 16.245 ;
      RECT 21.95 3.665 22.65 13.725 ;
      RECT 15.355 16.745 16.055 26.805 ;
      RECT 21.95 16.745 22.65 26.805 ;
      RECT 28.545 3.665 29.245 13.725 ;
      RECT 28.545 16.745 29.245 26.805 ;
      RECT 15.355 26.805 29.245 27.505 ;
      RECT 10.9 2.965 29.245 3.135 ;
      RECT 15.1 14.425 15.27 16.045 ;
      RECT 15.1 16.045 29.245 16.245 ;
      RECT 15.355 16.415 29.245 16.745 ;
      RECT 10.9 16.245 29.245 16.415 ;
      RECT 15.1 3.665 16.055 13.725 ;
      RECT 15.1 13.725 29.245 14.425 ;
      RECT 15.1 3.135 29.245 3.665 ;
      RECT 11.83 3.905 14.34 4.075 ;
      RECT 14.17 4.075 14.34 15.315 ;
      RECT 11.83 15.315 14.34 15.485 ;
      RECT 11.83 4.075 12 15.315 ;
      RECT 12.635 4.315 13.535 4.485 ;
      RECT 12.75 4.485 13.42 14.905 ;
      RECT 12.635 14.905 13.945 15.075 ;
      RECT 18.335 5.42 19.66 5.83 ;
      RECT 16.815 5.135 17.515 12.265 ;
      RECT 16.815 4.425 21.19 5.135 ;
      RECT 16.815 12.265 21.19 12.965 ;
      RECT 20.49 5.135 21.19 12.265 ;
      RECT 17.99 6 18.53 11.395 ;
      RECT 19.465 6 20.005 11.395 ;
      RECT 24.94 5.42 26.265 5.83 ;
      RECT 23.41 5.135 24.11 12.265 ;
      RECT 23.41 4.425 27.785 5.135 ;
      RECT 23.41 12.265 27.785 12.965 ;
      RECT 27.085 5.135 27.785 12.265 ;
      RECT 24.595 6 25.135 11.395 ;
      RECT 43.2 5.415 43.37 28.375 ;
      RECT 31.3 28.375 70.68 28.555 ;
      RECT 47.335 4.01 70.68 4.19 ;
      RECT 31.3 5.235 47.515 5.415 ;
      RECT 31.3 15.485 31.5 16.91 ;
      RECT 31.3 16.91 31.48 28.375 ;
      RECT 47.615 28.555 70.645 28.565 ;
      RECT 47.805 21.685 69.605 21.695 ;
      RECT 47.805 21.165 69.605 21.175 ;
      RECT 69.95 11.865 70.68 12.535 ;
      RECT 69.95 19.635 70.68 20.305 ;
      RECT 47.335 11.865 48.28 12.535 ;
      RECT 47.335 10.99 47.515 11.865 ;
      RECT 70.5 12.535 70.68 19.635 ;
      RECT 70.5 10.99 70.68 11.865 ;
      RECT 70.5 4.19 70.68 10.48 ;
      RECT 47.335 12.535 47.515 19.635 ;
      RECT 70.5 21.685 70.68 28.375 ;
      RECT 70.5 20.305 70.68 21.175 ;
      RECT 47.335 21.175 70.68 21.685 ;
      RECT 47.335 20.305 47.515 21.175 ;
      RECT 47.335 5.415 47.515 10.48 ;
      RECT 31.3 5.415 31.48 15.485 ;
      RECT 47.335 4.19 47.515 5.235 ;
      RECT 47.335 21.685 47.515 28.375 ;
      RECT 47.335 19.635 48.28 20.305 ;
      RECT 47.335 10.48 70.68 10.99 ;
      RECT 26.07 6 26.61 11.395 ;
      RECT 326.745 54.67 326.955 58.76 ;
      RECT 63.05 54.67 63.26 58.76 ;
      RECT 36.145 54.67 36.355 58.79 ;
      RECT 276.595 54.66 276.765 55.565 ;
      RECT 113.24 54.66 113.41 55.565 ;
      RECT 326.745 54.46 353.86 54.67 ;
      RECT 36.145 54.46 63.26 54.67 ;
      RECT 276.235 54.385 276.765 54.66 ;
      RECT 274.115 54.385 275.44 54.66 ;
      RECT 278.07 54.385 278.24 55.575 ;
      RECT 113.24 54.385 113.77 54.66 ;
      RECT 114.565 54.385 115.89 54.66 ;
      RECT 111.765 54.385 111.935 55.575 ;
      RECT 274.115 54.055 278.24 54.385 ;
      RECT 111.765 54.055 115.89 54.385 ;
      RECT 275.275 53.935 278.24 54.055 ;
      RECT 111.765 53.935 114.73 54.055 ;
      RECT 274.115 53.77 274.645 54.055 ;
      RECT 276.235 53.77 278.24 53.935 ;
      RECT 115.36 53.77 115.89 54.055 ;
      RECT 111.765 53.77 113.77 53.935 ;
      RECT 279.285 53.6 295.115 54.78 ;
      RECT 276.415 53.6 278.24 53.77 ;
      RECT 94.89 53.6 110.72 54.78 ;
      RECT 111.765 53.6 113.59 53.77 ;
      RECT 274.115 52.775 274.565 53.77 ;
      RECT 275.275 52.875 275.485 53.935 ;
      RECT 115.44 52.775 115.89 53.77 ;
      RECT 114.52 52.875 114.73 53.935 ;
      RECT 274.115 51.91 274.3 52.775 ;
      RECT 115.705 51.91 115.89 52.775 ;
      RECT 275.275 51.885 275.475 52.875 ;
      RECT 114.53 51.885 114.73 52.875 ;
      RECT 274.115 51.74 274.645 51.91 ;
      RECT 306.855 51.72 307.025 54.78 ;
      RECT 308.615 51.72 308.785 54.78 ;
      RECT 310.375 51.72 310.545 54.78 ;
      RECT 312.135 51.72 312.305 54.78 ;
      RECT 313.895 51.72 314.065 54.78 ;
      RECT 320.935 51.72 321.105 54.78 ;
      RECT 319.175 51.72 319.345 54.78 ;
      RECT 317.415 51.72 317.585 54.78 ;
      RECT 315.655 51.72 315.825 54.78 ;
      RECT 322.695 51.72 322.865 54.78 ;
      RECT 296.405 51.72 296.575 54.78 ;
      RECT 298.715 51.72 298.885 54.78 ;
      RECT 300.475 51.72 300.645 54.78 ;
      RECT 302.235 51.72 302.405 54.78 ;
      RECT 115.36 51.74 115.89 51.91 ;
      RECT 89.36 51.72 89.53 54.78 ;
      RECT 87.6 51.72 87.77 54.78 ;
      RECT 93.43 51.72 93.6 54.78 ;
      RECT 91.12 51.72 91.29 54.78 ;
      RECT 67.14 51.72 67.31 54.78 ;
      RECT 68.9 51.72 69.07 54.78 ;
      RECT 70.66 51.72 70.83 54.78 ;
      RECT 72.42 51.72 72.59 54.78 ;
      RECT 77.7 51.72 77.87 54.78 ;
      RECT 75.94 51.72 76.11 54.78 ;
      RECT 74.18 51.72 74.35 54.78 ;
      RECT 82.98 51.72 83.15 54.78 ;
      RECT 81.22 51.72 81.39 54.78 ;
      RECT 79.46 51.72 79.63 54.78 ;
      RECT 276.415 51.555 295.115 53.6 ;
      RECT 323.275 51.41 325.845 54.78 ;
      RECT 94.89 51.555 113.59 53.6 ;
      RECT 64.16 51.41 66.73 54.78 ;
      RECT 345.3 51.195 353.86 54.46 ;
      RECT 36.145 51.195 44.705 54.46 ;
      RECT 275.275 50.875 275.485 51.885 ;
      RECT 274.115 50.875 274.565 51.74 ;
      RECT 114.52 50.875 114.73 51.885 ;
      RECT 115.44 50.875 115.89 51.74 ;
      RECT 276.41 50.6 295.115 51.555 ;
      RECT 94.89 50.6 113.595 51.555 ;
      RECT 276.41 50.405 293.435 50.6 ;
      RECT 96.57 50.405 113.595 50.6 ;
      RECT 276.095 49.975 293.435 50.405 ;
      RECT 96.57 49.975 113.91 50.405 ;
      RECT 276.095 49.76 281.95 49.79 ;
      RECT 276.095 49.79 290.205 49.975 ;
      RECT 276.095 49.735 278.505 49.76 ;
      RECT 108.055 49.76 113.91 49.79 ;
      RECT 99.8 49.79 113.91 49.975 ;
      RECT 111.5 49.735 113.91 49.76 ;
      RECT 276.325 49.28 278.505 49.735 ;
      RECT 111.5 49.28 113.68 49.735 ;
      RECT 345.3 46.875 346.795 51.195 ;
      RECT 326.745 46.875 326.955 54.46 ;
      RECT 43.21 46.875 44.705 51.195 ;
      RECT 63.05 46.875 63.26 54.46 ;
      RECT 326.745 46.705 355.51 46.875 ;
      RECT 326.745 46.61 327.37 46.705 ;
      RECT 34.495 46.705 63.26 46.875 ;
      RECT 62.635 46.61 63.26 46.705 ;
      RECT 355.05 46.165 355.51 46.705 ;
      RECT 327.065 46.165 327.37 46.61 ;
      RECT 34.495 46.165 34.955 46.705 ;
      RECT 62.635 46.165 62.94 46.61 ;
      RECT 327.065 45.835 348.06 46.165 ;
      RECT 353.8 45.835 355.51 46.165 ;
      RECT 41.945 45.835 62.94 46.165 ;
      RECT 34.495 45.835 36.205 46.165 ;
      RECT 355.05 44.15 355.51 45.835 ;
      RECT 34.495 44.15 34.955 45.835 ;
      RECT 355.05 44.145 363.915 44.15 ;
      RECT 26.09 44.145 34.955 44.15 ;
      RECT 355.05 43.98 364.06 44.145 ;
      RECT 25.945 43.98 34.955 44.145 ;
      RECT 327.065 43.52 327.37 45.835 ;
      RECT 62.635 43.52 62.94 45.835 ;
      RECT 309.295 43.35 327.37 43.52 ;
      RECT 62.635 43.35 80.71 43.52 ;
      RECT 363.745 39.745 364.06 43.98 ;
      RECT 25.945 39.745 26.26 43.98 ;
      RECT 336.66 39.575 364.06 39.745 ;
      RECT 25.945 39.575 53.345 39.745 ;
      RECT 177.32 37.11 212.685 88.63 ;
      RECT 183.94 0.33 205.86 37.11 ;
      RECT 336.66 36.61 336.945 39.575 ;
      RECT 309.295 36.44 336.945 36.61 ;
      RECT 309.295 36.61 309.465 43.35 ;
      RECT 53.06 36.61 53.345 39.575 ;
      RECT 53.06 36.44 80.71 36.61 ;
      RECT 80.54 36.61 80.71 43.35 ;
      RECT 29.945 0.75 71.625 0.93 ;
      RECT 26.44 28.185 30.125 28.365 ;
      RECT 29.145 125.5 30.035 127.655 ;
      RECT 29.165 122.7 30.015 125.5 ;
      RECT 29.145 117.405 30.035 122.7 ;
      RECT 29.165 115.48 30.015 117.405 ;
      RECT 29.145 112.835 30.035 115.48 ;
      RECT 29.165 108.215 30.015 112.835 ;
      RECT 29.145 103.775 30.035 108.215 ;
      RECT 29.165 99.415 30.015 103.775 ;
      RECT 29.145 97.085 30.035 99.415 ;
      RECT 29.165 94.985 30.015 97.085 ;
      RECT 29.145 89.825 30.035 94.985 ;
      RECT 29.165 88.205 30.015 89.825 ;
      RECT 29.145 86.645 30.035 88.205 ;
      RECT 29.165 84.41 30.015 86.645 ;
      RECT 1.13 40.64 7.13 187.555 ;
      RECT 1.13 17.505 10.44 40.64 ;
      RECT 1.12 0.335 9.38 17.505 ;
      RECT 176.755 175.1 213.25 253.24 ;
      RECT 90.45 102.115 116.88 107.805 ;
      RECT 273.125 102.115 299.555 107.805 ;
      RECT 191.735 95.265 198.365 175.1 ;
      RECT 236.555 95.265 299.555 102.115 ;
      RECT 90.45 95.265 153.45 102.115 ;
      RECT 90.45 93.98 299.555 95.265 ;
      RECT 90.435 93.07 299.57 93.98 ;
      RECT 291.18 92.01 299.57 93.07 ;
      RECT 90.435 92.01 98.825 93.07 ;
      RECT 146.79 88.63 243.215 93.07 ;
      RECT 291.18 88.625 299.555 92.01 ;
      RECT 90.45 88.625 98.825 92.01 ;
      RECT 291.185 85.3 299.555 88.625 ;
      RECT 90.45 85.3 98.82 88.625 ;
      RECT 291.185 75.535 297.14 85.3 ;
      RECT 290.14 74.525 297.14 75.535 ;
      RECT 92.865 75.535 98.82 85.3 ;
      RECT 92.865 74.525 99.865 75.535 ;
      RECT 362.36 72.42 372.185 72.73 ;
      RECT 17.82 72.42 27.645 72.73 ;
      RECT 305.42 71.83 372.185 72.42 ;
      RECT 305.42 71.56 372.12 71.83 ;
      RECT 17.82 71.83 84.585 72.42 ;
      RECT 17.885 71.56 84.585 71.83 ;
      RECT 305.42 71.04 363.05 71.56 ;
      RECT 292.035 71.04 297.14 74.525 ;
      RECT 26.955 71.04 84.585 71.56 ;
      RECT 92.865 71.04 97.97 74.525 ;
      RECT 292.035 70.42 363.05 71.04 ;
      RECT 26.955 70.42 97.97 71.04 ;
      RECT 311.675 69.665 324.515 69.835 ;
      RECT 65.49 69.665 78.33 69.835 ;
      RECT 292.035 69.04 307.42 70.42 ;
      RECT 82.585 69.04 97.97 70.42 ;
      RECT 325.96 68.33 363.05 70.42 ;
      RECT 26.955 68.33 64.045 70.42 ;
      RECT 325.93 68.1 363.05 68.33 ;
      RECT 26.955 68.1 64.075 68.33 ;
      RECT 345.065 66.305 363.05 68.1 ;
      RECT 26.955 66.305 44.94 68.1 ;
      RECT 311.675 63.645 314.475 69.665 ;
      RECT 75.53 63.645 78.33 69.665 ;
      RECT 345.065 63.565 355.47 66.305 ;
      RECT 34.535 63.565 44.94 66.305 ;
      RECT 345.065 63.355 355.455 63.565 ;
      RECT 34.55 63.355 44.94 63.565 ;
      RECT 292.035 63.07 293.175 69.04 ;
      RECT 96.83 63.07 97.97 69.04 ;
      RECT 290.14 62.78 294.5 63.07 ;
      RECT 95.505 62.78 99.865 63.07 ;
      RECT 345.065 62.505 345.235 63.355 ;
      RECT 355.245 62.505 355.455 63.355 ;
      RECT 44.77 62.505 44.94 63.355 ;
      RECT 34.55 62.505 34.76 63.355 ;
      RECT 345.065 60.035 355.455 62.505 ;
      RECT 290.14 60.605 294.515 62.78 ;
      RECT 34.55 60.035 44.94 62.505 ;
      RECT 95.49 60.605 99.865 62.78 ;
      RECT 345.065 59.885 345.235 60.035 ;
      RECT 343.965 59.885 344.175 59.925 ;
      RECT 44.77 59.885 44.94 60.035 ;
      RECT 45.83 59.885 46.04 59.925 ;
      RECT 345.955 59.795 346.125 60.035 ;
      RECT 354.515 59.795 354.685 60.035 ;
      RECT 350.235 59.795 350.405 60.035 ;
      RECT 343.965 59.595 344.175 59.635 ;
      RECT 343.885 59.635 345.235 59.885 ;
      RECT 35.32 59.795 35.49 60.035 ;
      RECT 39.6 59.795 39.77 60.035 ;
      RECT 43.88 59.795 44.05 60.035 ;
      RECT 45.83 59.595 46.04 59.635 ;
      RECT 44.77 59.635 46.12 59.885 ;
      RECT 279.285 59.255 294.515 60.605 ;
      RECT 95.49 59.255 110.72 60.605 ;
      RECT 355.245 59 355.455 60.035 ;
      RECT 345.065 59 345.235 59.635 ;
      RECT 34.55 59 34.76 60.035 ;
      RECT 44.77 59 44.94 59.635 ;
      RECT 325.93 58.99 326.16 68.1 ;
      RECT 63.845 58.99 64.075 68.1 ;
      RECT 345.065 58.96 355.455 59 ;
      RECT 325.93 58.96 336.675 58.99 ;
      RECT 34.55 58.96 44.94 59 ;
      RECT 53.33 58.96 64.075 58.99 ;
      RECT 279.285 58.725 294.625 59.255 ;
      RECT 325.93 58.76 336.675 58.79 ;
      RECT 325.93 58.79 355.455 58.96 ;
      RECT 95.38 58.725 110.72 59.255 ;
      RECT 53.33 58.76 64.075 58.79 ;
      RECT 34.55 58.79 64.075 58.96 ;
      RECT 324.345 58.085 324.515 69.665 ;
      RECT 65.49 58.085 65.66 69.665 ;
      RECT 279.285 56.715 294.515 58.725 ;
      RECT 95.49 56.715 110.72 58.725 ;
      RECT 279.285 56.185 294.59 56.715 ;
      RECT 95.415 56.185 110.72 56.715 ;
      RECT 312.725 56.075 314.475 63.645 ;
      RECT 324.345 56.075 325.845 58.085 ;
      RECT 75.53 56.075 77.28 63.645 ;
      RECT 64.16 56.075 65.66 58.085 ;
      RECT 312.725 55.645 325.845 56.075 ;
      RECT 64.16 55.645 77.28 56.075 ;
      RECT 279.285 55.295 294.515 56.185 ;
      RECT 297.72 55.295 325.845 55.645 ;
      RECT 95.49 55.295 110.72 56.185 ;
      RECT 64.16 55.295 92.285 55.645 ;
      RECT 279.285 54.78 325.845 55.295 ;
      RECT 64.16 54.78 110.72 55.295 ;
      RECT 353.65 54.67 353.86 58.79 ;
      RECT 467.82 244.115 470.48 253.385 ;
      RECT 450.085 242.39 470.48 244.115 ;
      RECT 450.64 240.72 451.22 242.39 ;
      RECT 455.955 240.72 456.535 242.39 ;
      RECT 452.715 240.72 454.605 242.39 ;
      RECT 419.1 240.29 420.68 243.86 ;
      RECT 385 240.29 408.075 240.32 ;
      RECT 450.085 240.12 450.255 242.39 ;
      RECT 384.15 240.09 408.075 240.12 ;
      RECT 384.15 240.12 420.68 240.29 ;
      RECT 467.48 235.18 470.48 242.39 ;
      RECT 444.37 234.95 470.48 235.18 ;
      RECT 444.37 232.32 444.6 234.95 ;
      RECT 444.4 229.655 444.57 232.32 ;
      RECT 416.87 229.405 444.57 229.655 ;
      RECT 384.15 217.09 385.01 240.09 ;
      RECT 441.02 217.09 441.25 229.405 ;
      RECT 384.15 216.23 444.6 217.09 ;
      RECT 443.71 215.23 444.6 216.23 ;
      RECT 443.71 211.91 444.57 215.23 ;
      RECT 443.71 209.62 444.6 211.91 ;
      RECT 467.45 198.88 470.48 234.95 ;
      RECT 443.71 198.88 444.57 209.62 ;
      RECT 457.585 197.915 470.48 198.88 ;
      RECT 467.85 88.84 470.48 197.915 ;
      RECT 443.71 193.22 444.6 198.88 ;
      RECT 467.98 88.77 470.48 88.84 ;
      RECT 457.585 193.22 458.545 197.915 ;
      RECT 443.71 192.1 458.545 193.22 ;
      RECT 386.205 199.94 428.415 200.145 ;
      RECT 393.445 199.58 393.675 199.94 ;
      RECT 428.235 188.345 428.415 199.94 ;
      RECT 428.235 182.415 428.48 188.345 ;
      RECT 428.235 182.19 428.475 182.415 ;
      RECT 393.445 182.19 393.625 199.58 ;
      RECT 393.445 182.01 428.475 182.19 ;
      RECT 406.625 156.1 406.805 182.01 ;
      RECT 393.445 156.1 393.625 182.01 ;
      RECT 419.805 156.1 419.985 182.01 ;
      RECT 393.445 155.92 419.985 156.1 ;
      RECT 393.45 154.95 393.62 155.23 ;
      RECT 406.625 147.89 406.805 155.92 ;
      RECT 393.445 147.89 393.625 154.95 ;
      RECT 392.495 147.71 406.805 147.89 ;
      RECT 396.105 147.14 396.285 147.71 ;
      RECT 386.205 147.14 386.385 199.94 ;
      RECT 392.495 147.14 392.675 147.71 ;
      RECT 384.775 146.96 396.285 147.14 ;
      RECT 419.805 145.715 419.985 155.92 ;
      RECT 406.625 145.715 406.805 147.71 ;
      RECT 396.105 145.715 396.285 146.96 ;
      RECT 396.105 145.535 397.305 145.715 ;
      RECT 398.945 145.535 419.985 145.715 ;
      RECT 384.775 136.24 384.955 146.96 ;
      RECT 396.105 121.915 396.285 145.535 ;
      RECT 407.78 121.915 408.31 145.535 ;
      RECT 419.805 121.915 419.985 145.535 ;
      RECT 396.105 121.735 419.985 121.915 ;
      RECT 418.095 109.84 418.885 121.735 ;
      RECT 407.955 109.66 408.135 121.735 ;
      RECT 397.205 109.66 397.99 121.735 ;
      RECT 418.095 109.66 425.725 109.84 ;
      RECT 418.095 109.47 418.885 109.66 ;
      RECT 397.205 63.185 397.385 109.66 ;
      RECT 425.545 63.185 425.725 109.66 ;
      RECT 397.205 63.005 425.725 63.185 ;
      RECT 425.545 48.6 425.725 63.005 ;
      RECT 445.155 48.6 445.335 51.285 ;
      RECT 425.545 48.42 445.335 48.6 ;
      RECT 397.205 39.145 397.385 63.005 ;
      RECT 418.705 39.145 418.885 63.005 ;
      RECT 396.105 38.465 396.285 121.735 ;
      RECT 397.205 38.965 418.885 39.145 ;
      RECT 418.71 38.465 418.88 38.965 ;
      RECT 396.105 38.145 418.88 38.465 ;
      RECT 1.175 250.14 40.82 253.385 ;
      RECT 1.175 227.215 24.38 250.14 ;
      RECT 1.175 202.71 16.405 227.215 ;
      RECT 1.175 195.58 40.82 202.71 ;
      RECT 20.06 193.23 20.23 195.58 ;
      RECT 34.045 192.515 40.82 195.58 ;
      RECT 20.005 190.495 20.255 193.23 ;
      RECT 1.175 187.555 19.475 195.58 ;
      RECT 18.06 186.695 19.475 187.555 ;
      RECT 36.08 186.695 40.82 192.515 ;
      RECT 18.06 186.105 40.82 186.695 ;
      RECT 18.06 185.455 22.205 186.105 ;
      RECT 27.95 184.215 40.82 186.105 ;
      RECT 18.06 181.365 22.49 185.455 ;
      RECT 18.06 178.695 21.78 181.365 ;
      RECT 34.8 178.605 34.97 183.39 ;
      RECT 42.75 178.605 42.92 183.39 ;
      RECT 18.06 177.695 22.28 178.695 ;
      RECT 34.68 178.435 35.21 178.605 ;
      RECT 42.51 178.435 43.04 178.605 ;
      RECT 18.06 176.43 21.78 177.695 ;
      RECT 34.8 176.43 34.97 178.435 ;
      RECT 42.75 176.43 42.92 178.435 ;
      RECT 18.06 174.835 48.865 176.43 ;
      RECT 42.82 174.055 48.865 174.835 ;
      RECT 18.06 173.75 18.965 174.835 ;
      RECT 45.73 173.485 48.865 174.055 ;
      RECT 18.06 172.935 18.68 173.75 ;
      RECT 42.82 172.905 48.865 173.485 ;
      RECT 46.535 171.515 48.865 172.905 ;
      RECT 42.82 171.345 48.865 171.515 ;
      RECT 46.535 169.955 48.865 171.345 ;
      RECT 42.82 169.785 48.865 169.955 ;
      RECT 46.535 168.395 48.865 169.785 ;
      RECT 42.82 168.225 48.865 168.395 ;
      RECT 46.535 167.875 48.865 168.225 ;
      RECT 45.99 167.705 60.94 167.875 ;
      RECT 60.77 165.785 60.94 167.705 ;
      RECT 55.785 165.455 60.94 165.785 ;
      RECT 60.77 163.625 60.94 165.455 ;
      RECT 55.785 163.295 60.94 163.625 ;
      RECT 60.77 162.385 60.94 163.295 ;
      RECT 17.645 162.215 18.775 164.565 ;
      RECT 38.55 162.215 60.94 162.385 ;
      RECT 17.645 161.195 60.94 162.215 ;
      RECT 17.645 141.545 19.675 161.195 ;
      RECT 17.645 134.865 30.945 141.545 ;
      RECT 29.165 134.385 30.015 134.865 ;
      RECT 29.145 130.805 30.035 134.385 ;
      RECT 29.165 129.725 30.015 130.805 ;
      RECT 29.145 128.425 30.035 129.725 ;
      RECT 29.165 127.655 30.015 128.425 ;
      RECT 442.15 139.805 444.415 185.105 ;
      RECT 442.725 136.27 444.415 136.615 ;
      RECT 433.98 136.685 444.415 139.805 ;
      RECT 442.745 135.87 444.415 136.27 ;
      RECT 438.62 135.84 444.415 135.87 ;
      RECT 429.155 135.84 437.515 135.87 ;
      RECT 429.155 135.64 437.515 135.67 ;
      RECT 429.155 135.67 444.415 135.84 ;
      RECT 438.535 135.64 444.415 135.67 ;
      RECT 382.77 134.915 383.97 148.03 ;
      RECT 385.72 134.915 386.09 146.015 ;
      RECT 359.06 134.865 372.36 141.545 ;
      RECT 359.99 134.385 360.84 134.865 ;
      RECT 359.97 130.805 360.86 134.385 ;
      RECT 359.99 129.725 360.84 130.805 ;
      RECT 359.97 128.425 360.86 129.725 ;
      RECT 359.99 127.655 360.84 128.425 ;
      RECT 359.97 125.5 360.86 127.655 ;
      RECT 359.99 122.7 360.84 125.5 ;
      RECT 359.97 117.405 360.86 122.7 ;
      RECT 438.535 114.97 439.035 135.64 ;
      RECT 432.705 114.97 433.205 135.64 ;
      RECT 359.99 115.48 360.84 117.405 ;
      RECT 359.97 112.835 360.86 115.48 ;
      RECT 359.99 108.215 360.84 112.835 ;
      RECT 359.97 103.775 360.86 108.215 ;
      RECT 359.99 99.415 360.84 103.775 ;
      RECT 359.97 97.085 360.86 99.415 ;
      RECT 359.99 94.985 360.84 97.085 ;
      RECT 436.225 93.535 436.725 135.64 ;
      RECT 435.015 93.535 435.515 135.64 ;
      RECT 359.97 89.825 360.86 94.985 ;
      RECT 471.245 88.295 477.515 253.585 ;
      RECT 359.99 88.205 360.84 89.825 ;
      RECT 442.385 88.065 444.415 135.64 ;
      RECT 463.22 87.055 466.74 185.105 ;
      RECT 359.97 86.645 360.86 88.205 ;
      RECT 359.99 84.41 360.84 86.645 ;
      RECT 435.785 66.66 435.955 135.64 ;
      RECT 442.385 61.065 450.13 88.065 ;
      RECT 444.86 61.055 450.13 61.065 ;
      RECT 448.6 52.425 450.13 61.055 ;
      RECT 435.755 49.95 435.985 66.66 ;
      RECT 435.785 49.54 435.955 49.95 ;
      RECT 442.385 49.54 442.555 61.065 ;
      RECT 429.185 49.54 429.355 135.64 ;
      RECT 429.185 49.37 442.555 49.54 ;
      RECT 464.36 47.345 466.13 87.055 ;
      RECT 464.36 46.88 467.36 47.345 ;
      RECT 472.255 45.815 477.515 88.295 ;
      RECT 465.56 45.815 467.36 46.88 ;
      RECT 382.77 41.12 386.09 134.915 ;
      RECT 447.71 39.285 450.13 52.425 ;
      RECT 395.16 35.665 395.34 146.015 ;
      RECT 395.16 35.485 396.18 35.665 ;
      RECT 396.85 35.485 400.38 35.665 ;
      RECT 465.56 29 477.515 45.815 ;
      RECT 445.32 29 450.13 39.285 ;
      RECT 447.725 24.75 477.515 24.755 ;
      RECT 445.32 24.755 477.515 29 ;
      RECT 467.085 11.24 477.515 24.75 ;
      RECT 445.32 11.24 447.42 24.755 ;
      RECT 445.32 11.235 477.515 11.24 ;
      RECT 400.2 9.25 400.38 35.485 ;
      RECT 380.1 9.25 386.09 41.12 ;
      RECT 380.1 8.5 400.38 9.25 ;
      RECT 444.51 6.6 477.515 11.235 ;
      RECT 386.575 0.3 477.515 1.97 ;
      RECT 467.085 0.13 477.515 0.3 ;
      RECT 405.89 1.97 477.515 6.6 ;
      RECT 380.1 0.415 385.64 8.5 ;
      RECT 445.425 183.68 447.49 183.685 ;
      RECT 445.425 182.82 462.11 183.68 ;
      RECT 445.425 146.46 446.29 182.82 ;
      RECT 461.25 146.46 462.11 182.82 ;
      RECT 445.425 145.465 462.11 146.46 ;
      RECT 461.25 140.225 462.11 145.465 ;
      RECT 457.385 140.185 462.11 140.225 ;
      RECT 457.385 139.975 462.11 140.015 ;
      RECT 457.025 140.015 462.11 140.185 ;
      RECT 461.25 136.945 462.11 139.975 ;
      RECT 457.385 136.905 462.11 136.945 ;
      RECT 457.385 136.695 462.11 136.735 ;
      RECT 457.025 136.735 462.11 136.905 ;
      RECT 461.25 126.715 462.11 136.695 ;
      RECT 457.385 126.675 462.11 126.715 ;
      RECT 457.385 126.465 462.11 126.505 ;
      RECT 457.025 126.505 462.11 126.675 ;
      RECT 461.25 123.435 462.11 126.465 ;
      RECT 445.425 113.455 446.29 145.465 ;
      RECT 457.385 123.395 462.11 123.435 ;
      RECT 457.385 123.185 462.11 123.225 ;
      RECT 457.025 123.225 462.11 123.395 ;
      RECT 461.25 113.205 462.11 123.185 ;
      RECT 457.385 113.165 462.11 113.205 ;
      RECT 457.385 112.955 462.11 112.995 ;
      RECT 457.025 112.995 462.11 113.165 ;
      RECT 461.25 109.925 462.11 112.955 ;
      RECT 457.385 109.885 462.11 109.925 ;
      RECT 457.385 109.675 462.11 109.715 ;
      RECT 457.025 109.715 462.11 109.885 ;
      RECT 461.25 99.695 462.11 109.675 ;
      RECT 457.385 99.655 462.11 99.695 ;
      RECT 457.385 99.445 462.11 99.485 ;
      RECT 457.025 99.485 462.11 99.655 ;
      RECT 461.25 96.415 462.11 99.445 ;
      RECT 457.385 96.375 462.11 96.415 ;
      RECT 457.385 96.165 462.11 96.205 ;
      RECT 457.025 96.205 462.11 96.375 ;
      RECT 461.25 90.055 462.11 96.165 ;
      RECT 445.43 90.055 446.29 113.455 ;
      RECT 445.43 89.195 462.11 90.055 ;
      RECT 451.4 86.845 460.915 89.195 ;
      RECT 451.4 78.92 452.62 86.845 ;
      RECT 460.515 78.92 460.915 86.845 ;
      RECT 451.4 78.42 460.915 78.92 ;
      RECT 451.4 62.975 452.62 78.42 ;
      RECT 460.515 62.975 460.915 78.42 ;
      RECT 451.4 62.475 460.915 62.975 ;
      RECT 460.515 62.47 460.915 62.475 ;
      RECT 460.515 46.655 460.685 62.47 ;
      RECT 451.9 46.655 452.07 62.475 ;
      RECT 451.9 46.485 460.685 46.655 ;
      RECT 451.9 30.405 452.07 46.485 ;
      RECT 464.155 43.095 464.8 45.865 ;
      RECT 464.63 30.405 464.8 43.095 ;
      RECT 451.9 30.235 464.8 30.405 ;
      RECT 7.78 41.925 8.01 184.54 ;
      RECT 7.78 184.54 17.24 184.77 ;
      RECT 17.01 82.505 17.24 184.54 ;
      RECT 15.1 53.7 17.21 53.87 ;
      RECT 14.31 42.79 15.27 42.96 ;
      RECT 15.1 42.96 15.27 53.7 ;
      RECT 7.78 41.725 14.48 41.895 ;
      RECT 7.78 41.895 11.68 41.925 ;
      RECT 7.78 41.695 11.68 41.725 ;
      RECT 17.04 53.87 17.21 82.505 ;
      RECT 14.31 41.895 14.48 42.79 ;
      RECT 381.995 41.925 382.225 184.54 ;
      RECT 372.765 184.54 382.225 184.77 ;
      RECT 372.765 82.505 372.995 184.54 ;
      RECT 372.795 53.7 374.905 53.87 ;
      RECT 374.735 42.79 375.695 42.96 ;
      RECT 374.735 42.96 374.905 53.7 ;
      RECT 375.525 41.725 382.225 41.895 ;
      RECT 378.325 41.895 382.225 41.925 ;
      RECT 378.325 41.695 382.225 41.725 ;
      RECT 372.795 53.87 372.965 82.505 ;
      RECT 375.525 41.895 375.695 42.79 ;
      RECT 349.185 250.14 382.945 253.385 ;
      RECT 365.625 227.215 382.945 250.14 ;
      RECT 441.925 215.425 443.295 215.44 ;
      RECT 371.945 214.88 382.945 227.215 ;
      RECT 386.77 214.88 443.295 215.425 ;
      RECT 371.945 211.275 443.295 214.88 ;
      RECT 371.945 206.365 387.62 211.275 ;
      RECT 394.64 206.365 395.49 211.275 ;
      RECT 402.7 206.365 405.25 211.275 ;
      RECT 412.575 206.365 413.425 211.275 ;
      RECT 420.985 206.365 422.855 211.275 ;
      RECT 430.485 206.365 431.335 211.275 ;
      RECT 439.13 206.365 443.295 211.275 ;
      RECT 371.945 202.71 443.295 206.365 ;
      RECT 349.185 202.215 443.295 202.71 ;
      RECT 349.185 195.58 385.37 202.215 ;
      RECT 369.775 193.23 369.945 195.58 ;
      RECT 349.185 192.515 355.96 195.58 ;
      RECT 442.15 190.715 443.295 202.215 ;
      RECT 460.09 190.715 466.74 196.79 ;
      RECT 369.75 190.495 370 193.23 ;
      RECT 370.53 186.695 385.37 195.58 ;
      RECT 349.185 186.695 353.925 192.515 ;
      RECT 349.185 186.105 385.37 186.695 ;
      RECT 367.8 185.835 385.37 186.105 ;
      RECT 367.8 185.455 371.945 185.835 ;
      RECT 442.15 185.105 466.74 190.715 ;
      RECT 349.185 184.215 362.055 186.105 ;
      RECT 367.515 181.365 371.945 185.455 ;
      RECT 368.225 178.695 371.945 181.365 ;
      RECT 347.085 178.605 347.255 183.39 ;
      RECT 355.035 178.605 355.205 183.39 ;
      RECT 367.725 177.695 371.945 178.695 ;
      RECT 346.965 178.435 347.495 178.605 ;
      RECT 354.795 178.435 355.325 178.605 ;
      RECT 368.225 176.43 371.945 177.695 ;
      RECT 347.085 176.43 347.255 178.435 ;
      RECT 355.035 176.43 355.205 178.435 ;
      RECT 341.14 174.835 371.945 176.43 ;
      RECT 341.14 174.055 347.185 174.835 ;
      RECT 371.04 173.75 371.945 174.835 ;
      RECT 341.14 173.485 344.275 174.055 ;
      RECT 371.325 172.935 371.945 173.75 ;
      RECT 341.14 172.905 347.185 173.485 ;
      RECT 341.14 171.515 343.47 172.905 ;
      RECT 341.14 171.345 347.185 171.515 ;
      RECT 341.14 169.955 343.47 171.345 ;
      RECT 341.14 169.785 347.185 169.955 ;
      RECT 341.14 168.395 343.47 169.785 ;
      RECT 341.14 168.225 347.185 168.395 ;
      RECT 341.14 167.875 343.47 168.225 ;
      RECT 329.065 167.705 344.015 167.875 ;
      RECT 329.065 165.785 329.235 167.705 ;
      RECT 329.065 165.455 334.22 165.785 ;
      RECT 329.065 163.625 329.235 165.455 ;
      RECT 329.065 163.295 334.22 163.625 ;
      RECT 329.065 162.385 329.235 163.295 ;
      RECT 371.23 162.215 372.36 164.565 ;
      RECT 329.065 162.215 351.455 162.385 ;
      RECT 329.065 161.195 372.36 162.215 ;
      RECT 382.77 148.03 385.37 185.835 ;
      RECT 385.72 146.015 395.34 146.325 ;
      RECT 370.33 141.545 372.36 161.195 ;
      RECT 442.705 136.615 444.415 136.685 ;
    LAYER met5 ;
      RECT 0 0 480 55.05 ;
      RECT 278.015 124.875 459.455 131.875 ;
      RECT 285.015 131.875 446.62 144.71 ;
      RECT 171.99 194.875 225.015 201.875 ;
      RECT 164.99 124.875 218.015 131.875 ;
      RECT 171.99 131.875 218.015 194.875 ;
      RECT 51.79 145.105 104.99 145.595 ;
      RECT 51.79 145.595 104.99 148.75 ;
      RECT 39.28 132.55 104.99 133.085 ;
      RECT 39.28 133.085 104.99 145.105 ;
      RECT 31.07 124.875 104.99 131.875 ;
      RECT 38.07 131.875 104.99 132.55 ;
      RECT 54.945 194.875 107.38 197.27 ;
      RECT 0 149.515 28.46 159.715 ;
      RECT 54.945 197.27 111.99 201.875 ;
      RECT 54.945 148.75 104.99 194.875 ;
      RECT 0 159.715 28.46 207.655 ;
      RECT 285.015 194.875 389.455 201.875 ;
      RECT 59.55 201.875 387.64 203.69 ;
      RECT 285.015 150.95 439.89 151.44 ;
      RECT 285.015 151.44 396.455 194.875 ;
      RECT 285.015 144.71 446.09 145.24 ;
      RECT 285.015 145.24 440.38 150.95 ;
      RECT 29.145 122.95 466.455 124.875 ;
      RECT 478.815 149.5 480 228.7 ;
      RECT 0 207.655 49.505 228.7 ;
      RECT 285.015 138.275 452.655 138.675 ;
      RECT 285.015 138.675 452.255 139.075 ;
      RECT 285.015 139.075 451.855 139.475 ;
      RECT 285.015 139.475 451.455 139.875 ;
      RECT 285.015 139.875 451.055 140.275 ;
      RECT 285.015 140.275 450.655 140.675 ;
      RECT 285.015 140.675 450.255 141.075 ;
      RECT 285.015 141.075 449.855 141.475 ;
      RECT 285.015 141.475 449.455 141.875 ;
      RECT 285.015 141.875 449.055 142.275 ;
      RECT 285.015 142.275 448.655 142.675 ;
      RECT 285.015 142.675 448.255 143.075 ;
      RECT 285.015 143.075 447.855 143.475 ;
      RECT 285.015 143.475 447.455 143.875 ;
      RECT 285.015 143.875 447.055 144.275 ;
      RECT 285.015 144.275 446.655 144.675 ;
      RECT 285.015 144.675 446.62 144.71 ;
      RECT 55.345 197.27 107.38 197.67 ;
      RECT 55.745 197.67 107.785 198.07 ;
      RECT 56.145 198.07 108.185 198.47 ;
      RECT 56.545 198.47 108.585 198.87 ;
      RECT 56.945 198.87 108.985 199.27 ;
      RECT 57.345 199.27 109.385 199.67 ;
      RECT 57.745 199.67 109.785 200.07 ;
      RECT 58.145 200.07 110.185 200.47 ;
      RECT 58.545 200.47 110.585 200.87 ;
      RECT 58.945 200.87 110.985 201.27 ;
      RECT 59.345 201.27 111.385 201.67 ;
      RECT 59.55 201.67 111.785 201.875 ;
      RECT 52.19 145.595 104.99 145.995 ;
      RECT 52.59 145.995 104.99 146.395 ;
      RECT 52.99 146.395 104.99 146.795 ;
      RECT 53.39 146.795 104.99 147.195 ;
      RECT 53.79 147.195 104.99 147.595 ;
      RECT 54.19 147.595 104.99 147.995 ;
      RECT 54.59 147.995 104.99 148.395 ;
      RECT 54.945 148.395 104.99 148.75 ;
      RECT 54.945 194.875 104.99 195.275 ;
      RECT 54.945 195.275 105.39 195.675 ;
      RECT 54.945 195.675 105.79 196.075 ;
      RECT 54.945 196.075 106.19 196.475 ;
      RECT 54.945 196.475 106.59 196.875 ;
      RECT 54.945 196.875 106.99 197.27 ;
      RECT 39.68 133.085 104.99 133.485 ;
      RECT 40.08 133.485 104.99 133.885 ;
      RECT 40.48 133.885 104.99 134.285 ;
      RECT 40.88 134.285 104.99 134.685 ;
      RECT 41.28 134.685 104.99 135.085 ;
      RECT 41.68 135.085 104.99 135.485 ;
      RECT 42.08 135.485 104.99 135.885 ;
      RECT 42.48 135.885 104.99 136.285 ;
      RECT 42.88 136.285 104.99 136.685 ;
      RECT 43.28 136.685 104.99 137.085 ;
      RECT 43.68 137.085 104.99 137.485 ;
      RECT 44.08 137.485 104.99 137.885 ;
      RECT 44.48 137.885 104.99 138.285 ;
      RECT 44.88 138.285 104.99 138.685 ;
      RECT 45.28 138.685 104.99 139.085 ;
      RECT 45.68 139.085 104.99 139.485 ;
      RECT 46.08 139.485 104.99 139.885 ;
      RECT 46.48 139.885 104.99 140.285 ;
      RECT 46.88 140.285 104.99 140.685 ;
      RECT 47.28 140.685 104.99 141.085 ;
      RECT 47.68 141.085 104.99 141.485 ;
      RECT 48.08 141.485 104.99 141.885 ;
      RECT 48.48 141.885 104.99 142.285 ;
      RECT 48.88 142.285 104.99 142.685 ;
      RECT 49.28 142.685 104.99 143.085 ;
      RECT 49.68 143.085 104.99 143.485 ;
      RECT 50.08 143.485 104.99 143.885 ;
      RECT 50.48 143.885 104.99 144.285 ;
      RECT 50.88 144.285 104.99 144.685 ;
      RECT 51.28 144.685 104.99 145.085 ;
      RECT 51.3 145.085 104.99 145.105 ;
      RECT 31.47 124.875 111.59 125.275 ;
      RECT 31.87 125.275 111.19 125.675 ;
      RECT 32.27 125.675 110.79 126.075 ;
      RECT 32.67 126.075 110.39 126.475 ;
      RECT 33.07 126.475 109.99 126.875 ;
      RECT 33.47 126.875 109.59 127.275 ;
      RECT 33.87 127.275 109.19 127.675 ;
      RECT 34.27 127.675 108.79 128.075 ;
      RECT 34.67 128.075 108.39 128.475 ;
      RECT 35.07 128.475 107.99 128.875 ;
      RECT 35.47 128.875 107.59 129.275 ;
      RECT 35.87 129.275 107.19 129.675 ;
      RECT 36.27 129.675 106.79 130.075 ;
      RECT 36.67 130.075 106.39 130.475 ;
      RECT 37.07 130.475 105.99 130.875 ;
      RECT 37.47 130.875 105.59 131.275 ;
      RECT 37.87 131.275 105.19 131.675 ;
      RECT 38.07 131.675 104.99 131.875 ;
      RECT 38.405 131.875 104.99 132.21 ;
      RECT 38.745 132.21 104.99 132.55 ;
      RECT 285.015 164.64 426.29 165.04 ;
      RECT 285.015 164.24 426.69 164.64 ;
      RECT 285.015 163.84 427.09 164.24 ;
      RECT 285.015 163.44 427.49 163.84 ;
      RECT 285.015 163.04 427.89 163.44 ;
      RECT 285.015 162.64 428.29 163.04 ;
      RECT 285.015 162.24 428.69 162.64 ;
      RECT 285.015 161.84 429.09 162.24 ;
      RECT 285.015 161.44 429.49 161.84 ;
      RECT 285.015 161.04 429.89 161.44 ;
      RECT 285.015 160.64 430.29 161.04 ;
      RECT 285.015 160.24 430.69 160.64 ;
      RECT 285.015 159.84 431.09 160.24 ;
      RECT 285.015 159.44 431.49 159.84 ;
      RECT 285.015 159.04 431.89 159.44 ;
      RECT 285.015 158.64 432.29 159.04 ;
      RECT 285.015 158.24 432.69 158.64 ;
      RECT 285.015 157.84 433.09 158.24 ;
      RECT 285.015 157.44 433.49 157.84 ;
      RECT 285.015 157.04 433.89 157.44 ;
      RECT 285.015 156.64 434.29 157.04 ;
      RECT 285.015 156.24 434.69 156.64 ;
      RECT 285.015 155.84 435.09 156.24 ;
      RECT 285.015 155.44 435.49 155.84 ;
      RECT 285.015 155.04 435.89 155.44 ;
      RECT 285.015 154.64 436.29 155.04 ;
      RECT 285.015 154.24 436.69 154.64 ;
      RECT 285.015 153.84 437.09 154.24 ;
      RECT 285.015 153.44 437.49 153.84 ;
      RECT 285.015 153.04 437.89 153.44 ;
      RECT 285.015 152.64 438.29 153.04 ;
      RECT 285.015 152.24 438.69 152.64 ;
      RECT 285.015 151.84 439.09 152.24 ;
      RECT 285.015 151.44 439.49 151.84 ;
      RECT 171.99 194.875 218.015 195.275 ;
      RECT 171.59 195.275 218.415 195.675 ;
      RECT 171.19 195.675 218.815 196.075 ;
      RECT 170.79 196.075 219.215 196.475 ;
      RECT 170.39 196.475 219.615 196.875 ;
      RECT 169.99 196.875 220.015 197.275 ;
      RECT 169.59 197.275 220.415 197.675 ;
      RECT 169.19 197.675 220.815 198.075 ;
      RECT 168.79 198.075 221.215 198.475 ;
      RECT 168.39 198.475 221.615 198.875 ;
      RECT 167.99 198.875 222.015 199.275 ;
      RECT 167.59 199.275 222.415 199.675 ;
      RECT 167.19 199.675 222.815 200.075 ;
      RECT 166.79 200.075 223.215 200.475 ;
      RECT 166.39 200.475 223.615 200.875 ;
      RECT 165.99 200.875 224.015 201.275 ;
      RECT 165.59 201.275 224.415 201.675 ;
      RECT 165.19 201.675 224.815 201.875 ;
      RECT 285.015 194.875 396.055 195.275 ;
      RECT 284.615 195.275 395.655 195.675 ;
      RECT 284.215 195.675 395.255 196.075 ;
      RECT 283.815 196.075 394.855 196.475 ;
      RECT 283.415 196.475 394.455 196.875 ;
      RECT 283.015 196.875 394.055 197.275 ;
      RECT 282.615 197.275 393.655 197.675 ;
      RECT 282.215 197.675 393.255 198.075 ;
      RECT 281.815 198.075 392.855 198.475 ;
      RECT 281.415 198.475 392.455 198.875 ;
      RECT 281.015 198.875 392.055 199.275 ;
      RECT 280.615 199.275 391.655 199.675 ;
      RECT 280.215 199.675 391.255 200.075 ;
      RECT 279.815 200.075 390.855 200.475 ;
      RECT 279.415 200.475 390.455 200.875 ;
      RECT 279.015 200.875 390.055 201.275 ;
      RECT 278.615 201.275 389.655 201.675 ;
      RECT 278.215 201.675 389.455 201.875 ;
      RECT 165.39 124.875 224.615 125.275 ;
      RECT 165.79 125.275 224.215 125.675 ;
      RECT 166.19 125.675 223.815 126.075 ;
      RECT 166.59 126.075 223.415 126.475 ;
      RECT 166.99 126.475 223.015 126.875 ;
      RECT 167.39 126.875 222.615 127.275 ;
      RECT 167.79 127.275 222.215 127.675 ;
      RECT 168.19 127.675 221.815 128.075 ;
      RECT 168.59 128.075 221.415 128.475 ;
      RECT 168.99 128.475 221.015 128.875 ;
      RECT 169.39 128.875 220.615 129.275 ;
      RECT 169.79 129.275 220.215 129.675 ;
      RECT 170.19 129.675 219.815 130.075 ;
      RECT 170.59 130.075 219.415 130.475 ;
      RECT 170.99 130.475 219.015 130.875 ;
      RECT 171.39 130.875 218.615 131.275 ;
      RECT 171.79 131.275 218.215 131.675 ;
      RECT 171.99 131.675 218.015 131.875 ;
      RECT 278.415 124.875 466.055 125.275 ;
      RECT 278.815 125.275 465.655 125.675 ;
      RECT 279.215 125.675 465.255 126.075 ;
      RECT 279.615 126.075 464.855 126.475 ;
      RECT 280.015 126.475 464.455 126.875 ;
      RECT 280.415 126.875 464.055 127.275 ;
      RECT 280.815 127.275 463.655 127.675 ;
      RECT 281.215 127.675 463.255 128.075 ;
      RECT 281.615 128.075 462.855 128.475 ;
      RECT 282.015 128.475 462.455 128.875 ;
      RECT 282.415 128.875 462.055 129.275 ;
      RECT 282.815 129.275 461.655 129.675 ;
      RECT 283.215 129.675 461.255 130.075 ;
      RECT 283.615 130.075 460.855 130.475 ;
      RECT 284.015 130.475 460.455 130.875 ;
      RECT 284.415 130.875 460.055 131.275 ;
      RECT 284.815 131.275 459.655 131.675 ;
      RECT 285.015 131.675 459.455 131.875 ;
      RECT 29.545 122.95 467.98 123.35 ;
      RECT 29.945 123.35 467.58 123.75 ;
      RECT 30.345 123.75 467.18 124.15 ;
      RECT 30.745 124.15 466.78 124.55 ;
      RECT 31.07 124.55 466.455 124.875 ;
      RECT 285.015 131.875 459.055 132.275 ;
      RECT 285.015 132.275 458.655 132.675 ;
      RECT 285.015 132.675 458.255 133.075 ;
      RECT 285.015 133.075 457.855 133.475 ;
      RECT 285.015 133.475 457.455 133.875 ;
      RECT 285.015 133.875 457.055 134.275 ;
      RECT 285.015 134.275 456.655 134.675 ;
      RECT 285.015 134.675 456.255 135.075 ;
      RECT 285.015 135.075 455.855 135.475 ;
      RECT 285.015 135.475 455.455 135.875 ;
      RECT 285.015 135.875 455.055 136.275 ;
      RECT 285.015 136.275 454.655 136.675 ;
      RECT 285.015 136.675 454.255 137.075 ;
      RECT 285.015 137.075 453.855 137.475 ;
      RECT 285.015 137.475 453.455 137.875 ;
      RECT 285.015 137.875 453.055 138.275 ;
      RECT 0 226.855 47.66 227.255 ;
      RECT 0 227.255 48.06 227.655 ;
      RECT 0 227.655 48.46 228.055 ;
      RECT 0 228.055 48.86 228.455 ;
      RECT 0 228.455 49.26 228.7 ;
      RECT 0 149.515 18.26 149.915 ;
      RECT 0 149.915 18.66 150.315 ;
      RECT 0 150.315 19.06 150.715 ;
      RECT 0 150.715 19.46 151.115 ;
      RECT 0 151.115 19.86 151.515 ;
      RECT 0 151.515 20.26 151.915 ;
      RECT 0 151.915 20.66 152.315 ;
      RECT 0 152.315 21.06 152.715 ;
      RECT 0 152.715 21.46 153.115 ;
      RECT 0 153.115 21.86 153.515 ;
      RECT 0 153.515 22.26 153.915 ;
      RECT 0 153.915 22.66 154.315 ;
      RECT 0 154.315 23.06 154.715 ;
      RECT 0 154.715 23.46 155.115 ;
      RECT 0 155.115 23.86 155.515 ;
      RECT 0 155.515 24.26 155.915 ;
      RECT 0 155.915 24.66 156.315 ;
      RECT 0 156.315 25.06 156.715 ;
      RECT 0 156.715 25.46 157.115 ;
      RECT 0 157.115 25.86 157.515 ;
      RECT 0 157.515 26.26 157.915 ;
      RECT 0 157.915 26.66 158.315 ;
      RECT 0 158.315 27.06 158.715 ;
      RECT 0 158.715 27.46 159.115 ;
      RECT 0 159.115 27.86 159.515 ;
      RECT 0 159.515 28.26 159.715 ;
      RECT 59.95 201.875 389.055 202.275 ;
      RECT 60.35 202.275 388.655 202.675 ;
      RECT 60.75 202.675 388.255 203.075 ;
      RECT 61.15 203.075 387.855 203.475 ;
      RECT 61.365 203.475 387.64 203.69 ;
      RECT 285.015 145.24 445.69 145.64 ;
      RECT 285.015 145.64 445.29 146.04 ;
      RECT 285.015 146.04 444.89 146.44 ;
      RECT 285.015 146.44 444.49 146.84 ;
      RECT 285.015 146.84 444.09 147.24 ;
      RECT 285.015 147.24 443.69 147.64 ;
      RECT 285.015 147.64 443.29 148.04 ;
      RECT 285.015 148.04 442.89 148.44 ;
      RECT 285.015 148.44 442.49 148.84 ;
      RECT 285.015 148.84 442.09 149.24 ;
      RECT 285.015 149.24 441.69 149.64 ;
      RECT 285.015 149.64 441.29 150.04 ;
      RECT 285.015 150.04 440.89 150.44 ;
      RECT 285.015 150.44 440.49 150.84 ;
      RECT 285.015 150.84 440.38 150.95 ;
      RECT 285.015 194.64 396.455 194.875 ;
      RECT 285.015 194.24 396.69 194.64 ;
      RECT 285.015 193.84 397.09 194.24 ;
      RECT 285.015 193.44 397.49 193.84 ;
      RECT 285.015 193.04 397.89 193.44 ;
      RECT 285.015 192.64 398.29 193.04 ;
      RECT 285.015 192.24 398.69 192.64 ;
      RECT 285.015 191.84 399.09 192.24 ;
      RECT 285.015 191.44 399.49 191.84 ;
      RECT 285.015 191.04 399.89 191.44 ;
      RECT 285.015 190.64 400.29 191.04 ;
      RECT 285.015 190.24 400.69 190.64 ;
      RECT 285.015 189.84 401.09 190.24 ;
      RECT 285.015 189.44 401.49 189.84 ;
      RECT 285.015 189.04 401.89 189.44 ;
      RECT 285.015 188.64 402.29 189.04 ;
      RECT 285.015 188.24 402.69 188.64 ;
      RECT 285.015 187.84 403.09 188.24 ;
      RECT 285.015 187.44 403.49 187.84 ;
      RECT 285.015 187.04 403.89 187.44 ;
      RECT 285.015 186.64 404.29 187.04 ;
      RECT 285.015 186.24 404.69 186.64 ;
      RECT 285.015 185.84 405.09 186.24 ;
      RECT 285.015 185.44 405.49 185.84 ;
      RECT 285.015 185.04 405.89 185.44 ;
      RECT 285.015 184.64 406.29 185.04 ;
      RECT 285.015 184.24 406.69 184.64 ;
      RECT 285.015 183.84 407.09 184.24 ;
      RECT 285.015 183.44 407.49 183.84 ;
      RECT 285.015 183.04 407.89 183.44 ;
      RECT 285.015 182.64 408.29 183.04 ;
      RECT 285.015 182.24 408.69 182.64 ;
      RECT 285.015 181.84 409.09 182.24 ;
      RECT 285.015 181.44 409.49 181.84 ;
      RECT 285.015 181.04 409.89 181.44 ;
      RECT 285.015 180.64 410.29 181.04 ;
      RECT 285.015 180.24 410.69 180.64 ;
      RECT 285.015 179.84 411.09 180.24 ;
      RECT 285.015 179.44 411.49 179.84 ;
      RECT 285.015 179.04 411.89 179.44 ;
      RECT 285.015 178.64 412.29 179.04 ;
      RECT 285.015 178.24 412.69 178.64 ;
      RECT 285.015 177.84 413.09 178.24 ;
      RECT 285.015 177.44 413.49 177.84 ;
      RECT 285.015 177.04 413.89 177.44 ;
      RECT 285.015 176.64 414.29 177.04 ;
      RECT 285.015 176.24 414.69 176.64 ;
      RECT 285.015 175.84 415.09 176.24 ;
      RECT 285.015 175.44 415.49 175.84 ;
      RECT 285.015 175.04 415.89 175.44 ;
      RECT 285.015 174.64 416.29 175.04 ;
      RECT 285.015 174.24 416.69 174.64 ;
      RECT 285.015 173.84 417.09 174.24 ;
      RECT 285.015 173.44 417.49 173.84 ;
      RECT 285.015 173.04 417.89 173.44 ;
      RECT 285.015 172.64 418.29 173.04 ;
      RECT 285.015 172.24 418.69 172.64 ;
      RECT 285.015 171.84 419.09 172.24 ;
      RECT 285.015 171.44 419.49 171.84 ;
      RECT 285.015 171.04 419.89 171.44 ;
      RECT 285.015 170.64 420.29 171.04 ;
      RECT 285.015 170.24 420.69 170.64 ;
      RECT 285.015 169.84 421.09 170.24 ;
      RECT 285.015 169.44 421.49 169.84 ;
      RECT 285.015 169.04 421.89 169.44 ;
      RECT 285.015 168.64 422.29 169.04 ;
      RECT 285.015 168.24 422.69 168.64 ;
      RECT 285.015 167.84 423.09 168.24 ;
      RECT 285.015 167.44 423.49 167.84 ;
      RECT 285.015 167.04 423.89 167.44 ;
      RECT 285.015 166.64 424.29 167.04 ;
      RECT 285.015 166.24 424.69 166.64 ;
      RECT 285.015 165.84 425.09 166.24 ;
      RECT 285.015 165.44 425.49 165.84 ;
      RECT 285.015 165.04 425.89 165.44 ;
      RECT 447.615 180.7 480 181.1 ;
      RECT 448.015 180.3 480 180.7 ;
      RECT 448.415 179.9 480 180.3 ;
      RECT 448.815 179.5 480 179.9 ;
      RECT 449.215 179.1 480 179.5 ;
      RECT 449.615 178.7 480 179.1 ;
      RECT 450.015 178.3 480 178.7 ;
      RECT 450.415 177.9 480 178.3 ;
      RECT 450.815 177.5 480 177.9 ;
      RECT 451.215 177.1 480 177.5 ;
      RECT 451.615 176.7 480 177.1 ;
      RECT 452.015 176.3 480 176.7 ;
      RECT 452.415 175.9 480 176.3 ;
      RECT 452.815 175.5 480 175.9 ;
      RECT 453.215 175.1 480 175.5 ;
      RECT 453.615 174.7 480 175.1 ;
      RECT 454.015 174.3 480 174.7 ;
      RECT 454.415 173.9 480 174.3 ;
      RECT 454.815 173.5 480 173.9 ;
      RECT 455.215 173.1 480 173.5 ;
      RECT 455.615 172.7 480 173.1 ;
      RECT 456.015 172.3 480 172.7 ;
      RECT 456.415 171.9 480 172.3 ;
      RECT 456.815 171.5 480 171.9 ;
      RECT 457.215 171.1 480 171.5 ;
      RECT 457.615 170.7 480 171.1 ;
      RECT 458.015 170.3 480 170.7 ;
      RECT 458.415 169.9 480 170.3 ;
      RECT 458.815 169.5 480 169.9 ;
      RECT 459.215 169.1 480 169.5 ;
      RECT 459.615 168.7 480 169.1 ;
      RECT 460.015 168.3 480 168.7 ;
      RECT 460.415 167.9 480 168.3 ;
      RECT 460.815 167.5 480 167.9 ;
      RECT 461.215 167.1 480 167.5 ;
      RECT 461.615 166.7 480 167.1 ;
      RECT 462.015 166.3 480 166.7 ;
      RECT 462.415 165.9 480 166.3 ;
      RECT 462.815 165.5 480 165.9 ;
      RECT 463.215 165.1 480 165.5 ;
      RECT 463.615 164.7 480 165.1 ;
      RECT 464.015 164.3 480 164.7 ;
      RECT 464.415 163.9 480 164.3 ;
      RECT 464.815 163.5 480 163.9 ;
      RECT 465.215 163.1 480 163.5 ;
      RECT 465.615 162.7 480 163.1 ;
      RECT 466.015 162.3 480 162.7 ;
      RECT 466.415 161.9 480 162.3 ;
      RECT 466.815 161.5 480 161.9 ;
      RECT 467.215 161.1 480 161.5 ;
      RECT 467.615 160.7 480 161.1 ;
      RECT 468.015 160.3 480 160.7 ;
      RECT 468.415 159.9 480 160.3 ;
      RECT 468.815 159.5 480 159.9 ;
      RECT 469.215 159.1 480 159.5 ;
      RECT 469.615 158.7 480 159.1 ;
      RECT 470.015 158.3 480 158.7 ;
      RECT 470.415 157.9 480 158.3 ;
      RECT 470.815 157.5 480 157.9 ;
      RECT 471.215 157.1 480 157.5 ;
      RECT 471.615 156.7 480 157.1 ;
      RECT 472.015 156.3 480 156.7 ;
      RECT 472.415 155.9 480 156.3 ;
      RECT 472.815 155.5 480 155.9 ;
      RECT 473.215 155.1 480 155.5 ;
      RECT 473.615 154.7 480 155.1 ;
      RECT 474.015 154.3 480 154.7 ;
      RECT 474.415 153.9 480 154.3 ;
      RECT 474.815 153.5 480 153.9 ;
      RECT 475.215 153.1 480 153.5 ;
      RECT 475.615 152.7 480 153.1 ;
      RECT 476.015 152.3 480 152.7 ;
      RECT 476.415 151.9 480 152.3 ;
      RECT 476.815 151.5 480 151.9 ;
      RECT 477.215 151.1 480 151.5 ;
      RECT 477.615 150.7 480 151.1 ;
      RECT 478.015 150.3 480 150.7 ;
      RECT 478.415 149.9 480 150.3 ;
      RECT 478.815 149.5 480 149.9 ;
      RECT 0 207.655 28.46 208.055 ;
      RECT 0 208.055 28.86 208.455 ;
      RECT 0 208.455 29.26 208.855 ;
      RECT 0 208.855 29.66 209.255 ;
      RECT 0 209.255 30.06 209.655 ;
      RECT 0 209.655 30.46 210.055 ;
      RECT 0 210.055 30.86 210.455 ;
      RECT 0 210.455 31.26 210.855 ;
      RECT 0 210.855 31.66 211.255 ;
      RECT 0 211.255 32.06 211.655 ;
      RECT 0 211.655 32.46 212.055 ;
      RECT 0 212.055 32.86 212.455 ;
      RECT 0 212.455 33.26 212.855 ;
      RECT 0 212.855 33.66 213.255 ;
      RECT 0 213.255 34.06 213.655 ;
      RECT 0 213.655 34.46 214.055 ;
      RECT 0 214.055 34.86 214.455 ;
      RECT 0 214.455 35.26 214.855 ;
      RECT 0 214.855 35.66 215.255 ;
      RECT 0 215.255 36.06 215.655 ;
      RECT 0 215.655 36.46 216.055 ;
      RECT 0 216.055 36.86 216.455 ;
      RECT 0 216.455 37.26 216.855 ;
      RECT 0 216.855 37.66 217.255 ;
      RECT 0 217.255 38.06 217.655 ;
      RECT 0 217.655 38.46 218.055 ;
      RECT 0 218.055 38.86 218.455 ;
      RECT 0 218.455 39.26 218.855 ;
      RECT 0 218.855 39.66 219.255 ;
      RECT 0 219.255 40.06 219.655 ;
      RECT 0 219.655 40.46 220.055 ;
      RECT 0 220.055 40.86 220.455 ;
      RECT 0 220.455 41.26 220.855 ;
      RECT 0 220.855 41.66 221.255 ;
      RECT 0 221.255 42.06 221.655 ;
      RECT 0 221.655 42.46 222.055 ;
      RECT 0 222.055 42.86 222.455 ;
      RECT 0 222.455 43.26 222.855 ;
      RECT 0 222.855 43.66 223.255 ;
      RECT 0 223.255 44.06 223.655 ;
      RECT 0 223.655 44.46 224.055 ;
      RECT 0 224.055 44.86 224.455 ;
      RECT 0 224.455 45.26 224.855 ;
      RECT 0 224.855 45.66 225.255 ;
      RECT 0 225.255 46.06 225.655 ;
      RECT 0 225.655 46.46 226.055 ;
      RECT 0 226.055 46.86 226.455 ;
      RECT 0 226.455 47.26 226.855 ;
      RECT 0 159.715 28.46 207.655 ;
      RECT 285.015 150.95 439.89 151.44 ;
      RECT 285.015 144.71 446.09 145.24 ;
      RECT 171.99 131.875 218.015 194.875 ;
      RECT 39.28 132.55 104.99 133.085 ;
      RECT 51.79 145.105 104.99 145.595 ;
      RECT 54.945 148.75 104.99 194.875 ;
      RECT 0 0 480 55.05 ;
      RECT 400.015 228.3 480 228.7 ;
      RECT 400.415 227.9 480 228.3 ;
      RECT 400.815 227.5 480 227.9 ;
      RECT 401.215 227.1 480 227.5 ;
      RECT 401.615 226.7 480 227.1 ;
      RECT 402.015 226.3 480 226.7 ;
      RECT 402.415 225.9 480 226.3 ;
      RECT 402.815 225.5 480 225.9 ;
      RECT 403.215 225.1 480 225.5 ;
      RECT 403.615 224.7 480 225.1 ;
      RECT 404.015 224.3 480 224.7 ;
      RECT 404.415 223.9 480 224.3 ;
      RECT 404.815 223.5 480 223.9 ;
      RECT 405.215 223.1 480 223.5 ;
      RECT 405.615 222.7 480 223.1 ;
      RECT 406.015 222.3 480 222.7 ;
      RECT 406.415 221.9 480 222.3 ;
      RECT 406.815 221.5 480 221.9 ;
      RECT 407.215 221.1 480 221.5 ;
      RECT 407.615 220.7 480 221.1 ;
      RECT 408.015 220.3 480 220.7 ;
      RECT 408.415 219.9 480 220.3 ;
      RECT 408.815 219.5 480 219.9 ;
      RECT 409.215 219.1 480 219.5 ;
      RECT 409.615 218.7 480 219.1 ;
      RECT 410.015 218.3 480 218.7 ;
      RECT 410.415 217.9 480 218.3 ;
      RECT 410.815 217.5 480 217.9 ;
      RECT 411.215 217.1 480 217.5 ;
      RECT 411.615 216.7 480 217.1 ;
      RECT 412.015 216.3 480 216.7 ;
      RECT 412.415 215.9 480 216.3 ;
      RECT 412.815 215.5 480 215.9 ;
      RECT 413.215 215.1 480 215.5 ;
      RECT 413.615 214.7 480 215.1 ;
      RECT 414.015 214.3 480 214.7 ;
      RECT 414.415 213.9 480 214.3 ;
      RECT 414.815 213.5 480 213.9 ;
      RECT 415.215 213.1 480 213.5 ;
      RECT 415.615 212.7 480 213.1 ;
      RECT 416.015 212.3 480 212.7 ;
      RECT 416.415 211.9 480 212.3 ;
      RECT 416.815 211.5 480 211.9 ;
      RECT 417.215 211.1 480 211.5 ;
      RECT 417.615 210.7 480 211.1 ;
      RECT 418.015 210.3 480 210.7 ;
      RECT 418.415 209.9 480 210.3 ;
      RECT 418.815 209.5 480 209.9 ;
      RECT 419.215 209.1 480 209.5 ;
      RECT 419.615 208.7 480 209.1 ;
      RECT 420.015 208.3 480 208.7 ;
      RECT 420.415 207.9 480 208.3 ;
      RECT 420.815 207.5 480 207.9 ;
      RECT 421.215 207.1 480 207.5 ;
      RECT 421.615 206.7 480 207.1 ;
      RECT 422.015 206.3 480 206.7 ;
      RECT 422.415 205.9 480 206.3 ;
      RECT 422.815 205.5 480 205.9 ;
      RECT 423.215 205.1 480 205.5 ;
      RECT 423.615 204.7 480 205.1 ;
      RECT 424.015 204.3 480 204.7 ;
      RECT 424.415 203.9 480 204.3 ;
      RECT 424.815 203.5 480 203.9 ;
      RECT 425.215 203.1 480 203.5 ;
      RECT 425.615 202.7 480 203.1 ;
      RECT 426.015 202.3 480 202.7 ;
      RECT 426.415 201.9 480 202.3 ;
      RECT 426.815 201.5 480 201.9 ;
      RECT 427.215 201.1 480 201.5 ;
      RECT 427.615 200.7 480 201.1 ;
      RECT 428.015 200.3 480 200.7 ;
      RECT 428.415 199.9 480 200.3 ;
      RECT 428.815 199.5 480 199.9 ;
      RECT 429.215 199.1 480 199.5 ;
      RECT 429.615 198.7 480 199.1 ;
      RECT 430.015 198.3 480 198.7 ;
      RECT 430.415 197.9 480 198.3 ;
      RECT 430.815 197.5 480 197.9 ;
      RECT 431.215 197.1 480 197.5 ;
      RECT 431.615 196.7 480 197.1 ;
      RECT 432.015 196.3 480 196.7 ;
      RECT 432.415 195.9 480 196.3 ;
      RECT 432.815 195.5 480 195.9 ;
      RECT 433.215 195.1 480 195.5 ;
      RECT 433.615 194.7 480 195.1 ;
      RECT 434.015 194.3 480 194.7 ;
      RECT 434.415 193.9 480 194.3 ;
      RECT 434.815 193.5 480 193.9 ;
      RECT 435.215 193.1 480 193.5 ;
      RECT 435.615 192.7 480 193.1 ;
      RECT 436.015 192.3 480 192.7 ;
      RECT 436.415 191.9 480 192.3 ;
      RECT 436.815 191.5 480 191.9 ;
      RECT 437.215 191.1 480 191.5 ;
      RECT 437.615 190.7 480 191.1 ;
      RECT 438.015 190.3 480 190.7 ;
      RECT 438.415 189.9 480 190.3 ;
      RECT 438.815 189.5 480 189.9 ;
      RECT 439.215 189.1 480 189.5 ;
      RECT 439.615 188.7 480 189.1 ;
      RECT 440.015 188.3 480 188.7 ;
      RECT 440.415 187.9 480 188.3 ;
      RECT 440.815 187.5 480 187.9 ;
      RECT 441.215 187.1 480 187.5 ;
      RECT 441.615 186.7 480 187.1 ;
      RECT 442.015 186.3 480 186.7 ;
      RECT 442.415 185.9 480 186.3 ;
      RECT 442.815 185.5 480 185.9 ;
      RECT 443.215 185.1 480 185.5 ;
      RECT 443.615 184.7 480 185.1 ;
      RECT 444.015 184.3 480 184.7 ;
      RECT 444.415 183.9 480 184.3 ;
      RECT 444.815 183.5 480 183.9 ;
      RECT 445.215 183.1 480 183.5 ;
      RECT 445.615 182.7 480 183.1 ;
      RECT 446.015 182.3 480 182.7 ;
      RECT 446.415 181.9 480 182.3 ;
      RECT 446.815 181.5 480 181.9 ;
      RECT 447.215 181.1 480 181.5 ;
    LAYER met4 ;
      RECT 0 116.8 480 117.4 ;
      RECT 0 110.75 480 111.55 ;
      RECT 0 84.6 480 85.2 ;
      RECT 0 94.3 480 94.9 ;
      RECT 0 89.45 480 90.05 ;
      RECT 0 0 480 55.35 ;
      RECT 0 67.65 480 68.25 ;
      RECT 0 61.6 480 62.2 ;
      RECT 0 100.35 480 101.15 ;
      RECT 0 78.45 480 79.15 ;
      RECT 458.05 73.115 480 73.2 ;
      RECT 0 72.5 480 73.115 ;
      RECT 0 228.2 480 229.1 ;
      RECT 29.23 123.55 468.31 123.74 ;
      RECT 28.94 123.45 468.5 123.55 ;
      RECT 0 122.65 480 123.45 ;
      RECT 478.595 149.015 480 228.2 ;
      RECT 29.23 123.74 443.095 148.955 ;
      RECT 54.445 148.955 394.575 197.475 ;
      RECT 0 73.115 9.455 73.2 ;
      RECT 0 207.45 49.71 228.2 ;
      RECT 0 149.015 28.96 159.51 ;
      RECT 0 159.51 28.96 207.45 ;
      RECT 54.445 197.475 387.845 204.205 ;
      RECT 0 154.965 24.275 155.115 ;
      RECT 0 154.815 24.125 154.965 ;
      RECT 0 154.665 23.975 154.815 ;
      RECT 0 154.515 23.825 154.665 ;
      RECT 0 154.365 23.675 154.515 ;
      RECT 0 154.215 23.525 154.365 ;
      RECT 0 154.065 23.375 154.215 ;
      RECT 0 153.915 23.225 154.065 ;
      RECT 0 153.765 23.075 153.915 ;
      RECT 0 153.615 22.925 153.765 ;
      RECT 0 153.465 22.775 153.615 ;
      RECT 0 153.315 22.625 153.465 ;
      RECT 0 153.165 22.475 153.315 ;
      RECT 0 153.015 22.325 153.165 ;
      RECT 0 152.865 22.175 153.015 ;
      RECT 0 152.715 22.025 152.865 ;
      RECT 0 152.565 21.875 152.715 ;
      RECT 0 152.415 21.725 152.565 ;
      RECT 0 152.265 21.575 152.415 ;
      RECT 0 152.115 21.425 152.265 ;
      RECT 0 151.965 21.275 152.115 ;
      RECT 0 151.815 21.125 151.965 ;
      RECT 0 151.665 20.975 151.815 ;
      RECT 0 151.515 20.825 151.665 ;
      RECT 0 151.365 20.675 151.515 ;
      RECT 0 151.215 20.525 151.365 ;
      RECT 0 151.065 20.375 151.215 ;
      RECT 0 150.915 20.225 151.065 ;
      RECT 0 150.765 20.075 150.915 ;
      RECT 0 150.615 19.925 150.765 ;
      RECT 0 150.465 19.775 150.615 ;
      RECT 0 150.315 19.625 150.465 ;
      RECT 0 150.165 19.475 150.315 ;
      RECT 0 150.015 19.325 150.165 ;
      RECT 0 149.865 19.175 150.015 ;
      RECT 0 149.715 19.025 149.865 ;
      RECT 0 149.565 18.875 149.715 ;
      RECT 0 149.415 18.725 149.565 ;
      RECT 0 149.265 18.575 149.415 ;
      RECT 0 149.115 18.425 149.265 ;
      RECT 0 221.74 43.11 221.89 ;
      RECT 0 221.59 42.96 221.74 ;
      RECT 0 221.44 42.81 221.59 ;
      RECT 0 221.29 42.66 221.44 ;
      RECT 0 221.14 42.51 221.29 ;
      RECT 0 220.99 42.36 221.14 ;
      RECT 0 220.84 42.21 220.99 ;
      RECT 0 220.69 42.06 220.84 ;
      RECT 0 220.54 41.91 220.69 ;
      RECT 0 220.39 41.76 220.54 ;
      RECT 0 220.24 41.61 220.39 ;
      RECT 0 220.09 41.46 220.24 ;
      RECT 0 219.94 41.31 220.09 ;
      RECT 0 219.79 41.16 219.94 ;
      RECT 0 219.64 41.01 219.79 ;
      RECT 0 219.49 40.86 219.64 ;
      RECT 0 219.34 40.71 219.49 ;
      RECT 0 219.19 40.56 219.34 ;
      RECT 0 219.04 40.41 219.19 ;
      RECT 0 218.89 40.26 219.04 ;
      RECT 0 218.74 40.11 218.89 ;
      RECT 0 218.59 39.96 218.74 ;
      RECT 0 218.44 39.81 218.59 ;
      RECT 0 218.29 39.66 218.44 ;
      RECT 0 218.14 39.51 218.29 ;
      RECT 0 217.99 39.36 218.14 ;
      RECT 0 217.84 39.21 217.99 ;
      RECT 0 217.69 39.06 217.84 ;
      RECT 0 217.54 38.91 217.69 ;
      RECT 0 217.39 38.76 217.54 ;
      RECT 0 217.24 38.61 217.39 ;
      RECT 0 217.09 38.46 217.24 ;
      RECT 0 216.94 38.31 217.09 ;
      RECT 0 216.79 38.16 216.94 ;
      RECT 0 216.64 38.01 216.79 ;
      RECT 0 216.49 37.86 216.64 ;
      RECT 0 216.34 37.71 216.49 ;
      RECT 0 216.19 37.56 216.34 ;
      RECT 0 216.04 37.41 216.19 ;
      RECT 0 215.89 37.26 216.04 ;
      RECT 0 215.74 37.11 215.89 ;
      RECT 0 215.59 36.96 215.74 ;
      RECT 0 215.44 36.81 215.59 ;
      RECT 0 215.29 36.66 215.44 ;
      RECT 0 215.14 36.51 215.29 ;
      RECT 0 214.99 36.36 215.14 ;
      RECT 0 214.84 36.21 214.99 ;
      RECT 0 214.69 36.06 214.84 ;
      RECT 0 214.54 35.91 214.69 ;
      RECT 0 214.39 35.76 214.54 ;
      RECT 0 214.24 35.61 214.39 ;
      RECT 0 214.09 35.46 214.24 ;
      RECT 0 213.94 35.31 214.09 ;
      RECT 0 213.79 35.16 213.94 ;
      RECT 0 213.64 35.01 213.79 ;
      RECT 0 213.49 34.86 213.64 ;
      RECT 0 213.34 34.71 213.49 ;
      RECT 0 213.19 34.56 213.34 ;
      RECT 0 213.04 34.41 213.19 ;
      RECT 0 212.89 34.26 213.04 ;
      RECT 0 212.74 34.11 212.89 ;
      RECT 0 212.59 33.96 212.74 ;
      RECT 0 212.44 33.81 212.59 ;
      RECT 0 212.29 33.66 212.44 ;
      RECT 0 212.14 33.51 212.29 ;
      RECT 0 211.99 33.36 212.14 ;
      RECT 0 211.84 33.21 211.99 ;
      RECT 0 211.69 33.06 211.84 ;
      RECT 0 211.54 32.91 211.69 ;
      RECT 0 211.39 32.76 211.54 ;
      RECT 0 211.24 32.61 211.39 ;
      RECT 0 211.09 32.46 211.24 ;
      RECT 0 210.94 32.31 211.09 ;
      RECT 0 210.79 32.16 210.94 ;
      RECT 0 210.64 32.01 210.79 ;
      RECT 0 210.49 31.86 210.64 ;
      RECT 0 210.34 31.71 210.49 ;
      RECT 0 210.19 31.56 210.34 ;
      RECT 0 210.04 31.41 210.19 ;
      RECT 0 209.89 31.26 210.04 ;
      RECT 0 209.74 31.11 209.89 ;
      RECT 0 209.59 30.96 209.74 ;
      RECT 0 209.44 30.81 209.59 ;
      RECT 0 209.29 30.66 209.44 ;
      RECT 0 209.14 30.51 209.29 ;
      RECT 0 208.99 30.36 209.14 ;
      RECT 0 208.84 30.21 208.99 ;
      RECT 0 208.69 30.06 208.84 ;
      RECT 0 208.54 29.91 208.69 ;
      RECT 0 208.39 29.76 208.54 ;
      RECT 0 208.24 29.61 208.39 ;
      RECT 0 208.09 29.46 208.24 ;
      RECT 0 207.94 29.31 208.09 ;
      RECT 0 207.79 29.16 207.94 ;
      RECT 0 207.64 29.01 207.79 ;
      RECT 0 207.49 28.86 207.64 ;
      RECT 0 159.465 28.775 159.55 ;
      RECT 0 159.315 28.625 159.465 ;
      RECT 0 159.165 28.475 159.315 ;
      RECT 0 159.015 28.325 159.165 ;
      RECT 0 158.865 28.175 159.015 ;
      RECT 0 158.715 28.025 158.865 ;
      RECT 0 158.565 27.875 158.715 ;
      RECT 0 158.415 27.725 158.565 ;
      RECT 0 158.265 27.575 158.415 ;
      RECT 0 158.115 27.425 158.265 ;
      RECT 0 157.965 27.275 158.115 ;
      RECT 0 157.815 27.125 157.965 ;
      RECT 0 157.665 26.975 157.815 ;
      RECT 0 157.515 26.825 157.665 ;
      RECT 0 157.365 26.675 157.515 ;
      RECT 0 157.215 26.525 157.365 ;
      RECT 0 157.065 26.375 157.215 ;
      RECT 0 156.915 26.225 157.065 ;
      RECT 0 156.765 26.075 156.915 ;
      RECT 0 156.615 25.925 156.765 ;
      RECT 0 156.465 25.775 156.615 ;
      RECT 0 156.315 25.625 156.465 ;
      RECT 0 156.165 25.475 156.315 ;
      RECT 0 156.015 25.325 156.165 ;
      RECT 0 155.865 25.175 156.015 ;
      RECT 0 155.715 25.025 155.865 ;
      RECT 0 155.565 24.875 155.715 ;
      RECT 0 155.415 24.725 155.565 ;
      RECT 0 155.265 24.575 155.415 ;
      RECT 0 155.115 24.425 155.265 ;
      RECT 468.45 159.3 480 159.45 ;
      RECT 468.6 159.15 480 159.3 ;
      RECT 468.75 159 480 159.15 ;
      RECT 468.9 158.85 480 159 ;
      RECT 469.05 158.7 480 158.85 ;
      RECT 469.2 158.55 480 158.7 ;
      RECT 469.35 158.4 480 158.55 ;
      RECT 469.5 158.25 480 158.4 ;
      RECT 469.65 158.1 480 158.25 ;
      RECT 469.8 157.95 480 158.1 ;
      RECT 469.95 157.8 480 157.95 ;
      RECT 470.1 157.65 480 157.8 ;
      RECT 470.25 157.5 480 157.65 ;
      RECT 470.4 157.35 480 157.5 ;
      RECT 470.55 157.2 480 157.35 ;
      RECT 470.7 157.05 480 157.2 ;
      RECT 470.85 156.9 480 157.05 ;
      RECT 471.0 156.75 480 156.9 ;
      RECT 471.15 156.6 480 156.75 ;
      RECT 471.3 156.45 480 156.6 ;
      RECT 471.45 156.3 480 156.45 ;
      RECT 471.6 156.15 480 156.3 ;
      RECT 471.75 156 480 156.15 ;
      RECT 471.9 155.85 480 156 ;
      RECT 472.05 155.7 480 155.85 ;
      RECT 472.2 155.55 480 155.7 ;
      RECT 472.35 155.4 480 155.55 ;
      RECT 472.5 155.25 480 155.4 ;
      RECT 472.65 155.1 480 155.25 ;
      RECT 472.8 154.95 480 155.1 ;
      RECT 472.95 154.8 480 154.95 ;
      RECT 473.1 154.65 480 154.8 ;
      RECT 473.25 154.5 480 154.65 ;
      RECT 473.4 154.35 480 154.5 ;
      RECT 473.55 154.2 480 154.35 ;
      RECT 473.7 154.05 480 154.2 ;
      RECT 473.85 153.9 480 154.05 ;
      RECT 474.0 153.75 480 153.9 ;
      RECT 474.15 153.6 480 153.75 ;
      RECT 474.3 153.45 480 153.6 ;
      RECT 474.45 153.3 480 153.45 ;
      RECT 474.6 153.15 480 153.3 ;
      RECT 474.75 153 480 153.15 ;
      RECT 474.9 152.85 480 153 ;
      RECT 475.05 152.7 480 152.85 ;
      RECT 475.2 152.55 480 152.7 ;
      RECT 475.35 152.4 480 152.55 ;
      RECT 475.5 152.25 480 152.4 ;
      RECT 475.65 152.1 480 152.25 ;
      RECT 475.8 151.95 480 152.1 ;
      RECT 475.95 151.8 480 151.95 ;
      RECT 476.1 151.65 480 151.8 ;
      RECT 476.25 151.5 480 151.65 ;
      RECT 476.4 151.35 480 151.5 ;
      RECT 476.55 151.2 480 151.35 ;
      RECT 476.7 151.05 480 151.2 ;
      RECT 476.85 150.9 480 151.05 ;
      RECT 477.0 150.75 480 150.9 ;
      RECT 477.15 150.6 480 150.75 ;
      RECT 477.3 150.45 480 150.6 ;
      RECT 477.45 150.3 480 150.45 ;
      RECT 477.6 150.15 480 150.3 ;
      RECT 477.75 150 480 150.15 ;
      RECT 477.9 149.85 480 150 ;
      RECT 478.05 149.7 480 149.85 ;
      RECT 478.2 149.55 480 149.7 ;
      RECT 478.35 149.4 480 149.55 ;
      RECT 478.5 149.25 480 149.4 ;
      RECT 478.65 149.1 480 149.25 ;
      RECT 478.8 148.95 480 149.1 ;
      RECT 478.95 148.8 480 148.95 ;
      RECT 479.1 148.65 480 148.8 ;
      RECT 479.25 148.5 480 148.65 ;
      RECT 479.4 148.35 480 148.5 ;
      RECT 479.55 148.2 480 148.35 ;
      RECT 479.7 148.05 480 148.2 ;
      RECT 479.85 147.9 480 148.05 ;
      RECT 0 229.09 50.46 229.1 ;
      RECT 0 228.94 50.31 229.09 ;
      RECT 0 228.79 50.16 228.94 ;
      RECT 0 228.64 50.01 228.79 ;
      RECT 0 228.49 49.86 228.64 ;
      RECT 0 228.34 49.71 228.49 ;
      RECT 0 228.19 49.56 228.34 ;
      RECT 0 228.04 49.41 228.19 ;
      RECT 0 227.89 49.26 228.04 ;
      RECT 0 227.74 49.11 227.89 ;
      RECT 0 227.59 48.96 227.74 ;
      RECT 0 227.44 48.81 227.59 ;
      RECT 0 227.29 48.66 227.44 ;
      RECT 0 227.14 48.51 227.29 ;
      RECT 0 226.99 48.36 227.14 ;
      RECT 0 226.84 48.21 226.99 ;
      RECT 0 226.69 48.06 226.84 ;
      RECT 0 226.54 47.91 226.69 ;
      RECT 0 226.39 47.76 226.54 ;
      RECT 0 226.24 47.61 226.39 ;
      RECT 0 226.09 47.46 226.24 ;
      RECT 0 225.94 47.31 226.09 ;
      RECT 0 225.79 47.16 225.94 ;
      RECT 0 225.64 47.01 225.79 ;
      RECT 0 225.49 46.86 225.64 ;
      RECT 0 225.34 46.71 225.49 ;
      RECT 0 225.19 46.56 225.34 ;
      RECT 0 225.04 46.41 225.19 ;
      RECT 0 224.89 46.26 225.04 ;
      RECT 0 224.74 46.11 224.89 ;
      RECT 0 224.59 45.96 224.74 ;
      RECT 0 224.44 45.81 224.59 ;
      RECT 0 224.29 45.66 224.44 ;
      RECT 0 224.14 45.51 224.29 ;
      RECT 0 223.99 45.36 224.14 ;
      RECT 0 223.84 45.21 223.99 ;
      RECT 0 223.69 45.06 223.84 ;
      RECT 0 223.54 44.91 223.69 ;
      RECT 0 223.39 44.76 223.54 ;
      RECT 0 223.24 44.61 223.39 ;
      RECT 0 223.09 44.46 223.24 ;
      RECT 0 222.94 44.31 223.09 ;
      RECT 0 222.79 44.16 222.94 ;
      RECT 0 222.64 44.01 222.79 ;
      RECT 0 222.49 43.86 222.64 ;
      RECT 0 222.34 43.71 222.49 ;
      RECT 0 222.19 43.56 222.34 ;
      RECT 0 222.04 43.41 222.19 ;
      RECT 0 221.89 43.26 222.04 ;
      RECT 449.4 178.35 480 178.5 ;
      RECT 449.55 178.2 480 178.35 ;
      RECT 449.7 178.05 480 178.2 ;
      RECT 449.85 177.9 480 178.05 ;
      RECT 450.0 177.75 480 177.9 ;
      RECT 450.15 177.6 480 177.75 ;
      RECT 450.3 177.45 480 177.6 ;
      RECT 450.45 177.3 480 177.45 ;
      RECT 450.6 177.15 480 177.3 ;
      RECT 450.75 177 480 177.15 ;
      RECT 450.9 176.85 480 177 ;
      RECT 451.05 176.7 480 176.85 ;
      RECT 451.2 176.55 480 176.7 ;
      RECT 451.35 176.4 480 176.55 ;
      RECT 451.5 176.25 480 176.4 ;
      RECT 451.65 176.1 480 176.25 ;
      RECT 451.8 175.95 480 176.1 ;
      RECT 451.95 175.8 480 175.95 ;
      RECT 452.1 175.65 480 175.8 ;
      RECT 452.25 175.5 480 175.65 ;
      RECT 452.4 175.35 480 175.5 ;
      RECT 452.55 175.2 480 175.35 ;
      RECT 452.7 175.05 480 175.2 ;
      RECT 452.85 174.9 480 175.05 ;
      RECT 453.0 174.75 480 174.9 ;
      RECT 453.15 174.6 480 174.75 ;
      RECT 453.3 174.45 480 174.6 ;
      RECT 453.45 174.3 480 174.45 ;
      RECT 453.6 174.15 480 174.3 ;
      RECT 453.75 174 480 174.15 ;
      RECT 453.9 173.85 480 174 ;
      RECT 454.05 173.7 480 173.85 ;
      RECT 454.2 173.55 480 173.7 ;
      RECT 454.35 173.4 480 173.55 ;
      RECT 454.5 173.25 480 173.4 ;
      RECT 454.65 173.1 480 173.25 ;
      RECT 454.8 172.95 480 173.1 ;
      RECT 454.95 172.8 480 172.95 ;
      RECT 455.1 172.65 480 172.8 ;
      RECT 455.25 172.5 480 172.65 ;
      RECT 455.4 172.35 480 172.5 ;
      RECT 455.55 172.2 480 172.35 ;
      RECT 455.7 172.05 480 172.2 ;
      RECT 455.85 171.9 480 172.05 ;
      RECT 456.0 171.75 480 171.9 ;
      RECT 456.15 171.6 480 171.75 ;
      RECT 456.3 171.45 480 171.6 ;
      RECT 456.45 171.3 480 171.45 ;
      RECT 456.6 171.15 480 171.3 ;
      RECT 456.75 171 480 171.15 ;
      RECT 456.9 170.85 480 171 ;
      RECT 457.05 170.7 480 170.85 ;
      RECT 457.2 170.55 480 170.7 ;
      RECT 457.35 170.4 480 170.55 ;
      RECT 457.5 170.25 480 170.4 ;
      RECT 457.65 170.1 480 170.25 ;
      RECT 457.8 169.95 480 170.1 ;
      RECT 457.95 169.8 480 169.95 ;
      RECT 458.1 169.65 480 169.8 ;
      RECT 458.25 169.5 480 169.65 ;
      RECT 458.4 169.35 480 169.5 ;
      RECT 458.55 169.2 480 169.35 ;
      RECT 458.7 169.05 480 169.2 ;
      RECT 458.85 168.9 480 169.05 ;
      RECT 459.0 168.75 480 168.9 ;
      RECT 459.15 168.6 480 168.75 ;
      RECT 459.3 168.45 480 168.6 ;
      RECT 459.45 168.3 480 168.45 ;
      RECT 459.6 168.15 480 168.3 ;
      RECT 459.75 168 480 168.15 ;
      RECT 459.9 167.85 480 168 ;
      RECT 460.05 167.7 480 167.85 ;
      RECT 460.2 167.55 480 167.7 ;
      RECT 460.35 167.4 480 167.55 ;
      RECT 460.5 167.25 480 167.4 ;
      RECT 460.65 167.1 480 167.25 ;
      RECT 460.8 166.95 480 167.1 ;
      RECT 460.95 166.8 480 166.95 ;
      RECT 461.1 166.65 480 166.8 ;
      RECT 461.25 166.5 480 166.65 ;
      RECT 461.4 166.35 480 166.5 ;
      RECT 461.55 166.2 480 166.35 ;
      RECT 461.7 166.05 480 166.2 ;
      RECT 461.85 165.9 480 166.05 ;
      RECT 462.0 165.75 480 165.9 ;
      RECT 462.15 165.6 480 165.75 ;
      RECT 462.3 165.45 480 165.6 ;
      RECT 462.45 165.3 480 165.45 ;
      RECT 462.6 165.15 480 165.3 ;
      RECT 462.75 165 480 165.15 ;
      RECT 462.9 164.85 480 165 ;
      RECT 463.05 164.7 480 164.85 ;
      RECT 463.2 164.55 480 164.7 ;
      RECT 463.35 164.4 480 164.55 ;
      RECT 463.5 164.25 480 164.4 ;
      RECT 463.65 164.1 480 164.25 ;
      RECT 463.8 163.95 480 164.1 ;
      RECT 463.95 163.8 480 163.95 ;
      RECT 464.1 163.65 480 163.8 ;
      RECT 464.25 163.5 480 163.65 ;
      RECT 464.4 163.35 480 163.5 ;
      RECT 464.55 163.2 480 163.35 ;
      RECT 464.7 163.05 480 163.2 ;
      RECT 464.85 162.9 480 163.05 ;
      RECT 465.0 162.75 480 162.9 ;
      RECT 465.15 162.6 480 162.75 ;
      RECT 465.3 162.45 480 162.6 ;
      RECT 465.45 162.3 480 162.45 ;
      RECT 465.6 162.15 480 162.3 ;
      RECT 465.75 162 480 162.15 ;
      RECT 465.9 161.85 480 162 ;
      RECT 466.05 161.7 480 161.85 ;
      RECT 466.2 161.55 480 161.7 ;
      RECT 466.35 161.4 480 161.55 ;
      RECT 466.5 161.25 480 161.4 ;
      RECT 466.65 161.1 480 161.25 ;
      RECT 466.8 160.95 480 161.1 ;
      RECT 466.95 160.8 480 160.95 ;
      RECT 467.1 160.65 480 160.8 ;
      RECT 467.25 160.5 480 160.65 ;
      RECT 467.4 160.35 480 160.5 ;
      RECT 467.55 160.2 480 160.35 ;
      RECT 467.7 160.05 480 160.2 ;
      RECT 467.85 159.9 480 160.05 ;
      RECT 468.0 159.75 480 159.9 ;
      RECT 468.15 159.6 480 159.75 ;
      RECT 468.3 159.45 480 159.6 ;
      RECT 430.35 197.4 480 197.55 ;
      RECT 430.5 197.25 480 197.4 ;
      RECT 430.65 197.1 480 197.25 ;
      RECT 430.8 196.95 480 197.1 ;
      RECT 430.95 196.8 480 196.95 ;
      RECT 431.1 196.65 480 196.8 ;
      RECT 431.25 196.5 480 196.65 ;
      RECT 431.4 196.35 480 196.5 ;
      RECT 431.55 196.2 480 196.35 ;
      RECT 431.7 196.05 480 196.2 ;
      RECT 431.85 195.9 480 196.05 ;
      RECT 432.0 195.75 480 195.9 ;
      RECT 432.15 195.6 480 195.75 ;
      RECT 432.3 195.45 480 195.6 ;
      RECT 432.45 195.3 480 195.45 ;
      RECT 432.6 195.15 480 195.3 ;
      RECT 432.75 195 480 195.15 ;
      RECT 432.9 194.85 480 195 ;
      RECT 433.05 194.7 480 194.85 ;
      RECT 433.2 194.55 480 194.7 ;
      RECT 433.35 194.4 480 194.55 ;
      RECT 433.5 194.25 480 194.4 ;
      RECT 433.65 194.1 480 194.25 ;
      RECT 433.8 193.95 480 194.1 ;
      RECT 433.95 193.8 480 193.95 ;
      RECT 434.1 193.65 480 193.8 ;
      RECT 434.25 193.5 480 193.65 ;
      RECT 434.4 193.35 480 193.5 ;
      RECT 434.55 193.2 480 193.35 ;
      RECT 434.7 193.05 480 193.2 ;
      RECT 434.85 192.9 480 193.05 ;
      RECT 435.0 192.75 480 192.9 ;
      RECT 435.15 192.6 480 192.75 ;
      RECT 435.3 192.45 480 192.6 ;
      RECT 435.45 192.3 480 192.45 ;
      RECT 435.6 192.15 480 192.3 ;
      RECT 435.75 192 480 192.15 ;
      RECT 435.9 191.85 480 192 ;
      RECT 436.05 191.7 480 191.85 ;
      RECT 436.2 191.55 480 191.7 ;
      RECT 436.35 191.4 480 191.55 ;
      RECT 436.5 191.25 480 191.4 ;
      RECT 436.65 191.1 480 191.25 ;
      RECT 436.8 190.95 480 191.1 ;
      RECT 436.95 190.8 480 190.95 ;
      RECT 437.1 190.65 480 190.8 ;
      RECT 437.25 190.5 480 190.65 ;
      RECT 437.4 190.35 480 190.5 ;
      RECT 437.55 190.2 480 190.35 ;
      RECT 437.7 190.05 480 190.2 ;
      RECT 437.85 189.9 480 190.05 ;
      RECT 438.0 189.75 480 189.9 ;
      RECT 438.15 189.6 480 189.75 ;
      RECT 438.3 189.45 480 189.6 ;
      RECT 438.45 189.3 480 189.45 ;
      RECT 438.6 189.15 480 189.3 ;
      RECT 438.75 189 480 189.15 ;
      RECT 438.9 188.85 480 189 ;
      RECT 439.05 188.7 480 188.85 ;
      RECT 439.2 188.55 480 188.7 ;
      RECT 439.35 188.4 480 188.55 ;
      RECT 439.5 188.25 480 188.4 ;
      RECT 439.65 188.1 480 188.25 ;
      RECT 439.8 187.95 480 188.1 ;
      RECT 439.95 187.8 480 187.95 ;
      RECT 440.1 187.65 480 187.8 ;
      RECT 440.25 187.5 480 187.65 ;
      RECT 440.4 187.35 480 187.5 ;
      RECT 440.55 187.2 480 187.35 ;
      RECT 440.7 187.05 480 187.2 ;
      RECT 440.85 186.9 480 187.05 ;
      RECT 441.0 186.75 480 186.9 ;
      RECT 441.15 186.6 480 186.75 ;
      RECT 441.3 186.45 480 186.6 ;
      RECT 441.45 186.3 480 186.45 ;
      RECT 441.6 186.15 480 186.3 ;
      RECT 441.75 186 480 186.15 ;
      RECT 441.9 185.85 480 186 ;
      RECT 442.05 185.7 480 185.85 ;
      RECT 442.2 185.55 480 185.7 ;
      RECT 442.35 185.4 480 185.55 ;
      RECT 442.5 185.25 480 185.4 ;
      RECT 442.65 185.1 480 185.25 ;
      RECT 442.8 184.95 480 185.1 ;
      RECT 442.95 184.8 480 184.95 ;
      RECT 443.1 184.65 480 184.8 ;
      RECT 443.25 184.5 480 184.65 ;
      RECT 443.4 184.35 480 184.5 ;
      RECT 443.55 184.2 480 184.35 ;
      RECT 443.7 184.05 480 184.2 ;
      RECT 443.85 183.9 480 184.05 ;
      RECT 444.0 183.75 480 183.9 ;
      RECT 444.15 183.6 480 183.75 ;
      RECT 444.3 183.45 480 183.6 ;
      RECT 444.45 183.3 480 183.45 ;
      RECT 444.6 183.15 480 183.3 ;
      RECT 444.75 183 480 183.15 ;
      RECT 444.9 182.85 480 183 ;
      RECT 445.05 182.7 480 182.85 ;
      RECT 445.2 182.55 480 182.7 ;
      RECT 445.35 182.4 480 182.55 ;
      RECT 445.5 182.25 480 182.4 ;
      RECT 445.65 182.1 480 182.25 ;
      RECT 445.8 181.95 480 182.1 ;
      RECT 445.95 181.8 480 181.95 ;
      RECT 446.1 181.65 480 181.8 ;
      RECT 446.25 181.5 480 181.65 ;
      RECT 446.4 181.35 480 181.5 ;
      RECT 446.55 181.2 480 181.35 ;
      RECT 446.7 181.05 480 181.2 ;
      RECT 446.85 180.9 480 181.05 ;
      RECT 447.0 180.75 480 180.9 ;
      RECT 447.15 180.6 480 180.75 ;
      RECT 447.3 180.45 480 180.6 ;
      RECT 447.45 180.3 480 180.45 ;
      RECT 447.6 180.15 480 180.3 ;
      RECT 447.75 180 480 180.15 ;
      RECT 447.9 179.85 480 180 ;
      RECT 448.05 179.7 480 179.85 ;
      RECT 448.2 179.55 480 179.7 ;
      RECT 448.35 179.4 480 179.55 ;
      RECT 448.5 179.25 480 179.4 ;
      RECT 448.65 179.1 480 179.25 ;
      RECT 448.8 178.95 480 179.1 ;
      RECT 448.95 178.8 480 178.95 ;
      RECT 449.1 178.65 480 178.8 ;
      RECT 449.25 178.5 480 178.65 ;
      RECT 411.3 216.45 480 216.6 ;
      RECT 411.45 216.3 480 216.45 ;
      RECT 411.6 216.15 480 216.3 ;
      RECT 411.75 216 480 216.15 ;
      RECT 411.9 215.85 480 216 ;
      RECT 412.05 215.7 480 215.85 ;
      RECT 412.2 215.55 480 215.7 ;
      RECT 412.35 215.4 480 215.55 ;
      RECT 412.5 215.25 480 215.4 ;
      RECT 412.65 215.1 480 215.25 ;
      RECT 412.8 214.95 480 215.1 ;
      RECT 412.95 214.8 480 214.95 ;
      RECT 413.1 214.65 480 214.8 ;
      RECT 413.25 214.5 480 214.65 ;
      RECT 413.4 214.35 480 214.5 ;
      RECT 413.55 214.2 480 214.35 ;
      RECT 413.7 214.05 480 214.2 ;
      RECT 413.85 213.9 480 214.05 ;
      RECT 414.0 213.75 480 213.9 ;
      RECT 414.15 213.6 480 213.75 ;
      RECT 414.3 213.45 480 213.6 ;
      RECT 414.45 213.3 480 213.45 ;
      RECT 414.6 213.15 480 213.3 ;
      RECT 414.75 213 480 213.15 ;
      RECT 414.9 212.85 480 213 ;
      RECT 415.05 212.7 480 212.85 ;
      RECT 415.2 212.55 480 212.7 ;
      RECT 415.35 212.4 480 212.55 ;
      RECT 415.5 212.25 480 212.4 ;
      RECT 415.65 212.1 480 212.25 ;
      RECT 415.8 211.95 480 212.1 ;
      RECT 415.95 211.8 480 211.95 ;
      RECT 416.1 211.65 480 211.8 ;
      RECT 416.25 211.5 480 211.65 ;
      RECT 416.4 211.35 480 211.5 ;
      RECT 416.55 211.2 480 211.35 ;
      RECT 416.7 211.05 480 211.2 ;
      RECT 416.85 210.9 480 211.05 ;
      RECT 417.0 210.75 480 210.9 ;
      RECT 417.15 210.6 480 210.75 ;
      RECT 417.3 210.45 480 210.6 ;
      RECT 417.45 210.3 480 210.45 ;
      RECT 417.6 210.15 480 210.3 ;
      RECT 417.75 210 480 210.15 ;
      RECT 417.9 209.85 480 210 ;
      RECT 418.05 209.7 480 209.85 ;
      RECT 418.2 209.55 480 209.7 ;
      RECT 418.35 209.4 480 209.55 ;
      RECT 418.5 209.25 480 209.4 ;
      RECT 418.65 209.1 480 209.25 ;
      RECT 418.8 208.95 480 209.1 ;
      RECT 418.95 208.8 480 208.95 ;
      RECT 419.1 208.65 480 208.8 ;
      RECT 419.25 208.5 480 208.65 ;
      RECT 419.4 208.35 480 208.5 ;
      RECT 419.55 208.2 480 208.35 ;
      RECT 419.7 208.05 480 208.2 ;
      RECT 419.85 207.9 480 208.05 ;
      RECT 420.0 207.75 480 207.9 ;
      RECT 420.15 207.6 480 207.75 ;
      RECT 420.3 207.45 480 207.6 ;
      RECT 420.45 207.3 480 207.45 ;
      RECT 420.6 207.15 480 207.3 ;
      RECT 420.75 207 480 207.15 ;
      RECT 420.9 206.85 480 207 ;
      RECT 421.05 206.7 480 206.85 ;
      RECT 421.2 206.55 480 206.7 ;
      RECT 421.35 206.4 480 206.55 ;
      RECT 421.5 206.25 480 206.4 ;
      RECT 421.65 206.1 480 206.25 ;
      RECT 421.8 205.95 480 206.1 ;
      RECT 421.95 205.8 480 205.95 ;
      RECT 422.1 205.65 480 205.8 ;
      RECT 422.25 205.5 480 205.65 ;
      RECT 422.4 205.35 480 205.5 ;
      RECT 422.55 205.2 480 205.35 ;
      RECT 422.7 205.05 480 205.2 ;
      RECT 422.85 204.9 480 205.05 ;
      RECT 423.0 204.75 480 204.9 ;
      RECT 423.15 204.6 480 204.75 ;
      RECT 423.3 204.45 480 204.6 ;
      RECT 423.45 204.3 480 204.45 ;
      RECT 423.6 204.15 480 204.3 ;
      RECT 423.75 204 480 204.15 ;
      RECT 423.9 203.85 480 204 ;
      RECT 424.05 203.7 480 203.85 ;
      RECT 424.2 203.55 480 203.7 ;
      RECT 424.35 203.4 480 203.55 ;
      RECT 424.5 203.25 480 203.4 ;
      RECT 424.65 203.1 480 203.25 ;
      RECT 424.8 202.95 480 203.1 ;
      RECT 424.95 202.8 480 202.95 ;
      RECT 425.1 202.65 480 202.8 ;
      RECT 425.25 202.5 480 202.65 ;
      RECT 425.4 202.35 480 202.5 ;
      RECT 425.55 202.2 480 202.35 ;
      RECT 425.7 202.05 480 202.2 ;
      RECT 425.85 201.9 480 202.05 ;
      RECT 426.0 201.75 480 201.9 ;
      RECT 426.15 201.6 480 201.75 ;
      RECT 426.3 201.45 480 201.6 ;
      RECT 426.45 201.3 480 201.45 ;
      RECT 426.6 201.15 480 201.3 ;
      RECT 426.75 201 480 201.15 ;
      RECT 426.9 200.85 480 201 ;
      RECT 427.05 200.7 480 200.85 ;
      RECT 427.2 200.55 480 200.7 ;
      RECT 427.35 200.4 480 200.55 ;
      RECT 427.5 200.25 480 200.4 ;
      RECT 427.65 200.1 480 200.25 ;
      RECT 427.8 199.95 480 200.1 ;
      RECT 427.95 199.8 480 199.95 ;
      RECT 428.1 199.65 480 199.8 ;
      RECT 428.25 199.5 480 199.65 ;
      RECT 428.4 199.35 480 199.5 ;
      RECT 428.55 199.2 480 199.35 ;
      RECT 428.7 199.05 480 199.2 ;
      RECT 428.85 198.9 480 199.05 ;
      RECT 429.0 198.75 480 198.9 ;
      RECT 429.15 198.6 480 198.75 ;
      RECT 429.3 198.45 480 198.6 ;
      RECT 429.45 198.3 480 198.45 ;
      RECT 429.6 198.15 480 198.3 ;
      RECT 429.75 198 480 198.15 ;
      RECT 429.9 197.85 480 198 ;
      RECT 430.05 197.7 480 197.85 ;
      RECT 430.2 197.55 480 197.7 ;
      RECT 0 154.515 23.825 154.665 ;
      RECT 0 154.365 23.675 154.515 ;
      RECT 0 154.215 23.525 154.365 ;
      RECT 0 154.065 23.375 154.215 ;
      RECT 0 153.915 23.225 154.065 ;
      RECT 0 153.765 23.075 153.915 ;
      RECT 0 153.615 22.925 153.765 ;
      RECT 0 153.465 22.775 153.615 ;
      RECT 0 153.315 22.625 153.465 ;
      RECT 0 153.165 22.475 153.315 ;
      RECT 0 153.015 22.325 153.165 ;
      RECT 0 152.865 22.175 153.015 ;
      RECT 0 152.715 22.025 152.865 ;
      RECT 0 152.565 21.875 152.715 ;
      RECT 0 152.415 21.725 152.565 ;
      RECT 0 152.265 21.575 152.415 ;
      RECT 0 152.115 21.425 152.265 ;
      RECT 0 151.965 21.275 152.115 ;
      RECT 0 151.815 21.125 151.965 ;
      RECT 0 151.665 20.975 151.815 ;
      RECT 0 151.515 20.825 151.665 ;
      RECT 0 151.365 20.675 151.515 ;
      RECT 0 151.215 20.525 151.365 ;
      RECT 0 151.065 20.375 151.215 ;
      RECT 0 150.915 20.225 151.065 ;
      RECT 0 150.765 20.075 150.915 ;
      RECT 0 150.615 19.925 150.765 ;
      RECT 0 150.465 19.775 150.615 ;
      RECT 0 150.315 19.625 150.465 ;
      RECT 0 150.165 19.475 150.315 ;
      RECT 0 150.015 19.325 150.165 ;
      RECT 0 149.865 19.175 150.015 ;
      RECT 0 149.715 19.025 149.865 ;
      RECT 0 149.565 18.875 149.715 ;
      RECT 0 149.415 18.725 149.565 ;
      RECT 0 149.265 18.575 149.415 ;
      RECT 0 149.115 18.425 149.265 ;
      RECT 49.82 228.3 399.3 228.45 ;
      RECT 49.97 228.45 399.15 228.6 ;
      RECT 50.12 228.6 399.0 228.75 ;
      RECT 50.27 228.75 398.85 228.9 ;
      RECT 50.42 228.9 398.7 229.05 ;
      RECT 50.47 229.05 398.65 229.1 ;
      RECT 398.7 229.05 480 229.1 ;
      RECT 398.85 228.9 480 229.05 ;
      RECT 399.0 228.75 480 228.9 ;
      RECT 399.15 228.6 480 228.75 ;
      RECT 399.3 228.45 480 228.6 ;
      RECT 399.45 228.3 480 228.45 ;
      RECT 399.6 228.15 480 228.3 ;
      RECT 399.75 228 480 228.15 ;
      RECT 399.9 227.85 480 228 ;
      RECT 400.05 227.7 480 227.85 ;
      RECT 400.2 227.55 480 227.7 ;
      RECT 400.35 227.4 480 227.55 ;
      RECT 400.5 227.25 480 227.4 ;
      RECT 400.65 227.1 480 227.25 ;
      RECT 400.8 226.95 480 227.1 ;
      RECT 400.95 226.8 480 226.95 ;
      RECT 401.1 226.65 480 226.8 ;
      RECT 401.25 226.5 480 226.65 ;
      RECT 401.4 226.35 480 226.5 ;
      RECT 401.55 226.2 480 226.35 ;
      RECT 401.7 226.05 480 226.2 ;
      RECT 401.85 225.9 480 226.05 ;
      RECT 402.0 225.75 480 225.9 ;
      RECT 402.15 225.6 480 225.75 ;
      RECT 402.3 225.45 480 225.6 ;
      RECT 402.45 225.3 480 225.45 ;
      RECT 402.6 225.15 480 225.3 ;
      RECT 402.75 225 480 225.15 ;
      RECT 402.9 224.85 480 225 ;
      RECT 403.05 224.7 480 224.85 ;
      RECT 403.2 224.55 480 224.7 ;
      RECT 403.35 224.4 480 224.55 ;
      RECT 403.5 224.25 480 224.4 ;
      RECT 403.65 224.1 480 224.25 ;
      RECT 403.8 223.95 480 224.1 ;
      RECT 403.95 223.8 480 223.95 ;
      RECT 404.1 223.65 480 223.8 ;
      RECT 404.25 223.5 480 223.65 ;
      RECT 404.4 223.35 480 223.5 ;
      RECT 404.55 223.2 480 223.35 ;
      RECT 404.7 223.05 480 223.2 ;
      RECT 404.85 222.9 480 223.05 ;
      RECT 405.0 222.75 480 222.9 ;
      RECT 405.15 222.6 480 222.75 ;
      RECT 405.3 222.45 480 222.6 ;
      RECT 405.45 222.3 480 222.45 ;
      RECT 405.6 222.15 480 222.3 ;
      RECT 405.75 222 480 222.15 ;
      RECT 405.9 221.85 480 222 ;
      RECT 406.05 221.7 480 221.85 ;
      RECT 406.2 221.55 480 221.7 ;
      RECT 406.35 221.4 480 221.55 ;
      RECT 406.5 221.25 480 221.4 ;
      RECT 406.65 221.1 480 221.25 ;
      RECT 406.8 220.95 480 221.1 ;
      RECT 406.95 220.8 480 220.95 ;
      RECT 407.1 220.65 480 220.8 ;
      RECT 407.25 220.5 480 220.65 ;
      RECT 407.4 220.35 480 220.5 ;
      RECT 407.55 220.2 480 220.35 ;
      RECT 407.7 220.05 480 220.2 ;
      RECT 407.85 219.9 480 220.05 ;
      RECT 408.0 219.75 480 219.9 ;
      RECT 408.15 219.6 480 219.75 ;
      RECT 408.3 219.45 480 219.6 ;
      RECT 408.45 219.3 480 219.45 ;
      RECT 408.6 219.15 480 219.3 ;
      RECT 408.75 219 480 219.15 ;
      RECT 408.9 218.85 480 219 ;
      RECT 409.05 218.7 480 218.85 ;
      RECT 409.2 218.55 480 218.7 ;
      RECT 409.35 218.4 480 218.55 ;
      RECT 409.5 218.25 480 218.4 ;
      RECT 409.65 218.1 480 218.25 ;
      RECT 409.8 217.95 480 218.1 ;
      RECT 409.95 217.8 480 217.95 ;
      RECT 410.1 217.65 480 217.8 ;
      RECT 410.25 217.5 480 217.65 ;
      RECT 410.4 217.35 480 217.5 ;
      RECT 410.55 217.2 480 217.35 ;
      RECT 410.7 217.05 480 217.2 ;
      RECT 410.85 216.9 480 217.05 ;
      RECT 411.0 216.75 480 216.9 ;
      RECT 411.15 216.6 480 216.75 ;
      RECT 0 221.29 42.66 221.44 ;
      RECT 0 221.14 42.51 221.29 ;
      RECT 0 220.99 42.36 221.14 ;
      RECT 0 220.84 42.21 220.99 ;
      RECT 0 220.69 42.06 220.84 ;
      RECT 0 220.54 41.91 220.69 ;
      RECT 0 220.39 41.76 220.54 ;
      RECT 0 220.24 41.61 220.39 ;
      RECT 0 220.09 41.46 220.24 ;
      RECT 0 219.94 41.31 220.09 ;
      RECT 0 219.79 41.16 219.94 ;
      RECT 0 219.64 41.01 219.79 ;
      RECT 0 219.49 40.86 219.64 ;
      RECT 0 219.34 40.71 219.49 ;
      RECT 0 219.19 40.56 219.34 ;
      RECT 0 219.04 40.41 219.19 ;
      RECT 0 218.89 40.26 219.04 ;
      RECT 0 218.74 40.11 218.89 ;
      RECT 0 218.59 39.96 218.74 ;
      RECT 0 218.44 39.81 218.59 ;
      RECT 0 218.29 39.66 218.44 ;
      RECT 0 218.14 39.51 218.29 ;
      RECT 0 217.99 39.36 218.14 ;
      RECT 0 217.84 39.21 217.99 ;
      RECT 0 217.69 39.06 217.84 ;
      RECT 0 217.54 38.91 217.69 ;
      RECT 0 217.39 38.76 217.54 ;
      RECT 0 217.24 38.61 217.39 ;
      RECT 0 217.09 38.46 217.24 ;
      RECT 0 216.94 38.31 217.09 ;
      RECT 0 216.79 38.16 216.94 ;
      RECT 0 216.64 38.01 216.79 ;
      RECT 0 216.49 37.86 216.64 ;
      RECT 0 216.34 37.71 216.49 ;
      RECT 0 216.19 37.56 216.34 ;
      RECT 0 216.04 37.41 216.19 ;
      RECT 0 215.89 37.26 216.04 ;
      RECT 0 215.74 37.11 215.89 ;
      RECT 0 215.59 36.96 215.74 ;
      RECT 0 215.44 36.81 215.59 ;
      RECT 0 215.29 36.66 215.44 ;
      RECT 0 215.14 36.51 215.29 ;
      RECT 0 214.99 36.36 215.14 ;
      RECT 0 214.84 36.21 214.99 ;
      RECT 0 214.69 36.06 214.84 ;
      RECT 0 214.54 35.91 214.69 ;
      RECT 0 214.39 35.76 214.54 ;
      RECT 0 214.24 35.61 214.39 ;
      RECT 0 214.09 35.46 214.24 ;
      RECT 0 213.94 35.31 214.09 ;
      RECT 0 213.79 35.16 213.94 ;
      RECT 0 213.64 35.01 213.79 ;
      RECT 0 213.49 34.86 213.64 ;
      RECT 0 213.34 34.71 213.49 ;
      RECT 0 213.19 34.56 213.34 ;
      RECT 0 213.04 34.41 213.19 ;
      RECT 0 212.89 34.26 213.04 ;
      RECT 0 212.74 34.11 212.89 ;
      RECT 0 212.59 33.96 212.74 ;
      RECT 0 212.44 33.81 212.59 ;
      RECT 0 212.29 33.66 212.44 ;
      RECT 0 212.14 33.51 212.29 ;
      RECT 0 211.99 33.36 212.14 ;
      RECT 0 211.84 33.21 211.99 ;
      RECT 0 211.69 33.06 211.84 ;
      RECT 0 211.54 32.91 211.69 ;
      RECT 0 211.39 32.76 211.54 ;
      RECT 0 211.24 32.61 211.39 ;
      RECT 0 211.09 32.46 211.24 ;
      RECT 0 210.94 32.31 211.09 ;
      RECT 0 210.79 32.16 210.94 ;
      RECT 0 210.64 32.01 210.79 ;
      RECT 0 210.49 31.86 210.64 ;
      RECT 0 210.34 31.71 210.49 ;
      RECT 0 210.19 31.56 210.34 ;
      RECT 0 210.04 31.41 210.19 ;
      RECT 0 209.89 31.26 210.04 ;
      RECT 0 209.74 31.11 209.89 ;
      RECT 0 209.59 30.96 209.74 ;
      RECT 0 209.44 30.81 209.59 ;
      RECT 0 209.29 30.66 209.44 ;
      RECT 0 209.14 30.51 209.29 ;
      RECT 0 208.99 30.36 209.14 ;
      RECT 0 208.84 30.21 208.99 ;
      RECT 0 208.69 30.06 208.84 ;
      RECT 0 208.54 29.91 208.69 ;
      RECT 0 208.39 29.76 208.54 ;
      RECT 0 208.24 29.61 208.39 ;
      RECT 0 208.09 29.46 208.24 ;
      RECT 0 207.94 29.31 208.09 ;
      RECT 0 207.79 29.16 207.94 ;
      RECT 0 207.64 29.01 207.79 ;
      RECT 0 207.49 28.86 207.64 ;
      RECT 0 159.465 28.775 159.55 ;
      RECT 0 159.315 28.625 159.465 ;
      RECT 0 159.165 28.475 159.315 ;
      RECT 0 159.015 28.325 159.165 ;
      RECT 0 158.865 28.175 159.015 ;
      RECT 0 158.715 28.025 158.865 ;
      RECT 0 158.565 27.875 158.715 ;
      RECT 0 158.415 27.725 158.565 ;
      RECT 0 158.265 27.575 158.415 ;
      RECT 0 158.115 27.425 158.265 ;
      RECT 0 157.965 27.275 158.115 ;
      RECT 0 157.815 27.125 157.965 ;
      RECT 0 157.665 26.975 157.815 ;
      RECT 0 157.515 26.825 157.665 ;
      RECT 0 157.365 26.675 157.515 ;
      RECT 0 157.215 26.525 157.365 ;
      RECT 0 157.065 26.375 157.215 ;
      RECT 0 156.915 26.225 157.065 ;
      RECT 0 156.765 26.075 156.915 ;
      RECT 0 156.615 25.925 156.765 ;
      RECT 0 156.465 25.775 156.615 ;
      RECT 0 156.315 25.625 156.465 ;
      RECT 0 156.165 25.475 156.315 ;
      RECT 0 156.015 25.325 156.165 ;
      RECT 0 155.865 25.175 156.015 ;
      RECT 0 155.715 25.025 155.865 ;
      RECT 0 155.565 24.875 155.715 ;
      RECT 0 155.415 24.725 155.565 ;
      RECT 0 155.265 24.575 155.415 ;
      RECT 0 155.115 24.425 155.265 ;
      RECT 0 154.965 24.275 155.115 ;
      RECT 0 154.815 24.125 154.965 ;
      RECT 0 154.665 23.975 154.815 ;
      RECT 468.9 158.85 480 159 ;
      RECT 469.05 158.7 480 158.85 ;
      RECT 469.2 158.55 480 158.7 ;
      RECT 469.35 158.4 480 158.55 ;
      RECT 469.5 158.25 480 158.4 ;
      RECT 469.65 158.1 480 158.25 ;
      RECT 469.8 157.95 480 158.1 ;
      RECT 469.95 157.8 480 157.95 ;
      RECT 470.1 157.65 480 157.8 ;
      RECT 470.25 157.5 480 157.65 ;
      RECT 470.4 157.35 480 157.5 ;
      RECT 470.55 157.2 480 157.35 ;
      RECT 470.7 157.05 480 157.2 ;
      RECT 470.85 156.9 480 157.05 ;
      RECT 471.0 156.75 480 156.9 ;
      RECT 471.15 156.6 480 156.75 ;
      RECT 471.3 156.45 480 156.6 ;
      RECT 471.45 156.3 480 156.45 ;
      RECT 471.6 156.15 480 156.3 ;
      RECT 471.75 156 480 156.15 ;
      RECT 471.9 155.85 480 156 ;
      RECT 472.05 155.7 480 155.85 ;
      RECT 472.2 155.55 480 155.7 ;
      RECT 472.35 155.4 480 155.55 ;
      RECT 472.5 155.25 480 155.4 ;
      RECT 472.65 155.1 480 155.25 ;
      RECT 472.8 154.95 480 155.1 ;
      RECT 472.95 154.8 480 154.95 ;
      RECT 473.1 154.65 480 154.8 ;
      RECT 473.25 154.5 480 154.65 ;
      RECT 473.4 154.35 480 154.5 ;
      RECT 473.55 154.2 480 154.35 ;
      RECT 473.7 154.05 480 154.2 ;
      RECT 473.85 153.9 480 154.05 ;
      RECT 474.0 153.75 480 153.9 ;
      RECT 474.15 153.6 480 153.75 ;
      RECT 474.3 153.45 480 153.6 ;
      RECT 474.45 153.3 480 153.45 ;
      RECT 474.6 153.15 480 153.3 ;
      RECT 474.75 153 480 153.15 ;
      RECT 474.9 152.85 480 153 ;
      RECT 475.05 152.7 480 152.85 ;
      RECT 475.2 152.55 480 152.7 ;
      RECT 475.35 152.4 480 152.55 ;
      RECT 475.5 152.25 480 152.4 ;
      RECT 475.65 152.1 480 152.25 ;
      RECT 475.8 151.95 480 152.1 ;
      RECT 475.95 151.8 480 151.95 ;
      RECT 476.1 151.65 480 151.8 ;
      RECT 476.25 151.5 480 151.65 ;
      RECT 476.4 151.35 480 151.5 ;
      RECT 476.55 151.2 480 151.35 ;
      RECT 476.7 151.05 480 151.2 ;
      RECT 476.85 150.9 480 151.05 ;
      RECT 477.0 150.75 480 150.9 ;
      RECT 477.15 150.6 480 150.75 ;
      RECT 477.3 150.45 480 150.6 ;
      RECT 477.45 150.3 480 150.45 ;
      RECT 477.6 150.15 480 150.3 ;
      RECT 477.75 150 480 150.15 ;
      RECT 477.9 149.85 480 150 ;
      RECT 478.05 149.7 480 149.85 ;
      RECT 478.2 149.55 480 149.7 ;
      RECT 478.35 149.4 480 149.55 ;
      RECT 478.5 149.25 480 149.4 ;
      RECT 478.65 149.1 480 149.25 ;
      RECT 478.8 148.95 480 149.1 ;
      RECT 478.95 148.8 480 148.95 ;
      RECT 479.1 148.65 480 148.8 ;
      RECT 479.25 148.5 480 148.65 ;
      RECT 479.4 148.35 480 148.5 ;
      RECT 479.55 148.2 480 148.35 ;
      RECT 479.7 148.05 480 148.2 ;
      RECT 479.85 147.9 480 148.05 ;
      RECT 0 229.09 50.46 229.1 ;
      RECT 0 228.94 50.31 229.09 ;
      RECT 0 228.79 50.16 228.94 ;
      RECT 0 228.64 50.01 228.79 ;
      RECT 0 228.49 49.86 228.64 ;
      RECT 0 228.34 49.71 228.49 ;
      RECT 0 228.19 49.56 228.34 ;
      RECT 0 228.04 49.41 228.19 ;
      RECT 0 227.89 49.26 228.04 ;
      RECT 0 227.74 49.11 227.89 ;
      RECT 0 227.59 48.96 227.74 ;
      RECT 0 227.44 48.81 227.59 ;
      RECT 0 227.29 48.66 227.44 ;
      RECT 0 227.14 48.51 227.29 ;
      RECT 0 226.99 48.36 227.14 ;
      RECT 0 226.84 48.21 226.99 ;
      RECT 0 226.69 48.06 226.84 ;
      RECT 0 226.54 47.91 226.69 ;
      RECT 0 226.39 47.76 226.54 ;
      RECT 0 226.24 47.61 226.39 ;
      RECT 0 226.09 47.46 226.24 ;
      RECT 0 225.94 47.31 226.09 ;
      RECT 0 225.79 47.16 225.94 ;
      RECT 0 225.64 47.01 225.79 ;
      RECT 0 225.49 46.86 225.64 ;
      RECT 0 225.34 46.71 225.49 ;
      RECT 0 225.19 46.56 225.34 ;
      RECT 0 225.04 46.41 225.19 ;
      RECT 0 224.89 46.26 225.04 ;
      RECT 0 224.74 46.11 224.89 ;
      RECT 0 224.59 45.96 224.74 ;
      RECT 0 224.44 45.81 224.59 ;
      RECT 0 224.29 45.66 224.44 ;
      RECT 0 224.14 45.51 224.29 ;
      RECT 0 223.99 45.36 224.14 ;
      RECT 0 223.84 45.21 223.99 ;
      RECT 0 223.69 45.06 223.84 ;
      RECT 0 223.54 44.91 223.69 ;
      RECT 0 223.39 44.76 223.54 ;
      RECT 0 223.24 44.61 223.39 ;
      RECT 0 223.09 44.46 223.24 ;
      RECT 0 222.94 44.31 223.09 ;
      RECT 0 222.79 44.16 222.94 ;
      RECT 0 222.64 44.01 222.79 ;
      RECT 0 222.49 43.86 222.64 ;
      RECT 0 222.34 43.71 222.49 ;
      RECT 0 222.19 43.56 222.34 ;
      RECT 0 222.04 43.41 222.19 ;
      RECT 0 221.89 43.26 222.04 ;
      RECT 0 221.74 43.11 221.89 ;
      RECT 0 221.59 42.96 221.74 ;
      RECT 0 221.44 42.81 221.59 ;
      RECT 449.85 177.9 480 178.05 ;
      RECT 450.0 177.75 480 177.9 ;
      RECT 450.15 177.6 480 177.75 ;
      RECT 450.3 177.45 480 177.6 ;
      RECT 450.45 177.3 480 177.45 ;
      RECT 450.6 177.15 480 177.3 ;
      RECT 450.75 177 480 177.15 ;
      RECT 450.9 176.85 480 177 ;
      RECT 451.05 176.7 480 176.85 ;
      RECT 451.2 176.55 480 176.7 ;
      RECT 451.35 176.4 480 176.55 ;
      RECT 451.5 176.25 480 176.4 ;
      RECT 451.65 176.1 480 176.25 ;
      RECT 451.8 175.95 480 176.1 ;
      RECT 451.95 175.8 480 175.95 ;
      RECT 452.1 175.65 480 175.8 ;
      RECT 452.25 175.5 480 175.65 ;
      RECT 452.4 175.35 480 175.5 ;
      RECT 452.55 175.2 480 175.35 ;
      RECT 452.7 175.05 480 175.2 ;
      RECT 452.85 174.9 480 175.05 ;
      RECT 453.0 174.75 480 174.9 ;
      RECT 453.15 174.6 480 174.75 ;
      RECT 453.3 174.45 480 174.6 ;
      RECT 453.45 174.3 480 174.45 ;
      RECT 453.6 174.15 480 174.3 ;
      RECT 453.75 174 480 174.15 ;
      RECT 453.9 173.85 480 174 ;
      RECT 454.05 173.7 480 173.85 ;
      RECT 454.2 173.55 480 173.7 ;
      RECT 454.35 173.4 480 173.55 ;
      RECT 454.5 173.25 480 173.4 ;
      RECT 454.65 173.1 480 173.25 ;
      RECT 454.8 172.95 480 173.1 ;
      RECT 454.95 172.8 480 172.95 ;
      RECT 455.1 172.65 480 172.8 ;
      RECT 455.25 172.5 480 172.65 ;
      RECT 455.4 172.35 480 172.5 ;
      RECT 455.55 172.2 480 172.35 ;
      RECT 455.7 172.05 480 172.2 ;
      RECT 455.85 171.9 480 172.05 ;
      RECT 456.0 171.75 480 171.9 ;
      RECT 456.15 171.6 480 171.75 ;
      RECT 456.3 171.45 480 171.6 ;
      RECT 456.45 171.3 480 171.45 ;
      RECT 456.6 171.15 480 171.3 ;
      RECT 456.75 171 480 171.15 ;
      RECT 456.9 170.85 480 171 ;
      RECT 457.05 170.7 480 170.85 ;
      RECT 457.2 170.55 480 170.7 ;
      RECT 457.35 170.4 480 170.55 ;
      RECT 457.5 170.25 480 170.4 ;
      RECT 457.65 170.1 480 170.25 ;
      RECT 457.8 169.95 480 170.1 ;
      RECT 457.95 169.8 480 169.95 ;
      RECT 458.1 169.65 480 169.8 ;
      RECT 458.25 169.5 480 169.65 ;
      RECT 458.4 169.35 480 169.5 ;
      RECT 458.55 169.2 480 169.35 ;
      RECT 458.7 169.05 480 169.2 ;
      RECT 458.85 168.9 480 169.05 ;
      RECT 459.0 168.75 480 168.9 ;
      RECT 459.15 168.6 480 168.75 ;
      RECT 459.3 168.45 480 168.6 ;
      RECT 459.45 168.3 480 168.45 ;
      RECT 459.6 168.15 480 168.3 ;
      RECT 459.75 168 480 168.15 ;
      RECT 459.9 167.85 480 168 ;
      RECT 460.05 167.7 480 167.85 ;
      RECT 460.2 167.55 480 167.7 ;
      RECT 460.35 167.4 480 167.55 ;
      RECT 460.5 167.25 480 167.4 ;
      RECT 460.65 167.1 480 167.25 ;
      RECT 460.8 166.95 480 167.1 ;
      RECT 460.95 166.8 480 166.95 ;
      RECT 461.1 166.65 480 166.8 ;
      RECT 461.25 166.5 480 166.65 ;
      RECT 461.4 166.35 480 166.5 ;
      RECT 461.55 166.2 480 166.35 ;
      RECT 461.7 166.05 480 166.2 ;
      RECT 461.85 165.9 480 166.05 ;
      RECT 462.0 165.75 480 165.9 ;
      RECT 462.15 165.6 480 165.75 ;
      RECT 462.3 165.45 480 165.6 ;
      RECT 462.45 165.3 480 165.45 ;
      RECT 462.6 165.15 480 165.3 ;
      RECT 462.75 165 480 165.15 ;
      RECT 462.9 164.85 480 165 ;
      RECT 463.05 164.7 480 164.85 ;
      RECT 463.2 164.55 480 164.7 ;
      RECT 463.35 164.4 480 164.55 ;
      RECT 463.5 164.25 480 164.4 ;
      RECT 463.65 164.1 480 164.25 ;
      RECT 463.8 163.95 480 164.1 ;
      RECT 463.95 163.8 480 163.95 ;
      RECT 464.1 163.65 480 163.8 ;
      RECT 464.25 163.5 480 163.65 ;
      RECT 464.4 163.35 480 163.5 ;
      RECT 464.55 163.2 480 163.35 ;
      RECT 464.7 163.05 480 163.2 ;
      RECT 464.85 162.9 480 163.05 ;
      RECT 465.0 162.75 480 162.9 ;
      RECT 465.15 162.6 480 162.75 ;
      RECT 465.3 162.45 480 162.6 ;
      RECT 465.45 162.3 480 162.45 ;
      RECT 465.6 162.15 480 162.3 ;
      RECT 465.75 162 480 162.15 ;
      RECT 465.9 161.85 480 162 ;
      RECT 466.05 161.7 480 161.85 ;
      RECT 466.2 161.55 480 161.7 ;
      RECT 466.35 161.4 480 161.55 ;
      RECT 466.5 161.25 480 161.4 ;
      RECT 466.65 161.1 480 161.25 ;
      RECT 466.8 160.95 480 161.1 ;
      RECT 466.95 160.8 480 160.95 ;
      RECT 467.1 160.65 480 160.8 ;
      RECT 467.25 160.5 480 160.65 ;
      RECT 467.4 160.35 480 160.5 ;
      RECT 467.55 160.2 480 160.35 ;
      RECT 467.7 160.05 480 160.2 ;
      RECT 467.85 159.9 480 160.05 ;
      RECT 468.0 159.75 480 159.9 ;
      RECT 468.15 159.6 480 159.75 ;
      RECT 468.3 159.45 480 159.6 ;
      RECT 468.45 159.3 480 159.45 ;
      RECT 468.6 159.15 480 159.3 ;
      RECT 468.75 159 480 159.15 ;
      RECT 430.8 196.95 480 197.1 ;
      RECT 430.95 196.8 480 196.95 ;
      RECT 431.1 196.65 480 196.8 ;
      RECT 431.25 196.5 480 196.65 ;
      RECT 431.4 196.35 480 196.5 ;
      RECT 431.55 196.2 480 196.35 ;
      RECT 431.7 196.05 480 196.2 ;
      RECT 431.85 195.9 480 196.05 ;
      RECT 432.0 195.75 480 195.9 ;
      RECT 432.15 195.6 480 195.75 ;
      RECT 432.3 195.45 480 195.6 ;
      RECT 432.45 195.3 480 195.45 ;
      RECT 432.6 195.15 480 195.3 ;
      RECT 432.75 195 480 195.15 ;
      RECT 432.9 194.85 480 195 ;
      RECT 433.05 194.7 480 194.85 ;
      RECT 433.2 194.55 480 194.7 ;
      RECT 433.35 194.4 480 194.55 ;
      RECT 433.5 194.25 480 194.4 ;
      RECT 433.65 194.1 480 194.25 ;
      RECT 433.8 193.95 480 194.1 ;
      RECT 433.95 193.8 480 193.95 ;
      RECT 434.1 193.65 480 193.8 ;
      RECT 434.25 193.5 480 193.65 ;
      RECT 434.4 193.35 480 193.5 ;
      RECT 434.55 193.2 480 193.35 ;
      RECT 434.7 193.05 480 193.2 ;
      RECT 434.85 192.9 480 193.05 ;
      RECT 435.0 192.75 480 192.9 ;
      RECT 435.15 192.6 480 192.75 ;
      RECT 435.3 192.45 480 192.6 ;
      RECT 435.45 192.3 480 192.45 ;
      RECT 435.6 192.15 480 192.3 ;
      RECT 435.75 192 480 192.15 ;
      RECT 435.9 191.85 480 192 ;
      RECT 436.05 191.7 480 191.85 ;
      RECT 436.2 191.55 480 191.7 ;
      RECT 436.35 191.4 480 191.55 ;
      RECT 436.5 191.25 480 191.4 ;
      RECT 436.65 191.1 480 191.25 ;
      RECT 436.8 190.95 480 191.1 ;
      RECT 436.95 190.8 480 190.95 ;
      RECT 437.1 190.65 480 190.8 ;
      RECT 437.25 190.5 480 190.65 ;
      RECT 437.4 190.35 480 190.5 ;
      RECT 437.55 190.2 480 190.35 ;
      RECT 437.7 190.05 480 190.2 ;
      RECT 437.85 189.9 480 190.05 ;
      RECT 438.0 189.75 480 189.9 ;
      RECT 438.15 189.6 480 189.75 ;
      RECT 438.3 189.45 480 189.6 ;
      RECT 438.45 189.3 480 189.45 ;
      RECT 438.6 189.15 480 189.3 ;
      RECT 438.75 189 480 189.15 ;
      RECT 438.9 188.85 480 189 ;
      RECT 439.05 188.7 480 188.85 ;
      RECT 439.2 188.55 480 188.7 ;
      RECT 439.35 188.4 480 188.55 ;
      RECT 439.5 188.25 480 188.4 ;
      RECT 439.65 188.1 480 188.25 ;
      RECT 439.8 187.95 480 188.1 ;
      RECT 439.95 187.8 480 187.95 ;
      RECT 440.1 187.65 480 187.8 ;
      RECT 440.25 187.5 480 187.65 ;
      RECT 440.4 187.35 480 187.5 ;
      RECT 440.55 187.2 480 187.35 ;
      RECT 440.7 187.05 480 187.2 ;
      RECT 440.85 186.9 480 187.05 ;
      RECT 441.0 186.75 480 186.9 ;
      RECT 441.15 186.6 480 186.75 ;
      RECT 441.3 186.45 480 186.6 ;
      RECT 441.45 186.3 480 186.45 ;
      RECT 441.6 186.15 480 186.3 ;
      RECT 441.75 186 480 186.15 ;
      RECT 441.9 185.85 480 186 ;
      RECT 442.05 185.7 480 185.85 ;
      RECT 442.2 185.55 480 185.7 ;
      RECT 442.35 185.4 480 185.55 ;
      RECT 442.5 185.25 480 185.4 ;
      RECT 442.65 185.1 480 185.25 ;
      RECT 442.8 184.95 480 185.1 ;
      RECT 442.95 184.8 480 184.95 ;
      RECT 443.1 184.65 480 184.8 ;
      RECT 443.25 184.5 480 184.65 ;
      RECT 443.4 184.35 480 184.5 ;
      RECT 443.55 184.2 480 184.35 ;
      RECT 443.7 184.05 480 184.2 ;
      RECT 443.85 183.9 480 184.05 ;
      RECT 444.0 183.75 480 183.9 ;
      RECT 444.15 183.6 480 183.75 ;
      RECT 444.3 183.45 480 183.6 ;
      RECT 444.45 183.3 480 183.45 ;
      RECT 444.6 183.15 480 183.3 ;
      RECT 444.75 183 480 183.15 ;
      RECT 444.9 182.85 480 183 ;
      RECT 445.05 182.7 480 182.85 ;
      RECT 445.2 182.55 480 182.7 ;
      RECT 445.35 182.4 480 182.55 ;
      RECT 445.5 182.25 480 182.4 ;
      RECT 445.65 182.1 480 182.25 ;
      RECT 445.8 181.95 480 182.1 ;
      RECT 445.95 181.8 480 181.95 ;
      RECT 446.1 181.65 480 181.8 ;
      RECT 446.25 181.5 480 181.65 ;
      RECT 446.4 181.35 480 181.5 ;
      RECT 446.55 181.2 480 181.35 ;
      RECT 446.7 181.05 480 181.2 ;
      RECT 446.85 180.9 480 181.05 ;
      RECT 447.0 180.75 480 180.9 ;
      RECT 447.15 180.6 480 180.75 ;
      RECT 447.3 180.45 480 180.6 ;
      RECT 447.45 180.3 480 180.45 ;
      RECT 447.6 180.15 480 180.3 ;
      RECT 447.75 180 480 180.15 ;
      RECT 447.9 179.85 480 180 ;
      RECT 448.05 179.7 480 179.85 ;
      RECT 448.2 179.55 480 179.7 ;
      RECT 448.35 179.4 480 179.55 ;
      RECT 448.5 179.25 480 179.4 ;
      RECT 448.65 179.1 480 179.25 ;
      RECT 448.8 178.95 480 179.1 ;
      RECT 448.95 178.8 480 178.95 ;
      RECT 449.1 178.65 480 178.8 ;
      RECT 449.25 178.5 480 178.65 ;
      RECT 449.4 178.35 480 178.5 ;
      RECT 449.55 178.2 480 178.35 ;
      RECT 449.7 178.05 480 178.2 ;
      RECT 411.75 216 480 216.15 ;
      RECT 411.9 215.85 480 216 ;
      RECT 412.05 215.7 480 215.85 ;
      RECT 412.2 215.55 480 215.7 ;
      RECT 412.35 215.4 480 215.55 ;
      RECT 412.5 215.25 480 215.4 ;
      RECT 412.65 215.1 480 215.25 ;
      RECT 412.8 214.95 480 215.1 ;
      RECT 412.95 214.8 480 214.95 ;
      RECT 413.1 214.65 480 214.8 ;
      RECT 413.25 214.5 480 214.65 ;
      RECT 413.4 214.35 480 214.5 ;
      RECT 413.55 214.2 480 214.35 ;
      RECT 413.7 214.05 480 214.2 ;
      RECT 413.85 213.9 480 214.05 ;
      RECT 414.0 213.75 480 213.9 ;
      RECT 414.15 213.6 480 213.75 ;
      RECT 414.3 213.45 480 213.6 ;
      RECT 414.45 213.3 480 213.45 ;
      RECT 414.6 213.15 480 213.3 ;
      RECT 414.75 213 480 213.15 ;
      RECT 414.9 212.85 480 213 ;
      RECT 415.05 212.7 480 212.85 ;
      RECT 415.2 212.55 480 212.7 ;
      RECT 415.35 212.4 480 212.55 ;
      RECT 415.5 212.25 480 212.4 ;
      RECT 415.65 212.1 480 212.25 ;
      RECT 415.8 211.95 480 212.1 ;
      RECT 415.95 211.8 480 211.95 ;
      RECT 416.1 211.65 480 211.8 ;
      RECT 416.25 211.5 480 211.65 ;
      RECT 416.4 211.35 480 211.5 ;
      RECT 416.55 211.2 480 211.35 ;
      RECT 416.7 211.05 480 211.2 ;
      RECT 416.85 210.9 480 211.05 ;
      RECT 417.0 210.75 480 210.9 ;
      RECT 417.15 210.6 480 210.75 ;
      RECT 417.3 210.45 480 210.6 ;
      RECT 417.45 210.3 480 210.45 ;
      RECT 417.6 210.15 480 210.3 ;
      RECT 417.75 210 480 210.15 ;
      RECT 417.9 209.85 480 210 ;
      RECT 418.05 209.7 480 209.85 ;
      RECT 418.2 209.55 480 209.7 ;
      RECT 418.35 209.4 480 209.55 ;
      RECT 418.5 209.25 480 209.4 ;
      RECT 418.65 209.1 480 209.25 ;
      RECT 418.8 208.95 480 209.1 ;
      RECT 418.95 208.8 480 208.95 ;
      RECT 419.1 208.65 480 208.8 ;
      RECT 419.25 208.5 480 208.65 ;
      RECT 419.4 208.35 480 208.5 ;
      RECT 419.55 208.2 480 208.35 ;
      RECT 419.7 208.05 480 208.2 ;
      RECT 419.85 207.9 480 208.05 ;
      RECT 420.0 207.75 480 207.9 ;
      RECT 420.15 207.6 480 207.75 ;
      RECT 420.3 207.45 480 207.6 ;
      RECT 420.45 207.3 480 207.45 ;
      RECT 420.6 207.15 480 207.3 ;
      RECT 420.75 207 480 207.15 ;
      RECT 420.9 206.85 480 207 ;
      RECT 421.05 206.7 480 206.85 ;
      RECT 421.2 206.55 480 206.7 ;
      RECT 421.35 206.4 480 206.55 ;
      RECT 421.5 206.25 480 206.4 ;
      RECT 421.65 206.1 480 206.25 ;
      RECT 421.8 205.95 480 206.1 ;
      RECT 421.95 205.8 480 205.95 ;
      RECT 422.1 205.65 480 205.8 ;
      RECT 422.25 205.5 480 205.65 ;
      RECT 422.4 205.35 480 205.5 ;
      RECT 422.55 205.2 480 205.35 ;
      RECT 422.7 205.05 480 205.2 ;
      RECT 422.85 204.9 480 205.05 ;
      RECT 423.0 204.75 480 204.9 ;
      RECT 423.15 204.6 480 204.75 ;
      RECT 423.3 204.45 480 204.6 ;
      RECT 423.45 204.3 480 204.45 ;
      RECT 423.6 204.15 480 204.3 ;
      RECT 423.75 204 480 204.15 ;
      RECT 423.9 203.85 480 204 ;
      RECT 424.05 203.7 480 203.85 ;
      RECT 424.2 203.55 480 203.7 ;
      RECT 424.35 203.4 480 203.55 ;
      RECT 424.5 203.25 480 203.4 ;
      RECT 424.65 203.1 480 203.25 ;
      RECT 424.8 202.95 480 203.1 ;
      RECT 424.95 202.8 480 202.95 ;
      RECT 425.1 202.65 480 202.8 ;
      RECT 425.25 202.5 480 202.65 ;
      RECT 425.4 202.35 480 202.5 ;
      RECT 425.55 202.2 480 202.35 ;
      RECT 425.7 202.05 480 202.2 ;
      RECT 425.85 201.9 480 202.05 ;
      RECT 426.0 201.75 480 201.9 ;
      RECT 426.15 201.6 480 201.75 ;
      RECT 426.3 201.45 480 201.6 ;
      RECT 426.45 201.3 480 201.45 ;
      RECT 426.6 201.15 480 201.3 ;
      RECT 426.75 201 480 201.15 ;
      RECT 426.9 200.85 480 201 ;
      RECT 427.05 200.7 480 200.85 ;
      RECT 427.2 200.55 480 200.7 ;
      RECT 427.35 200.4 480 200.55 ;
      RECT 427.5 200.25 480 200.4 ;
      RECT 427.65 200.1 480 200.25 ;
      RECT 427.8 199.95 480 200.1 ;
      RECT 427.95 199.8 480 199.95 ;
      RECT 428.1 199.65 480 199.8 ;
      RECT 428.25 199.5 480 199.65 ;
      RECT 428.4 199.35 480 199.5 ;
      RECT 428.55 199.2 480 199.35 ;
      RECT 428.7 199.05 480 199.2 ;
      RECT 428.85 198.9 480 199.05 ;
      RECT 429.0 198.75 480 198.9 ;
      RECT 429.15 198.6 480 198.75 ;
      RECT 429.3 198.45 480 198.6 ;
      RECT 429.45 198.3 480 198.45 ;
      RECT 429.6 198.15 480 198.3 ;
      RECT 429.75 198 480 198.15 ;
      RECT 429.9 197.85 480 198 ;
      RECT 430.05 197.7 480 197.85 ;
      RECT 430.2 197.55 480 197.7 ;
      RECT 430.35 197.4 480 197.55 ;
      RECT 430.5 197.25 480 197.4 ;
      RECT 430.65 197.1 480 197.25 ;
      RECT 473.235 154.515 480 154.665 ;
      RECT 473.385 154.365 480 154.515 ;
      RECT 473.535 154.215 480 154.365 ;
      RECT 473.685 154.065 480 154.215 ;
      RECT 473.835 153.915 480 154.065 ;
      RECT 473.985 153.765 480 153.915 ;
      RECT 474.135 153.615 480 153.765 ;
      RECT 474.285 153.465 480 153.615 ;
      RECT 474.435 153.315 480 153.465 ;
      RECT 474.585 153.165 480 153.315 ;
      RECT 474.735 153.015 480 153.165 ;
      RECT 474.885 152.865 480 153.015 ;
      RECT 475.035 152.715 480 152.865 ;
      RECT 475.185 152.565 480 152.715 ;
      RECT 475.335 152.415 480 152.565 ;
      RECT 475.485 152.265 480 152.415 ;
      RECT 475.635 152.115 480 152.265 ;
      RECT 475.785 151.965 480 152.115 ;
      RECT 475.935 151.815 480 151.965 ;
      RECT 476.085 151.665 480 151.815 ;
      RECT 476.235 151.515 480 151.665 ;
      RECT 476.385 151.365 480 151.515 ;
      RECT 476.535 151.215 480 151.365 ;
      RECT 476.685 151.065 480 151.215 ;
      RECT 476.835 150.915 480 151.065 ;
      RECT 476.985 150.765 480 150.915 ;
      RECT 477.135 150.615 480 150.765 ;
      RECT 477.285 150.465 480 150.615 ;
      RECT 477.435 150.315 480 150.465 ;
      RECT 477.585 150.165 480 150.315 ;
      RECT 477.735 150.015 480 150.165 ;
      RECT 477.885 149.865 480 150.015 ;
      RECT 478.035 149.715 480 149.865 ;
      RECT 478.185 149.565 480 149.715 ;
      RECT 478.335 149.415 480 149.565 ;
      RECT 478.485 149.265 480 149.415 ;
      RECT 478.635 149.115 480 149.265 ;
      RECT 458.13 73.015 480 73.055 ;
      RECT 458.17 73.055 480 73.095 ;
      RECT 458.175 73.095 480 73.1 ;
      RECT 398.7 229.05 480 229.1 ;
      RECT 398.85 228.9 480 229.05 ;
      RECT 399.0 228.75 480 228.9 ;
      RECT 399.15 228.6 480 228.75 ;
      RECT 399.3 228.45 480 228.6 ;
      RECT 399.45 228.3 480 228.45 ;
      RECT 399.6 228.15 480 228.3 ;
      RECT 399.75 228 480 228.15 ;
      RECT 399.9 227.85 480 228 ;
      RECT 400.05 227.7 480 227.85 ;
      RECT 400.2 227.55 480 227.7 ;
      RECT 400.35 227.4 480 227.55 ;
      RECT 400.5 227.25 480 227.4 ;
      RECT 400.65 227.1 480 227.25 ;
      RECT 400.8 226.95 480 227.1 ;
      RECT 400.95 226.8 480 226.95 ;
      RECT 401.1 226.65 480 226.8 ;
      RECT 401.25 226.5 480 226.65 ;
      RECT 401.4 226.35 480 226.5 ;
      RECT 401.55 226.2 480 226.35 ;
      RECT 401.7 226.05 480 226.2 ;
      RECT 401.85 225.9 480 226.05 ;
      RECT 402.0 225.75 480 225.9 ;
      RECT 402.15 225.6 480 225.75 ;
      RECT 402.3 225.45 480 225.6 ;
      RECT 402.45 225.3 480 225.45 ;
      RECT 402.6 225.15 480 225.3 ;
      RECT 402.75 225 480 225.15 ;
      RECT 402.9 224.85 480 225 ;
      RECT 403.05 224.7 480 224.85 ;
      RECT 403.2 224.55 480 224.7 ;
      RECT 403.35 224.4 480 224.55 ;
      RECT 403.5 224.25 480 224.4 ;
      RECT 403.65 224.1 480 224.25 ;
      RECT 403.8 223.95 480 224.1 ;
      RECT 403.95 223.8 480 223.95 ;
      RECT 404.1 223.65 480 223.8 ;
      RECT 404.25 223.5 480 223.65 ;
      RECT 404.4 223.35 480 223.5 ;
      RECT 404.55 223.2 480 223.35 ;
      RECT 404.7 223.05 480 223.2 ;
      RECT 404.85 222.9 480 223.05 ;
      RECT 405.0 222.75 480 222.9 ;
      RECT 405.15 222.6 480 222.75 ;
      RECT 405.3 222.45 480 222.6 ;
      RECT 405.45 222.3 480 222.45 ;
      RECT 405.6 222.15 480 222.3 ;
      RECT 405.75 222 480 222.15 ;
      RECT 405.9 221.85 480 222 ;
      RECT 406.05 221.7 480 221.85 ;
      RECT 406.2 221.55 480 221.7 ;
      RECT 406.35 221.4 480 221.55 ;
      RECT 406.5 221.25 480 221.4 ;
      RECT 406.65 221.1 480 221.25 ;
      RECT 406.8 220.95 480 221.1 ;
      RECT 406.95 220.8 480 220.95 ;
      RECT 407.1 220.65 480 220.8 ;
      RECT 407.25 220.5 480 220.65 ;
      RECT 407.4 220.35 480 220.5 ;
      RECT 407.55 220.2 480 220.35 ;
      RECT 407.7 220.05 480 220.2 ;
      RECT 407.85 219.9 480 220.05 ;
      RECT 408.0 219.75 480 219.9 ;
      RECT 408.15 219.6 480 219.75 ;
      RECT 408.3 219.45 480 219.6 ;
      RECT 408.45 219.3 480 219.45 ;
      RECT 408.6 219.15 480 219.3 ;
      RECT 408.75 219 480 219.15 ;
      RECT 408.9 218.85 480 219 ;
      RECT 409.05 218.7 480 218.85 ;
      RECT 409.2 218.55 480 218.7 ;
      RECT 409.35 218.4 480 218.55 ;
      RECT 409.5 218.25 480 218.4 ;
      RECT 409.65 218.1 480 218.25 ;
      RECT 409.8 217.95 480 218.1 ;
      RECT 409.95 217.8 480 217.95 ;
      RECT 410.1 217.65 480 217.8 ;
      RECT 410.25 217.5 480 217.65 ;
      RECT 410.4 217.35 480 217.5 ;
      RECT 410.55 217.2 480 217.35 ;
      RECT 410.7 217.05 480 217.2 ;
      RECT 410.85 216.9 480 217.05 ;
      RECT 411.0 216.75 480 216.9 ;
      RECT 411.15 216.6 480 216.75 ;
      RECT 411.3 216.45 480 216.6 ;
      RECT 411.45 216.3 480 216.45 ;
      RECT 411.6 216.15 480 216.3 ;
      RECT 454.185 173.565 480 173.715 ;
      RECT 454.335 173.415 480 173.565 ;
      RECT 454.485 173.265 480 173.415 ;
      RECT 454.635 173.115 480 173.265 ;
      RECT 454.785 172.965 480 173.115 ;
      RECT 454.935 172.815 480 172.965 ;
      RECT 455.085 172.665 480 172.815 ;
      RECT 455.235 172.515 480 172.665 ;
      RECT 455.385 172.365 480 172.515 ;
      RECT 455.535 172.215 480 172.365 ;
      RECT 455.685 172.065 480 172.215 ;
      RECT 455.835 171.915 480 172.065 ;
      RECT 455.985 171.765 480 171.915 ;
      RECT 456.135 171.615 480 171.765 ;
      RECT 456.285 171.465 480 171.615 ;
      RECT 456.435 171.315 480 171.465 ;
      RECT 456.585 171.165 480 171.315 ;
      RECT 456.735 171.015 480 171.165 ;
      RECT 456.885 170.865 480 171.015 ;
      RECT 457.035 170.715 480 170.865 ;
      RECT 457.185 170.565 480 170.715 ;
      RECT 457.335 170.415 480 170.565 ;
      RECT 457.485 170.265 480 170.415 ;
      RECT 457.635 170.115 480 170.265 ;
      RECT 457.785 169.965 480 170.115 ;
      RECT 457.935 169.815 480 169.965 ;
      RECT 458.085 169.665 480 169.815 ;
      RECT 458.235 169.515 480 169.665 ;
      RECT 458.385 169.365 480 169.515 ;
      RECT 458.535 169.215 480 169.365 ;
      RECT 458.685 169.065 480 169.215 ;
      RECT 458.835 168.915 480 169.065 ;
      RECT 458.985 168.765 480 168.915 ;
      RECT 459.135 168.615 480 168.765 ;
      RECT 459.285 168.465 480 168.615 ;
      RECT 459.435 168.315 480 168.465 ;
      RECT 459.585 168.165 480 168.315 ;
      RECT 459.735 168.015 480 168.165 ;
      RECT 459.885 167.865 480 168.015 ;
      RECT 460.035 167.715 480 167.865 ;
      RECT 460.185 167.565 480 167.715 ;
      RECT 460.335 167.415 480 167.565 ;
      RECT 460.485 167.265 480 167.415 ;
      RECT 460.635 167.115 480 167.265 ;
      RECT 460.785 166.965 480 167.115 ;
      RECT 460.935 166.815 480 166.965 ;
      RECT 461.085 166.665 480 166.815 ;
      RECT 461.235 166.515 480 166.665 ;
      RECT 461.385 166.365 480 166.515 ;
      RECT 461.535 166.215 480 166.365 ;
      RECT 461.685 166.065 480 166.215 ;
      RECT 461.835 165.915 480 166.065 ;
      RECT 461.985 165.765 480 165.915 ;
      RECT 462.135 165.615 480 165.765 ;
      RECT 462.285 165.465 480 165.615 ;
      RECT 462.435 165.315 480 165.465 ;
      RECT 462.585 165.165 480 165.315 ;
      RECT 462.735 165.015 480 165.165 ;
      RECT 462.885 164.865 480 165.015 ;
      RECT 463.035 164.715 480 164.865 ;
      RECT 463.185 164.565 480 164.715 ;
      RECT 463.335 164.415 480 164.565 ;
      RECT 463.485 164.265 480 164.415 ;
      RECT 463.635 164.115 480 164.265 ;
      RECT 463.785 163.965 480 164.115 ;
      RECT 463.935 163.815 480 163.965 ;
      RECT 464.085 163.665 480 163.815 ;
      RECT 464.235 163.515 480 163.665 ;
      RECT 464.385 163.365 480 163.515 ;
      RECT 464.535 163.215 480 163.365 ;
      RECT 464.685 163.065 480 163.215 ;
      RECT 464.835 162.915 480 163.065 ;
      RECT 464.985 162.765 480 162.915 ;
      RECT 465.135 162.615 480 162.765 ;
      RECT 465.285 162.465 480 162.615 ;
      RECT 465.435 162.315 480 162.465 ;
      RECT 465.585 162.165 480 162.315 ;
      RECT 465.735 162.015 480 162.165 ;
      RECT 465.885 161.865 480 162.015 ;
      RECT 466.035 161.715 480 161.865 ;
      RECT 466.185 161.565 480 161.715 ;
      RECT 466.335 161.415 480 161.565 ;
      RECT 466.485 161.265 480 161.415 ;
      RECT 466.635 161.115 480 161.265 ;
      RECT 466.785 160.965 480 161.115 ;
      RECT 466.935 160.815 480 160.965 ;
      RECT 467.085 160.665 480 160.815 ;
      RECT 467.235 160.515 480 160.665 ;
      RECT 467.385 160.365 480 160.515 ;
      RECT 467.535 160.215 480 160.365 ;
      RECT 467.685 160.065 480 160.215 ;
      RECT 467.835 159.915 480 160.065 ;
      RECT 467.985 159.765 480 159.915 ;
      RECT 468.135 159.615 480 159.765 ;
      RECT 468.285 159.465 480 159.615 ;
      RECT 468.435 159.315 480 159.465 ;
      RECT 468.585 159.165 480 159.315 ;
      RECT 468.735 159.015 480 159.165 ;
      RECT 468.885 158.865 480 159.015 ;
      RECT 469.035 158.715 480 158.865 ;
      RECT 469.185 158.565 480 158.715 ;
      RECT 469.335 158.415 480 158.565 ;
      RECT 469.485 158.265 480 158.415 ;
      RECT 469.635 158.115 480 158.265 ;
      RECT 469.785 157.965 480 158.115 ;
      RECT 469.935 157.815 480 157.965 ;
      RECT 470.085 157.665 480 157.815 ;
      RECT 470.235 157.515 480 157.665 ;
      RECT 470.385 157.365 480 157.515 ;
      RECT 470.535 157.215 480 157.365 ;
      RECT 470.685 157.065 480 157.215 ;
      RECT 470.835 156.915 480 157.065 ;
      RECT 470.985 156.765 480 156.915 ;
      RECT 471.135 156.615 480 156.765 ;
      RECT 471.285 156.465 480 156.615 ;
      RECT 471.435 156.315 480 156.465 ;
      RECT 471.585 156.165 480 156.315 ;
      RECT 471.735 156.015 480 156.165 ;
      RECT 471.885 155.865 480 156.015 ;
      RECT 472.035 155.715 480 155.865 ;
      RECT 472.185 155.565 480 155.715 ;
      RECT 472.335 155.415 480 155.565 ;
      RECT 472.485 155.265 480 155.415 ;
      RECT 472.635 155.115 480 155.265 ;
      RECT 472.785 154.965 480 155.115 ;
      RECT 472.935 154.815 480 154.965 ;
      RECT 473.085 154.665 480 154.815 ;
      RECT 435.135 192.615 480 192.765 ;
      RECT 435.285 192.465 480 192.615 ;
      RECT 435.435 192.315 480 192.465 ;
      RECT 435.585 192.165 480 192.315 ;
      RECT 435.735 192.015 480 192.165 ;
      RECT 435.885 191.865 480 192.015 ;
      RECT 436.035 191.715 480 191.865 ;
      RECT 436.185 191.565 480 191.715 ;
      RECT 436.335 191.415 480 191.565 ;
      RECT 436.485 191.265 480 191.415 ;
      RECT 436.635 191.115 480 191.265 ;
      RECT 436.785 190.965 480 191.115 ;
      RECT 436.935 190.815 480 190.965 ;
      RECT 437.085 190.665 480 190.815 ;
      RECT 437.235 190.515 480 190.665 ;
      RECT 437.385 190.365 480 190.515 ;
      RECT 437.535 190.215 480 190.365 ;
      RECT 437.685 190.065 480 190.215 ;
      RECT 437.835 189.915 480 190.065 ;
      RECT 437.985 189.765 480 189.915 ;
      RECT 438.135 189.615 480 189.765 ;
      RECT 438.285 189.465 480 189.615 ;
      RECT 438.435 189.315 480 189.465 ;
      RECT 438.585 189.165 480 189.315 ;
      RECT 438.735 189.015 480 189.165 ;
      RECT 438.885 188.865 480 189.015 ;
      RECT 439.035 188.715 480 188.865 ;
      RECT 439.185 188.565 480 188.715 ;
      RECT 439.335 188.415 480 188.565 ;
      RECT 439.485 188.265 480 188.415 ;
      RECT 439.635 188.115 480 188.265 ;
      RECT 439.785 187.965 480 188.115 ;
      RECT 439.935 187.815 480 187.965 ;
      RECT 440.085 187.665 480 187.815 ;
      RECT 440.235 187.515 480 187.665 ;
      RECT 440.385 187.365 480 187.515 ;
      RECT 440.535 187.215 480 187.365 ;
      RECT 440.685 187.065 480 187.215 ;
      RECT 440.835 186.915 480 187.065 ;
      RECT 440.985 186.765 480 186.915 ;
      RECT 441.135 186.615 480 186.765 ;
      RECT 441.285 186.465 480 186.615 ;
      RECT 441.435 186.315 480 186.465 ;
      RECT 441.585 186.165 480 186.315 ;
      RECT 441.735 186.015 480 186.165 ;
      RECT 441.885 185.865 480 186.015 ;
      RECT 442.035 185.715 480 185.865 ;
      RECT 442.185 185.565 480 185.715 ;
      RECT 442.335 185.415 480 185.565 ;
      RECT 442.485 185.265 480 185.415 ;
      RECT 442.635 185.115 480 185.265 ;
      RECT 442.785 184.965 480 185.115 ;
      RECT 442.935 184.815 480 184.965 ;
      RECT 443.085 184.665 480 184.815 ;
      RECT 443.235 184.515 480 184.665 ;
      RECT 443.385 184.365 480 184.515 ;
      RECT 443.535 184.215 480 184.365 ;
      RECT 443.685 184.065 480 184.215 ;
      RECT 443.835 183.915 480 184.065 ;
      RECT 443.985 183.765 480 183.915 ;
      RECT 444.135 183.615 480 183.765 ;
      RECT 444.285 183.465 480 183.615 ;
      RECT 444.435 183.315 480 183.465 ;
      RECT 444.585 183.165 480 183.315 ;
      RECT 444.735 183.015 480 183.165 ;
      RECT 444.885 182.865 480 183.015 ;
      RECT 445.035 182.715 480 182.865 ;
      RECT 445.185 182.565 480 182.715 ;
      RECT 445.335 182.415 480 182.565 ;
      RECT 445.485 182.265 480 182.415 ;
      RECT 445.635 182.115 480 182.265 ;
      RECT 445.785 181.965 480 182.115 ;
      RECT 445.935 181.815 480 181.965 ;
      RECT 446.085 181.665 480 181.815 ;
      RECT 446.235 181.515 480 181.665 ;
      RECT 446.385 181.365 480 181.515 ;
      RECT 446.535 181.215 480 181.365 ;
      RECT 446.685 181.065 480 181.215 ;
      RECT 446.835 180.915 480 181.065 ;
      RECT 446.985 180.765 480 180.915 ;
      RECT 447.135 180.615 480 180.765 ;
      RECT 447.285 180.465 480 180.615 ;
      RECT 447.435 180.315 480 180.465 ;
      RECT 447.585 180.165 480 180.315 ;
      RECT 447.735 180.015 480 180.165 ;
      RECT 447.885 179.865 480 180.015 ;
      RECT 448.035 179.715 480 179.865 ;
      RECT 448.185 179.565 480 179.715 ;
      RECT 448.335 179.415 480 179.565 ;
      RECT 448.485 179.265 480 179.415 ;
      RECT 448.635 179.115 480 179.265 ;
      RECT 448.785 178.965 480 179.115 ;
      RECT 448.935 178.815 480 178.965 ;
      RECT 449.085 178.665 480 178.815 ;
      RECT 449.235 178.515 480 178.665 ;
      RECT 449.385 178.365 480 178.515 ;
      RECT 449.535 178.215 480 178.365 ;
      RECT 449.685 178.065 480 178.215 ;
      RECT 449.835 177.915 480 178.065 ;
      RECT 449.985 177.765 480 177.915 ;
      RECT 450.135 177.615 480 177.765 ;
      RECT 450.285 177.465 480 177.615 ;
      RECT 450.435 177.315 480 177.465 ;
      RECT 450.585 177.165 480 177.315 ;
      RECT 450.735 177.015 480 177.165 ;
      RECT 450.885 176.865 480 177.015 ;
      RECT 451.035 176.715 480 176.865 ;
      RECT 451.185 176.565 480 176.715 ;
      RECT 451.335 176.415 480 176.565 ;
      RECT 451.485 176.265 480 176.415 ;
      RECT 451.635 176.115 480 176.265 ;
      RECT 451.785 175.965 480 176.115 ;
      RECT 451.935 175.815 480 175.965 ;
      RECT 452.085 175.665 480 175.815 ;
      RECT 452.235 175.515 480 175.665 ;
      RECT 452.385 175.365 480 175.515 ;
      RECT 452.535 175.215 480 175.365 ;
      RECT 452.685 175.065 480 175.215 ;
      RECT 452.835 174.915 480 175.065 ;
      RECT 452.985 174.765 480 174.915 ;
      RECT 453.135 174.615 480 174.765 ;
      RECT 453.285 174.465 480 174.615 ;
      RECT 453.435 174.315 480 174.465 ;
      RECT 453.585 174.165 480 174.315 ;
      RECT 453.735 174.015 480 174.165 ;
      RECT 453.885 173.865 480 174.015 ;
      RECT 454.035 173.715 480 173.865 ;
      RECT 416.085 211.665 480 211.815 ;
      RECT 416.235 211.515 480 211.665 ;
      RECT 416.385 211.365 480 211.515 ;
      RECT 416.535 211.215 480 211.365 ;
      RECT 416.685 211.065 480 211.215 ;
      RECT 416.835 210.915 480 211.065 ;
      RECT 416.985 210.765 480 210.915 ;
      RECT 417.135 210.615 480 210.765 ;
      RECT 417.285 210.465 480 210.615 ;
      RECT 417.435 210.315 480 210.465 ;
      RECT 417.585 210.165 480 210.315 ;
      RECT 417.735 210.015 480 210.165 ;
      RECT 417.885 209.865 480 210.015 ;
      RECT 418.035 209.715 480 209.865 ;
      RECT 418.185 209.565 480 209.715 ;
      RECT 418.335 209.415 480 209.565 ;
      RECT 418.485 209.265 480 209.415 ;
      RECT 418.635 209.115 480 209.265 ;
      RECT 418.785 208.965 480 209.115 ;
      RECT 418.935 208.815 480 208.965 ;
      RECT 419.085 208.665 480 208.815 ;
      RECT 419.235 208.515 480 208.665 ;
      RECT 419.385 208.365 480 208.515 ;
      RECT 419.535 208.215 480 208.365 ;
      RECT 419.685 208.065 480 208.215 ;
      RECT 419.835 207.915 480 208.065 ;
      RECT 419.985 207.765 480 207.915 ;
      RECT 420.135 207.615 480 207.765 ;
      RECT 420.285 207.465 480 207.615 ;
      RECT 420.435 207.315 480 207.465 ;
      RECT 420.585 207.165 480 207.315 ;
      RECT 420.735 207.015 480 207.165 ;
      RECT 420.885 206.865 480 207.015 ;
      RECT 421.035 206.715 480 206.865 ;
      RECT 421.185 206.565 480 206.715 ;
      RECT 421.335 206.415 480 206.565 ;
      RECT 421.485 206.265 480 206.415 ;
      RECT 421.635 206.115 480 206.265 ;
      RECT 421.785 205.965 480 206.115 ;
      RECT 421.935 205.815 480 205.965 ;
      RECT 422.085 205.665 480 205.815 ;
      RECT 422.235 205.515 480 205.665 ;
      RECT 422.385 205.365 480 205.515 ;
      RECT 422.535 205.215 480 205.365 ;
      RECT 422.685 205.065 480 205.215 ;
      RECT 422.835 204.915 480 205.065 ;
      RECT 422.985 204.765 480 204.915 ;
      RECT 423.135 204.615 480 204.765 ;
      RECT 423.285 204.465 480 204.615 ;
      RECT 423.435 204.315 480 204.465 ;
      RECT 423.585 204.165 480 204.315 ;
      RECT 423.735 204.015 480 204.165 ;
      RECT 423.885 203.865 480 204.015 ;
      RECT 424.035 203.715 480 203.865 ;
      RECT 424.185 203.565 480 203.715 ;
      RECT 424.335 203.415 480 203.565 ;
      RECT 424.485 203.265 480 203.415 ;
      RECT 424.635 203.115 480 203.265 ;
      RECT 424.785 202.965 480 203.115 ;
      RECT 424.935 202.815 480 202.965 ;
      RECT 425.085 202.665 480 202.815 ;
      RECT 425.235 202.515 480 202.665 ;
      RECT 425.385 202.365 480 202.515 ;
      RECT 425.535 202.215 480 202.365 ;
      RECT 425.685 202.065 480 202.215 ;
      RECT 425.835 201.915 480 202.065 ;
      RECT 425.985 201.765 480 201.915 ;
      RECT 426.135 201.615 480 201.765 ;
      RECT 426.285 201.465 480 201.615 ;
      RECT 426.435 201.315 480 201.465 ;
      RECT 426.585 201.165 480 201.315 ;
      RECT 426.735 201.015 480 201.165 ;
      RECT 426.885 200.865 480 201.015 ;
      RECT 427.035 200.715 480 200.865 ;
      RECT 427.185 200.565 480 200.715 ;
      RECT 427.335 200.415 480 200.565 ;
      RECT 427.485 200.265 480 200.415 ;
      RECT 427.635 200.115 480 200.265 ;
      RECT 427.785 199.965 480 200.115 ;
      RECT 427.935 199.815 480 199.965 ;
      RECT 428.085 199.665 480 199.815 ;
      RECT 428.235 199.515 480 199.665 ;
      RECT 428.385 199.365 480 199.515 ;
      RECT 428.535 199.215 480 199.365 ;
      RECT 428.685 199.065 480 199.215 ;
      RECT 428.835 198.915 480 199.065 ;
      RECT 428.985 198.765 480 198.915 ;
      RECT 429.135 198.615 480 198.765 ;
      RECT 429.285 198.465 480 198.615 ;
      RECT 429.435 198.315 480 198.465 ;
      RECT 429.585 198.165 480 198.315 ;
      RECT 429.735 198.015 480 198.165 ;
      RECT 429.885 197.865 480 198.015 ;
      RECT 430.035 197.715 480 197.865 ;
      RECT 430.185 197.565 480 197.715 ;
      RECT 430.335 197.415 480 197.565 ;
      RECT 430.485 197.265 480 197.415 ;
      RECT 430.635 197.115 480 197.265 ;
      RECT 430.785 196.965 480 197.115 ;
      RECT 430.935 196.815 480 196.965 ;
      RECT 431.085 196.665 480 196.815 ;
      RECT 431.235 196.515 480 196.665 ;
      RECT 431.385 196.365 480 196.515 ;
      RECT 431.535 196.215 480 196.365 ;
      RECT 431.685 196.065 480 196.215 ;
      RECT 431.835 195.915 480 196.065 ;
      RECT 431.985 195.765 480 195.915 ;
      RECT 432.135 195.615 480 195.765 ;
      RECT 432.285 195.465 480 195.615 ;
      RECT 432.435 195.315 480 195.465 ;
      RECT 432.585 195.165 480 195.315 ;
      RECT 432.735 195.015 480 195.165 ;
      RECT 432.885 194.865 480 195.015 ;
      RECT 433.035 194.715 480 194.865 ;
      RECT 433.185 194.565 480 194.715 ;
      RECT 433.335 194.415 480 194.565 ;
      RECT 433.485 194.265 480 194.415 ;
      RECT 433.635 194.115 480 194.265 ;
      RECT 433.785 193.965 480 194.115 ;
      RECT 433.935 193.815 480 193.965 ;
      RECT 434.085 193.665 480 193.815 ;
      RECT 434.235 193.515 480 193.665 ;
      RECT 434.385 193.365 480 193.515 ;
      RECT 434.535 193.215 480 193.365 ;
      RECT 434.685 193.065 480 193.215 ;
      RECT 434.835 192.915 480 193.065 ;
      RECT 434.985 192.765 480 192.915 ;
      RECT 58.895 201.635 390.125 201.785 ;
      RECT 59.045 201.785 389.975 201.935 ;
      RECT 59.195 201.935 389.825 202.085 ;
      RECT 59.345 202.085 389.675 202.235 ;
      RECT 59.495 202.235 389.525 202.385 ;
      RECT 59.645 202.385 389.375 202.535 ;
      RECT 59.795 202.535 389.225 202.685 ;
      RECT 59.945 202.685 389.075 202.835 ;
      RECT 60.095 202.835 388.925 202.985 ;
      RECT 60.245 202.985 388.775 203.135 ;
      RECT 60.395 203.135 388.625 203.285 ;
      RECT 60.545 203.285 388.475 203.435 ;
      RECT 60.695 203.435 388.325 203.585 ;
      RECT 60.845 203.585 388.175 203.735 ;
      RECT 60.995 203.735 388.025 203.885 ;
      RECT 61.145 203.885 387.875 204.035 ;
      RECT 61.215 204.035 387.805 204.105 ;
      RECT 399.585 228.165 480 228.3 ;
      RECT 399.735 228.015 480 228.165 ;
      RECT 399.885 227.865 480 228.015 ;
      RECT 400.035 227.715 480 227.865 ;
      RECT 400.185 227.565 480 227.715 ;
      RECT 400.335 227.415 480 227.565 ;
      RECT 400.485 227.265 480 227.415 ;
      RECT 400.635 227.115 480 227.265 ;
      RECT 400.785 226.965 480 227.115 ;
      RECT 400.935 226.815 480 226.965 ;
      RECT 401.085 226.665 480 226.815 ;
      RECT 401.235 226.515 480 226.665 ;
      RECT 401.385 226.365 480 226.515 ;
      RECT 401.535 226.215 480 226.365 ;
      RECT 401.685 226.065 480 226.215 ;
      RECT 401.835 225.915 480 226.065 ;
      RECT 401.985 225.765 480 225.915 ;
      RECT 402.135 225.615 480 225.765 ;
      RECT 402.285 225.465 480 225.615 ;
      RECT 402.435 225.315 480 225.465 ;
      RECT 402.585 225.165 480 225.315 ;
      RECT 402.735 225.015 480 225.165 ;
      RECT 402.885 224.865 480 225.015 ;
      RECT 403.035 224.715 480 224.865 ;
      RECT 403.185 224.565 480 224.715 ;
      RECT 403.335 224.415 480 224.565 ;
      RECT 403.485 224.265 480 224.415 ;
      RECT 403.635 224.115 480 224.265 ;
      RECT 403.785 223.965 480 224.115 ;
      RECT 403.935 223.815 480 223.965 ;
      RECT 404.085 223.665 480 223.815 ;
      RECT 404.235 223.515 480 223.665 ;
      RECT 404.385 223.365 480 223.515 ;
      RECT 404.535 223.215 480 223.365 ;
      RECT 404.685 223.065 480 223.215 ;
      RECT 404.835 222.915 480 223.065 ;
      RECT 404.985 222.765 480 222.915 ;
      RECT 405.135 222.615 480 222.765 ;
      RECT 405.285 222.465 480 222.615 ;
      RECT 405.435 222.315 480 222.465 ;
      RECT 405.585 222.165 480 222.315 ;
      RECT 405.735 222.015 480 222.165 ;
      RECT 405.885 221.865 480 222.015 ;
      RECT 406.035 221.715 480 221.865 ;
      RECT 406.185 221.565 480 221.715 ;
      RECT 406.335 221.415 480 221.565 ;
      RECT 406.485 221.265 480 221.415 ;
      RECT 406.635 221.115 480 221.265 ;
      RECT 406.785 220.965 480 221.115 ;
      RECT 406.935 220.815 480 220.965 ;
      RECT 407.085 220.665 480 220.815 ;
      RECT 407.235 220.515 480 220.665 ;
      RECT 407.385 220.365 480 220.515 ;
      RECT 407.535 220.215 480 220.365 ;
      RECT 407.685 220.065 480 220.215 ;
      RECT 407.835 219.915 480 220.065 ;
      RECT 407.985 219.765 480 219.915 ;
      RECT 408.135 219.615 480 219.765 ;
      RECT 408.285 219.465 480 219.615 ;
      RECT 408.435 219.315 480 219.465 ;
      RECT 408.585 219.165 480 219.315 ;
      RECT 408.735 219.015 480 219.165 ;
      RECT 408.885 218.865 480 219.015 ;
      RECT 409.035 218.715 480 218.865 ;
      RECT 409.185 218.565 480 218.715 ;
      RECT 409.335 218.415 480 218.565 ;
      RECT 409.485 218.265 480 218.415 ;
      RECT 409.635 218.115 480 218.265 ;
      RECT 409.785 217.965 480 218.115 ;
      RECT 409.935 217.815 480 217.965 ;
      RECT 410.085 217.665 480 217.815 ;
      RECT 410.235 217.515 480 217.665 ;
      RECT 410.385 217.365 480 217.515 ;
      RECT 410.535 217.215 480 217.365 ;
      RECT 410.685 217.065 480 217.215 ;
      RECT 410.835 216.915 480 217.065 ;
      RECT 410.985 216.765 480 216.915 ;
      RECT 411.135 216.615 480 216.765 ;
      RECT 411.285 216.465 480 216.615 ;
      RECT 411.435 216.315 480 216.465 ;
      RECT 411.585 216.165 480 216.315 ;
      RECT 411.735 216.015 480 216.165 ;
      RECT 411.885 215.865 480 216.015 ;
      RECT 412.035 215.715 480 215.865 ;
      RECT 412.185 215.565 480 215.715 ;
      RECT 412.335 215.415 480 215.565 ;
      RECT 412.485 215.265 480 215.415 ;
      RECT 412.635 215.115 480 215.265 ;
      RECT 412.785 214.965 480 215.115 ;
      RECT 412.935 214.815 480 214.965 ;
      RECT 413.085 214.665 480 214.815 ;
      RECT 413.235 214.515 480 214.665 ;
      RECT 413.385 214.365 480 214.515 ;
      RECT 413.535 214.215 480 214.365 ;
      RECT 413.685 214.065 480 214.215 ;
      RECT 413.835 213.915 480 214.065 ;
      RECT 413.985 213.765 480 213.915 ;
      RECT 414.135 213.615 480 213.765 ;
      RECT 414.285 213.465 480 213.615 ;
      RECT 414.435 213.315 480 213.465 ;
      RECT 414.585 213.165 480 213.315 ;
      RECT 414.735 213.015 480 213.165 ;
      RECT 414.885 212.865 480 213.015 ;
      RECT 415.035 212.715 480 212.865 ;
      RECT 415.185 212.565 480 212.715 ;
      RECT 415.335 212.415 480 212.565 ;
      RECT 415.485 212.265 480 212.415 ;
      RECT 415.635 212.115 480 212.265 ;
      RECT 415.785 211.965 480 212.115 ;
      RECT 415.935 211.815 480 211.965 ;
      RECT 54.545 163.615 428.145 163.765 ;
      RECT 54.545 163.465 428.295 163.615 ;
      RECT 54.545 163.315 428.445 163.465 ;
      RECT 54.545 163.165 428.595 163.315 ;
      RECT 54.545 163.015 428.745 163.165 ;
      RECT 54.545 162.865 428.895 163.015 ;
      RECT 54.545 162.715 429.045 162.865 ;
      RECT 54.545 162.565 429.195 162.715 ;
      RECT 54.545 162.415 429.345 162.565 ;
      RECT 54.545 162.265 429.495 162.415 ;
      RECT 54.545 162.115 429.645 162.265 ;
      RECT 54.545 161.965 429.795 162.115 ;
      RECT 54.545 161.815 429.945 161.965 ;
      RECT 54.545 161.665 430.095 161.815 ;
      RECT 54.545 161.515 430.245 161.665 ;
      RECT 54.545 161.365 430.395 161.515 ;
      RECT 54.545 161.215 430.545 161.365 ;
      RECT 54.545 161.065 430.695 161.215 ;
      RECT 54.545 160.915 430.845 161.065 ;
      RECT 54.545 160.765 430.995 160.915 ;
      RECT 54.545 160.615 431.145 160.765 ;
      RECT 54.545 160.465 431.295 160.615 ;
      RECT 54.545 160.315 431.445 160.465 ;
      RECT 54.545 160.165 431.595 160.315 ;
      RECT 54.545 160.015 431.745 160.165 ;
      RECT 54.545 159.865 431.895 160.015 ;
      RECT 54.545 159.715 432.045 159.865 ;
      RECT 54.545 159.565 432.195 159.715 ;
      RECT 54.545 159.415 432.345 159.565 ;
      RECT 54.545 159.265 432.495 159.415 ;
      RECT 54.545 159.115 432.645 159.265 ;
      RECT 54.545 158.965 432.795 159.115 ;
      RECT 54.545 158.815 432.945 158.965 ;
      RECT 54.545 158.665 433.095 158.815 ;
      RECT 54.545 158.515 433.245 158.665 ;
      RECT 54.545 158.365 433.395 158.515 ;
      RECT 54.545 158.215 433.545 158.365 ;
      RECT 54.545 158.065 433.695 158.215 ;
      RECT 54.545 157.915 433.845 158.065 ;
      RECT 54.545 157.765 433.995 157.915 ;
      RECT 54.545 157.615 434.145 157.765 ;
      RECT 54.545 157.465 434.295 157.615 ;
      RECT 54.545 157.315 434.445 157.465 ;
      RECT 54.545 157.165 434.595 157.315 ;
      RECT 54.545 157.015 434.745 157.165 ;
      RECT 54.545 156.865 434.895 157.015 ;
      RECT 54.545 156.715 435.045 156.865 ;
      RECT 54.545 156.565 435.195 156.715 ;
      RECT 54.545 156.415 435.345 156.565 ;
      RECT 54.545 156.265 435.495 156.415 ;
      RECT 54.545 156.115 435.645 156.265 ;
      RECT 54.545 155.965 435.795 156.115 ;
      RECT 54.545 155.815 435.945 155.965 ;
      RECT 54.545 155.665 436.095 155.815 ;
      RECT 54.545 155.515 436.245 155.665 ;
      RECT 54.545 155.365 436.395 155.515 ;
      RECT 54.545 155.215 436.545 155.365 ;
      RECT 54.545 155.065 436.695 155.215 ;
      RECT 54.545 154.915 436.845 155.065 ;
      RECT 54.545 154.765 436.995 154.915 ;
      RECT 54.545 154.615 437.145 154.765 ;
      RECT 54.545 154.465 437.295 154.615 ;
      RECT 54.545 154.315 437.445 154.465 ;
      RECT 54.545 154.165 437.595 154.315 ;
      RECT 54.545 154.015 437.745 154.165 ;
      RECT 54.545 153.865 437.895 154.015 ;
      RECT 54.545 153.715 438.045 153.865 ;
      RECT 54.545 153.565 438.195 153.715 ;
      RECT 54.545 153.415 438.345 153.565 ;
      RECT 54.545 153.265 438.495 153.415 ;
      RECT 54.545 153.115 438.645 153.265 ;
      RECT 54.545 152.965 438.795 153.115 ;
      RECT 54.545 152.815 438.945 152.965 ;
      RECT 54.545 152.665 439.095 152.815 ;
      RECT 54.545 152.515 439.245 152.665 ;
      RECT 54.545 152.365 439.395 152.515 ;
      RECT 54.545 152.215 439.545 152.365 ;
      RECT 54.545 152.065 439.695 152.215 ;
      RECT 54.545 151.915 439.845 152.065 ;
      RECT 54.545 151.765 439.995 151.915 ;
      RECT 54.545 151.615 440.145 151.765 ;
      RECT 54.545 151.465 440.295 151.615 ;
      RECT 54.545 151.315 440.445 151.465 ;
      RECT 54.545 151.165 440.595 151.315 ;
      RECT 54.545 151.015 440.745 151.165 ;
      RECT 54.545 150.865 440.895 151.015 ;
      RECT 54.545 150.715 441.045 150.865 ;
      RECT 54.545 150.565 441.195 150.715 ;
      RECT 54.545 150.415 441.345 150.565 ;
      RECT 54.545 150.265 441.495 150.415 ;
      RECT 54.545 150.115 441.645 150.265 ;
      RECT 54.545 149.965 441.795 150.115 ;
      RECT 54.545 149.815 441.945 149.965 ;
      RECT 54.545 149.665 442.095 149.815 ;
      RECT 54.545 149.515 442.245 149.665 ;
      RECT 54.545 149.365 442.395 149.515 ;
      RECT 54.545 149.215 442.545 149.365 ;
      RECT 54.545 149.065 442.695 149.215 ;
      RECT 54.545 148.915 442.845 149.065 ;
      RECT 54.695 197.435 394.325 197.585 ;
      RECT 54.845 197.585 394.175 197.735 ;
      RECT 54.995 197.735 394.025 197.885 ;
      RECT 55.145 197.885 393.875 198.035 ;
      RECT 55.295 198.035 393.725 198.185 ;
      RECT 55.445 198.185 393.575 198.335 ;
      RECT 55.595 198.335 393.425 198.485 ;
      RECT 55.745 198.485 393.275 198.635 ;
      RECT 55.895 198.635 393.125 198.785 ;
      RECT 56.045 198.785 392.975 198.935 ;
      RECT 56.195 198.935 392.825 199.085 ;
      RECT 56.345 199.085 392.675 199.235 ;
      RECT 56.495 199.235 392.525 199.385 ;
      RECT 56.645 199.385 392.375 199.535 ;
      RECT 56.795 199.535 392.225 199.685 ;
      RECT 56.945 199.685 392.075 199.835 ;
      RECT 57.095 199.835 391.925 199.985 ;
      RECT 57.245 199.985 391.775 200.135 ;
      RECT 57.395 200.135 391.625 200.285 ;
      RECT 57.545 200.285 391.475 200.435 ;
      RECT 57.695 200.435 391.325 200.585 ;
      RECT 57.845 200.585 391.175 200.735 ;
      RECT 57.995 200.735 391.025 200.885 ;
      RECT 58.145 200.885 390.875 201.035 ;
      RECT 58.295 201.035 390.725 201.185 ;
      RECT 58.445 201.185 390.575 201.335 ;
      RECT 58.595 201.335 390.425 201.485 ;
      RECT 58.745 201.485 390.275 201.635 ;
      RECT 54.545 182.665 409.095 182.815 ;
      RECT 54.545 182.515 409.245 182.665 ;
      RECT 54.545 182.365 409.395 182.515 ;
      RECT 54.545 182.215 409.545 182.365 ;
      RECT 54.545 182.065 409.695 182.215 ;
      RECT 54.545 181.915 409.845 182.065 ;
      RECT 54.545 181.765 409.995 181.915 ;
      RECT 54.545 181.615 410.145 181.765 ;
      RECT 54.545 181.465 410.295 181.615 ;
      RECT 54.545 181.315 410.445 181.465 ;
      RECT 54.545 181.165 410.595 181.315 ;
      RECT 54.545 181.015 410.745 181.165 ;
      RECT 54.545 180.865 410.895 181.015 ;
      RECT 54.545 180.715 411.045 180.865 ;
      RECT 54.545 180.565 411.195 180.715 ;
      RECT 54.545 180.415 411.345 180.565 ;
      RECT 54.545 180.265 411.495 180.415 ;
      RECT 54.545 180.115 411.645 180.265 ;
      RECT 54.545 179.965 411.795 180.115 ;
      RECT 54.545 179.815 411.945 179.965 ;
      RECT 54.545 179.665 412.095 179.815 ;
      RECT 54.545 179.515 412.245 179.665 ;
      RECT 54.545 179.365 412.395 179.515 ;
      RECT 54.545 179.215 412.545 179.365 ;
      RECT 54.545 179.065 412.695 179.215 ;
      RECT 54.545 178.915 412.845 179.065 ;
      RECT 54.545 178.765 412.995 178.915 ;
      RECT 54.545 178.615 413.145 178.765 ;
      RECT 54.545 178.465 413.295 178.615 ;
      RECT 54.545 178.315 413.445 178.465 ;
      RECT 54.545 178.165 413.595 178.315 ;
      RECT 54.545 178.015 413.745 178.165 ;
      RECT 54.545 177.865 413.895 178.015 ;
      RECT 54.545 177.715 414.045 177.865 ;
      RECT 54.545 177.565 414.195 177.715 ;
      RECT 54.545 177.415 414.345 177.565 ;
      RECT 54.545 177.265 414.495 177.415 ;
      RECT 54.545 177.115 414.645 177.265 ;
      RECT 54.545 176.965 414.795 177.115 ;
      RECT 54.545 176.815 414.945 176.965 ;
      RECT 54.545 176.665 415.095 176.815 ;
      RECT 54.545 176.515 415.245 176.665 ;
      RECT 54.545 176.365 415.395 176.515 ;
      RECT 54.545 176.215 415.545 176.365 ;
      RECT 54.545 176.065 415.695 176.215 ;
      RECT 54.545 175.915 415.845 176.065 ;
      RECT 54.545 175.765 415.995 175.915 ;
      RECT 54.545 175.615 416.145 175.765 ;
      RECT 54.545 175.465 416.295 175.615 ;
      RECT 54.545 175.315 416.445 175.465 ;
      RECT 54.545 175.165 416.595 175.315 ;
      RECT 54.545 175.015 416.745 175.165 ;
      RECT 54.545 174.865 416.895 175.015 ;
      RECT 54.545 174.715 417.045 174.865 ;
      RECT 54.545 174.565 417.195 174.715 ;
      RECT 54.545 174.415 417.345 174.565 ;
      RECT 54.545 174.265 417.495 174.415 ;
      RECT 54.545 174.115 417.645 174.265 ;
      RECT 54.545 173.965 417.795 174.115 ;
      RECT 54.545 173.815 417.945 173.965 ;
      RECT 54.545 173.665 418.095 173.815 ;
      RECT 54.545 173.515 418.245 173.665 ;
      RECT 54.545 173.365 418.395 173.515 ;
      RECT 54.545 173.215 418.545 173.365 ;
      RECT 54.545 173.065 418.695 173.215 ;
      RECT 54.545 172.915 418.845 173.065 ;
      RECT 54.545 172.765 418.995 172.915 ;
      RECT 54.545 172.615 419.145 172.765 ;
      RECT 54.545 172.465 419.295 172.615 ;
      RECT 54.545 172.315 419.445 172.465 ;
      RECT 54.545 172.165 419.595 172.315 ;
      RECT 54.545 172.015 419.745 172.165 ;
      RECT 54.545 171.865 419.895 172.015 ;
      RECT 54.545 171.715 420.045 171.865 ;
      RECT 54.545 171.565 420.195 171.715 ;
      RECT 54.545 171.415 420.345 171.565 ;
      RECT 54.545 171.265 420.495 171.415 ;
      RECT 54.545 171.115 420.645 171.265 ;
      RECT 54.545 170.965 420.795 171.115 ;
      RECT 54.545 170.815 420.945 170.965 ;
      RECT 54.545 170.665 421.095 170.815 ;
      RECT 54.545 170.515 421.245 170.665 ;
      RECT 54.545 170.365 421.395 170.515 ;
      RECT 54.545 170.215 421.545 170.365 ;
      RECT 54.545 170.065 421.695 170.215 ;
      RECT 54.545 169.915 421.845 170.065 ;
      RECT 54.545 169.765 421.995 169.915 ;
      RECT 54.545 169.615 422.145 169.765 ;
      RECT 54.545 169.465 422.295 169.615 ;
      RECT 54.545 169.315 422.445 169.465 ;
      RECT 54.545 169.165 422.595 169.315 ;
      RECT 54.545 169.015 422.745 169.165 ;
      RECT 54.545 168.865 422.895 169.015 ;
      RECT 54.545 168.715 423.045 168.865 ;
      RECT 54.545 168.565 423.195 168.715 ;
      RECT 54.545 168.415 423.345 168.565 ;
      RECT 54.545 168.265 423.495 168.415 ;
      RECT 54.545 168.115 423.645 168.265 ;
      RECT 54.545 167.965 423.795 168.115 ;
      RECT 54.545 167.815 423.945 167.965 ;
      RECT 54.545 167.665 424.095 167.815 ;
      RECT 54.545 167.515 424.245 167.665 ;
      RECT 54.545 167.365 424.395 167.515 ;
      RECT 54.545 167.215 424.545 167.365 ;
      RECT 54.545 167.065 424.695 167.215 ;
      RECT 54.545 166.915 424.845 167.065 ;
      RECT 54.545 166.765 424.995 166.915 ;
      RECT 54.545 166.615 425.145 166.765 ;
      RECT 54.545 166.465 425.295 166.615 ;
      RECT 54.545 166.315 425.445 166.465 ;
      RECT 54.545 166.165 425.595 166.315 ;
      RECT 54.545 166.015 425.745 166.165 ;
      RECT 54.545 165.865 425.895 166.015 ;
      RECT 54.545 165.715 426.045 165.865 ;
      RECT 54.545 165.565 426.195 165.715 ;
      RECT 54.545 165.415 426.345 165.565 ;
      RECT 54.545 165.265 426.495 165.415 ;
      RECT 54.545 165.115 426.645 165.265 ;
      RECT 54.545 164.965 426.795 165.115 ;
      RECT 54.545 164.815 426.945 164.965 ;
      RECT 54.545 164.665 427.095 164.815 ;
      RECT 54.545 164.515 427.245 164.665 ;
      RECT 54.545 164.365 427.395 164.515 ;
      RECT 54.545 164.215 427.545 164.365 ;
      RECT 54.545 164.065 427.695 164.215 ;
      RECT 54.545 163.915 427.845 164.065 ;
      RECT 54.545 163.765 427.995 163.915 ;
      RECT 33.68 127.9 463.86 128.05 ;
      RECT 33.53 127.75 464.01 127.9 ;
      RECT 33.38 127.6 464.16 127.75 ;
      RECT 33.23 127.45 464.31 127.6 ;
      RECT 33.08 127.3 464.46 127.45 ;
      RECT 32.93 127.15 464.61 127.3 ;
      RECT 32.78 127 464.76 127.15 ;
      RECT 32.63 126.85 464.91 127 ;
      RECT 32.48 126.7 465.06 126.85 ;
      RECT 32.33 126.55 465.21 126.7 ;
      RECT 32.18 126.4 465.36 126.55 ;
      RECT 32.03 126.25 465.51 126.4 ;
      RECT 31.88 126.1 465.66 126.25 ;
      RECT 31.73 125.95 465.81 126.1 ;
      RECT 31.58 125.8 465.96 125.95 ;
      RECT 31.43 125.65 466.11 125.8 ;
      RECT 31.28 125.5 466.26 125.65 ;
      RECT 31.13 125.35 466.41 125.5 ;
      RECT 30.98 125.2 466.56 125.35 ;
      RECT 30.83 125.05 466.71 125.2 ;
      RECT 30.68 124.9 466.86 125.05 ;
      RECT 30.53 124.75 467.01 124.9 ;
      RECT 30.38 124.6 467.16 124.75 ;
      RECT 30.23 124.45 467.31 124.6 ;
      RECT 30.08 124.3 467.46 124.45 ;
      RECT 29.93 124.15 467.61 124.3 ;
      RECT 29.78 124 467.76 124.15 ;
      RECT 29.63 123.85 467.91 124 ;
      RECT 29.48 123.7 468.06 123.85 ;
      RECT 54.545 197.365 394.475 197.435 ;
      RECT 54.545 197.215 394.545 197.365 ;
      RECT 54.545 197.065 394.695 197.215 ;
      RECT 54.545 196.915 394.845 197.065 ;
      RECT 54.545 196.765 394.995 196.915 ;
      RECT 54.545 196.615 395.145 196.765 ;
      RECT 54.545 196.465 395.295 196.615 ;
      RECT 54.545 196.315 395.445 196.465 ;
      RECT 54.545 196.165 395.595 196.315 ;
      RECT 54.545 196.015 395.745 196.165 ;
      RECT 54.545 195.865 395.895 196.015 ;
      RECT 54.545 195.715 396.045 195.865 ;
      RECT 54.545 195.565 396.195 195.715 ;
      RECT 54.545 195.415 396.345 195.565 ;
      RECT 54.545 195.265 396.495 195.415 ;
      RECT 54.545 195.115 396.645 195.265 ;
      RECT 54.545 194.965 396.795 195.115 ;
      RECT 54.545 194.815 396.945 194.965 ;
      RECT 54.545 194.665 397.095 194.815 ;
      RECT 54.545 194.515 397.245 194.665 ;
      RECT 54.545 194.365 397.395 194.515 ;
      RECT 54.545 194.215 397.545 194.365 ;
      RECT 54.545 194.065 397.695 194.215 ;
      RECT 54.545 193.915 397.845 194.065 ;
      RECT 54.545 193.765 397.995 193.915 ;
      RECT 54.545 193.615 398.145 193.765 ;
      RECT 54.545 193.465 398.295 193.615 ;
      RECT 54.545 193.315 398.445 193.465 ;
      RECT 54.545 193.165 398.595 193.315 ;
      RECT 54.545 193.015 398.745 193.165 ;
      RECT 54.545 192.865 398.895 193.015 ;
      RECT 54.545 192.715 399.045 192.865 ;
      RECT 54.545 192.565 399.195 192.715 ;
      RECT 54.545 192.415 399.345 192.565 ;
      RECT 54.545 192.265 399.495 192.415 ;
      RECT 54.545 192.115 399.645 192.265 ;
      RECT 54.545 191.965 399.795 192.115 ;
      RECT 54.545 191.815 399.945 191.965 ;
      RECT 54.545 191.665 400.095 191.815 ;
      RECT 54.545 191.515 400.245 191.665 ;
      RECT 54.545 191.365 400.395 191.515 ;
      RECT 54.545 191.215 400.545 191.365 ;
      RECT 54.545 191.065 400.695 191.215 ;
      RECT 54.545 190.915 400.845 191.065 ;
      RECT 54.545 190.765 400.995 190.915 ;
      RECT 54.545 190.615 401.145 190.765 ;
      RECT 54.545 190.465 401.295 190.615 ;
      RECT 54.545 190.315 401.445 190.465 ;
      RECT 54.545 190.165 401.595 190.315 ;
      RECT 54.545 190.015 401.745 190.165 ;
      RECT 54.545 189.865 401.895 190.015 ;
      RECT 54.545 189.715 402.045 189.865 ;
      RECT 54.545 189.565 402.195 189.715 ;
      RECT 54.545 189.415 402.345 189.565 ;
      RECT 54.545 189.265 402.495 189.415 ;
      RECT 54.545 189.115 402.645 189.265 ;
      RECT 54.545 188.965 402.795 189.115 ;
      RECT 54.545 188.815 402.945 188.965 ;
      RECT 54.545 188.665 403.095 188.815 ;
      RECT 54.545 188.515 403.245 188.665 ;
      RECT 54.545 188.365 403.395 188.515 ;
      RECT 54.545 188.215 403.545 188.365 ;
      RECT 54.545 188.065 403.695 188.215 ;
      RECT 54.545 187.915 403.845 188.065 ;
      RECT 54.545 187.765 403.995 187.915 ;
      RECT 54.545 187.615 404.145 187.765 ;
      RECT 54.545 187.465 404.295 187.615 ;
      RECT 54.545 187.315 404.445 187.465 ;
      RECT 54.545 187.165 404.595 187.315 ;
      RECT 54.545 187.015 404.745 187.165 ;
      RECT 54.545 186.865 404.895 187.015 ;
      RECT 54.545 186.715 405.045 186.865 ;
      RECT 54.545 186.565 405.195 186.715 ;
      RECT 54.545 186.415 405.345 186.565 ;
      RECT 54.545 186.265 405.495 186.415 ;
      RECT 54.545 186.115 405.645 186.265 ;
      RECT 54.545 185.965 405.795 186.115 ;
      RECT 54.545 185.815 405.945 185.965 ;
      RECT 54.545 185.665 406.095 185.815 ;
      RECT 54.545 185.515 406.245 185.665 ;
      RECT 54.545 185.365 406.395 185.515 ;
      RECT 54.545 185.215 406.545 185.365 ;
      RECT 54.545 185.065 406.695 185.215 ;
      RECT 54.545 184.915 406.845 185.065 ;
      RECT 54.545 184.765 406.995 184.915 ;
      RECT 54.545 184.615 407.145 184.765 ;
      RECT 54.545 184.465 407.295 184.615 ;
      RECT 54.545 184.315 407.445 184.465 ;
      RECT 54.545 184.165 407.595 184.315 ;
      RECT 54.545 184.015 407.745 184.165 ;
      RECT 54.545 183.865 407.895 184.015 ;
      RECT 54.545 183.715 408.045 183.865 ;
      RECT 54.545 183.565 408.195 183.715 ;
      RECT 54.545 183.415 408.345 183.565 ;
      RECT 54.545 183.265 408.495 183.415 ;
      RECT 54.545 183.115 408.645 183.265 ;
      RECT 54.545 182.965 408.795 183.115 ;
      RECT 54.545 182.815 408.945 182.965 ;
      RECT 52.73 146.95 444.81 147.1 ;
      RECT 52.58 146.8 444.96 146.95 ;
      RECT 52.43 146.65 445.11 146.8 ;
      RECT 52.28 146.5 445.26 146.65 ;
      RECT 52.13 146.35 445.41 146.5 ;
      RECT 51.98 146.2 445.56 146.35 ;
      RECT 51.83 146.05 445.71 146.2 ;
      RECT 51.68 145.9 445.86 146.05 ;
      RECT 51.53 145.75 446.01 145.9 ;
      RECT 51.38 145.6 446.16 145.75 ;
      RECT 51.23 145.45 446.31 145.6 ;
      RECT 51.08 145.3 446.46 145.45 ;
      RECT 50.93 145.15 446.61 145.3 ;
      RECT 50.78 145 446.76 145.15 ;
      RECT 50.63 144.85 446.91 145 ;
      RECT 50.48 144.7 447.06 144.85 ;
      RECT 50.33 144.55 447.21 144.7 ;
      RECT 50.18 144.4 447.36 144.55 ;
      RECT 50.03 144.25 447.51 144.4 ;
      RECT 49.88 144.1 447.66 144.25 ;
      RECT 49.73 143.95 447.81 144.1 ;
      RECT 49.58 143.8 447.96 143.95 ;
      RECT 49.43 143.65 448.11 143.8 ;
      RECT 49.28 143.5 448.26 143.65 ;
      RECT 49.13 143.35 448.41 143.5 ;
      RECT 48.98 143.2 448.56 143.35 ;
      RECT 48.83 143.05 448.71 143.2 ;
      RECT 48.68 142.9 448.86 143.05 ;
      RECT 48.53 142.75 449.01 142.9 ;
      RECT 48.38 142.6 449.16 142.75 ;
      RECT 48.23 142.45 449.31 142.6 ;
      RECT 48.08 142.3 449.46 142.45 ;
      RECT 47.93 142.15 449.61 142.3 ;
      RECT 47.78 142 449.76 142.15 ;
      RECT 47.63 141.85 449.91 142 ;
      RECT 47.48 141.7 450.06 141.85 ;
      RECT 47.33 141.55 450.21 141.7 ;
      RECT 47.18 141.4 450.36 141.55 ;
      RECT 47.03 141.25 450.51 141.4 ;
      RECT 46.88 141.1 450.66 141.25 ;
      RECT 46.73 140.95 450.81 141.1 ;
      RECT 46.58 140.8 450.96 140.95 ;
      RECT 46.43 140.65 451.11 140.8 ;
      RECT 46.28 140.5 451.26 140.65 ;
      RECT 46.13 140.35 451.41 140.5 ;
      RECT 45.98 140.2 451.56 140.35 ;
      RECT 45.83 140.05 451.71 140.2 ;
      RECT 45.68 139.9 451.86 140.05 ;
      RECT 45.53 139.75 452.01 139.9 ;
      RECT 45.38 139.6 452.16 139.75 ;
      RECT 45.23 139.45 452.31 139.6 ;
      RECT 45.08 139.3 452.46 139.45 ;
      RECT 44.93 139.15 452.61 139.3 ;
      RECT 44.78 139 452.76 139.15 ;
      RECT 44.63 138.85 452.91 139 ;
      RECT 44.48 138.7 453.06 138.85 ;
      RECT 44.33 138.55 453.21 138.7 ;
      RECT 44.18 138.4 453.36 138.55 ;
      RECT 44.03 138.25 453.51 138.4 ;
      RECT 43.88 138.1 453.66 138.25 ;
      RECT 43.73 137.95 453.81 138.1 ;
      RECT 43.58 137.8 453.96 137.95 ;
      RECT 43.43 137.65 454.11 137.8 ;
      RECT 43.28 137.5 454.26 137.65 ;
      RECT 43.13 137.35 454.41 137.5 ;
      RECT 42.98 137.2 454.56 137.35 ;
      RECT 42.83 137.05 454.71 137.2 ;
      RECT 42.68 136.9 454.86 137.05 ;
      RECT 42.53 136.75 455.01 136.9 ;
      RECT 42.38 136.6 455.16 136.75 ;
      RECT 42.23 136.45 455.31 136.6 ;
      RECT 42.08 136.3 455.46 136.45 ;
      RECT 41.93 136.15 455.61 136.3 ;
      RECT 41.78 136 455.76 136.15 ;
      RECT 41.63 135.85 455.91 136 ;
      RECT 41.48 135.7 456.06 135.85 ;
      RECT 41.33 135.55 456.21 135.7 ;
      RECT 41.18 135.4 456.36 135.55 ;
      RECT 41.03 135.25 456.51 135.4 ;
      RECT 40.88 135.1 456.66 135.25 ;
      RECT 40.73 134.95 456.81 135.1 ;
      RECT 40.58 134.8 456.96 134.95 ;
      RECT 40.43 134.65 457.11 134.8 ;
      RECT 40.28 134.5 457.26 134.65 ;
      RECT 40.13 134.35 457.41 134.5 ;
      RECT 39.98 134.2 457.56 134.35 ;
      RECT 39.83 134.05 457.71 134.2 ;
      RECT 39.68 133.9 457.86 134.05 ;
      RECT 39.53 133.75 458.01 133.9 ;
      RECT 39.38 133.6 458.16 133.75 ;
      RECT 39.23 133.45 458.31 133.6 ;
      RECT 39.08 133.3 458.46 133.45 ;
      RECT 38.93 133.15 458.61 133.3 ;
      RECT 38.78 133 458.76 133.15 ;
      RECT 38.63 132.85 458.91 133 ;
      RECT 38.48 132.7 459.06 132.85 ;
      RECT 38.33 132.55 459.21 132.7 ;
      RECT 38.18 132.4 459.36 132.55 ;
      RECT 38.03 132.25 459.51 132.4 ;
      RECT 37.88 132.1 459.66 132.25 ;
      RECT 37.73 131.95 459.81 132.1 ;
      RECT 37.58 131.8 459.96 131.95 ;
      RECT 37.43 131.65 460.11 131.8 ;
      RECT 37.28 131.5 460.26 131.65 ;
      RECT 37.13 131.35 460.41 131.5 ;
      RECT 36.98 131.2 460.56 131.35 ;
      RECT 36.83 131.05 460.71 131.2 ;
      RECT 36.68 130.9 460.86 131.05 ;
      RECT 36.53 130.75 461.01 130.9 ;
      RECT 36.38 130.6 461.16 130.75 ;
      RECT 36.23 130.45 461.31 130.6 ;
      RECT 36.08 130.3 461.46 130.45 ;
      RECT 35.93 130.15 461.61 130.3 ;
      RECT 35.78 130 461.76 130.15 ;
      RECT 35.63 129.85 461.91 130 ;
      RECT 35.48 129.7 462.06 129.85 ;
      RECT 35.33 129.55 462.21 129.7 ;
      RECT 35.18 129.4 462.36 129.55 ;
      RECT 35.03 129.25 462.51 129.4 ;
      RECT 34.88 129.1 462.66 129.25 ;
      RECT 34.73 128.95 462.81 129.1 ;
      RECT 34.58 128.8 462.96 128.95 ;
      RECT 34.43 128.65 463.11 128.8 ;
      RECT 34.28 128.5 463.26 128.65 ;
      RECT 34.13 128.35 463.41 128.5 ;
      RECT 33.98 128.2 463.56 128.35 ;
      RECT 33.83 128.05 463.71 128.2 ;
      RECT 0 61.6 480 62.2 ;
      RECT 0 67.65 480 68.25 ;
      RECT 0 72.5 480 73.015 ;
      RECT 0 116.8 480 117.4 ;
      RECT 0 122.65 480 123.35 ;
      RECT 0 0 480 55.35 ;
      RECT 0 84.6 480 85.2 ;
      RECT 0 89.45 480 90.05 ;
      RECT 0 94.3 480 94.9 ;
      RECT 0 100.35 480 101.05 ;
      RECT 0 78.55 480 79.15 ;
      RECT 0 110.85 480 111.55 ;
      RECT 0 159.55 28.86 207.49 ;
      RECT 0 73.015 9.46 73.055 ;
      RECT 0 73.055 9.42 73.095 ;
      RECT 0 73.095 9.415 73.1 ;
      RECT 29.03 123.35 468.51 123.4 ;
      RECT 29.08 123.4 468.46 123.45 ;
      RECT 29.33 123.45 468.335 123.575 ;
      RECT 29.33 123.575 468.21 123.7 ;
      RECT 54.545 148.9 442.995 148.915 ;
      RECT 54.53 148.75 443.01 148.9 ;
      RECT 54.38 148.6 443.16 148.75 ;
      RECT 54.23 148.45 443.31 148.6 ;
      RECT 54.08 148.3 443.46 148.45 ;
      RECT 53.93 148.15 443.61 148.3 ;
      RECT 53.78 148 443.76 148.15 ;
      RECT 53.63 147.85 443.91 148 ;
      RECT 53.48 147.7 444.06 147.85 ;
      RECT 53.33 147.55 444.21 147.7 ;
      RECT 53.18 147.4 444.36 147.55 ;
      RECT 53.03 147.25 444.51 147.4 ;
      RECT 52.88 147.1 444.66 147.25 ;
    LAYER met1 ;
      RECT 0 0 480 253.715 ;
    LAYER met3 ;
      RECT 0 0 480 253.715 ;
  END
END sky130_fd_io__top_sio_macro

END LIBRARY
