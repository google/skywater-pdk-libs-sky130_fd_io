# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__overlay_gpiov2
  CLASS COVER ;
  FOREIGN sky130_fd_io__overlay_gpiov2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  80.00000 BY  200.0000 ;
  SYMMETRY X Y ;
  PIN AMUXBUS_A
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 80.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 80.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN PAD
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 11.100000 104.395000 73.800000 166.960000 ;
    END
  END PAD
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 80.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 80.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 80.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 80.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 80.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 80.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 80.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 80.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 80.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 80.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met4 ;
      RECT 0.000000  2.035000 80.000000  47.965000 ;
      RECT 0.000000 51.745000 80.000000  52.725000 ;
      RECT 0.000000 56.505000 80.000000 200.000000 ;
    LAYER met5 ;
      RECT  0.000000  19.885000 80.000000  24.335000 ;
      RECT  0.000000  36.835000 80.000000  40.085000 ;
      RECT  0.000000  96.585000 80.000000 102.795000 ;
      RECT  0.000000 102.795000  9.500000 168.560000 ;
      RECT  0.000000 168.560000 80.000000 200.000000 ;
      RECT 75.400000 102.795000 80.000000 168.560000 ;
  END
END sky130_fd_io__overlay_gpiov2
END LIBRARY
