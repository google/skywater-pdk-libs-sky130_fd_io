# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sky130_fd_io__top_analog_pad
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 75 BY 198 ;
  SYMMETRY R90 ;

  PIN pad_core
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 9.43 146.45 10.39 169.22 ;
        RECT 4.955 141.825 10.39 141.975 ;
        RECT 5.105 141.975 10.39 142.125 ;
        RECT 5.255 142.125 10.39 142.275 ;
        RECT 5.405 142.275 10.39 142.425 ;
        RECT 5.555 142.425 10.39 142.575 ;
        RECT 5.705 142.575 10.39 142.725 ;
        RECT 5.855 142.725 10.39 142.875 ;
        RECT 6.005 142.875 10.39 143.025 ;
        RECT 6.155 143.025 10.39 143.175 ;
        RECT 6.305 143.175 10.39 143.325 ;
        RECT 6.455 143.325 10.39 143.475 ;
        RECT 6.605 143.475 10.39 143.625 ;
        RECT 6.755 143.625 10.39 143.775 ;
        RECT 6.905 143.775 10.39 143.925 ;
        RECT 7.055 143.925 10.39 144.075 ;
        RECT 7.205 144.075 10.39 144.225 ;
        RECT 7.355 144.225 10.39 144.375 ;
        RECT 7.505 144.375 10.39 144.525 ;
        RECT 7.655 144.525 10.39 144.675 ;
        RECT 7.805 144.675 10.39 144.825 ;
        RECT 7.955 144.825 10.39 144.975 ;
        RECT 8.105 144.975 10.39 145.125 ;
        RECT 8.255 145.125 10.39 145.275 ;
        RECT 8.405 145.275 10.39 145.425 ;
        RECT 8.555 145.425 10.39 145.575 ;
        RECT 8.705 145.575 10.39 145.725 ;
        RECT 8.855 145.725 10.39 145.875 ;
        RECT 9.005 145.875 10.39 146.025 ;
        RECT 9.155 146.025 10.39 146.175 ;
        RECT 9.305 146.175 10.39 146.325 ;
        RECT 9.43 146.325 10.39 146.45 ;
        RECT 24.31 135.995 25.27 171.125 ;
        RECT 34.23 135.975 35.21 171.125 ;
        RECT 29.27 135.975 30.23 171.125 ;
        RECT 39.19 135.975 40.15 171.125 ;
        RECT 19.35 135.975 20.31 171.125 ;
        RECT 34.23 135.505 35.53 135.655 ;
        RECT 34.23 135.655 35.38 135.805 ;
        RECT 34.23 135.805 35.23 135.955 ;
        RECT 34.23 135.955 35.21 135.975 ;
        RECT 39.19 135.505 40.47 135.655 ;
        RECT 39.19 135.655 40.32 135.805 ;
        RECT 39.19 135.805 40.17 135.955 ;
        RECT 39.19 135.955 40.15 135.975 ;
        RECT 24.31 135.505 25.61 135.655 ;
        RECT 24.31 135.655 25.46 135.805 ;
        RECT 24.31 135.805 25.31 135.955 ;
        RECT 24.31 135.955 25.27 135.995 ;
        RECT 19.35 135.505 20.63 135.655 ;
        RECT 19.35 135.655 20.48 135.805 ;
        RECT 19.35 135.805 20.33 135.955 ;
        RECT 19.35 135.955 20.31 135.975 ;
        RECT 29.27 135.485 30.57 135.635 ;
        RECT 29.27 135.635 30.42 135.785 ;
        RECT 29.27 135.785 30.27 135.935 ;
        RECT 29.27 135.935 30.23 135.975 ;
        RECT 14.39 134.76 15.35 171.125 ;
        RECT 14.39 134.29 15.67 134.44 ;
        RECT 14.39 134.44 15.52 134.59 ;
        RECT 14.39 134.59 15.37 134.74 ;
        RECT 14.39 134.74 15.35 134.76 ;
        RECT 34.23 133.65 35.68 135.505 ;
        RECT 24.31 133.65 25.76 135.505 ;
        RECT 39.19 133.63 40.62 135.505 ;
        RECT 29.27 133.63 30.72 135.485 ;
        RECT 19.35 133.63 20.78 135.505 ;
        RECT 34.72 133.16 35.68 133.31 ;
        RECT 34.57 133.31 35.68 133.46 ;
        RECT 34.42 133.46 35.68 133.61 ;
        RECT 34.27 133.61 35.68 133.65 ;
        RECT 24.8 133.16 25.76 133.31 ;
        RECT 24.65 133.31 25.76 133.46 ;
        RECT 24.5 133.46 25.76 133.61 ;
        RECT 24.35 133.61 25.76 133.65 ;
        RECT 29.76 133.14 30.72 133.29 ;
        RECT 29.61 133.29 30.72 133.44 ;
        RECT 29.46 133.44 30.72 133.59 ;
        RECT 29.31 133.59 30.72 133.63 ;
        RECT 39.7 133.12 40.62 133.27 ;
        RECT 39.55 133.27 40.62 133.42 ;
        RECT 39.4 133.42 40.62 133.57 ;
        RECT 39.25 133.57 40.62 133.63 ;
        RECT 19.86 133.12 20.78 133.27 ;
        RECT 19.71 133.27 20.78 133.42 ;
        RECT 19.56 133.42 20.78 133.57 ;
        RECT 19.41 133.57 20.78 133.63 ;
        RECT 14.39 132.83 15.82 134.29 ;
        RECT 14.9 132.32 15.82 132.47 ;
        RECT 14.75 132.47 15.82 132.62 ;
        RECT 14.6 132.62 15.82 132.77 ;
        RECT 14.45 132.77 15.82 132.83 ;
        RECT 4.805 124.405 10.39 141.825 ;
        RECT 6.125 123.09 10.39 123.24 ;
        RECT 5.975 123.24 10.39 123.39 ;
        RECT 5.825 123.39 10.39 123.54 ;
        RECT 5.675 123.54 10.39 123.69 ;
        RECT 5.525 123.69 10.39 123.84 ;
        RECT 5.375 123.84 10.39 123.99 ;
        RECT 5.225 123.99 10.39 124.14 ;
        RECT 5.075 124.14 10.39 124.29 ;
        RECT 4.925 124.29 10.39 124.405 ;
        RECT 6.595 122.62 10.71 122.77 ;
        RECT 6.445 122.77 10.56 122.92 ;
        RECT 6.295 122.92 10.41 123.07 ;
        RECT 6.145 123.07 10.39 123.09 ;
        RECT 9.91 119.305 10.86 119.455 ;
        RECT 9.76 119.455 10.86 119.605 ;
        RECT 9.61 119.605 10.86 119.755 ;
        RECT 9.46 119.755 10.86 119.905 ;
        RECT 9.31 119.905 10.86 120.055 ;
        RECT 9.16 120.055 10.86 120.205 ;
        RECT 9.01 120.205 10.86 120.355 ;
        RECT 8.86 120.355 10.86 120.505 ;
        RECT 8.71 120.505 10.86 120.655 ;
        RECT 8.56 120.655 10.86 120.805 ;
        RECT 8.41 120.805 10.86 120.955 ;
        RECT 8.26 120.955 10.86 121.105 ;
        RECT 8.11 121.105 10.86 121.255 ;
        RECT 7.96 121.255 10.86 121.405 ;
        RECT 7.81 121.405 10.86 121.555 ;
        RECT 7.66 121.555 10.86 121.705 ;
        RECT 7.51 121.705 10.86 121.855 ;
        RECT 7.36 121.855 10.86 122.005 ;
        RECT 7.21 122.005 10.86 122.155 ;
        RECT 7.06 122.155 10.86 122.305 ;
        RECT 6.91 122.305 10.86 122.455 ;
        RECT 6.76 122.455 10.86 122.605 ;
        RECT 6.61 122.605 10.86 122.62 ;
        RECT 29.76 65.32 30.72 133.14 ;
        RECT 34.72 65.32 35.68 133.16 ;
        RECT 39.7 65.32 40.62 133.12 ;
        RECT 24.8 65.32 25.76 133.16 ;
        RECT 19.86 65.32 20.78 133.12 ;
        RECT 14.9 65.32 15.82 132.32 ;
        RECT 24.79 65.3 25.76 65.31 ;
        RECT 24.8 65.31 25.76 65.32 ;
        RECT 9.91 65.29 10.86 119.305 ;
        RECT 14.885 65.29 15.82 65.305 ;
        RECT 14.9 65.305 15.82 65.32 ;
        RECT 24.065 64.435 26.475 64.585 ;
        RECT 24.215 64.585 26.325 64.735 ;
        RECT 24.365 64.735 26.175 64.885 ;
        RECT 24.515 64.885 26.025 65.035 ;
        RECT 24.665 65.035 25.875 65.185 ;
        RECT 24.78 65.185 25.76 65.3 ;
        RECT 29.025 64.435 31.455 64.585 ;
        RECT 29.175 64.585 31.305 64.735 ;
        RECT 29.325 64.735 31.155 64.885 ;
        RECT 29.475 64.885 31.005 65.035 ;
        RECT 29.625 65.035 30.855 65.185 ;
        RECT 29.76 65.185 30.72 65.32 ;
        RECT 33.985 64.435 36.415 64.585 ;
        RECT 34.135 64.585 36.265 64.735 ;
        RECT 34.285 64.735 36.115 64.885 ;
        RECT 34.435 64.885 35.965 65.035 ;
        RECT 34.585 65.035 35.815 65.185 ;
        RECT 34.72 65.185 35.68 65.32 ;
        RECT 38.965 64.435 40.62 64.585 ;
        RECT 39.115 64.585 40.62 64.735 ;
        RECT 39.265 64.735 40.62 64.885 ;
        RECT 39.415 64.885 40.62 65.035 ;
        RECT 39.565 65.035 40.62 65.185 ;
        RECT 39.7 65.185 40.62 65.32 ;
        RECT 19.125 64.435 21.515 64.585 ;
        RECT 19.275 64.585 21.365 64.735 ;
        RECT 19.425 64.735 21.215 64.885 ;
        RECT 19.575 64.885 21.065 65.035 ;
        RECT 19.725 65.035 20.915 65.185 ;
        RECT 19.86 65.185 20.78 65.32 ;
        RECT 9.91 64.435 11.565 64.585 ;
        RECT 9.91 64.585 11.415 64.735 ;
        RECT 9.91 64.735 11.265 64.885 ;
        RECT 9.91 64.885 11.115 65.035 ;
        RECT 9.91 65.035 10.965 65.185 ;
        RECT 9.91 65.185 10.86 65.29 ;
        RECT 14.165 64.435 16.525 64.585 ;
        RECT 14.315 64.585 16.375 64.735 ;
        RECT 14.465 64.735 16.225 64.885 ;
        RECT 14.615 64.885 16.075 65.035 ;
        RECT 14.765 65.035 15.925 65.185 ;
        RECT 14.87 65.185 15.82 65.29 ;
        RECT 9.91 61.99 40.62 64.435 ;
        RECT 11.25 60.65 40.62 60.8 ;
        RECT 11.1 60.8 40.62 60.95 ;
        RECT 10.95 60.95 40.62 61.1 ;
        RECT 10.8 61.1 40.62 61.25 ;
        RECT 10.65 61.25 40.62 61.4 ;
        RECT 10.5 61.4 40.62 61.55 ;
        RECT 10.35 61.55 40.62 61.7 ;
        RECT 10.2 61.7 40.62 61.85 ;
        RECT 10.05 61.85 40.62 61.99 ;
        RECT 19.475 52.425 32.395 52.575 ;
        RECT 19.325 52.575 32.545 52.725 ;
        RECT 19.175 52.725 32.695 52.875 ;
        RECT 19.025 52.875 32.845 53.025 ;
        RECT 18.875 53.025 32.995 53.175 ;
        RECT 18.725 53.175 33.145 53.325 ;
        RECT 18.575 53.325 33.295 53.475 ;
        RECT 18.425 53.475 33.445 53.625 ;
        RECT 18.275 53.625 33.595 53.775 ;
        RECT 18.125 53.775 33.745 53.925 ;
        RECT 17.975 53.925 33.895 54.075 ;
        RECT 17.825 54.075 34.045 54.225 ;
        RECT 17.675 54.225 34.195 54.375 ;
        RECT 17.525 54.375 34.345 54.525 ;
        RECT 17.375 54.525 34.495 54.675 ;
        RECT 17.225 54.675 34.645 54.825 ;
        RECT 17.075 54.825 34.795 54.975 ;
        RECT 16.925 54.975 34.945 55.125 ;
        RECT 16.775 55.125 35.095 55.275 ;
        RECT 16.625 55.275 35.245 55.425 ;
        RECT 16.475 55.425 35.395 55.575 ;
        RECT 16.325 55.575 35.545 55.725 ;
        RECT 16.175 55.725 35.695 55.875 ;
        RECT 16.025 55.875 35.845 56.025 ;
        RECT 15.875 56.025 35.995 56.175 ;
        RECT 15.725 56.175 36.145 56.325 ;
        RECT 15.575 56.325 36.295 56.475 ;
        RECT 15.425 56.475 36.445 56.625 ;
        RECT 15.275 56.625 36.595 56.775 ;
        RECT 15.125 56.775 36.745 56.925 ;
        RECT 14.975 56.925 36.895 57.075 ;
        RECT 14.825 57.075 37.045 57.225 ;
        RECT 14.675 57.225 37.195 57.375 ;
        RECT 14.525 57.375 37.345 57.525 ;
        RECT 14.375 57.525 37.495 57.675 ;
        RECT 14.225 57.675 37.645 57.825 ;
        RECT 14.075 57.825 37.795 57.975 ;
        RECT 13.925 57.975 37.945 58.125 ;
        RECT 13.775 58.125 38.095 58.275 ;
        RECT 13.625 58.275 38.245 58.425 ;
        RECT 13.475 58.425 38.395 58.575 ;
        RECT 13.325 58.575 38.545 58.725 ;
        RECT 13.175 58.725 38.695 58.875 ;
        RECT 13.025 58.875 38.845 59.025 ;
        RECT 12.875 59.025 38.995 59.175 ;
        RECT 12.725 59.175 39.145 59.325 ;
        RECT 12.575 59.325 39.295 59.475 ;
        RECT 12.425 59.475 39.445 59.625 ;
        RECT 12.275 59.625 39.595 59.775 ;
        RECT 12.125 59.775 39.745 59.925 ;
        RECT 11.975 59.925 39.895 60.075 ;
        RECT 11.825 60.075 40.045 60.225 ;
        RECT 11.675 60.225 40.195 60.375 ;
        RECT 11.525 60.375 40.345 60.525 ;
        RECT 11.375 60.525 40.495 60.65 ;
        RECT 20.835 51.065 32.395 51.215 ;
        RECT 20.685 51.215 32.395 51.365 ;
        RECT 20.535 51.365 32.395 51.515 ;
        RECT 20.385 51.515 32.395 51.665 ;
        RECT 20.235 51.665 32.395 51.815 ;
        RECT 20.085 51.815 32.395 51.965 ;
        RECT 19.935 51.965 32.395 52.115 ;
        RECT 19.785 52.115 32.395 52.265 ;
        RECT 19.635 52.265 32.395 52.415 ;
        RECT 19.485 52.415 32.395 52.425 ;
        RECT 20.835 35.455 32.395 51.065 ;
        RECT 20.835 34.315 33.385 34.465 ;
        RECT 20.835 34.465 33.235 34.615 ;
        RECT 20.835 34.615 33.085 34.765 ;
        RECT 20.835 34.765 32.935 34.915 ;
        RECT 20.835 34.915 32.785 35.065 ;
        RECT 20.835 35.065 32.635 35.215 ;
        RECT 20.835 35.215 32.485 35.365 ;
        RECT 20.835 35.365 32.395 35.455 ;
        RECT 20.86 34.29 33.535 34.315 ;
        RECT 21.01 34.14 33.56 34.29 ;
        RECT 21.16 33.99 33.71 34.14 ;
        RECT 21.31 33.84 33.86 33.99 ;
        RECT 21.46 33.69 34.01 33.84 ;
        RECT 21.61 33.54 34.16 33.69 ;
        RECT 21.76 33.39 34.31 33.54 ;
        RECT 21.91 33.24 34.46 33.39 ;
        RECT 22.06 33.09 34.61 33.24 ;
        RECT 22.21 32.94 34.76 33.09 ;
        RECT 22.36 32.79 34.91 32.94 ;
        RECT 22.51 32.64 35.06 32.79 ;
        RECT 22.66 32.49 35.21 32.64 ;
        RECT 22.81 32.34 35.36 32.49 ;
        RECT 22.96 32.19 35.51 32.34 ;
        RECT 23.11 32.04 35.66 32.19 ;
        RECT 23.26 31.89 35.81 32.04 ;
        RECT 23.41 31.74 35.96 31.89 ;
        RECT 23.56 31.59 36.11 31.74 ;
        RECT 23.71 31.44 36.26 31.59 ;
        RECT 23.86 31.29 36.41 31.44 ;
        RECT 24.01 31.14 36.56 31.29 ;
        RECT 24.16 30.99 36.71 31.14 ;
        RECT 24.31 30.84 36.86 30.99 ;
        RECT 24.46 30.69 37.01 30.84 ;
        RECT 24.61 30.54 37.16 30.69 ;
        RECT 24.76 30.39 37.31 30.54 ;
        RECT 24.91 30.24 37.46 30.39 ;
        RECT 25.06 30.09 37.61 30.24 ;
        RECT 25.21 29.94 37.76 30.09 ;
        RECT 25.36 29.79 37.91 29.94 ;
        RECT 25.51 29.64 38.06 29.79 ;
        RECT 25.66 29.49 38.21 29.64 ;
        RECT 25.81 29.34 38.36 29.49 ;
        RECT 25.96 29.19 38.51 29.34 ;
        RECT 26.11 29.04 38.66 29.19 ;
        RECT 26.26 28.89 38.81 29.04 ;
        RECT 26.41 28.74 38.96 28.89 ;
        RECT 26.56 28.59 39.11 28.74 ;
        RECT 26.71 28.44 39.26 28.59 ;
        RECT 26.86 28.29 39.41 28.44 ;
        RECT 27.01 28.14 39.56 28.29 ;
        RECT 27.16 27.99 39.71 28.14 ;
        RECT 27.31 27.84 39.86 27.99 ;
        RECT 27.46 27.69 40.01 27.84 ;
        RECT 27.61 27.54 40.16 27.69 ;
        RECT 27.76 27.39 40.31 27.54 ;
        RECT 27.91 27.24 40.46 27.39 ;
        RECT 28.06 27.09 40.61 27.24 ;
        RECT 28.21 26.94 40.76 27.09 ;
        RECT 28.36 26.79 40.91 26.94 ;
        RECT 28.51 26.64 41.06 26.79 ;
        RECT 28.66 26.49 41.21 26.64 ;
        RECT 28.81 26.34 41.36 26.49 ;
        RECT 28.96 26.19 41.51 26.34 ;
        RECT 29.11 26.04 41.66 26.19 ;
        RECT 29.26 25.89 41.81 26.04 ;
        RECT 29.41 25.74 41.96 25.89 ;
        RECT 29.56 25.59 42.11 25.74 ;
        RECT 29.71 25.44 42.26 25.59 ;
        RECT 29.86 25.29 42.41 25.44 ;
        RECT 30.01 25.14 42.56 25.29 ;
        RECT 30.16 24.99 42.71 25.14 ;
        RECT 30.31 24.84 42.86 24.99 ;
        RECT 30.46 24.69 43.01 24.84 ;
        RECT 30.61 24.54 43.16 24.69 ;
        RECT 30.76 24.39 43.31 24.54 ;
        RECT 30.91 24.24 43.46 24.39 ;
        RECT 31.06 24.09 43.61 24.24 ;
        RECT 31.21 23.94 43.76 24.09 ;
        RECT 31.36 23.79 43.91 23.94 ;
        RECT 31.51 23.64 44.06 23.79 ;
        RECT 31.66 23.49 44.21 23.64 ;
        RECT 31.81 23.34 44.36 23.49 ;
        RECT 31.96 23.19 44.51 23.34 ;
        RECT 32.11 23.04 44.66 23.19 ;
        RECT 32.26 22.89 44.81 23.04 ;
        RECT 32.41 22.74 44.96 22.89 ;
        RECT 32.56 22.59 45.11 22.74 ;
        RECT 32.71 22.44 45.26 22.59 ;
        RECT 32.86 22.29 45.41 22.44 ;
        RECT 33.01 22.14 45.56 22.29 ;
        RECT 33.16 21.99 45.71 22.14 ;
        RECT 33.31 21.84 45.86 21.99 ;
        RECT 33.46 21.69 46.01 21.84 ;
        RECT 33.61 21.54 46.16 21.69 ;
        RECT 33.76 21.39 46.31 21.54 ;
        RECT 33.91 21.24 46.46 21.39 ;
        RECT 34.06 21.09 46.61 21.24 ;
        RECT 34.21 20.94 46.76 21.09 ;
        RECT 34.36 20.79 46.91 20.94 ;
        RECT 34.51 20.64 47.06 20.79 ;
        RECT 34.66 20.49 47.21 20.64 ;
        RECT 34.81 20.34 47.36 20.49 ;
        RECT 34.96 20.19 47.51 20.34 ;
        RECT 35.11 20.04 47.66 20.19 ;
        RECT 38.83 16.32 47.81 16.47 ;
        RECT 38.68 16.47 47.81 16.62 ;
        RECT 38.53 16.62 47.81 16.77 ;
        RECT 38.38 16.77 47.81 16.92 ;
        RECT 38.23 16.92 47.81 17.07 ;
        RECT 38.08 17.07 47.81 17.22 ;
        RECT 37.93 17.22 47.81 17.37 ;
        RECT 37.78 17.37 47.81 17.52 ;
        RECT 37.63 17.52 47.81 17.67 ;
        RECT 37.48 17.67 47.81 17.82 ;
        RECT 37.33 17.82 47.81 17.97 ;
        RECT 37.18 17.97 47.81 18.12 ;
        RECT 37.03 18.12 47.81 18.27 ;
        RECT 36.88 18.27 47.81 18.42 ;
        RECT 36.73 18.42 47.81 18.57 ;
        RECT 36.58 18.57 47.81 18.72 ;
        RECT 36.43 18.72 47.81 18.87 ;
        RECT 36.28 18.87 47.81 19.02 ;
        RECT 36.13 19.02 47.81 19.17 ;
        RECT 35.98 19.17 47.81 19.32 ;
        RECT 35.83 19.32 47.81 19.47 ;
        RECT 35.68 19.47 47.81 19.62 ;
        RECT 35.53 19.62 47.81 19.77 ;
        RECT 35.38 19.77 47.81 19.92 ;
        RECT 35.23 19.92 47.81 20.04 ;
        RECT 38.83 0 47.81 16.32 ;
    END
    ANTENNAPARTIALMETALSIDEAREA 14.856 LAYER met3 ;
  END pad_core

  PIN amuxbus_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0 46.365 75 49.345 ;
    END
    ANTENNAPARTIALMETALSIDEAREA 111.168 LAYER met4 ;
  END amuxbus_b

  PIN amuxbus_a
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0 51.125 75 54.105 ;
    END
    ANTENNAPARTIALMETALSIDEAREA 111.168 LAYER met4 ;
  END amuxbus_a

  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 6.985 75 11.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 6.885 75 11.535 ;
    END
  END vccd

  PIN vddio_q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 62.185 75 66.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 62.085 75 66.535 ;
    END
  END vddio_q

  PIN vssa
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 34.835 75 38.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0 45.735 75 54.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 34.735 75 38.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 45.735 75 46.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 49.645 75 50.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 54.405 75 54.735 ;
    END
  END vssa

  PIN vddio
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 17.885 75 22.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 0 68.035 75 92.985 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 17.785 75 22.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 68.035 75 93 ;
    END
  END vddio

  PIN vcchib
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 0.135 75 5.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 0.035 75 5.485 ;
    END
  END vcchib

  PIN vswitch
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 29.985 75 33.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 29.885 75 33.335 ;
    END
  END vswitch

  PIN vssio_q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 56.335 75 60.585 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 56.235 75 60.685 ;
    END
  END vssio_q

  PIN vdda
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 13.035 75 16.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 12.935 75 16.385 ;
    END
  END vdda

  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 39.685 75 44.135 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 39.585 75 44.235 ;
    END
  END vssd

  PIN pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 4.8 102.23 70.2 164.57 ;
        RECT 5.6 164.57 69.4 165.37 ;
        RECT 6.4 165.37 68.6 166.17 ;
        RECT 7.2 166.17 67.8 166.97 ;
        RECT 8 166.97 67 167.77 ;
        RECT 8.8 167.77 66.2 168.57 ;
        RECT 9.6 168.57 65.4 169.37 ;
        RECT 10.4 169.37 64.6 170.17 ;
        RECT 11.2 170.17 63.8 170.97 ;
        RECT 11.33 170.97 63.67 171.1 ;
        RECT 11.33 95.7 63.67 96.5 ;
        RECT 10.53 96.5 64.47 97.3 ;
        RECT 9.73 97.3 65.27 98.1 ;
        RECT 8.93 98.1 66.07 98.9 ;
        RECT 8.13 98.9 66.87 99.7 ;
        RECT 7.33 99.7 67.67 100.5 ;
        RECT 6.53 100.5 68.47 101.3 ;
        RECT 5.73 101.3 69.27 102.1 ;
        RECT 4.93 102.1 70.07 102.23 ;
    END
    ANTENNADIFFAREA 426.8 LAYER met1 ;
    ANTENNADIFFAREA 426.8 LAYER met2 ;
    ANTENNADIFFAREA 426.8 LAYER met3 ;
    ANTENNADIFFAREA 426.8 LAYER met4 ;
    ANTENNADIFFAREA 426.8 LAYER met5 ;
    ANTENNAPARTIALMETALSIDEAREA 245.627 LAYER met5 ;
  END pad

  PIN vssio
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 23.935 75 28.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0 173.785 75 198 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 23.835 75 28.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 173.785 75 198 ;
    END
  END vssio
  OBS
    LAYER met3 ;
      RECT 11.34 65.235 14.43 65.415 ;
      RECT 11.88 64.835 14.25 65.235 ;
      RECT 0 61.825 9.51 65.235 ;
      RECT 41.02 60.485 75 65.235 ;
      RECT 32.795 52.26 75 60.485 ;
      RECT 0 50.9 9.51 61.825 ;
      RECT 32.795 35.62 75 52.26 ;
      RECT 48.21 20.205 75 35.62 ;
      RECT 0 16.155 20.435 34.15 ;
      RECT 48.21 0 75 20.205 ;
      RECT 0 0 38.43 16.155 ;
      RECT 0 34.15 20.435 50.9 ;
      RECT 0 171.425 75 198 ;
      RECT 0 169.52 14.09 171.425 ;
      RECT 10.69 148.94 14.09 169.52 ;
      RECT 10.69 148.84 10.79 148.94 ;
      RECT 0 147.28 9.13 169.52 ;
      RECT 0 147.18 9.13 147.28 ;
      RECT 0 146.615 9.03 147.18 ;
      RECT 0 141.99 9.03 146.615 ;
      RECT 25.57 136.12 28.97 171.425 ;
      RECT 35.51 136.1 38.89 171.425 ;
      RECT 40.45 136.1 75 171.425 ;
      RECT 20.61 136.1 24.01 171.425 ;
      RECT 30.53 136.1 33.93 171.425 ;
      RECT 35.98 135.63 38.89 136.1 ;
      RECT 40.92 135.63 75 136.1 ;
      RECT 26.06 135.63 28.97 136.12 ;
      RECT 21.08 135.63 24.01 136.1 ;
      RECT 31.02 135.61 33.93 136.1 ;
      RECT 15.65 134.885 19.05 171.425 ;
      RECT 16.12 134.415 19.05 134.885 ;
      RECT 21.08 133.525 24.01 135.63 ;
      RECT 31.02 133.525 33.93 135.61 ;
      RECT 35.98 133.505 38.89 135.63 ;
      RECT 26.06 133.505 28.97 135.63 ;
      RECT 16.12 133.505 19.05 134.415 ;
      RECT 21.08 133.035 24.01 133.525 ;
      RECT 31.02 133.035 33.93 133.525 ;
      RECT 26.06 133.015 28.97 133.505 ;
      RECT 35.98 132.995 38.89 133.505 ;
      RECT 16.12 132.995 19.05 133.505 ;
      RECT 10.79 132.705 14.09 148.94 ;
      RECT 10.79 132.195 14.09 132.705 ;
      RECT 0 124.005 4.405 141.99 ;
      RECT 10.79 123.255 14.6 132.195 ;
      RECT 11.26 122.785 14.6 123.255 ;
      RECT 0 119.14 4.645 124.005 ;
      RECT 0 118.57 9.51 119.14 ;
      RECT 0 118.475 9.51 118.57 ;
      RECT 11.26 116.82 14.6 122.785 ;
      RECT 35.98 66.15 39.4 132.995 ;
      RECT 21.08 66.15 24.5 133.035 ;
      RECT 31.02 66.15 34.42 133.035 ;
      RECT 26.06 66.15 29.46 133.015 ;
      RECT 16.12 66.15 19.56 132.995 ;
      RECT 11.16 66.15 14.6 116.82 ;
      RECT 26.06 66.13 29.46 66.15 ;
      RECT 16.12 66.12 19.56 66.15 ;
      RECT 36.08 66.05 39.4 66.15 ;
      RECT 11.16 66.05 14.6 66.15 ;
      RECT 21.18 66.05 24.5 66.15 ;
      RECT 31.12 66.05 34.42 66.15 ;
      RECT 26.14 66.05 29.44 66.13 ;
      RECT 16.19 66.05 19.53 66.12 ;
      RECT 26.16 66.03 29.36 66.05 ;
      RECT 16.22 66.02 19.46 66.05 ;
      RECT 36.08 65.485 39.4 66.05 ;
      RECT 11.16 65.485 14.5 66.05 ;
      RECT 21.18 65.485 24.4 66.05 ;
      RECT 31.12 65.485 34.32 66.05 ;
      RECT 26.16 65.485 29.36 66.03 ;
      RECT 16.22 65.485 19.46 66.02 ;
      RECT 26.16 65.465 29.36 65.485 ;
      RECT 16.22 65.455 19.46 65.485 ;
      RECT 36.12 65.445 39.4 65.485 ;
      RECT 11.16 65.415 14.5 65.485 ;
      RECT 36.33 65.235 39.4 65.445 ;
      RECT 36.73 64.835 39.05 65.235 ;
      RECT 40.92 65.235 75 135.63 ;
      RECT 0 65.235 9.61 118.475 ;
      RECT 21.83 64.835 24.4 65.485 ;
      RECT 31.77 64.835 34.32 65.485 ;
      RECT 26.79 64.835 29.34 65.465 ;
      RECT 16.84 64.835 19.43 65.455 ;
      RECT 36.28 65.285 39.1 65.435 ;
      RECT 36.13 65.435 39.25 65.485 ;
      RECT 26.16 132.975 29.21 133.125 ;
      RECT 26.16 133.125 29.06 133.275 ;
      RECT 26.16 133.275 28.91 133.425 ;
      RECT 26.16 133.425 28.87 133.465 ;
      RECT 26.16 65.465 29.34 65.475 ;
      RECT 26.16 65.475 29.35 65.485 ;
      RECT 16.22 134.455 18.95 134.605 ;
      RECT 16.07 134.605 18.95 134.755 ;
      RECT 15.92 134.755 18.95 134.905 ;
      RECT 15.77 134.905 18.95 134.925 ;
      RECT 0 146.49 8.905 146.615 ;
      RECT 0 146.34 8.755 146.49 ;
      RECT 0 146.19 8.605 146.34 ;
      RECT 0 146.04 8.455 146.19 ;
      RECT 0 145.89 8.305 146.04 ;
      RECT 0 145.74 8.155 145.89 ;
      RECT 0 145.59 8.005 145.74 ;
      RECT 0 145.44 7.855 145.59 ;
      RECT 0 145.29 7.705 145.44 ;
      RECT 0 145.14 7.555 145.29 ;
      RECT 0 144.99 7.405 145.14 ;
      RECT 0 144.84 7.255 144.99 ;
      RECT 0 144.69 7.105 144.84 ;
      RECT 0 144.54 6.955 144.69 ;
      RECT 0 144.39 6.805 144.54 ;
      RECT 0 144.24 6.655 144.39 ;
      RECT 0 144.09 6.505 144.24 ;
      RECT 0 143.94 6.355 144.09 ;
      RECT 0 143.79 6.205 143.94 ;
      RECT 0 143.64 6.055 143.79 ;
      RECT 0 143.49 5.905 143.64 ;
      RECT 0 143.34 5.755 143.49 ;
      RECT 0 143.19 5.605 143.34 ;
      RECT 0 143.04 5.455 143.19 ;
      RECT 0 142.89 5.305 143.04 ;
      RECT 0 142.74 5.155 142.89 ;
      RECT 0 142.59 5.005 142.74 ;
      RECT 0 142.44 4.855 142.59 ;
      RECT 0 142.29 4.705 142.44 ;
      RECT 0 142.14 4.555 142.29 ;
      RECT 0 141.99 4.405 142.14 ;
      RECT 32.945 52.26 75 52.41 ;
      RECT 33.095 52.41 75 52.56 ;
      RECT 33.245 52.56 75 52.71 ;
      RECT 33.395 52.71 75 52.86 ;
      RECT 33.545 52.86 75 53.01 ;
      RECT 33.695 53.01 75 53.16 ;
      RECT 33.845 53.16 75 53.31 ;
      RECT 33.995 53.31 75 53.46 ;
      RECT 34.145 53.46 75 53.61 ;
      RECT 34.295 53.61 75 53.76 ;
      RECT 34.445 53.76 75 53.91 ;
      RECT 34.595 53.91 75 54.06 ;
      RECT 34.745 54.06 75 54.21 ;
      RECT 34.895 54.21 75 54.36 ;
      RECT 35.045 54.36 75 54.51 ;
      RECT 35.195 54.51 75 54.66 ;
      RECT 35.345 54.66 75 54.81 ;
      RECT 35.495 54.81 75 54.96 ;
      RECT 35.645 54.96 75 55.11 ;
      RECT 35.795 55.11 75 55.26 ;
      RECT 35.945 55.26 75 55.41 ;
      RECT 36.095 55.41 75 55.56 ;
      RECT 36.245 55.56 75 55.71 ;
      RECT 36.395 55.71 75 55.86 ;
      RECT 36.545 55.86 75 56.01 ;
      RECT 36.695 56.01 75 56.16 ;
      RECT 36.845 56.16 75 56.31 ;
      RECT 36.995 56.31 75 56.46 ;
      RECT 37.145 56.46 75 56.61 ;
      RECT 37.295 56.61 75 56.76 ;
      RECT 37.445 56.76 75 56.91 ;
      RECT 37.595 56.91 75 57.06 ;
      RECT 37.745 57.06 75 57.21 ;
      RECT 37.895 57.21 75 57.36 ;
      RECT 38.045 57.36 75 57.51 ;
      RECT 38.195 57.51 75 57.66 ;
      RECT 38.345 57.66 75 57.81 ;
      RECT 38.495 57.81 75 57.96 ;
      RECT 38.645 57.96 75 58.11 ;
      RECT 38.795 58.11 75 58.26 ;
      RECT 38.945 58.26 75 58.41 ;
      RECT 39.095 58.41 75 58.56 ;
      RECT 39.245 58.56 75 58.71 ;
      RECT 39.395 58.71 75 58.86 ;
      RECT 39.545 58.86 75 59.01 ;
      RECT 39.695 59.01 75 59.16 ;
      RECT 39.845 59.16 75 59.31 ;
      RECT 39.995 59.31 75 59.46 ;
      RECT 40.145 59.46 75 59.61 ;
      RECT 40.295 59.61 75 59.76 ;
      RECT 40.445 59.76 75 59.91 ;
      RECT 40.595 59.91 75 60.06 ;
      RECT 40.745 60.06 75 60.21 ;
      RECT 40.895 60.21 75 60.36 ;
      RECT 41.02 60.36 75 60.485 ;
      RECT 41.02 135.67 75 135.82 ;
      RECT 40.87 135.82 75 135.97 ;
      RECT 40.72 135.97 75 136.12 ;
      RECT 40.57 136.12 75 136.14 ;
      RECT 10.79 132.155 14.35 132.305 ;
      RECT 10.79 132.305 14.2 132.455 ;
      RECT 10.79 132.455 14.05 132.605 ;
      RECT 10.79 132.605 13.99 132.665 ;
      RECT 11.26 122.785 14.5 122.935 ;
      RECT 11.11 122.935 14.5 123.085 ;
      RECT 10.96 123.085 14.5 123.235 ;
      RECT 10.81 123.235 14.5 123.255 ;
      RECT 34.41 34.005 75 34.155 ;
      RECT 34.56 33.855 75 34.005 ;
      RECT 34.71 33.705 75 33.855 ;
      RECT 34.86 33.555 75 33.705 ;
      RECT 35.01 33.405 75 33.555 ;
      RECT 35.16 33.255 75 33.405 ;
      RECT 35.31 33.105 75 33.255 ;
      RECT 35.46 32.955 75 33.105 ;
      RECT 35.61 32.805 75 32.955 ;
      RECT 35.76 32.655 75 32.805 ;
      RECT 35.91 32.505 75 32.655 ;
      RECT 36.06 32.355 75 32.505 ;
      RECT 36.21 32.205 75 32.355 ;
      RECT 36.36 32.055 75 32.205 ;
      RECT 36.51 31.905 75 32.055 ;
      RECT 36.66 31.755 75 31.905 ;
      RECT 36.81 31.605 75 31.755 ;
      RECT 36.96 31.455 75 31.605 ;
      RECT 37.11 31.305 75 31.455 ;
      RECT 37.26 31.155 75 31.305 ;
      RECT 37.41 31.005 75 31.155 ;
      RECT 37.56 30.855 75 31.005 ;
      RECT 37.71 30.705 75 30.855 ;
      RECT 37.86 30.555 75 30.705 ;
      RECT 38.01 30.405 75 30.555 ;
      RECT 38.16 30.255 75 30.405 ;
      RECT 38.31 30.105 75 30.255 ;
      RECT 38.46 29.955 75 30.105 ;
      RECT 38.61 29.805 75 29.955 ;
      RECT 38.76 29.655 75 29.805 ;
      RECT 38.91 29.505 75 29.655 ;
      RECT 39.06 29.355 75 29.505 ;
      RECT 39.21 29.205 75 29.355 ;
      RECT 39.36 29.055 75 29.205 ;
      RECT 39.51 28.905 75 29.055 ;
      RECT 39.66 28.755 75 28.905 ;
      RECT 39.81 28.605 75 28.755 ;
      RECT 39.96 28.455 75 28.605 ;
      RECT 40.11 28.305 75 28.455 ;
      RECT 40.26 28.155 75 28.305 ;
      RECT 40.41 28.005 75 28.155 ;
      RECT 40.56 27.855 75 28.005 ;
      RECT 40.71 27.705 75 27.855 ;
      RECT 40.86 27.555 75 27.705 ;
      RECT 41.01 27.405 75 27.555 ;
      RECT 41.16 27.255 75 27.405 ;
      RECT 41.31 27.105 75 27.255 ;
      RECT 41.46 26.955 75 27.105 ;
      RECT 41.61 26.805 75 26.955 ;
      RECT 41.76 26.655 75 26.805 ;
      RECT 41.91 26.505 75 26.655 ;
      RECT 42.06 26.355 75 26.505 ;
      RECT 42.21 26.205 75 26.355 ;
      RECT 42.36 26.055 75 26.205 ;
      RECT 42.51 25.905 75 26.055 ;
      RECT 42.66 25.755 75 25.905 ;
      RECT 42.81 25.605 75 25.755 ;
      RECT 42.96 25.455 75 25.605 ;
      RECT 43.11 25.305 75 25.455 ;
      RECT 43.26 25.155 75 25.305 ;
      RECT 43.41 25.005 75 25.155 ;
      RECT 43.56 24.855 75 25.005 ;
      RECT 43.71 24.705 75 24.855 ;
      RECT 43.86 24.555 75 24.705 ;
      RECT 44.01 24.405 75 24.555 ;
      RECT 44.16 24.255 75 24.405 ;
      RECT 44.31 24.105 75 24.255 ;
      RECT 44.46 23.955 75 24.105 ;
      RECT 44.61 23.805 75 23.955 ;
      RECT 44.76 23.655 75 23.805 ;
      RECT 44.91 23.505 75 23.655 ;
      RECT 45.06 23.355 75 23.505 ;
      RECT 45.21 23.205 75 23.355 ;
      RECT 45.36 23.055 75 23.205 ;
      RECT 45.51 22.905 75 23.055 ;
      RECT 45.66 22.755 75 22.905 ;
      RECT 45.81 22.605 75 22.755 ;
      RECT 45.96 22.455 75 22.605 ;
      RECT 46.11 22.305 75 22.455 ;
      RECT 46.26 22.155 75 22.305 ;
      RECT 46.41 22.005 75 22.155 ;
      RECT 46.56 21.855 75 22.005 ;
      RECT 46.71 21.705 75 21.855 ;
      RECT 46.86 21.555 75 21.705 ;
      RECT 47.01 21.405 75 21.555 ;
      RECT 47.16 21.255 75 21.405 ;
      RECT 47.31 21.105 75 21.255 ;
      RECT 47.46 20.955 75 21.105 ;
      RECT 47.61 20.805 75 20.955 ;
      RECT 47.76 20.655 75 20.805 ;
      RECT 47.91 20.505 75 20.655 ;
      RECT 48.06 20.355 75 20.505 ;
      RECT 48.21 20.205 75 20.355 ;
      RECT 21.18 132.995 24.25 133.145 ;
      RECT 21.18 133.145 24.1 133.295 ;
      RECT 21.18 133.295 23.95 133.445 ;
      RECT 21.18 133.445 23.91 133.485 ;
      RECT 21.83 64.835 23.75 64.985 ;
      RECT 21.68 64.985 23.9 65.135 ;
      RECT 21.53 65.135 24.05 65.285 ;
      RECT 21.38 65.285 24.2 65.435 ;
      RECT 21.23 65.435 24.35 65.485 ;
      RECT 31.12 132.995 34.17 133.145 ;
      RECT 31.12 133.145 34.02 133.295 ;
      RECT 31.12 133.295 33.87 133.445 ;
      RECT 31.12 133.445 33.83 133.485 ;
      RECT 31.77 64.835 33.67 64.985 ;
      RECT 31.62 64.985 33.82 65.135 ;
      RECT 31.47 65.135 33.97 65.285 ;
      RECT 31.32 65.285 34.12 65.435 ;
      RECT 31.17 65.435 34.27 65.485 ;
      RECT 16.22 132.955 19.31 133.105 ;
      RECT 16.22 133.105 19.16 133.255 ;
      RECT 16.22 133.255 19.01 133.405 ;
      RECT 16.22 133.405 18.95 133.465 ;
      RECT 16.22 65.455 19.43 65.47 ;
      RECT 16.22 65.47 19.445 65.485 ;
      RECT 36.08 132.955 39.15 133.105 ;
      RECT 36.08 133.105 39.0 133.255 ;
      RECT 36.08 133.255 38.85 133.405 ;
      RECT 36.08 133.405 38.79 133.465 ;
      RECT 36.73 64.835 38.65 64.985 ;
      RECT 36.58 64.985 38.8 65.135 ;
      RECT 36.43 65.135 38.95 65.285 ;
      RECT 0 33.405 21.03 33.555 ;
      RECT 0 33.255 21.18 33.405 ;
      RECT 0 33.105 21.33 33.255 ;
      RECT 0 32.955 21.48 33.105 ;
      RECT 0 32.805 21.63 32.955 ;
      RECT 0 32.655 21.78 32.805 ;
      RECT 0 32.505 21.93 32.655 ;
      RECT 0 32.355 22.08 32.505 ;
      RECT 0 32.205 22.23 32.355 ;
      RECT 0 32.055 22.38 32.205 ;
      RECT 0 31.905 22.53 32.055 ;
      RECT 0 31.755 22.68 31.905 ;
      RECT 0 31.605 22.83 31.755 ;
      RECT 0 31.455 22.98 31.605 ;
      RECT 0 31.305 23.13 31.455 ;
      RECT 0 31.155 23.28 31.305 ;
      RECT 0 31.005 23.43 31.155 ;
      RECT 0 30.855 23.58 31.005 ;
      RECT 0 30.705 23.73 30.855 ;
      RECT 0 30.555 23.88 30.705 ;
      RECT 0 30.405 24.03 30.555 ;
      RECT 0 30.255 24.18 30.405 ;
      RECT 0 30.105 24.33 30.255 ;
      RECT 0 29.955 24.48 30.105 ;
      RECT 0 29.805 24.63 29.955 ;
      RECT 0 29.655 24.78 29.805 ;
      RECT 0 29.505 24.93 29.655 ;
      RECT 0 29.355 25.08 29.505 ;
      RECT 0 29.205 25.23 29.355 ;
      RECT 0 29.055 25.38 29.205 ;
      RECT 0 28.905 25.53 29.055 ;
      RECT 0 28.755 25.68 28.905 ;
      RECT 0 28.605 25.83 28.755 ;
      RECT 0 28.455 25.98 28.605 ;
      RECT 0 28.305 26.13 28.455 ;
      RECT 0 28.155 26.28 28.305 ;
      RECT 0 28.005 26.43 28.155 ;
      RECT 0 27.855 26.58 28.005 ;
      RECT 0 27.705 26.73 27.855 ;
      RECT 0 27.555 26.88 27.705 ;
      RECT 0 27.405 27.03 27.555 ;
      RECT 0 27.255 27.18 27.405 ;
      RECT 0 27.105 27.33 27.255 ;
      RECT 0 26.955 27.48 27.105 ;
      RECT 0 26.805 27.63 26.955 ;
      RECT 0 26.655 27.78 26.805 ;
      RECT 0 26.505 27.93 26.655 ;
      RECT 0 26.355 28.08 26.505 ;
      RECT 0 26.205 28.23 26.355 ;
      RECT 0 26.055 28.38 26.205 ;
      RECT 0 25.905 28.53 26.055 ;
      RECT 0 25.755 28.68 25.905 ;
      RECT 0 25.605 28.83 25.755 ;
      RECT 0 25.455 28.98 25.605 ;
      RECT 0 25.305 29.13 25.455 ;
      RECT 0 25.155 29.28 25.305 ;
      RECT 0 25.005 29.43 25.155 ;
      RECT 0 24.855 29.58 25.005 ;
      RECT 0 24.705 29.73 24.855 ;
      RECT 0 24.555 29.88 24.705 ;
      RECT 0 24.405 30.03 24.555 ;
      RECT 0 24.255 30.18 24.405 ;
      RECT 0 24.105 30.33 24.255 ;
      RECT 0 23.955 30.48 24.105 ;
      RECT 0 23.805 30.63 23.955 ;
      RECT 0 23.655 30.78 23.805 ;
      RECT 0 23.505 30.93 23.655 ;
      RECT 0 23.355 31.08 23.505 ;
      RECT 0 23.205 31.23 23.355 ;
      RECT 0 23.055 31.38 23.205 ;
      RECT 0 22.905 31.53 23.055 ;
      RECT 0 22.755 31.68 22.905 ;
      RECT 0 22.605 31.83 22.755 ;
      RECT 0 22.455 31.98 22.605 ;
      RECT 0 22.305 32.13 22.455 ;
      RECT 0 22.155 32.28 22.305 ;
      RECT 0 22.005 32.43 22.155 ;
      RECT 0 21.855 32.58 22.005 ;
      RECT 0 21.705 32.73 21.855 ;
      RECT 0 21.555 32.88 21.705 ;
      RECT 0 21.405 33.03 21.555 ;
      RECT 0 21.255 33.18 21.405 ;
      RECT 0 21.105 33.33 21.255 ;
      RECT 0 20.955 33.48 21.105 ;
      RECT 0 20.805 33.63 20.955 ;
      RECT 0 20.655 33.78 20.805 ;
      RECT 0 20.505 33.93 20.655 ;
      RECT 0 20.355 34.08 20.505 ;
      RECT 0 20.205 34.23 20.355 ;
      RECT 0 20.055 34.38 20.205 ;
      RECT 0 19.905 34.53 20.055 ;
      RECT 0 19.755 34.68 19.905 ;
      RECT 0 19.605 34.83 19.755 ;
      RECT 0 19.455 34.98 19.605 ;
      RECT 0 19.305 35.13 19.455 ;
      RECT 0 19.155 35.28 19.305 ;
      RECT 0 19.005 35.43 19.155 ;
      RECT 0 18.855 35.58 19.005 ;
      RECT 0 18.705 35.73 18.855 ;
      RECT 0 18.555 35.88 18.705 ;
      RECT 0 18.405 36.03 18.555 ;
      RECT 0 18.255 36.18 18.405 ;
      RECT 0 18.105 36.33 18.255 ;
      RECT 0 17.955 36.48 18.105 ;
      RECT 0 17.805 36.63 17.955 ;
      RECT 0 17.655 36.78 17.805 ;
      RECT 0 17.505 36.93 17.655 ;
      RECT 0 17.355 37.08 17.505 ;
      RECT 0 17.205 37.23 17.355 ;
      RECT 0 17.055 37.38 17.205 ;
      RECT 0 16.905 37.53 17.055 ;
      RECT 0 16.755 37.68 16.905 ;
      RECT 0 16.605 37.83 16.755 ;
      RECT 0 16.455 37.98 16.605 ;
      RECT 0 16.305 38.13 16.455 ;
      RECT 0 16.155 38.28 16.305 ;
      RECT 32.91 35.505 75 35.62 ;
      RECT 33.06 35.355 75 35.505 ;
      RECT 33.21 35.205 75 35.355 ;
      RECT 33.36 35.055 75 35.205 ;
      RECT 33.51 34.905 75 35.055 ;
      RECT 33.66 34.755 75 34.905 ;
      RECT 33.81 34.605 75 34.755 ;
      RECT 33.96 34.455 75 34.605 ;
      RECT 34.11 34.305 75 34.455 ;
      RECT 34.26 34.155 75 34.305 ;
      RECT 21.03 135.82 23.91 135.97 ;
      RECT 20.88 135.97 23.91 136.12 ;
      RECT 20.73 136.12 23.91 136.14 ;
      RECT 31.12 135.65 33.83 135.8 ;
      RECT 30.97 135.8 33.83 135.95 ;
      RECT 30.82 135.95 33.83 136.1 ;
      RECT 30.67 136.1 33.83 136.14 ;
      RECT 36.08 135.67 38.79 135.82 ;
      RECT 35.93 135.82 38.79 135.97 ;
      RECT 35.78 135.97 38.79 136.12 ;
      RECT 35.63 136.12 38.79 136.14 ;
      RECT 11.26 65.455 14.47 65.47 ;
      RECT 11.26 65.47 14.485 65.485 ;
      RECT 0 119.14 9.36 119.29 ;
      RECT 0 119.29 9.21 119.44 ;
      RECT 0 119.44 9.06 119.59 ;
      RECT 0 119.59 8.91 119.74 ;
      RECT 0 119.74 8.76 119.89 ;
      RECT 0 119.89 8.61 120.04 ;
      RECT 0 120.04 8.46 120.19 ;
      RECT 0 120.19 8.31 120.34 ;
      RECT 0 120.34 8.16 120.49 ;
      RECT 0 120.49 8.01 120.64 ;
      RECT 0 120.64 7.86 120.79 ;
      RECT 0 120.79 7.71 120.94 ;
      RECT 0 120.94 7.56 121.09 ;
      RECT 0 121.09 7.41 121.24 ;
      RECT 0 121.24 7.26 121.39 ;
      RECT 0 121.39 7.11 121.54 ;
      RECT 0 121.54 6.96 121.69 ;
      RECT 0 121.69 6.81 121.84 ;
      RECT 0 121.84 6.66 121.99 ;
      RECT 0 121.99 6.51 122.14 ;
      RECT 0 122.14 6.36 122.29 ;
      RECT 0 122.29 6.21 122.44 ;
      RECT 0 122.44 6.06 122.59 ;
      RECT 0 122.59 5.91 122.74 ;
      RECT 0 122.74 5.76 122.89 ;
      RECT 0 122.89 5.61 123.04 ;
      RECT 0 123.04 5.46 123.19 ;
      RECT 0 123.19 5.31 123.34 ;
      RECT 0 123.34 5.16 123.49 ;
      RECT 0 123.49 5.01 123.64 ;
      RECT 0 123.64 4.86 123.79 ;
      RECT 0 123.79 4.71 123.94 ;
      RECT 0 123.94 4.645 124.005 ;
      RECT 0 61.7 9.51 61.825 ;
      RECT 0 61.55 9.635 61.7 ;
      RECT 0 61.4 9.785 61.55 ;
      RECT 0 61.25 9.935 61.4 ;
      RECT 0 61.1 10.085 61.25 ;
      RECT 0 60.95 10.235 61.1 ;
      RECT 0 60.8 10.385 60.95 ;
      RECT 0 60.65 10.535 60.8 ;
      RECT 0 60.5 10.685 60.65 ;
      RECT 0 60.35 10.835 60.5 ;
      RECT 0 60.2 10.985 60.35 ;
      RECT 0 60.05 11.135 60.2 ;
      RECT 0 59.9 11.285 60.05 ;
      RECT 0 59.75 11.435 59.9 ;
      RECT 0 59.6 11.585 59.75 ;
      RECT 0 59.45 11.735 59.6 ;
      RECT 0 59.3 11.885 59.45 ;
      RECT 0 59.15 12.035 59.3 ;
      RECT 0 59 12.185 59.15 ;
      RECT 0 58.85 12.335 59 ;
      RECT 0 58.7 12.485 58.85 ;
      RECT 0 58.55 12.635 58.7 ;
      RECT 0 58.4 12.785 58.55 ;
      RECT 0 58.25 12.935 58.4 ;
      RECT 0 58.1 13.085 58.25 ;
      RECT 0 57.95 13.235 58.1 ;
      RECT 0 57.8 13.385 57.95 ;
      RECT 0 57.65 13.535 57.8 ;
      RECT 0 57.5 13.685 57.65 ;
      RECT 0 57.35 13.835 57.5 ;
      RECT 0 57.2 13.985 57.35 ;
      RECT 0 57.05 14.135 57.2 ;
      RECT 0 56.9 14.285 57.05 ;
      RECT 0 56.75 14.435 56.9 ;
      RECT 0 56.6 14.585 56.75 ;
      RECT 0 56.45 14.735 56.6 ;
      RECT 0 56.3 14.885 56.45 ;
      RECT 0 56.15 15.035 56.3 ;
      RECT 0 56 15.185 56.15 ;
      RECT 0 55.85 15.335 56 ;
      RECT 0 55.7 15.485 55.85 ;
      RECT 0 55.55 15.635 55.7 ;
      RECT 0 55.4 15.785 55.55 ;
      RECT 0 55.25 15.935 55.4 ;
      RECT 0 55.1 16.085 55.25 ;
      RECT 0 54.95 16.235 55.1 ;
      RECT 0 54.8 16.385 54.95 ;
      RECT 0 54.65 16.535 54.8 ;
      RECT 0 54.5 16.685 54.65 ;
      RECT 0 54.35 16.835 54.5 ;
      RECT 0 54.2 16.985 54.35 ;
      RECT 0 54.05 17.135 54.2 ;
      RECT 0 53.9 17.285 54.05 ;
      RECT 0 53.75 17.435 53.9 ;
      RECT 0 53.6 17.585 53.75 ;
      RECT 0 53.45 17.735 53.6 ;
      RECT 0 53.3 17.885 53.45 ;
      RECT 0 53.15 18.035 53.3 ;
      RECT 0 53 18.185 53.15 ;
      RECT 0 52.85 18.335 53 ;
      RECT 0 52.7 18.485 52.85 ;
      RECT 0 52.55 18.635 52.7 ;
      RECT 0 52.4 18.785 52.55 ;
      RECT 0 52.25 18.935 52.4 ;
      RECT 0 52.1 19.085 52.25 ;
      RECT 0 51.95 19.235 52.1 ;
      RECT 0 51.8 19.385 51.95 ;
      RECT 0 51.65 19.535 51.8 ;
      RECT 0 51.5 19.685 51.65 ;
      RECT 0 51.35 19.835 51.5 ;
      RECT 0 51.2 19.985 51.35 ;
      RECT 0 51.05 20.135 51.2 ;
      RECT 0 50.9 20.285 51.05 ;
      RECT 0 34.005 20.435 34.15 ;
      RECT 0 33.855 20.58 34.005 ;
      RECT 0 33.705 20.73 33.855 ;
      RECT 0 33.555 20.88 33.705 ;
      RECT 0 19.305 35.13 19.455 ;
      RECT 0 19.155 35.28 19.305 ;
      RECT 0 19.005 35.43 19.155 ;
      RECT 0 18.855 35.58 19.005 ;
      RECT 0 18.705 35.73 18.855 ;
      RECT 0 18.555 35.88 18.705 ;
      RECT 0 18.405 36.03 18.555 ;
      RECT 0 18.255 36.18 18.405 ;
      RECT 0 18.105 36.33 18.255 ;
      RECT 0 17.955 36.48 18.105 ;
      RECT 0 17.805 36.63 17.955 ;
      RECT 0 17.655 36.78 17.805 ;
      RECT 0 17.505 36.93 17.655 ;
      RECT 0 17.355 37.08 17.505 ;
      RECT 0 17.205 37.23 17.355 ;
      RECT 0 17.055 37.38 17.205 ;
      RECT 0 16.905 37.53 17.055 ;
      RECT 0 16.755 37.68 16.905 ;
      RECT 0 16.605 37.83 16.755 ;
      RECT 0 16.455 37.98 16.605 ;
      RECT 0 16.305 38.13 16.455 ;
      RECT 0 16.155 38.28 16.305 ;
      RECT 21.83 64.835 23.75 64.985 ;
      RECT 21.68 64.985 23.9 65.135 ;
      RECT 21.53 65.135 24.05 65.285 ;
      RECT 21.38 65.285 24.2 65.435 ;
      RECT 21.23 65.435 24.35 65.485 ;
      RECT 31.77 64.835 33.67 64.985 ;
      RECT 31.62 64.985 33.82 65.135 ;
      RECT 31.47 65.135 33.97 65.285 ;
      RECT 31.32 65.285 34.12 65.435 ;
      RECT 31.17 65.435 34.27 65.485 ;
      RECT 16.22 65.455 19.43 65.47 ;
      RECT 16.22 65.47 19.445 65.485 ;
      RECT 16.84 64.835 18.81 64.985 ;
      RECT 16.69 64.985 18.96 65.135 ;
      RECT 16.54 65.135 19.11 65.285 ;
      RECT 16.39 65.285 19.26 65.435 ;
      RECT 16.24 65.435 19.41 65.455 ;
      RECT 36.73 64.835 38.65 64.985 ;
      RECT 36.58 64.985 38.8 65.135 ;
      RECT 36.43 65.135 38.95 65.285 ;
      RECT 36.28 65.285 39.1 65.435 ;
      RECT 36.13 65.435 39.25 65.485 ;
      RECT 26.16 65.465 29.34 65.475 ;
      RECT 26.16 65.475 29.35 65.485 ;
      RECT 26.79 64.835 28.71 64.985 ;
      RECT 26.64 64.985 28.86 65.135 ;
      RECT 26.49 65.135 29.01 65.285 ;
      RECT 26.34 65.285 29.16 65.435 ;
      RECT 26.19 65.435 29.31 65.465 ;
      RECT 36.08 135.67 38.79 135.82 ;
      RECT 35.93 135.82 38.79 135.97 ;
      RECT 35.78 135.97 38.79 136.12 ;
      RECT 35.63 136.12 38.79 136.14 ;
      RECT 36.08 132.955 39.15 133.105 ;
      RECT 36.08 133.105 39.0 133.255 ;
      RECT 36.08 133.255 38.85 133.405 ;
      RECT 36.08 133.405 38.79 133.465 ;
      RECT 26.16 135.67 28.87 135.82 ;
      RECT 26.01 135.82 28.87 135.97 ;
      RECT 25.86 135.97 28.87 136.12 ;
      RECT 25.71 136.12 28.87 136.16 ;
      RECT 26.16 132.975 29.21 133.125 ;
      RECT 26.16 133.125 29.06 133.275 ;
      RECT 26.16 133.275 28.91 133.425 ;
      RECT 26.16 133.425 28.87 133.465 ;
      RECT 21.18 135.67 23.91 135.82 ;
      RECT 21.03 135.82 23.91 135.97 ;
      RECT 20.88 135.97 23.91 136.12 ;
      RECT 20.73 136.12 23.91 136.14 ;
      RECT 21.18 132.995 24.25 133.145 ;
      RECT 21.18 133.145 24.1 133.295 ;
      RECT 21.18 133.295 23.95 133.445 ;
      RECT 21.18 133.445 23.91 133.485 ;
      RECT 31.12 135.65 33.83 135.8 ;
      RECT 30.97 135.8 33.83 135.95 ;
      RECT 30.82 135.95 33.83 136.1 ;
      RECT 30.67 136.1 33.83 136.14 ;
      RECT 31.12 132.995 34.17 133.145 ;
      RECT 31.12 133.145 34.02 133.295 ;
      RECT 31.12 133.295 33.87 133.445 ;
      RECT 31.12 133.445 33.83 133.485 ;
      RECT 16.22 134.455 18.95 134.605 ;
      RECT 16.07 134.605 18.95 134.755 ;
      RECT 15.92 134.755 18.95 134.905 ;
      RECT 15.77 134.905 18.95 134.925 ;
      RECT 16.22 132.955 19.31 133.105 ;
      RECT 16.22 133.105 19.16 133.255 ;
      RECT 16.22 133.255 19.01 133.405 ;
      RECT 16.22 133.405 18.95 133.465 ;
      RECT 11.88 64.835 13.85 64.985 ;
      RECT 11.73 64.985 14.0 65.135 ;
      RECT 11.58 65.135 14.15 65.285 ;
      RECT 11.43 65.285 14.3 65.435 ;
      RECT 11.28 65.435 14.45 65.455 ;
      RECT 16.84 64.835 18.81 64.985 ;
      RECT 16.69 64.985 18.96 65.135 ;
      RECT 16.54 65.135 19.11 65.285 ;
      RECT 16.39 65.285 19.26 65.435 ;
      RECT 16.24 65.435 19.41 65.455 ;
      RECT 26.79 64.835 28.71 64.985 ;
      RECT 26.64 64.985 28.86 65.135 ;
      RECT 26.49 65.135 29.01 65.285 ;
      RECT 26.34 65.285 29.16 65.435 ;
      RECT 26.19 65.435 29.31 65.465 ;
      RECT 26.16 135.67 28.87 135.82 ;
      RECT 26.01 135.82 28.87 135.97 ;
      RECT 25.86 135.97 28.87 136.12 ;
      RECT 25.71 136.12 28.87 136.16 ;
      RECT 21.18 135.67 23.91 135.82 ;
      RECT 44.01 24.405 75 24.555 ;
      RECT 44.16 24.255 75 24.405 ;
      RECT 44.31 24.105 75 24.255 ;
      RECT 44.46 23.955 75 24.105 ;
      RECT 44.61 23.805 75 23.955 ;
      RECT 44.76 23.655 75 23.805 ;
      RECT 44.91 23.505 75 23.655 ;
      RECT 45.06 23.355 75 23.505 ;
      RECT 45.21 23.205 75 23.355 ;
      RECT 45.36 23.055 75 23.205 ;
      RECT 45.51 22.905 75 23.055 ;
      RECT 45.66 22.755 75 22.905 ;
      RECT 45.81 22.605 75 22.755 ;
      RECT 45.96 22.455 75 22.605 ;
      RECT 46.11 22.305 75 22.455 ;
      RECT 46.26 22.155 75 22.305 ;
      RECT 46.41 22.005 75 22.155 ;
      RECT 46.56 21.855 75 22.005 ;
      RECT 46.71 21.705 75 21.855 ;
      RECT 46.86 21.555 75 21.705 ;
      RECT 47.01 21.405 75 21.555 ;
      RECT 47.16 21.255 75 21.405 ;
      RECT 47.31 21.105 75 21.255 ;
      RECT 47.46 20.955 75 21.105 ;
      RECT 47.61 20.805 75 20.955 ;
      RECT 47.76 20.655 75 20.805 ;
      RECT 47.91 20.505 75 20.655 ;
      RECT 48.06 20.355 75 20.505 ;
      RECT 48.21 20.205 75 20.355 ;
      RECT 0 34.005 20.435 34.15 ;
      RECT 0 33.855 20.58 34.005 ;
      RECT 0 33.705 20.73 33.855 ;
      RECT 0 33.555 20.88 33.705 ;
      RECT 0 33.405 21.03 33.555 ;
      RECT 0 33.255 21.18 33.405 ;
      RECT 0 33.105 21.33 33.255 ;
      RECT 0 32.955 21.48 33.105 ;
      RECT 0 32.805 21.63 32.955 ;
      RECT 0 32.655 21.78 32.805 ;
      RECT 0 32.505 21.93 32.655 ;
      RECT 0 32.355 22.08 32.505 ;
      RECT 0 32.205 22.23 32.355 ;
      RECT 0 32.055 22.38 32.205 ;
      RECT 0 31.905 22.53 32.055 ;
      RECT 0 31.755 22.68 31.905 ;
      RECT 0 31.605 22.83 31.755 ;
      RECT 0 31.455 22.98 31.605 ;
      RECT 0 31.305 23.13 31.455 ;
      RECT 0 31.155 23.28 31.305 ;
      RECT 0 31.005 23.43 31.155 ;
      RECT 0 30.855 23.58 31.005 ;
      RECT 0 30.705 23.73 30.855 ;
      RECT 0 30.555 23.88 30.705 ;
      RECT 0 30.405 24.03 30.555 ;
      RECT 0 30.255 24.18 30.405 ;
      RECT 0 30.105 24.33 30.255 ;
      RECT 0 29.955 24.48 30.105 ;
      RECT 0 29.805 24.63 29.955 ;
      RECT 0 29.655 24.78 29.805 ;
      RECT 0 29.505 24.93 29.655 ;
      RECT 0 29.355 25.08 29.505 ;
      RECT 0 29.205 25.23 29.355 ;
      RECT 0 29.055 25.38 29.205 ;
      RECT 0 28.905 25.53 29.055 ;
      RECT 0 28.755 25.68 28.905 ;
      RECT 0 28.605 25.83 28.755 ;
      RECT 0 28.455 25.98 28.605 ;
      RECT 0 28.305 26.13 28.455 ;
      RECT 0 28.155 26.28 28.305 ;
      RECT 0 28.005 26.43 28.155 ;
      RECT 0 27.855 26.58 28.005 ;
      RECT 0 27.705 26.73 27.855 ;
      RECT 0 27.555 26.88 27.705 ;
      RECT 0 27.405 27.03 27.555 ;
      RECT 0 27.255 27.18 27.405 ;
      RECT 0 27.105 27.33 27.255 ;
      RECT 0 26.955 27.48 27.105 ;
      RECT 0 26.805 27.63 26.955 ;
      RECT 0 26.655 27.78 26.805 ;
      RECT 0 26.505 27.93 26.655 ;
      RECT 0 26.355 28.08 26.505 ;
      RECT 0 26.205 28.23 26.355 ;
      RECT 0 26.055 28.38 26.205 ;
      RECT 0 25.905 28.53 26.055 ;
      RECT 0 25.755 28.68 25.905 ;
      RECT 0 25.605 28.83 25.755 ;
      RECT 0 25.455 28.98 25.605 ;
      RECT 0 25.305 29.13 25.455 ;
      RECT 0 25.155 29.28 25.305 ;
      RECT 0 25.005 29.43 25.155 ;
      RECT 0 24.855 29.58 25.005 ;
      RECT 0 24.705 29.73 24.855 ;
      RECT 0 24.555 29.88 24.705 ;
      RECT 0 24.405 30.03 24.555 ;
      RECT 0 24.255 30.18 24.405 ;
      RECT 0 24.105 30.33 24.255 ;
      RECT 0 23.955 30.48 24.105 ;
      RECT 0 23.805 30.63 23.955 ;
      RECT 0 23.655 30.78 23.805 ;
      RECT 0 23.505 30.93 23.655 ;
      RECT 0 23.355 31.08 23.505 ;
      RECT 0 23.205 31.23 23.355 ;
      RECT 0 23.055 31.38 23.205 ;
      RECT 0 22.905 31.53 23.055 ;
      RECT 0 22.755 31.68 22.905 ;
      RECT 0 22.605 31.83 22.755 ;
      RECT 0 22.455 31.98 22.605 ;
      RECT 0 22.305 32.13 22.455 ;
      RECT 0 22.155 32.28 22.305 ;
      RECT 0 22.005 32.43 22.155 ;
      RECT 0 21.855 32.58 22.005 ;
      RECT 0 21.705 32.73 21.855 ;
      RECT 0 21.555 32.88 21.705 ;
      RECT 0 21.405 33.03 21.555 ;
      RECT 0 21.255 33.18 21.405 ;
      RECT 0 21.105 33.33 21.255 ;
      RECT 0 20.955 33.48 21.105 ;
      RECT 0 20.805 33.63 20.955 ;
      RECT 0 20.655 33.78 20.805 ;
      RECT 0 20.505 33.93 20.655 ;
      RECT 0 20.355 34.08 20.505 ;
      RECT 0 20.205 34.23 20.355 ;
      RECT 0 20.055 34.38 20.205 ;
      RECT 0 19.905 34.53 20.055 ;
      RECT 0 19.755 34.68 19.905 ;
      RECT 0 19.605 34.83 19.755 ;
      RECT 0 19.455 34.98 19.605 ;
      RECT 0 58.55 12.635 58.7 ;
      RECT 0 58.4 12.785 58.55 ;
      RECT 0 58.25 12.935 58.4 ;
      RECT 0 58.1 13.085 58.25 ;
      RECT 0 57.95 13.235 58.1 ;
      RECT 0 57.8 13.385 57.95 ;
      RECT 0 57.65 13.535 57.8 ;
      RECT 0 57.5 13.685 57.65 ;
      RECT 0 57.35 13.835 57.5 ;
      RECT 0 57.2 13.985 57.35 ;
      RECT 0 57.05 14.135 57.2 ;
      RECT 0 56.9 14.285 57.05 ;
      RECT 0 56.75 14.435 56.9 ;
      RECT 0 56.6 14.585 56.75 ;
      RECT 0 56.45 14.735 56.6 ;
      RECT 0 56.3 14.885 56.45 ;
      RECT 0 56.15 15.035 56.3 ;
      RECT 0 56 15.185 56.15 ;
      RECT 0 55.85 15.335 56 ;
      RECT 0 55.7 15.485 55.85 ;
      RECT 0 55.55 15.635 55.7 ;
      RECT 0 55.4 15.785 55.55 ;
      RECT 0 55.25 15.935 55.4 ;
      RECT 0 55.1 16.085 55.25 ;
      RECT 0 54.95 16.235 55.1 ;
      RECT 0 54.8 16.385 54.95 ;
      RECT 0 54.65 16.535 54.8 ;
      RECT 0 54.5 16.685 54.65 ;
      RECT 0 54.35 16.835 54.5 ;
      RECT 0 54.2 16.985 54.35 ;
      RECT 0 54.05 17.135 54.2 ;
      RECT 0 53.9 17.285 54.05 ;
      RECT 0 53.75 17.435 53.9 ;
      RECT 0 53.6 17.585 53.75 ;
      RECT 0 53.45 17.735 53.6 ;
      RECT 0 53.3 17.885 53.45 ;
      RECT 0 53.15 18.035 53.3 ;
      RECT 0 53 18.185 53.15 ;
      RECT 0 52.85 18.335 53 ;
      RECT 0 52.7 18.485 52.85 ;
      RECT 0 52.55 18.635 52.7 ;
      RECT 0 52.4 18.785 52.55 ;
      RECT 0 52.25 18.935 52.4 ;
      RECT 0 52.1 19.085 52.25 ;
      RECT 0 51.95 19.235 52.1 ;
      RECT 0 51.8 19.385 51.95 ;
      RECT 0 51.65 19.535 51.8 ;
      RECT 0 51.5 19.685 51.65 ;
      RECT 0 51.35 19.835 51.5 ;
      RECT 0 51.2 19.985 51.35 ;
      RECT 0 51.05 20.135 51.2 ;
      RECT 0 50.9 20.285 51.05 ;
      RECT 32.91 35.505 75 35.62 ;
      RECT 33.06 35.355 75 35.505 ;
      RECT 33.21 35.205 75 35.355 ;
      RECT 33.36 35.055 75 35.205 ;
      RECT 33.51 34.905 75 35.055 ;
      RECT 33.66 34.755 75 34.905 ;
      RECT 33.81 34.605 75 34.755 ;
      RECT 33.96 34.455 75 34.605 ;
      RECT 34.11 34.305 75 34.455 ;
      RECT 34.26 34.155 75 34.305 ;
      RECT 34.41 34.005 75 34.155 ;
      RECT 34.56 33.855 75 34.005 ;
      RECT 34.71 33.705 75 33.855 ;
      RECT 34.86 33.555 75 33.705 ;
      RECT 35.01 33.405 75 33.555 ;
      RECT 35.16 33.255 75 33.405 ;
      RECT 35.31 33.105 75 33.255 ;
      RECT 35.46 32.955 75 33.105 ;
      RECT 35.61 32.805 75 32.955 ;
      RECT 35.76 32.655 75 32.805 ;
      RECT 35.91 32.505 75 32.655 ;
      RECT 36.06 32.355 75 32.505 ;
      RECT 36.21 32.205 75 32.355 ;
      RECT 36.36 32.055 75 32.205 ;
      RECT 36.51 31.905 75 32.055 ;
      RECT 36.66 31.755 75 31.905 ;
      RECT 36.81 31.605 75 31.755 ;
      RECT 36.96 31.455 75 31.605 ;
      RECT 37.11 31.305 75 31.455 ;
      RECT 37.26 31.155 75 31.305 ;
      RECT 37.41 31.005 75 31.155 ;
      RECT 37.56 30.855 75 31.005 ;
      RECT 37.71 30.705 75 30.855 ;
      RECT 37.86 30.555 75 30.705 ;
      RECT 38.01 30.405 75 30.555 ;
      RECT 38.16 30.255 75 30.405 ;
      RECT 38.31 30.105 75 30.255 ;
      RECT 38.46 29.955 75 30.105 ;
      RECT 38.61 29.805 75 29.955 ;
      RECT 38.76 29.655 75 29.805 ;
      RECT 38.91 29.505 75 29.655 ;
      RECT 39.06 29.355 75 29.505 ;
      RECT 39.21 29.205 75 29.355 ;
      RECT 39.36 29.055 75 29.205 ;
      RECT 39.51 28.905 75 29.055 ;
      RECT 39.66 28.755 75 28.905 ;
      RECT 39.81 28.605 75 28.755 ;
      RECT 39.96 28.455 75 28.605 ;
      RECT 40.11 28.305 75 28.455 ;
      RECT 40.26 28.155 75 28.305 ;
      RECT 40.41 28.005 75 28.155 ;
      RECT 40.56 27.855 75 28.005 ;
      RECT 40.71 27.705 75 27.855 ;
      RECT 40.86 27.555 75 27.705 ;
      RECT 41.01 27.405 75 27.555 ;
      RECT 41.16 27.255 75 27.405 ;
      RECT 41.31 27.105 75 27.255 ;
      RECT 41.46 26.955 75 27.105 ;
      RECT 41.61 26.805 75 26.955 ;
      RECT 41.76 26.655 75 26.805 ;
      RECT 41.91 26.505 75 26.655 ;
      RECT 42.06 26.355 75 26.505 ;
      RECT 42.21 26.205 75 26.355 ;
      RECT 42.36 26.055 75 26.205 ;
      RECT 42.51 25.905 75 26.055 ;
      RECT 42.66 25.755 75 25.905 ;
      RECT 42.81 25.605 75 25.755 ;
      RECT 42.96 25.455 75 25.605 ;
      RECT 43.11 25.305 75 25.455 ;
      RECT 43.26 25.155 75 25.305 ;
      RECT 43.41 25.005 75 25.155 ;
      RECT 43.56 24.855 75 25.005 ;
      RECT 43.71 24.705 75 24.855 ;
      RECT 43.86 24.555 75 24.705 ;
      RECT 10.79 132.155 14.35 132.305 ;
      RECT 10.79 132.305 14.2 132.455 ;
      RECT 10.79 132.455 14.05 132.605 ;
      RECT 10.79 132.605 13.99 132.665 ;
      RECT 11.26 122.785 14.5 122.935 ;
      RECT 11.11 122.935 14.5 123.085 ;
      RECT 10.96 123.085 14.5 123.235 ;
      RECT 10.81 123.235 14.5 123.255 ;
      RECT 0 119.14 9.36 119.29 ;
      RECT 0 119.29 9.21 119.44 ;
      RECT 0 119.44 9.06 119.59 ;
      RECT 0 119.59 8.91 119.74 ;
      RECT 0 119.74 8.76 119.89 ;
      RECT 0 119.89 8.61 120.04 ;
      RECT 0 120.04 8.46 120.19 ;
      RECT 0 120.19 8.31 120.34 ;
      RECT 0 120.34 8.16 120.49 ;
      RECT 0 120.49 8.01 120.64 ;
      RECT 0 120.64 7.86 120.79 ;
      RECT 0 120.79 7.71 120.94 ;
      RECT 0 120.94 7.56 121.09 ;
      RECT 0 121.09 7.41 121.24 ;
      RECT 0 121.24 7.26 121.39 ;
      RECT 0 121.39 7.11 121.54 ;
      RECT 0 121.54 6.96 121.69 ;
      RECT 0 121.69 6.81 121.84 ;
      RECT 0 121.84 6.66 121.99 ;
      RECT 0 121.99 6.51 122.14 ;
      RECT 0 122.14 6.36 122.29 ;
      RECT 0 122.29 6.21 122.44 ;
      RECT 0 122.44 6.06 122.59 ;
      RECT 0 122.59 5.91 122.74 ;
      RECT 0 122.74 5.76 122.89 ;
      RECT 0 122.89 5.61 123.04 ;
      RECT 0 123.04 5.46 123.19 ;
      RECT 0 123.19 5.31 123.34 ;
      RECT 0 123.34 5.16 123.49 ;
      RECT 0 123.49 5.01 123.64 ;
      RECT 0 123.64 4.86 123.79 ;
      RECT 0 123.79 4.71 123.94 ;
      RECT 0 123.94 4.645 124.005 ;
      RECT 11.26 65.455 14.47 65.47 ;
      RECT 11.26 65.47 14.485 65.485 ;
      RECT 11.88 64.835 13.85 64.985 ;
      RECT 11.73 64.985 14.0 65.135 ;
      RECT 11.58 65.135 14.15 65.285 ;
      RECT 11.43 65.285 14.3 65.435 ;
      RECT 11.28 65.435 14.45 65.455 ;
      RECT 32.945 52.26 75 52.41 ;
      RECT 33.095 52.41 75 52.56 ;
      RECT 33.245 52.56 75 52.71 ;
      RECT 33.395 52.71 75 52.86 ;
      RECT 33.545 52.86 75 53.01 ;
      RECT 33.695 53.01 75 53.16 ;
      RECT 33.845 53.16 75 53.31 ;
      RECT 33.995 53.31 75 53.46 ;
      RECT 34.145 53.46 75 53.61 ;
      RECT 34.295 53.61 75 53.76 ;
      RECT 34.445 53.76 75 53.91 ;
      RECT 34.595 53.91 75 54.06 ;
      RECT 34.745 54.06 75 54.21 ;
      RECT 34.895 54.21 75 54.36 ;
      RECT 35.045 54.36 75 54.51 ;
      RECT 35.195 54.51 75 54.66 ;
      RECT 35.345 54.66 75 54.81 ;
      RECT 35.495 54.81 75 54.96 ;
      RECT 35.645 54.96 75 55.11 ;
      RECT 35.795 55.11 75 55.26 ;
      RECT 35.945 55.26 75 55.41 ;
      RECT 36.095 55.41 75 55.56 ;
      RECT 36.245 55.56 75 55.71 ;
      RECT 36.395 55.71 75 55.86 ;
      RECT 36.545 55.86 75 56.01 ;
      RECT 36.695 56.01 75 56.16 ;
      RECT 36.845 56.16 75 56.31 ;
      RECT 36.995 56.31 75 56.46 ;
      RECT 37.145 56.46 75 56.61 ;
      RECT 37.295 56.61 75 56.76 ;
      RECT 37.445 56.76 75 56.91 ;
      RECT 37.595 56.91 75 57.06 ;
      RECT 37.745 57.06 75 57.21 ;
      RECT 37.895 57.21 75 57.36 ;
      RECT 38.045 57.36 75 57.51 ;
      RECT 38.195 57.51 75 57.66 ;
      RECT 38.345 57.66 75 57.81 ;
      RECT 38.495 57.81 75 57.96 ;
      RECT 38.645 57.96 75 58.11 ;
      RECT 38.795 58.11 75 58.26 ;
      RECT 38.945 58.26 75 58.41 ;
      RECT 39.095 58.41 75 58.56 ;
      RECT 39.245 58.56 75 58.71 ;
      RECT 39.395 58.71 75 58.86 ;
      RECT 39.545 58.86 75 59.01 ;
      RECT 39.695 59.01 75 59.16 ;
      RECT 39.845 59.16 75 59.31 ;
      RECT 39.995 59.31 75 59.46 ;
      RECT 40.145 59.46 75 59.61 ;
      RECT 40.295 59.61 75 59.76 ;
      RECT 40.445 59.76 75 59.91 ;
      RECT 40.595 59.91 75 60.06 ;
      RECT 40.745 60.06 75 60.21 ;
      RECT 40.895 60.21 75 60.36 ;
      RECT 41.02 60.36 75 60.485 ;
      RECT 0 61.7 9.51 61.825 ;
      RECT 0 61.55 9.635 61.7 ;
      RECT 0 61.4 9.785 61.55 ;
      RECT 0 61.25 9.935 61.4 ;
      RECT 0 61.1 10.085 61.25 ;
      RECT 0 60.95 10.235 61.1 ;
      RECT 0 60.8 10.385 60.95 ;
      RECT 0 60.65 10.535 60.8 ;
      RECT 0 60.5 10.685 60.65 ;
      RECT 0 60.35 10.835 60.5 ;
      RECT 0 60.2 10.985 60.35 ;
      RECT 0 60.05 11.135 60.2 ;
      RECT 0 59.9 11.285 60.05 ;
      RECT 0 59.75 11.435 59.9 ;
      RECT 0 59.6 11.585 59.75 ;
      RECT 0 59.45 11.735 59.6 ;
      RECT 0 59.3 11.885 59.45 ;
      RECT 0 59.15 12.035 59.3 ;
      RECT 0 59 12.185 59.15 ;
      RECT 0 58.85 12.335 59 ;
      RECT 0 58.7 12.485 58.85 ;
      RECT 36.08 133.465 38.79 135.67 ;
      RECT 26.16 133.465 28.87 135.67 ;
      RECT 21.18 133.485 23.91 135.67 ;
      RECT 31.12 133.485 33.83 135.65 ;
      RECT 16.22 133.465 18.95 134.455 ;
      RECT 36.08 133.465 38.79 135.67 ;
      RECT 26.16 133.465 28.87 135.67 ;
      RECT 21.18 133.485 23.91 135.67 ;
      RECT 31.12 133.485 33.83 135.65 ;
      RECT 16.22 133.465 18.95 134.455 ;
      RECT 25.67 136.16 28.87 171.525 ;
      RECT 20.71 136.14 23.91 171.525 ;
      RECT 30.63 136.14 33.83 171.525 ;
      RECT 35.61 136.14 38.79 171.525 ;
      RECT 0 124.005 4.405 141.99 ;
      RECT 11.26 65.485 14.5 122.785 ;
      RECT 0 61.825 9.51 119.14 ;
      RECT 32.795 35.62 75 52.26 ;
      RECT 0 34.15 20.435 50.9 ;
      RECT 0 0 38.43 16.155 ;
      RECT 48.21 0 75 20.205 ;
      RECT 21.18 65.485 24.4 132.995 ;
      RECT 31.12 65.485 34.32 132.995 ;
      RECT 16.22 65.485 19.46 132.955 ;
      RECT 36.08 65.485 39.3 132.955 ;
      RECT 26.16 65.485 29.36 132.975 ;
      RECT 15.75 134.925 18.95 198 ;
      RECT 15.75 134.925 18.95 171.525 ;
      RECT 0 146.615 9.03 198 ;
      RECT 0 146.615 9.03 169.62 ;
      RECT 0 171.525 75 198 ;
      RECT 40.55 136.14 75 171.525 ;
      RECT 41.02 60.485 75 171.525 ;
      RECT 41.02 60.485 75 135.67 ;
      RECT 0 169.62 13.99 198 ;
      RECT 0 169.62 13.99 171.525 ;
      RECT 10.79 132.665 13.99 198 ;
      RECT 10.79 132.665 13.99 169.62 ;
      RECT 10.79 123.255 13.99 169.62 ;
      RECT 10.79 123.255 14.5 132.155 ;
      RECT 0 146.49 8.905 146.615 ;
      RECT 0 146.34 8.755 146.49 ;
      RECT 0 146.19 8.605 146.34 ;
      RECT 0 146.04 8.455 146.19 ;
      RECT 0 145.89 8.305 146.04 ;
      RECT 0 145.74 8.155 145.89 ;
      RECT 0 145.59 8.005 145.74 ;
      RECT 0 145.44 7.855 145.59 ;
      RECT 0 145.29 7.705 145.44 ;
      RECT 0 145.14 7.555 145.29 ;
      RECT 0 144.99 7.405 145.14 ;
      RECT 0 144.84 7.255 144.99 ;
      RECT 0 144.69 7.105 144.84 ;
      RECT 0 144.54 6.955 144.69 ;
      RECT 0 144.39 6.805 144.54 ;
      RECT 0 144.24 6.655 144.39 ;
      RECT 0 144.09 6.505 144.24 ;
      RECT 0 143.94 6.355 144.09 ;
      RECT 0 143.79 6.205 143.94 ;
      RECT 0 143.64 6.055 143.79 ;
      RECT 0 143.49 5.905 143.64 ;
      RECT 0 143.34 5.755 143.49 ;
      RECT 0 143.19 5.605 143.34 ;
      RECT 0 143.04 5.455 143.19 ;
      RECT 0 142.89 5.305 143.04 ;
      RECT 0 142.74 5.155 142.89 ;
      RECT 0 142.59 5.005 142.74 ;
      RECT 0 142.44 4.855 142.59 ;
      RECT 0 142.29 4.705 142.44 ;
      RECT 0 142.14 4.555 142.29 ;
      RECT 0 141.99 4.405 142.14 ;
      RECT 41.02 135.67 75 135.82 ;
      RECT 40.87 135.82 75 135.97 ;
      RECT 40.72 135.97 75 136.12 ;
      RECT 40.57 136.12 75 136.14 ;
    LAYER li1 ;
      RECT 34.46 147.22 34.99 147.32 ;
      RECT 38.31 146.19 38.91 162.235 ;
      RECT 40.46 146.19 41.06 161.705 ;
      RECT 40.46 161.705 41.1 162.235 ;
      RECT 39.235 147.32 40.135 160.075 ;
      RECT 39.42 147.22 39.95 147.32 ;
      RECT 43.27 146.19 43.87 162.235 ;
      RECT 45.42 146.19 46.02 162.235 ;
      RECT 44.195 147.32 45.095 160.075 ;
      RECT 44.38 147.22 44.91 147.32 ;
      RECT 41.57 147.085 42.76 160.075 ;
      RECT 48.23 146.19 48.83 162.235 ;
      RECT 46.53 147.085 47.72 160.075 ;
      RECT 49.155 147.32 50.055 160.075 ;
      RECT 49.34 147.22 49.87 147.32 ;
      RECT 50.38 146.19 50.98 162.235 ;
      RECT 53.19 146.19 53.79 162.235 ;
      RECT 51.49 147.085 52.68 160.075 ;
      RECT 55.34 146.19 55.94 162.235 ;
      RECT 56.45 147.085 57.64 160.075 ;
      RECT 54.115 147.32 55.015 160.075 ;
      RECT 54.3 147.22 54.83 147.32 ;
      RECT 58.15 146.19 58.75 162.235 ;
      RECT 60.3 146.19 60.9 162.235 ;
      RECT 61.41 147.085 62.6 160.075 ;
      RECT 59.075 147.32 59.975 160.075 ;
      RECT 59.26 147.22 59.79 147.32 ;
      RECT 65.26 146.19 65.86 162.235 ;
      RECT 63.11 146.19 63.71 162.235 ;
      RECT 66.37 147.085 67.56 160.075 ;
      RECT 64.035 147.32 64.935 160.075 ;
      RECT 64.22 147.22 64.75 147.32 ;
      RECT 70.22 146.19 70.82 162.235 ;
      RECT 68.07 146.19 68.67 162.235 ;
      RECT 68.995 147.32 69.895 160.075 ;
      RECT 69.18 147.22 69.71 147.32 ;
      RECT 0.295 137.815 74.41 141.445 ;
      RECT 0.27 143.105 1.12 166.005 ;
      RECT 73.51 143.105 74.91 166.005 ;
      RECT 0.27 142.215 74.91 143.105 ;
      RECT 0.27 166.005 74.91 166.895 ;
      RECT 0.985 89.275 73.86 92.945 ;
      RECT -0.205 125.9 41.52 127.225 ;
      RECT 62.04 125.9 74.915 127.22 ;
      RECT -0.205 94.575 58.735 96.65 ;
      RECT 62.04 127.22 74.41 127.225 ;
      RECT 72.3 94.575 74.915 96.65 ;
      RECT 0.265 100.32 1.305 122.315 ;
      RECT -0.085 99.395 74.915 99.42 ;
      RECT 73.695 100.32 74.915 122.315 ;
      RECT -0.205 92.945 74.915 94.575 ;
      RECT -0.205 123.24 74.915 125.9 ;
      RECT -0.205 96.65 74.915 99.395 ;
      RECT 0.265 99.42 74.915 100.32 ;
      RECT 0.265 122.315 74.915 123.24 ;
      RECT 59.12 95.42 60.135 95.65 ;
      RECT 59.12 95.65 60.13 95.75 ;
      RECT 70.17 95.295 71.18 95.935 ;
      RECT 2.07 120.09 72.925 121.09 ;
      RECT 2.07 101.16 72.925 102.16 ;
      RECT 2.07 102.16 3.56 120.09 ;
      RECT 71.44 102.16 72.925 120.09 ;
      RECT 6.215 103.545 6.815 119.445 ;
      RECT 4.99 105.565 5.89 118.315 ;
      RECT 4.065 103.545 4.665 119.445 ;
      RECT 7.325 105.505 8.515 118.415 ;
      RECT 9.025 103.545 9.625 119.445 ;
      RECT 11.175 103.545 11.775 119.445 ;
      RECT 9.95 105.565 10.85 118.315 ;
      RECT 13.985 103.545 14.585 119.445 ;
      RECT 16.135 103.545 16.735 119.445 ;
      RECT 12.285 105.505 13.475 118.415 ;
      RECT 14.91 105.565 15.81 118.315 ;
      RECT 18.945 103.545 19.545 119.445 ;
      RECT 17.245 105.505 18.435 118.415 ;
      RECT 19.87 105.565 20.77 118.315 ;
      RECT 23.905 103.545 24.505 119.445 ;
      RECT 21.095 103.545 21.695 119.445 ;
      RECT 22.205 105.505 23.395 118.415 ;
      RECT 26.055 103.545 26.655 119.445 ;
      RECT 28.865 103.545 29.465 119.445 ;
      RECT 27.165 105.505 28.355 118.415 ;
      RECT 24.83 105.565 25.73 118.315 ;
      RECT 31.015 103.545 31.615 119.445 ;
      RECT 32.125 105.505 33.315 118.415 ;
      RECT 29.79 105.565 30.69 118.315 ;
      RECT 33.825 103.545 34.425 119.445 ;
      RECT 35.975 103.545 36.575 119.445 ;
      RECT 34.75 105.565 35.65 118.315 ;
      RECT 37.085 105.505 38.275 118.415 ;
      RECT 38.785 103.545 39.385 119.445 ;
      RECT 40.935 103.545 41.535 119.445 ;
      RECT 39.71 105.565 40.61 118.315 ;
      RECT 43.745 103.545 44.345 119.445 ;
      RECT 44.67 105.565 45.57 118.32 ;
      RECT 42.045 105.505 43.235 118.415 ;
      RECT 48.705 103.545 49.305 119.445 ;
      RECT 45.895 103.545 46.495 119.445 ;
      RECT 49.63 105.565 50.53 118.415 ;
      RECT 47.005 105.505 48.195 118.415 ;
      RECT 53.665 103.545 54.265 119.445 ;
      RECT 50.855 103.545 51.455 119.445 ;
      RECT 51.965 105.505 53.155 118.475 ;
      RECT 55.815 103.545 56.415 119.445 ;
      RECT 54.59 105.565 55.49 118.315 ;
      RECT 56.925 105.505 58.115 118.415 ;
      RECT 58.625 103.545 59.225 119.445 ;
      RECT 60.775 103.545 61.375 119.445 ;
      RECT 59.55 105.565 60.45 118.315 ;
      RECT 61.885 105.505 63.075 118.415 ;
      RECT 65.735 103.545 66.335 119.445 ;
      RECT 63.585 103.545 64.185 119.445 ;
      RECT 64.51 105.565 65.41 118.315 ;
      RECT 68.545 103.545 69.145 119.445 ;
      RECT 70.335 103.545 70.935 119.445 ;
      RECT 69.655 105.565 69.825 118.315 ;
      RECT 66.845 105.505 68.035 118.415 ;
      RECT 1.25 134.585 2.265 134.815 ;
      RECT 1.25 134.815 2.26 134.865 ;
      RECT 1.25 134.535 2.26 134.585 ;
      RECT 0.245 133.97 0.755 135.43 ;
      RECT 14.11 133.97 74.81 135.43 ;
      RECT 0.245 127.995 74.81 133.97 ;
      RECT 0.285 135.43 74.81 137.05 ;
      RECT 12.3 134.815 13.31 134.865 ;
      RECT 12.295 134.245 13.31 134.815 ;
      RECT 2.105 144.655 72.665 145.505 ;
      RECT 2.105 163.695 72.665 164.545 ;
      RECT 71.26 145.505 72.665 163.695 ;
      RECT 2.105 145.505 3.51 163.695 ;
      RECT 3.95 146.19 4.55 162.235 ;
      RECT 5.74 146.19 6.34 162.235 ;
      RECT 6.85 147.085 8.04 160.075 ;
      RECT 5.06 147.22 5.23 160.075 ;
      RECT 10.7 146.19 11.3 162.235 ;
      RECT 8.55 146.19 9.15 162.235 ;
      RECT 9.475 147.32 10.375 160.075 ;
      RECT 11.81 147.085 13 160.075 ;
      RECT 13.51 146.19 14.11 162.235 ;
      RECT 15.66 146.19 16.26 162.235 ;
      RECT 14.435 147.32 15.335 160.075 ;
      RECT 14.62 147.22 15.15 147.32 ;
      RECT 18.47 146.19 19.07 162.235 ;
      RECT 16.77 147.085 17.96 160.075 ;
      RECT 19.395 147.32 20.295 160.075 ;
      RECT 19.58 147.22 20.11 147.32 ;
      RECT 23.43 146.19 24.03 162.235 ;
      RECT 20.62 146.19 21.22 162.235 ;
      RECT 21.73 147.085 22.92 160.075 ;
      RECT 24.355 147.32 25.255 160.075 ;
      RECT 24.54 147.22 25.07 147.32 ;
      RECT 28.39 146.19 28.99 162.235 ;
      RECT 25.58 146.19 26.18 162.235 ;
      RECT 26.69 147.085 27.88 160.075 ;
      RECT 30.54 146.19 31.14 162.235 ;
      RECT 31.65 147.085 32.84 160.075 ;
      RECT 29.315 147.32 30.215 160.075 ;
      RECT 29.5 147.22 30.03 147.32 ;
      RECT 33.35 146.19 33.95 162.235 ;
      RECT 35.5 146.19 36.1 162.235 ;
      RECT 36.61 147.085 37.8 160.075 ;
      RECT 34.275 147.32 35.175 160.075 ;
    LAYER met5 ;
      RECT 0 165.235 10.15 172.185 ;
      RECT 0 94.585 3.2 101.565 ;
      RECT 64.815 94.585 75 101.565 ;
      RECT 71.8 165.235 75 172.185 ;
      RECT 71.8 101.565 75 165.235 ;
      RECT 0 101.565 3.2 165.235 ;
      RECT 71.8 165.235 75 166.03 ;
      RECT 71.005 166.03 75 166.83 ;
      RECT 70.205 166.83 75 167.63 ;
      RECT 69.405 167.63 75 168.43 ;
      RECT 68.6 168.43 75 169.23 ;
      RECT 67.8 169.23 75 170.03 ;
      RECT 67.005 170.03 75 170.83 ;
      RECT 66.205 170.83 75 171.63 ;
      RECT 65.405 171.63 75 172.185 ;
      RECT 65.615 94.585 75 95.385 ;
      RECT 66.42 95.385 75 96.185 ;
      RECT 67.22 96.185 75 96.985 ;
      RECT 68.02 96.985 75 97.785 ;
      RECT 68.82 97.785 75 98.585 ;
      RECT 69.615 98.585 75 99.385 ;
      RECT 70.42 99.385 75 100.185 ;
      RECT 71.22 100.185 75 100.985 ;
      RECT 71.8 100.985 75 101.565 ;
      RECT 0 165.235 3.2 166.03 ;
      RECT 0 166.03 3.995 166.83 ;
      RECT 0 166.83 4.795 167.63 ;
      RECT 0 167.63 5.595 168.43 ;
      RECT 0 168.43 6.395 169.23 ;
      RECT 0 169.23 7.195 170.03 ;
      RECT 0 170.03 7.995 170.83 ;
      RECT 0 170.83 8.795 171.63 ;
      RECT 0 171.63 9.595 172.185 ;
      RECT 0 94.585 9.38 95.385 ;
      RECT 0 95.385 8.58 96.185 ;
      RECT 0 96.185 7.78 96.985 ;
      RECT 0 96.985 6.98 97.785 ;
      RECT 0 97.785 6.18 98.585 ;
      RECT 0 98.585 5.38 99.385 ;
      RECT 0 99.385 4.58 100.185 ;
      RECT 0 100.185 3.78 100.985 ;
      RECT 0 100.985 3.2 101.565 ;
    LAYER met4 ;
      RECT 0 55.035 75 55.835 ;
      RECT 0 44.635 75 45.435 ;
      RECT 0 5.885 75 6.485 ;
      RECT 0 16.785 75 17.385 ;
      RECT 0 11.935 75 12.535 ;
      RECT 0 55.135 75 55.835 ;
      RECT 0 44.635 75 45.335 ;
      RECT 0 22.835 75 23.435 ;
      RECT 0 66.935 75 67.635 ;
      RECT 0 61.085 75 61.685 ;
      RECT 0 38.585 75 39.185 ;
      RECT 0 33.735 75 34.335 ;
      RECT 0 28.885 75 29.485 ;
      RECT 0 93.4 75 173.385 ;
    LAYER met1 ;
      RECT 0 125.26 75 135.945 ;
      RECT 0 0 75 97.8 ;
      RECT -0.145 142.155 75.145 166.955 ;
      RECT -0.145 99.32 75.145 125.26 ;
      RECT -0.145 97.8 75 125.26 ;
      RECT -0.145 97.8 75 99.32 ;
      RECT 0 166.955 75 198 ;
      RECT 0 0 75 198 ;
      RECT 0 0 75 198 ;
      RECT 0 0 75 198 ;
      RECT 0 135.945 75.145 166.955 ;
      RECT 0 135.945 75.145 142.155 ;
    LAYER met2 ;
      RECT 0 0 75 198 ;
  END
END sky130_fd_io__top_analog_pad

END LIBRARY
