# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__top_ground_hvc_wpad
  CLASS PAD ;
  FOREIGN sky130_fd_io__top_ground_hvc_wpad ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  75.00000 BY  200.0000 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN G_PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 6.100000 104.010000 68.800000 166.625000 ;
    END
  END G_PAD
  PIN DRN_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 37.890000 0.000000 48.890000 96.150000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 100.105000 42.840000 100.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 100.215000 42.840000 102.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 102.135000 42.840000 102.285000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 102.285000 42.990000 102.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 102.435000 43.140000 102.585000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 102.585000 43.290000 102.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 102.735000 43.440000 102.885000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 102.885000 43.590000 103.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 103.035000 43.740000 103.185000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 103.185000 43.890000 103.335000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 103.335000 44.040000 103.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 103.485000 44.190000 103.635000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 103.635000 44.340000 103.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 103.785000 44.490000 103.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 103.935000 44.640000 104.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 104.085000 44.790000 104.235000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 104.235000 44.940000 104.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 104.535000 45.240000 104.685000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 104.685000 45.390000 104.835000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 104.835000 45.540000 104.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 104.985000 45.690000 105.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 105.135000 45.840000 105.285000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 105.285000 45.990000 105.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 105.435000 46.140000 105.585000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 105.585000 46.290000 105.655000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 105.655000 42.855000 110.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 96.150000 48.890000 96.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 96.300000 49.040000 96.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 96.450000 49.190000 96.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 96.600000 49.340000 96.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 96.750000 49.490000 96.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 96.900000 49.640000 97.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 97.050000 49.790000 97.200000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 97.200000 49.940000 97.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 97.350000 50.090000 97.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 97.500000 50.240000 97.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 97.650000 50.390000 97.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 97.800000 50.540000 97.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 97.950000 50.690000 98.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 98.100000 50.840000 98.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 98.300000 51.040000 99.505000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 99.505000 43.400000 99.655000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 99.655000 43.250000 99.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890000 99.805000 43.100000 99.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.965000 170.460000 42.855000 175.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.965000 175.350000 48.855000 190.020000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.040000 105.655000 46.360000 105.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.055000 175.260000 48.855000 175.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.190000 105.805000 46.510000 105.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.205000 175.110000 48.855000 175.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.355000 174.960000 48.855000 175.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.490000 106.105000 46.810000 106.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.505000 174.810000 48.855000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.640000 106.255000 46.960000 106.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.655000 174.660000 48.855000 174.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.790000 106.405000 47.110000 106.555000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.805000 174.510000 48.855000 174.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.940000 106.555000 47.260000 106.705000 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.955000 174.360000 48.855000 174.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.090000 106.705000 47.410000 106.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.105000 174.210000 48.855000 174.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.240000 106.855000 47.560000 107.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.255000 174.060000 48.855000 174.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.390000 107.005000 47.710000 107.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.405000 173.910000 48.855000 174.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.540000 107.155000 47.860000 107.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.555000 173.760000 48.855000 173.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.690000 107.305000 48.010000 107.455000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.705000 173.610000 48.855000 173.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.840000 107.455000 48.160000 107.605000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.855000 173.460000 48.855000 173.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.990000 107.605000 48.310000 107.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.005000 173.310000 48.855000 173.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.140000 107.755000 48.460000 107.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.155000 173.160000 48.855000 173.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.290000 107.905000 48.610000 108.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.305000 173.010000 48.855000 173.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.455000 172.860000 48.855000 173.010000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.535000 108.150000 48.855000 108.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.605000 172.710000 48.855000 172.860000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.685000 108.300000 48.855000 108.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.755000 172.560000 48.855000 172.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.835000 108.450000 48.855000 108.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.905000 172.410000 48.855000 172.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.985000 108.600000 48.855000 108.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.055000 172.260000 48.855000 172.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.135000 108.750000 48.855000 108.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.205000 172.110000 48.855000 172.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.285000 108.900000 48.855000 109.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.355000 171.960000 48.855000 172.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.435000 109.050000 48.855000 109.200000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.505000 171.810000 48.855000 171.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.585000 109.200000 48.855000 109.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.655000 171.660000 48.855000 171.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.735000 109.350000 48.855000 109.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.805000 171.510000 48.855000 171.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.885000 109.500000 48.855000 109.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.955000 171.360000 48.855000 171.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.035000 109.650000 48.855000 109.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.105000 171.210000 48.855000 171.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.185000 109.800000 48.855000 109.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.255000 171.060000 48.855000 171.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.335000 109.950000 48.855000 110.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.405000 170.910000 48.855000 171.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.485000 110.100000 48.855000 110.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.555000 170.760000 48.855000 170.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.635000 110.250000 48.855000 110.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.840000 102.135000 45.240000 104.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.840000 99.505000 43.550000 100.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.855000 108.150000 48.855000 110.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.855000 110.620000 48.855000 170.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.855000 170.460000 48.855000 170.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.550000 99.505000 45.260000 100.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.655000 99.505000 51.040000 99.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.760000 99.610000 51.040000 99.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.910000 99.715000 51.040000 99.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.060000 99.865000 51.190000 100.015000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.240000 104.535000 46.715000 106.010000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260000 100.165000 51.490000 100.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260000 100.215000 51.540000 100.365000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260000 100.365000 51.690000 100.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260000 100.515000 51.840000 100.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260000 100.665000 51.990000 100.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260000 100.815000 52.140000 100.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260000 100.965000 52.290000 101.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260000 101.115000 52.440000 101.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260000 101.265000 52.590000 101.415000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260000 101.415000 52.740000 101.565000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260000 101.565000 52.890000 101.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260000 101.715000 53.040000 101.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260000 101.865000 53.190000 102.015000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260000 102.015000 53.340000 102.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260000 102.165000 53.490000 102.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260000 102.315000 53.640000 102.415000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260000 102.415000 47.380000 104.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.410000 102.415000 53.740000 102.565000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.560000 102.565000 53.890000 102.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.710000 102.715000 54.040000 102.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.860000 102.865000 54.190000 103.015000 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.010000 103.015000 54.340000 103.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.160000 103.165000 54.490000 103.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.310000 103.315000 54.640000 103.465000 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.460000 103.465000 54.790000 103.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.610000 103.615000 54.940000 103.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.715000 106.010000 48.855000 108.150000 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.760000 103.765000 55.090000 103.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.910000 103.915000 55.240000 104.065000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.060000 104.065000 55.390000 104.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.210000 104.215000 55.540000 104.365000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.380000 104.535000 48.855000 106.010000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.510000 104.515000 55.840000 104.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.660000 104.665000 55.990000 104.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.810000 104.815000 56.140000 104.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.960000 104.965000 56.290000 105.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.110000 105.115000 56.440000 105.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.260000 105.265000 56.590000 105.415000 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.410000 105.415000 56.740000 105.565000 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.560000 105.565000 56.890000 105.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.855000 106.010000 50.995000 108.150000 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.860000 105.865000 57.190000 106.015000 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.890000 96.150000 51.040000 98.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.010000 106.015000 57.340000 106.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.160000 106.165000 57.490000 106.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.310000 106.315000 57.640000 106.465000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.460000 106.465000 57.790000 106.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.610000 106.615000 57.940000 106.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.760000 106.765000 58.090000 106.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775000 169.135000 53.285000 172.645000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775000 172.645000 59.285000 173.020000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775000 172.645000 59.285000 173.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775000 173.170000 59.435000 173.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775000 173.320000 59.585000 173.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775000 173.470000 59.735000 173.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775000 173.620000 59.885000 173.770000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775000 173.770000 60.035000 173.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775000 173.920000 60.185000 174.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775000 174.070000 60.335000 174.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775000 174.220000 60.485000 174.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775000 174.370000 60.635000 174.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775000 174.520000 60.785000 174.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775000 174.680000 60.945000 190.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.835000 172.585000 59.285000 172.645000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.910000 106.915000 58.240000 107.065000 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.985000 172.435000 59.285000 172.585000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.060000 107.065000 58.390000 107.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.135000 172.285000 59.285000 172.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.210000 107.215000 58.540000 107.365000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.285000 172.135000 59.285000 172.285000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.360000 107.365000 58.690000 107.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.435000 171.985000 59.285000 172.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.510000 107.515000 58.840000 107.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.585000 171.835000 59.285000 171.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.660000 107.665000 58.990000 107.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.735000 171.685000 59.285000 171.835000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.885000 171.535000 59.285000 171.685000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.995000 108.150000 53.285000 110.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.035000 171.385000 59.285000 171.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.040000 99.715000 59.285000 107.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.105000 108.110000 59.285000 108.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.185000 171.235000 59.285000 171.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255000 108.260000 59.285000 108.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.335000 171.085000 59.285000 171.235000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.405000 108.410000 59.285000 108.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.485000 170.935000 59.285000 171.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.555000 108.560000 59.285000 108.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.635000 170.785000 59.285000 170.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.705000 108.710000 59.285000 108.860000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.785000 170.635000 59.285000 170.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.855000 108.860000 59.285000 109.010000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.935000 170.485000 59.285000 170.635000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.005000 109.010000 59.285000 109.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.085000 170.335000 59.285000 170.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.155000 109.160000 59.285000 109.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.235000 170.185000 59.285000 170.335000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.305000 109.310000 59.285000 109.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.385000 170.035000 59.285000 170.185000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.455000 109.460000 59.285000 109.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.535000 169.885000 59.285000 170.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.605000 109.610000 59.285000 109.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.685000 169.735000 59.285000 169.885000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.755000 109.760000 59.285000 109.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 169.585000 59.285000 169.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.905000 109.910000 59.285000 110.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.985000 169.435000 59.285000 169.585000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.055000 110.060000 59.285000 110.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 107.960000 59.285000 110.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 110.440000 59.285000 169.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 169.135000 59.285000 169.285000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.285000 173.020000 60.945000 174.680000 ;
    END
  END DRN_HVC
  PIN G_CORE
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 50.390000 0.000000 74.290000 90.185000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000 90.185000 56.355000 96.150000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.540000 90.185000 74.290000 90.335000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.690000 90.335000 74.290000 90.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.840000 90.485000 74.290000 90.635000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.990000 90.635000 74.290000 90.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.140000 90.785000 74.290000 90.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.290000 90.935000 74.290000 91.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.440000 91.085000 74.290000 91.235000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.590000 91.235000 74.290000 91.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.740000 91.385000 74.290000 91.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.890000 91.535000 74.290000 91.685000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.040000 91.685000 74.290000 91.835000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.190000 91.835000 74.290000 91.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.340000 91.985000 74.290000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.490000 92.135000 74.290000 92.285000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.640000 92.285000 74.290000 92.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.790000 92.435000 74.290000 92.585000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940000 92.585000 74.290000 92.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.090000 92.735000 74.290000 92.885000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.240000 92.885000 74.290000 93.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.390000 93.035000 74.290000 93.185000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.540000 93.185000 74.290000 93.335000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 93.335000 74.290000 93.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.840000 93.485000 74.290000 93.635000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.990000 93.635000 74.290000 93.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.140000 93.785000 74.290000 93.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.290000 93.935000 74.290000 94.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.440000 94.085000 74.290000 94.235000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.590000 94.235000 74.290000 94.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.740000 94.385000 74.290000 94.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.890000 94.535000 74.290000 94.685000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.040000 94.685000 74.290000 94.835000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.190000 94.835000 74.290000 94.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.340000 94.985000 74.290000 95.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.490000 95.135000 74.290000 95.285000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.640000 95.285000 74.290000 95.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.790000 95.435000 74.290000 95.585000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.940000 95.585000 74.290000 95.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.090000 95.735000 74.290000 95.885000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.355000 96.150000 59.920000 99.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.390000 96.035000 74.290000 96.185000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.540000 96.185000 74.290000 96.335000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.690000 96.335000 74.290000 96.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840000 96.485000 74.290000 96.635000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990000 96.635000 74.290000 96.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.140000 96.785000 74.290000 96.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.290000 96.935000 74.290000 97.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.440000 97.085000 74.290000 97.235000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.590000 97.235000 74.290000 97.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 97.385000 74.290000 97.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.890000 97.535000 74.290000 97.685000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.040000 97.685000 74.290000 97.835000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.190000 97.835000 74.290000 97.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.340000 97.985000 74.290000 98.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.490000 98.135000 74.290000 98.285000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.640000 98.285000 74.290000 98.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.790000 98.435000 74.290000 98.585000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.940000 98.585000 74.290000 98.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.090000 98.735000 74.290000 98.885000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.240000 98.885000 74.290000 99.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.390000 99.035000 74.290000 99.185000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.540000 99.185000 74.290000 99.335000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.690000 99.335000 74.290000 99.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.920000 99.715000 61.500000 101.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.990000 99.635000 74.290000 99.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.140000 99.785000 74.290000 99.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.290000 99.935000 74.290000 100.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.440000 100.085000 74.290000 100.235000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.590000 100.235000 74.290000 100.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.740000 100.385000 74.290000 100.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.890000 100.535000 74.290000 100.685000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040000 100.685000 74.290000 100.835000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.190000 100.835000 74.290000 100.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.340000 100.985000 74.290000 101.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.500000 101.285000 74.290000 101.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.500000 101.295000 74.290000 173.320000 ;
    END
  END G_CORE
  PIN OGC_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 25.895000 0.000000 27.895000 0.535000 ;
    END
  END OGC_HVC
  PIN SRC_BDY_HVC
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 14.050000 171.305000 15.500000 172.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.050000 172.755000 25.010000 195.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.055000 172.750000 25.010000 172.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.110000 172.695000 25.010000 172.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.165000 172.640000 25.010000 172.695000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.300000 172.505000 24.875000 172.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.450000 172.355000 24.725000 172.505000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.600000 172.205000 24.575000 172.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.750000 172.055000 24.425000 172.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.900000 171.905000 24.275000 172.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.050000 171.755000 24.125000 171.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.200000 171.605000 23.975000 171.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 102.200000 23.830000 102.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 102.350000 23.680000 102.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 102.500000 23.530000 102.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 102.650000 23.380000 102.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 102.800000 23.230000 102.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 102.950000 23.080000 103.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 103.100000 22.930000 103.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 103.250000 22.780000 103.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 103.400000 22.630000 103.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 103.550000 22.480000 103.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 103.700000 22.330000 103.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 103.850000 22.180000 104.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 104.000000 22.030000 104.150000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 104.150000 21.880000 104.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 104.300000 21.730000 104.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 104.450000 21.580000 104.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 104.600000 21.500000 104.680000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 104.680000 21.500000 169.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 158.470000 21.500000 169.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 169.280000 21.650000 169.430000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 169.430000 21.800000 169.580000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 169.580000 21.950000 169.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 169.730000 22.100000 169.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 169.880000 22.250000 170.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 170.030000 22.400000 170.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 170.180000 22.550000 170.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 170.330000 22.700000 170.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 170.480000 22.850000 170.630000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 170.630000 23.000000 170.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 170.780000 23.150000 170.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 170.930000 23.300000 171.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 171.080000 23.450000 171.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 171.230000 23.600000 171.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500000 99.395000 18.305000 102.200000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645000 102.055000 23.980000 102.200000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.795000 101.905000 24.125000 102.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 101.755000 24.275000 101.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.095000 101.605000 24.425000 101.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.245000 101.455000 24.575000 101.605000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.395000 101.305000 24.725000 101.455000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.545000 101.155000 24.875000 101.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.695000 101.005000 25.025000 101.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.845000 100.855000 25.175000 101.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.995000 100.705000 25.325000 100.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.145000 100.555000 25.475000 100.705000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.295000 100.405000 25.625000 100.555000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.445000 100.255000 25.775000 100.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.745000 99.955000 26.075000 100.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.895000 99.805000 26.225000 99.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 99.655000 26.375000 99.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.305000 96.665000 21.035000 99.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.345000 99.355000 26.675000 99.505000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.495000 99.205000 26.825000 99.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.645000 99.055000 26.975000 99.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.795000 98.905000 27.125000 99.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.945000 98.755000 27.275000 98.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.095000 98.605000 27.425000 98.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.245000 98.455000 27.575000 98.605000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.395000 98.305000 27.725000 98.455000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.545000 98.155000 27.875000 98.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.845000 97.855000 28.175000 98.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 97.705000 28.325000 97.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.145000 97.555000 28.475000 97.705000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.295000 97.405000 28.625000 97.555000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.445000 97.255000 28.775000 97.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.595000 97.105000 28.925000 97.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.745000 96.955000 29.075000 97.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.035000 93.955000 23.745000 96.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.195000 96.505000 29.525000 96.655000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.345000 96.355000 29.525000 96.505000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.495000 96.205000 29.525000 96.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.500000 100.250000 25.930000 104.680000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.500000 169.130000 25.010000 172.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645000 96.055000 29.525000 96.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.795000 95.905000 29.525000 96.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.945000 95.755000 29.525000 95.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.095000 95.605000 29.525000 95.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.245000 95.455000 29.525000 95.605000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.395000 95.305000 29.525000 95.455000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.545000 95.155000 29.525000 95.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.695000 95.005000 29.525000 95.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845000 94.855000 29.525000 95.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.995000 94.705000 29.525000 94.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.145000 94.555000 29.525000 94.705000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.295000 94.405000 29.525000 94.555000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.445000 94.255000 29.525000 94.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 91.150000 25.135000 92.540000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 92.540000 29.525000 96.655000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 92.540000 29.935000 92.690000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 92.690000 29.785000 92.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 92.840000 29.635000 92.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 92.990000 29.525000 93.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 93.100000 29.525000 93.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.820000 92.465000 30.085000 92.540000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.945000 92.340000 36.895000 92.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.095000 92.190000 36.895000 92.340000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.245000 92.040000 36.895000 92.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.395000 91.890000 36.895000 92.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.545000 91.740000 36.895000 91.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.695000 91.590000 36.895000 91.740000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.845000 91.440000 36.895000 91.590000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.135000 90.390000 25.895000 91.150000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.145000 91.140000 36.895000 91.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.295000 90.990000 36.895000 91.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.445000 90.840000 36.895000 90.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.595000 90.690000 36.895000 90.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.895000 0.000000 36.895000 90.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.895000 90.390000 36.895000 90.540000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 100.250000 28.070000 102.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 102.390000 34.250000 102.540000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 102.540000 34.100000 102.690000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 102.690000 33.950000 102.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 102.840000 33.800000 102.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 102.990000 33.650000 103.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 103.140000 33.500000 103.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 103.290000 33.350000 103.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 103.440000 33.200000 103.590000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 103.590000 33.050000 103.740000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 103.740000 32.900000 103.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 103.890000 32.750000 104.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 104.040000 32.600000 104.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 104.190000 32.450000 104.340000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 104.340000 32.300000 104.490000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 104.490000 32.150000 104.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 104.640000 32.000000 104.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 104.790000 31.930000 104.860000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 104.860000 31.930000 170.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 158.470000 31.930000 170.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 170.610000 32.080000 170.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 170.760000 32.230000 170.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 170.910000 32.380000 171.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 171.060000 32.530000 171.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 171.210000 32.680000 171.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 171.360000 32.830000 171.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 171.510000 32.980000 171.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 171.660000 33.130000 171.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 171.810000 33.280000 171.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 171.960000 33.430000 172.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 172.110000 33.580000 172.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 172.260000 33.730000 172.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 172.410000 33.880000 172.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 172.560000 34.030000 172.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 172.860000 34.330000 173.010000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 173.010000 34.480000 173.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 173.160000 34.630000 173.310000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 173.460000 34.930000 173.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 173.610000 35.080000 173.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 173.760000 35.230000 173.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 173.910000 35.380000 174.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 174.210000 35.680000 174.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 174.360000 35.830000 174.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 174.510000 35.980000 174.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 174.810000 36.280000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 174.960000 36.430000 175.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 175.110000 36.580000 175.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 175.350000 36.820000 195.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930000 98.145000 28.035000 100.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.025000 102.295000 34.400000 102.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.175000 102.145000 34.495000 102.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.325000 101.995000 34.645000 102.145000 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.475000 101.845000 34.795000 101.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.625000 101.695000 34.945000 101.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.775000 101.545000 35.095000 101.695000 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.925000 101.395000 35.245000 101.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.075000 101.245000 35.395000 101.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.225000 101.095000 35.545000 101.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.375000 100.945000 35.695000 101.095000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.525000 100.795000 35.845000 100.945000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.675000 100.645000 35.995000 100.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.825000 100.495000 36.145000 100.645000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.035000 96.655000 29.525000 98.145000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.070000 98.145000 30.175000 100.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.125000 100.195000 36.445000 100.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.275000 100.045000 36.595000 100.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.495000 99.825000 36.895000 99.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.645000 99.675000 36.895000 99.825000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.795000 99.525000 36.895000 99.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.945000 99.375000 36.895000 99.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.095000 99.225000 36.895000 99.375000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.245000 99.075000 36.895000 99.225000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.395000 98.925000 36.895000 99.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.525000 92.390000 30.235000 93.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.545000 98.775000 36.895000 98.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.695000 98.625000 36.895000 98.775000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.845000 98.475000 36.895000 98.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.995000 98.325000 36.895000 98.475000 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.175000 96.375000 31.945000 98.145000 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.295000 98.025000 36.895000 98.175000 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.445000 97.875000 36.895000 98.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.595000 97.725000 36.895000 97.875000 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.745000 97.575000 36.895000 97.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.895000 97.425000 36.895000 97.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.045000 97.275000 36.895000 97.425000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.195000 97.125000 36.895000 97.275000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.235000 92.390000 31.945000 93.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.345000 96.975000 36.895000 97.125000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.385000 92.390000 36.895000 92.540000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.495000 96.825000 36.895000 96.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.535000 92.540000 36.895000 92.690000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.645000 96.675000 36.895000 96.825000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.685000 92.690000 36.895000 92.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.930000 170.460000 34.225000 172.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.930000 99.895000 36.895000 104.860000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.945000 89.470000 36.895000 99.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.945000 92.990000 36.895000 93.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.945000 93.100000 36.895000 96.375000 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.225000 172.755000 34.790000 173.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.790000 173.320000 35.540000 174.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.540000 174.070000 36.230000 174.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.230000 174.760000 36.820000 175.350000 ;
    END
  END SRC_BDY_HVC
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT 1.070000 1.000000 72.775000 199.695000 ;
    LAYER met1 ;
      RECT 0.185000 0.970000 73.620000 199.725000 ;
    LAYER met2 ;
      RECT  0.265000 0.000000 25.615000   0.815000 ;
      RECT  0.265000 0.815000 74.290000 195.075000 ;
      RECT 28.175000 0.000000 74.290000   0.815000 ;
    LAYER met3 ;
      RECT  0.240000   0.000000 25.495000  89.990000 ;
      RECT  0.240000  89.990000 24.735000  90.750000 ;
      RECT  0.240000  90.750000 23.345000  93.555000 ;
      RECT  0.240000  93.555000 20.635000  96.265000 ;
      RECT  0.240000  96.265000 17.905000  98.995000 ;
      RECT  0.240000  98.995000 15.100000 170.905000 ;
      RECT  0.240000 170.905000 13.650000 175.350000 ;
      RECT 21.900000 105.080000 25.530000 168.730000 ;
      RECT 25.410000 168.730000 25.530000 175.350000 ;
      RECT 29.925000  93.500000 31.545000  95.975000 ;
      RECT 30.635000  92.790000 30.835000  93.500000 ;
      RECT 32.330000 105.260000 37.490000 111.020000 ;
      RECT 32.330000 111.020000 42.455000 170.060000 ;
      RECT 34.625000 170.060000 37.565000 172.355000 ;
      RECT 35.190000 172.355000 37.565000 172.920000 ;
      RECT 35.940000 172.920000 37.565000 173.670000 ;
      RECT 36.630000 173.670000 37.565000 174.360000 ;
      RECT 37.220000 174.360000 37.565000 175.350000 ;
      RECT 37.295000   0.000000 37.490000 105.260000 ;
      RECT 43.240000 100.615000 44.860000 101.735000 ;
      RECT 43.950000  99.905000 44.150000 100.615000 ;
      RECT 49.255000 108.550000 50.595000 110.840000 ;
      RECT 49.255000 110.840000 52.885000 168.735000 ;
      RECT 49.255000 168.735000 49.375000 175.350000 ;
      RECT 49.290000   0.000000 49.990000  95.750000 ;
      RECT 51.440000  96.550000 55.955000  99.315000 ;
      RECT 59.685000 101.695000 61.100000 172.620000 ;
      RECT 61.345000 173.720000 74.290000 175.350000 ;
    LAYER met4 ;
      RECT 0.000000  2.035000 75.000000  47.965000 ;
      RECT 0.000000 51.745000 75.000000  52.725000 ;
      RECT 0.000000 56.505000 75.000000 200.000000 ;
    LAYER met5 ;
      RECT  0.000000   2.135000 72.130000  15.035000 ;
      RECT  0.000000  15.035000 72.435000  19.885000 ;
      RECT  0.000000  19.885000 75.000000  24.335000 ;
      RECT  0.000000  24.335000 72.130000  36.835000 ;
      RECT  0.000000  36.835000 75.000000  40.085000 ;
      RECT  0.000000  40.085000 72.130000  96.585000 ;
      RECT  0.000000  96.585000 75.000000 102.410000 ;
      RECT  0.000000 102.410000  4.500000 168.225000 ;
      RECT  0.000000 168.225000 75.000000 200.000000 ;
      RECT 70.400000 102.410000 75.000000 168.225000 ;
  END
END sky130_fd_io__top_ground_hvc_wpad
END LIBRARY
