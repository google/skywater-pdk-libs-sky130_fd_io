# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__top_ground_lvc_wpad
  CLASS PAD ;
  FOREIGN sky130_fd_io__top_ground_lvc_wpad ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  75.00000 BY  198.0000 ;
  SYMMETRY R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN G_PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 9.315000 100.140000 65.955000 167.570000 ;
    END
  END G_PAD
  PIN BDY2_B2B
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 34.440000 0.000000 44.440000 0.325000 ;
    END
  END BDY2_B2B
  PIN DRN_LVC1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 26.000000 0.000000 36.880000 20.220000 ;
    END
  END DRN_LVC1
  PIN DRN_LVC2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.380000 0.000000 49.255000 22.900000 ;
    END
  END DRN_LVC2
  PIN G_CORE
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 50.755000 0.000000 74.700000 84.465000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000 84.465000 51.100000 84.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.905000 84.465000 74.700000 84.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.100000 84.810000 54.665000 88.375000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.205000 84.765000 74.700000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.355000 84.915000 74.700000 85.065000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.505000 85.065000 74.700000 85.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655000 85.215000 74.700000 85.365000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.805000 85.365000 74.700000 85.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.955000 85.515000 74.700000 85.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.105000 85.665000 74.700000 85.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.255000 85.815000 74.700000 85.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 85.965000 74.700000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.555000 86.115000 74.700000 86.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.705000 86.265000 74.700000 86.415000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.855000 86.415000 74.700000 86.565000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.005000 86.565000 74.700000 86.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.155000 86.715000 74.700000 86.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305000 86.865000 74.700000 87.015000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.455000 87.015000 74.700000 87.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.605000 87.165000 74.700000 87.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.755000 87.315000 74.700000 87.465000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.905000 87.465000 74.700000 87.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 87.615000 74.700000 87.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.205000 87.765000 74.700000 87.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.355000 87.915000 74.700000 88.065000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.505000 88.065000 74.700000 88.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.665000 88.375000 58.310000 92.020000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.805000 88.365000 74.700000 88.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.955000 88.515000 74.700000 88.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.105000 88.665000 74.700000 88.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.255000 88.815000 74.700000 88.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.405000 88.965000 74.700000 89.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.555000 89.115000 74.700000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 89.265000 74.700000 89.415000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.855000 89.415000 74.700000 89.565000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.005000 89.565000 74.700000 89.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.155000 89.715000 74.700000 89.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.305000 89.865000 74.700000 90.015000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 90.015000 74.700000 90.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.605000 90.165000 74.700000 90.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.755000 90.315000 74.700000 90.465000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.905000 90.465000 74.700000 90.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.055000 90.615000 74.700000 90.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.205000 90.765000 74.700000 90.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355000 90.915000 74.700000 91.065000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.505000 91.065000 74.700000 91.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.655000 91.215000 74.700000 91.365000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.805000 91.365000 74.700000 91.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.955000 91.515000 74.700000 91.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 91.665000 74.700000 91.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.400000 92.110000 62.045000 95.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.405000 91.965000 74.700000 92.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.555000 92.115000 74.700000 92.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.705000 92.265000 74.700000 92.415000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.855000 92.415000 74.700000 92.565000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.005000 92.565000 74.700000 92.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.155000 92.715000 74.700000 92.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.305000 92.865000 74.700000 93.015000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.455000 93.015000 74.700000 93.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.605000 93.165000 74.700000 93.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755000 93.315000 74.700000 93.465000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.905000 93.465000 74.700000 93.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.055000 93.615000 74.700000 93.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.205000 93.765000 74.700000 93.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.355000 93.915000 74.700000 94.065000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 94.065000 74.700000 94.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.655000 94.215000 74.700000 94.365000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.805000 94.365000 74.700000 94.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.955000 94.515000 74.700000 94.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.105000 94.665000 74.700000 94.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.255000 94.815000 74.700000 94.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405000 94.965000 74.700000 95.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.555000 95.115000 74.700000 95.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.705000 95.265000 74.700000 95.415000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.855000 95.415000 74.700000 95.565000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.045000 0.000000 74.700000 95.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.045000 95.755000 74.700000 172.235000 ;
    END
  END G_CORE
  PIN OGC_LVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 26.210000 0.000000 27.700000 0.170000 ;
    END
  END OGC_LVC
  PIN SRC_BDY_LVC1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.500000 0.000000 20.495000 1.485000 ;
    END
  END SRC_BDY_LVC1
  PIN SRC_BDY_LVC2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 54.715000 0.000000 74.700000 3.660000 ;
    END
  END SRC_BDY_LVC2
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT 0.240000 1.020000 74.755000 197.780000 ;
    LAYER met1 ;
      RECT  0.120000 0.000000 25.930000   0.450000 ;
      RECT  0.120000 0.450000 74.785000 197.840000 ;
      RECT 27.980000 0.000000 74.785000   0.450000 ;
    LAYER met2 ;
      RECT  0.500000 1.765000 54.435000   3.940000 ;
      RECT  0.500000 3.940000 74.700000 194.430000 ;
      RECT 20.775000 0.000000 34.160000   0.605000 ;
      RECT 20.775000 0.605000 54.435000   1.765000 ;
      RECT 44.720000 0.000000 54.435000   0.605000 ;
    LAYER met3 ;
      RECT  0.500000   0.000000 25.600000  20.620000 ;
      RECT  0.500000  20.620000 37.980000  23.300000 ;
      RECT  0.500000  23.300000 50.355000  85.210000 ;
      RECT  0.500000  85.210000 50.700000  88.775000 ;
      RECT  0.500000  88.775000 54.265000  92.420000 ;
      RECT  0.500000  92.420000 58.000000  96.155000 ;
      RECT  0.500000  96.155000 61.645000 172.635000 ;
      RECT  0.500000 172.635000 62.045000 189.515000 ;
      RECT 37.280000   0.000000 37.980000  20.620000 ;
      RECT 49.655000   0.000000 50.355000  23.300000 ;
    LAYER met4 ;
      RECT 0.000000  0.035000 75.000000  45.965000 ;
      RECT 0.000000 49.745000 75.000000  50.725000 ;
      RECT 0.000000 54.505000 75.000000 198.000000 ;
    LAYER met5 ;
      RECT  0.000000   0.135000 72.130000  13.035000 ;
      RECT  0.000000  13.035000 72.435000  17.885000 ;
      RECT  0.000000  17.885000 75.000000  22.335000 ;
      RECT  0.000000  22.335000 72.130000  34.835000 ;
      RECT  0.000000  34.835000 75.000000  38.085000 ;
      RECT  0.000000  38.085000 72.130000  94.585000 ;
      RECT  0.000000  94.585000 75.000000  98.540000 ;
      RECT  0.000000  98.540000  7.715000 169.170000 ;
      RECT  0.000000 169.170000 75.000000 198.000000 ;
      RECT 67.555000  98.540000 75.000000 169.170000 ;
  END
END sky130_fd_io__top_ground_lvc_wpad
END LIBRARY
