# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_io__top_xres4v2
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 200 ;
  SYMMETRY R90 ;
  PIN AMUXBUS_A
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    ANTENNAPARTIALMETALSIDEAREA  111.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN DISABLE_PULLUP_H
    ANTENNAPARTIALCUTAREA  0.045000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 28.635000 28.540000 33.025000 28.580000 ;
        RECT 28.635000 28.580000 28.950000 28.650000 ;
        RECT 28.635000 28.650000 28.880000 28.720000 ;
        RECT 28.635000 28.720000 28.865000 28.735000 ;
        RECT 28.635000 28.735000 28.865000 32.435000 ;
        RECT 28.685000 28.490000 33.025000 28.540000 ;
        RECT 28.755000 28.420000 33.025000 28.490000 ;
        RECT 28.825000 28.350000 33.025000 28.420000 ;
        RECT 32.555000 28.340000 33.025000 28.350000 ;
        RECT 32.625000 28.270000 33.025000 28.340000 ;
        RECT 32.695000 28.200000 33.025000 28.270000 ;
        RECT 32.760000  0.000000 33.020000  8.720000 ;
        RECT 32.760000  8.720000 33.020000  8.725000 ;
        RECT 32.760000  8.725000 33.025000  8.830000 ;
        RECT 32.765000  8.830000 33.025000  8.835000 ;
        RECT 32.765000  8.835000 33.025000 28.130000 ;
        RECT 32.765000 28.130000 33.025000 28.200000 ;
    END
    PORT
      LAYER met2 ;
        RECT 32.760000 0.000000 33.020000 0.640000 ;
    END
  END DISABLE_PULLUP_H
  PIN ENABLE_H
    ANTENNAPARTIALCUTAREA  0.180000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 12.145000  6.635000 12.545000  6.665000 ;
        RECT 12.215000  6.565000 12.545000  6.635000 ;
        RECT 12.285000  0.000000 12.545000  6.495000 ;
        RECT 12.285000  6.495000 12.545000  6.565000 ;
        RECT 12.370000  6.665000 12.545000  6.775000 ;
        RECT 12.370000  6.775000 12.545000  6.845000 ;
        RECT 12.370000  6.845000 12.615000  6.915000 ;
        RECT 12.370000  6.915000 12.685000  6.925000 ;
        RECT 12.440000  6.925000 12.695000  6.995000 ;
        RECT 12.510000  6.995000 12.765000  7.065000 ;
        RECT 12.575000  7.065000 12.835000  7.130000 ;
        RECT 12.635000  7.130000 12.900000  7.190000 ;
        RECT 12.695000  7.190000 12.900000  7.250000 ;
        RECT 12.695000  7.250000 12.900000 10.230000 ;
        RECT 12.800000 10.230000 12.865000 10.265000 ;
        RECT 12.800000 10.265000 12.830000 10.300000 ;
        RECT 12.800000 10.300000 12.825000 10.305000 ;
    END
    PORT
      LAYER met2 ;
        RECT 12.285000 0.000000 12.545000 1.470000 ;
    END
  END ENABLE_H
  PIN ENABLE_VDDIO
    ANTENNAPARTIALCUTAREA  0.200000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.425000 0.000000 8.895000 1.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.775000 17.410000  7.400000 17.515000 ;
        RECT 6.775000 17.515000  7.295000 17.620000 ;
        RECT 6.775000 17.620000  7.295000 31.295000 ;
        RECT 6.775000 31.295000  7.295000 31.400000 ;
        RECT 6.775000 31.400000  7.400000 31.505000 ;
        RECT 6.840000 17.345000  7.505000 17.410000 ;
        RECT 6.925000 31.505000  7.505000 31.655000 ;
        RECT 6.990000 17.195000  7.570000 17.345000 ;
        RECT 7.075000 31.655000  7.655000 31.805000 ;
        RECT 7.140000 17.045000  7.720000 17.195000 ;
        RECT 7.225000 31.805000  7.805000 31.955000 ;
        RECT 7.290000 16.895000  7.870000 17.045000 ;
        RECT 7.375000 31.955000  7.955000 32.105000 ;
        RECT 7.440000 16.745000  8.020000 16.895000 ;
        RECT 7.525000 32.105000  8.105000 32.255000 ;
        RECT 7.590000 16.595000  8.170000 16.745000 ;
        RECT 7.675000 32.255000  8.255000 32.405000 ;
        RECT 7.740000 16.445000  8.320000 16.595000 ;
        RECT 7.825000 32.405000  8.405000 32.555000 ;
        RECT 7.890000 16.295000  8.470000 16.445000 ;
        RECT 7.975000 32.555000  8.555000 32.705000 ;
        RECT 8.040000 16.145000  8.620000 16.295000 ;
        RECT 8.125000 32.705000  8.705000 32.855000 ;
        RECT 8.190000 15.995000  8.770000 16.145000 ;
        RECT 8.275000 32.855000  8.855000 33.005000 ;
        RECT 8.295000 15.890000  8.920000 15.995000 ;
        RECT 8.400000  0.000000  8.920000 15.785000 ;
        RECT 8.400000 15.785000  8.920000 15.890000 ;
        RECT 8.425000 33.005000  9.005000 33.155000 ;
        RECT 8.575000 33.155000  9.155000 33.305000 ;
        RECT 8.665000 33.305000  9.305000 33.395000 ;
        RECT 8.815000 33.395000 22.275000 33.545000 ;
        RECT 8.965000 33.545000 22.275000 33.695000 ;
        RECT 9.115000 33.695000 22.275000 33.845000 ;
        RECT 9.265000 33.845000 22.275000 33.995000 ;
        RECT 9.395000 33.995000 22.275000 34.125000 ;
    END
  END ENABLE_VDDIO
  PIN EN_VDDIO_SIG_H
    ANTENNAPARTIALCUTAREA  0.157500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 22.360000 0.000000 22.660000 1.205000 ;
    END
    PORT
      LAYER met2 ;
        RECT  9.735000  4.520000 10.050000  4.575000 ;
        RECT  9.735000  4.575000  9.995000  4.630000 ;
        RECT  9.735000  4.630000  9.995000  8.860000 ;
        RECT  9.735000  8.860000  9.995000  8.915000 ;
        RECT  9.735000  8.915000 10.050000  8.970000 ;
        RECT  9.790000  4.465000 10.105000  4.520000 ;
        RECT  9.805000  8.970000 10.105000  9.040000 ;
        RECT  9.860000  4.395000 10.160000  4.465000 ;
        RECT  9.875000  9.040000 10.175000  9.110000 ;
        RECT  9.930000  4.325000 10.230000  4.395000 ;
        RECT  9.945000  9.110000 10.245000  9.180000 ;
        RECT 10.000000  4.255000 10.300000  4.325000 ;
        RECT 10.015000  9.180000 10.315000  9.250000 ;
        RECT 10.070000  4.185000 10.370000  4.255000 ;
        RECT 10.085000  9.250000 10.385000  9.320000 ;
        RECT 10.140000  4.115000 10.440000  4.185000 ;
        RECT 10.155000  9.320000 10.455000  9.390000 ;
        RECT 10.210000  4.045000 10.510000  4.115000 ;
        RECT 10.225000  9.390000 10.525000  9.460000 ;
        RECT 10.280000  3.975000 10.580000  4.045000 ;
        RECT 10.295000  9.460000 10.595000  9.530000 ;
        RECT 10.350000  3.905000 10.650000  3.975000 ;
        RECT 10.365000  9.530000 10.665000  9.600000 ;
        RECT 10.420000  3.835000 10.720000  3.905000 ;
        RECT 10.435000  9.600000 10.735000  9.670000 ;
        RECT 10.490000  3.765000 10.790000  3.835000 ;
        RECT 10.505000  9.670000 10.805000  9.740000 ;
        RECT 10.560000  3.695000 10.860000  3.765000 ;
        RECT 10.575000  9.740000 10.875000  9.810000 ;
        RECT 10.610000  3.645000 15.095000  3.695000 ;
        RECT 10.645000  9.810000 10.945000  9.880000 ;
        RECT 10.650000 26.825000 11.125000 27.085000 ;
        RECT 10.650000 27.085000 11.055000 27.155000 ;
        RECT 10.650000 27.155000 10.985000 27.225000 ;
        RECT 10.650000 27.225000 10.915000 27.295000 ;
        RECT 10.650000 27.295000 10.910000 27.300000 ;
        RECT 10.650000 27.300000 10.910000 27.935000 ;
        RECT 10.650000 27.935000 10.910000 28.005000 ;
        RECT 10.650000 28.005000 10.980000 28.075000 ;
        RECT 10.650000 28.075000 11.050000 28.145000 ;
        RECT 10.650000 28.145000 11.120000 28.150000 ;
        RECT 10.650000 28.150000 11.125000 28.410000 ;
        RECT 10.655000 26.820000 11.125000 26.825000 ;
        RECT 10.680000  3.575000 15.025000  3.645000 ;
        RECT 10.715000  9.880000 11.015000  9.950000 ;
        RECT 10.720000 28.410000 11.125000 28.480000 ;
        RECT 10.725000 26.750000 11.125000 26.820000 ;
        RECT 10.750000  3.505000 14.955000  3.575000 ;
        RECT 10.755000  9.950000 11.085000  9.990000 ;
        RECT 10.790000 28.480000 11.125000 28.550000 ;
        RECT 10.795000 26.680000 11.125000 26.750000 ;
        RECT 10.810000  9.990000 11.125000 10.045000 ;
        RECT 10.820000  3.435000 14.885000  3.505000 ;
        RECT 10.860000 28.550000 11.125000 28.620000 ;
        RECT 10.865000 10.045000 11.125000 10.100000 ;
        RECT 10.865000 10.100000 11.125000 26.610000 ;
        RECT 10.865000 26.610000 11.125000 26.680000 ;
        RECT 10.865000 28.620000 11.125000 28.625000 ;
        RECT 10.865000 28.625000 11.125000 31.085000 ;
        RECT 10.865000 31.085000 11.125000 31.140000 ;
        RECT 10.865000 31.140000 11.180000 31.195000 ;
        RECT 10.935000 31.195000 11.235000 31.265000 ;
        RECT 11.005000 31.265000 11.305000 31.335000 ;
        RECT 11.075000 31.335000 11.375000 31.405000 ;
        RECT 11.145000 31.405000 11.445000 31.475000 ;
        RECT 11.150000 31.475000 11.515000 31.480000 ;
        RECT 11.205000 31.480000 11.520000 31.535000 ;
        RECT 11.260000 31.535000 11.520000 31.590000 ;
        RECT 11.260000 31.590000 11.520000 36.020000 ;
        RECT 11.260000 36.020000 12.150000 36.280000 ;
        RECT 14.845000  3.695000 15.145000  3.765000 ;
        RECT 14.915000  3.765000 15.215000  3.835000 ;
        RECT 14.985000  3.835000 15.285000  3.905000 ;
        RECT 15.055000  3.905000 15.355000  3.975000 ;
        RECT 15.125000  3.975000 15.425000  4.045000 ;
        RECT 15.195000  4.045000 15.495000  4.115000 ;
        RECT 15.265000  4.115000 15.565000  4.185000 ;
        RECT 15.335000  4.185000 15.635000  4.255000 ;
        RECT 15.405000  4.255000 15.705000  4.325000 ;
        RECT 15.475000  4.325000 15.775000  4.395000 ;
        RECT 15.545000  4.395000 15.845000  4.465000 ;
        RECT 15.615000  4.465000 15.915000  4.535000 ;
        RECT 15.625000  4.535000 15.985000  4.545000 ;
        RECT 15.695000  4.545000 28.765000  4.615000 ;
        RECT 15.765000  4.615000 28.835000  4.685000 ;
        RECT 15.835000  4.685000 28.905000  4.755000 ;
        RECT 15.885000  4.755000 28.975000  4.805000 ;
        RECT 22.065000  4.540000 22.940000  4.545000 ;
        RECT 22.135000  4.470000 22.870000  4.540000 ;
        RECT 22.205000  4.400000 22.800000  4.470000 ;
        RECT 22.275000  4.330000 22.730000  4.400000 ;
        RECT 22.345000  4.260000 22.660000  4.330000 ;
        RECT 22.350000  4.255000 22.660000  4.260000 ;
        RECT 22.355000  4.250000 22.660000  4.255000 ;
        RECT 22.360000  0.000000 22.660000  4.245000 ;
        RECT 22.360000  4.245000 22.660000  4.250000 ;
        RECT 28.725000  4.805000 29.025000  4.875000 ;
        RECT 28.795000  4.875000 29.095000  4.945000 ;
        RECT 28.865000  4.945000 29.165000  5.015000 ;
        RECT 28.935000  5.015000 29.235000  5.085000 ;
        RECT 29.005000  5.085000 29.305000  5.155000 ;
        RECT 29.075000  5.155000 29.375000  5.225000 ;
        RECT 29.145000  5.225000 29.445000  5.295000 ;
        RECT 29.210000  5.295000 29.515000  5.360000 ;
        RECT 29.265000  5.360000 29.580000  5.415000 ;
        RECT 29.320000  5.415000 29.580000  5.470000 ;
        RECT 29.320000  5.470000 29.580000 10.975000 ;
        RECT 29.320000 10.975000 29.580000 11.030000 ;
        RECT 29.320000 11.030000 29.635000 11.085000 ;
        RECT 29.390000 11.085000 29.690000 11.155000 ;
        RECT 29.460000 11.155000 29.760000 11.225000 ;
        RECT 29.530000 11.225000 29.830000 11.295000 ;
        RECT 29.600000 11.295000 29.900000 11.365000 ;
        RECT 29.660000 11.365000 29.970000 11.425000 ;
        RECT 29.715000 11.425000 30.030000 11.480000 ;
        RECT 29.770000 11.480000 30.030000 11.535000 ;
        RECT 29.770000 11.535000 30.030000 15.645000 ;
        RECT 29.770000 15.645000 30.030000 15.700000 ;
        RECT 29.770000 15.700000 30.085000 15.755000 ;
        RECT 29.840000 15.755000 30.140000 15.825000 ;
        RECT 29.910000 15.825000 30.210000 15.895000 ;
        RECT 29.980000 15.895000 30.280000 15.965000 ;
        RECT 30.050000 15.965000 30.350000 16.035000 ;
        RECT 30.120000 16.035000 30.420000 16.105000 ;
        RECT 30.190000 16.105000 30.490000 16.175000 ;
        RECT 30.255000 16.175000 30.560000 16.240000 ;
        RECT 30.310000 16.240000 30.625000 16.295000 ;
        RECT 30.365000 16.295000 30.625000 16.350000 ;
        RECT 30.365000 16.350000 30.625000 20.495000 ;
    END
  END EN_VDDIO_SIG_H
  PIN FILT_IN_H
    ANTENNAPARTIALCUTAREA  0.960000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.075000 0.000000 21.225000 3.455000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.075000 0.000000 21.225000  6.670000 ;
        RECT 20.075000 6.670000 21.225000  6.820000 ;
        RECT 20.075000 6.820000 21.375000  6.970000 ;
        RECT 20.075000 6.970000 21.525000  7.120000 ;
        RECT 20.075000 7.120000 21.675000  7.150000 ;
        RECT 20.225000 7.150000 21.705000  7.300000 ;
        RECT 20.375000 7.300000 21.855000  7.450000 ;
        RECT 20.525000 7.450000 22.005000  7.600000 ;
        RECT 20.675000 7.600000 22.155000  7.750000 ;
        RECT 20.825000 7.750000 22.305000  7.900000 ;
        RECT 20.975000 7.900000 22.455000  8.050000 ;
        RECT 21.125000 8.050000 22.605000  8.200000 ;
        RECT 21.275000 8.200000 22.755000  8.350000 ;
        RECT 21.425000 8.350000 22.905000  8.500000 ;
        RECT 21.575000 8.500000 23.055000  8.650000 ;
        RECT 21.725000 8.650000 23.205000  8.800000 ;
        RECT 21.875000 8.800000 23.355000  8.950000 ;
        RECT 22.025000 8.950000 23.505000  9.100000 ;
        RECT 22.175000 9.100000 23.655000  9.250000 ;
        RECT 22.325000 9.250000 23.805000  9.400000 ;
        RECT 22.420000 9.400000 23.955000  9.495000 ;
        RECT 22.570000 9.495000 24.050000  9.645000 ;
        RECT 22.720000 9.645000 24.050000  9.795000 ;
        RECT 22.870000 9.795000 24.050000  9.945000 ;
        RECT 22.905000 9.945000 24.050000  9.980000 ;
        RECT 22.905000 9.980000 24.050000 12.265000 ;
    END
  END FILT_IN_H
  PIN INP_SEL_H
    ANTENNAGATEAREA  6.240000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.600000 11.420000 16.830000 12.310000 ;
        RECT 16.600000 12.310000 16.830000 12.360000 ;
        RECT 16.600000 12.360000 16.880000 12.410000 ;
        RECT 16.670000 12.410000 16.930000 12.480000 ;
        RECT 16.740000 12.480000 17.000000 12.550000 ;
        RECT 16.810000 12.550000 17.070000 12.620000 ;
        RECT 16.825000 12.620000 17.140000 12.635000 ;
        RECT 16.870000 12.635000 25.295000 12.680000 ;
        RECT 16.915000 12.680000 25.340000 12.725000 ;
        RECT 16.985000 12.725000 25.385000 12.795000 ;
        RECT 17.055000 12.795000 25.385000 12.865000 ;
        RECT 24.640000 12.615000 25.275000 12.635000 ;
        RECT 24.710000 12.545000 25.205000 12.615000 ;
        RECT 24.780000 12.475000 25.135000 12.545000 ;
        RECT 24.785000 12.470000 25.135000 12.475000 ;
        RECT 24.845000 12.410000 25.135000 12.470000 ;
        RECT 24.905000  0.000000 25.135000 12.350000 ;
        RECT 24.905000 12.350000 25.135000 12.410000 ;
        RECT 24.975000 12.865000 25.385000 12.935000 ;
        RECT 25.045000 12.935000 25.385000 13.005000 ;
        RECT 25.115000 13.005000 25.385000 13.075000 ;
        RECT 25.155000 13.075000 25.385000 13.115000 ;
        RECT 25.155000 13.115000 25.385000 15.035000 ;
        RECT 25.155000 15.035000 25.385000 15.085000 ;
        RECT 25.155000 15.085000 25.435000 15.135000 ;
        RECT 25.225000 15.135000 25.485000 15.205000 ;
        RECT 25.295000 15.205000 25.555000 15.275000 ;
        RECT 25.365000 15.275000 25.625000 15.345000 ;
        RECT 25.435000 15.345000 25.695000 15.415000 ;
        RECT 25.505000 15.415000 25.765000 15.485000 ;
        RECT 25.575000 15.485000 25.835000 15.555000 ;
        RECT 25.635000 15.555000 25.905000 15.615000 ;
        RECT 25.705000 15.615000 29.965000 15.685000 ;
        RECT 25.775000 15.685000 30.035000 15.755000 ;
        RECT 25.845000 15.755000 30.105000 15.825000 ;
        RECT 25.865000 15.825000 30.175000 15.845000 ;
        RECT 29.935000 15.845000 30.195000 15.915000 ;
        RECT 30.005000 15.915000 30.265000 15.985000 ;
        RECT 30.075000 15.985000 30.335000 16.055000 ;
        RECT 30.145000 16.055000 30.405000 16.125000 ;
        RECT 30.215000 16.125000 30.475000 16.195000 ;
        RECT 30.285000 16.195000 30.545000 16.265000 ;
        RECT 30.355000 16.265000 30.615000 16.335000 ;
        RECT 30.425000 16.335000 30.685000 16.405000 ;
        RECT 30.495000 16.405000 30.755000 16.475000 ;
        RECT 30.565000 16.475000 30.825000 16.545000 ;
        RECT 30.635000 16.545000 30.895000 16.615000 ;
        RECT 30.705000 16.615000 30.965000 16.685000 ;
        RECT 30.755000 16.685000 31.035000 16.735000 ;
        RECT 30.805000 16.735000 31.035000 16.785000 ;
        RECT 30.805000 16.785000 31.035000 19.345000 ;
    END
  END INP_SEL_H
  PIN PAD
    ANTENNAPARTIALMETALSIDEAREA  245.6270 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 29.695000 127.115000 41.990000 145.625000 ;
    END
  END PAD
  PIN PAD_A_ESD_H
    ANTENNAPARTIALCUTAREA  0.960000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.245000 0.000000 18.910000 3.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.245000 0.000000 18.910000 3.135000 ;
    END
  END PAD_A_ESD_H
  PIN PULLUP_H
    ANTENNAPARTIALCUTAREA  0.270000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  6.065000 43.285000 24.570000 43.355000 ;
        RECT  6.065000 43.355000 24.500000 43.425000 ;
        RECT  6.065000 43.425000 24.430000 43.495000 ;
        RECT  6.065000 43.495000 24.380000 43.545000 ;
        RECT 14.555000  0.000000 15.135000 12.210000 ;
        RECT 14.555000 12.210000 15.135000 12.275000 ;
        RECT 14.555000 12.275000 15.200000 12.340000 ;
        RECT 14.625000 12.340000 15.265000 12.410000 ;
        RECT 14.695000 12.410000 15.335000 12.480000 ;
        RECT 14.765000 12.480000 15.405000 12.550000 ;
        RECT 14.835000 12.550000 15.475000 12.620000 ;
        RECT 14.905000 12.620000 15.545000 12.690000 ;
        RECT 14.975000 12.690000 15.615000 12.760000 ;
        RECT 15.045000 12.760000 15.685000 12.830000 ;
        RECT 15.115000 12.830000 15.755000 12.900000 ;
        RECT 15.185000 12.900000 15.825000 12.970000 ;
        RECT 15.255000 12.970000 15.895000 13.040000 ;
        RECT 15.325000 13.040000 15.965000 13.110000 ;
        RECT 15.395000 13.110000 16.035000 13.180000 ;
        RECT 15.465000 13.180000 16.105000 13.250000 ;
        RECT 15.535000 13.250000 16.175000 13.320000 ;
        RECT 15.605000 13.320000 16.245000 13.390000 ;
        RECT 15.675000 13.390000 16.315000 13.460000 ;
        RECT 15.745000 13.460000 16.385000 13.530000 ;
        RECT 15.815000 13.530000 16.455000 13.600000 ;
        RECT 15.885000 13.600000 16.525000 13.670000 ;
        RECT 15.955000 13.670000 16.595000 13.740000 ;
        RECT 16.025000 13.740000 16.665000 13.810000 ;
        RECT 16.095000 13.810000 16.735000 13.880000 ;
        RECT 16.165000 13.880000 16.805000 13.950000 ;
        RECT 16.235000 13.950000 16.875000 14.020000 ;
        RECT 16.305000 14.020000 16.945000 14.090000 ;
        RECT 16.375000 14.090000 17.015000 14.160000 ;
        RECT 16.445000 14.160000 17.085000 14.230000 ;
        RECT 16.515000 14.230000 17.155000 14.300000 ;
        RECT 16.585000 14.300000 17.225000 14.370000 ;
        RECT 16.655000 14.370000 17.295000 14.440000 ;
        RECT 16.725000 14.440000 17.365000 14.510000 ;
        RECT 16.795000 14.510000 17.435000 14.580000 ;
        RECT 16.865000 14.580000 17.505000 14.650000 ;
        RECT 16.935000 14.650000 17.575000 14.720000 ;
        RECT 17.005000 14.720000 17.645000 14.790000 ;
        RECT 17.075000 14.790000 17.715000 14.860000 ;
        RECT 17.145000 14.860000 17.785000 14.930000 ;
        RECT 17.215000 14.930000 17.855000 15.000000 ;
        RECT 17.285000 15.000000 17.925000 15.070000 ;
        RECT 17.355000 15.070000 17.995000 15.140000 ;
        RECT 17.425000 15.140000 18.065000 15.210000 ;
        RECT 17.495000 15.210000 18.135000 15.280000 ;
        RECT 17.565000 15.280000 18.205000 15.350000 ;
        RECT 17.635000 15.350000 18.275000 15.420000 ;
        RECT 17.705000 15.420000 21.745000 15.490000 ;
        RECT 17.775000 15.490000 21.815000 15.560000 ;
        RECT 17.845000 15.560000 21.885000 15.630000 ;
        RECT 17.915000 15.630000 21.955000 15.700000 ;
        RECT 17.985000 15.700000 22.025000 15.770000 ;
        RECT 18.055000 15.770000 22.095000 15.840000 ;
        RECT 18.125000 15.840000 22.165000 15.910000 ;
        RECT 18.135000 15.910000 22.235000 15.920000 ;
        RECT 21.605000 15.920000 22.245000 15.990000 ;
        RECT 21.675000 15.990000 22.315000 16.060000 ;
        RECT 21.745000 16.060000 22.385000 16.130000 ;
        RECT 21.815000 16.130000 22.455000 16.200000 ;
        RECT 21.885000 16.200000 22.525000 16.270000 ;
        RECT 21.955000 16.270000 22.595000 16.340000 ;
        RECT 22.025000 16.340000 22.665000 16.410000 ;
        RECT 22.095000 16.410000 22.735000 16.480000 ;
        RECT 22.165000 16.480000 22.805000 16.550000 ;
        RECT 22.235000 16.550000 22.875000 16.620000 ;
        RECT 22.305000 16.620000 22.945000 16.690000 ;
        RECT 22.375000 16.690000 23.015000 16.760000 ;
        RECT 22.445000 16.760000 23.085000 16.830000 ;
        RECT 22.515000 16.830000 23.155000 16.900000 ;
        RECT 22.585000 16.900000 23.225000 16.970000 ;
        RECT 22.655000 16.970000 23.295000 17.040000 ;
        RECT 22.725000 17.040000 23.365000 17.110000 ;
        RECT 22.795000 17.110000 23.435000 17.180000 ;
        RECT 22.865000 17.180000 23.505000 17.250000 ;
        RECT 22.935000 17.250000 23.575000 17.320000 ;
        RECT 23.005000 17.320000 23.645000 17.390000 ;
        RECT 23.075000 17.390000 23.715000 17.460000 ;
        RECT 23.145000 17.460000 23.785000 17.530000 ;
        RECT 23.215000 17.530000 23.855000 17.600000 ;
        RECT 23.285000 17.600000 23.925000 17.670000 ;
        RECT 23.355000 17.670000 23.995000 17.740000 ;
        RECT 23.425000 17.740000 24.065000 17.810000 ;
        RECT 23.495000 17.810000 24.135000 17.880000 ;
        RECT 23.565000 17.880000 24.205000 17.950000 ;
        RECT 23.635000 17.950000 24.275000 18.020000 ;
        RECT 23.705000 18.020000 24.345000 18.090000 ;
        RECT 23.775000 18.090000 24.415000 18.160000 ;
        RECT 23.845000 18.160000 24.485000 18.230000 ;
        RECT 23.915000 18.230000 24.555000 18.300000 ;
        RECT 23.985000 18.300000 24.625000 18.370000 ;
        RECT 24.015000 18.370000 24.695000 18.400000 ;
        RECT 24.085000 18.400000 24.725000 18.470000 ;
        RECT 24.155000 18.470000 24.725000 18.540000 ;
        RECT 24.225000 18.540000 24.725000 18.610000 ;
        RECT 24.225000 18.610000 24.725000 25.145000 ;
        RECT 24.225000 25.145000 24.725000 25.215000 ;
        RECT 24.225000 25.215000 24.795000 25.285000 ;
        RECT 24.225000 25.285000 24.865000 25.355000 ;
        RECT 24.295000 25.355000 24.935000 25.425000 ;
        RECT 24.325000 43.230000 24.640000 43.285000 ;
        RECT 24.365000 25.425000 25.005000 25.495000 ;
        RECT 24.395000 43.160000 24.695000 43.230000 ;
        RECT 24.435000 25.495000 25.075000 25.565000 ;
        RECT 24.465000 43.090000 24.765000 43.160000 ;
        RECT 24.505000 25.565000 25.145000 25.635000 ;
        RECT 24.535000 43.020000 24.835000 43.090000 ;
        RECT 24.575000 25.635000 25.215000 25.705000 ;
        RECT 24.605000 25.705000 25.285000 25.735000 ;
        RECT 24.605000 42.950000 24.905000 43.020000 ;
        RECT 24.675000 25.735000 25.315000 25.805000 ;
        RECT 24.675000 42.880000 24.975000 42.950000 ;
        RECT 24.745000 25.805000 25.315000 25.875000 ;
        RECT 24.745000 42.810000 25.045000 42.880000 ;
        RECT 24.815000 25.875000 25.315000 25.945000 ;
        RECT 24.815000 25.945000 25.315000 42.610000 ;
        RECT 24.815000 42.610000 25.250000 42.675000 ;
        RECT 24.815000 42.675000 25.185000 42.740000 ;
        RECT 24.815000 42.740000 25.115000 42.810000 ;
    END
    PORT
      LAYER met2 ;
        RECT 14.555000 0.000000 15.135000 0.985000 ;
    END
  END PULLUP_H
  PIN TIE_HI_ESD
    ANTENNAPARTIALCUTAREA  0.045000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 28.185000 4.895000 30.220000 4.965000 ;
        RECT 28.185000 4.965000 30.150000 5.035000 ;
        RECT 28.185000 5.035000 30.080000 5.105000 ;
        RECT 28.185000 5.105000 30.010000 5.175000 ;
        RECT 28.185000 5.175000 29.940000 5.245000 ;
        RECT 28.185000 5.245000 29.870000 5.315000 ;
        RECT 28.185000 5.315000 29.800000 5.385000 ;
        RECT 28.185000 5.385000 29.730000 5.455000 ;
        RECT 28.185000 5.455000 29.660000 5.525000 ;
        RECT 28.185000 5.525000 29.640000 5.545000 ;
        RECT 29.395000 4.870000 30.290000 4.895000 ;
        RECT 29.465000 4.800000 30.315000 4.870000 ;
        RECT 29.535000 4.730000 30.385000 4.800000 ;
        RECT 29.605000 4.660000 30.455000 4.730000 ;
        RECT 29.675000 4.590000 30.525000 4.660000 ;
        RECT 29.745000 4.520000 30.595000 4.590000 ;
        RECT 29.815000 4.450000 30.665000 4.520000 ;
        RECT 29.885000 4.380000 30.735000 4.450000 ;
        RECT 29.955000 4.310000 30.805000 4.380000 ;
        RECT 30.025000 4.240000 30.875000 4.310000 ;
        RECT 30.095000 4.170000 30.945000 4.240000 ;
        RECT 30.165000 4.100000 31.015000 4.170000 ;
        RECT 30.235000 4.030000 31.085000 4.100000 ;
        RECT 30.295000 3.970000 31.155000 4.030000 ;
        RECT 30.365000 3.900000 31.155000 3.970000 ;
        RECT 30.435000 3.830000 31.155000 3.900000 ;
        RECT 30.505000 0.000000 31.155000 3.760000 ;
        RECT 30.505000 3.760000 31.155000 3.830000 ;
    END
    PORT
      LAYER met2 ;
        RECT 30.505000 0.000000 31.155000 0.330000 ;
    END
  END TIE_HI_ESD
  PIN TIE_LO_ESD
    ANTENNAPARTIALCUTAREA  0.045000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 27.580000 0.000000 28.230000 2.855000 ;
        RECT 27.580000 2.855000 28.230000 2.925000 ;
        RECT 27.580000 2.925000 28.300000 2.995000 ;
        RECT 27.580000 2.995000 28.370000 3.065000 ;
        RECT 27.580000 3.065000 28.440000 3.125000 ;
        RECT 27.650000 3.125000 28.500000 3.195000 ;
        RECT 27.720000 3.195000 28.570000 3.265000 ;
        RECT 27.790000 3.265000 28.640000 3.335000 ;
        RECT 27.860000 3.335000 28.710000 3.405000 ;
        RECT 27.915000 3.405000 28.780000 3.460000 ;
        RECT 27.985000 3.460000 28.835000 3.530000 ;
        RECT 28.055000 3.530000 28.835000 3.600000 ;
        RECT 28.125000 3.600000 28.835000 3.670000 ;
        RECT 28.185000 3.670000 28.835000 3.730000 ;
        RECT 28.185000 3.730000 28.835000 4.105000 ;
    END
    PORT
      LAYER met2 ;
        RECT 27.580000 0.000000 28.230000 0.330000 ;
    END
  END TIE_LO_ESD
  PIN TIE_WEAK_HI_H
    ANTENNAPARTIALCUTAREA  0.520000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.215000 0.000000 73.235000 0.770000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.860000 71.930000 66.310000 72.080000 ;
        RECT 64.860000 72.080000 66.160000 72.230000 ;
        RECT 64.860000 72.230000 66.010000 72.380000 ;
        RECT 64.860000 72.380000 65.990000 72.400000 ;
        RECT 64.860000 72.400000 65.990000 94.645000 ;
        RECT 64.990000 71.800000 66.460000 71.930000 ;
        RECT 65.140000 71.650000 66.590000 71.800000 ;
        RECT 65.290000 71.500000 66.740000 71.650000 ;
        RECT 65.440000 71.350000 66.890000 71.500000 ;
        RECT 65.590000 71.200000 67.040000 71.350000 ;
        RECT 65.740000 71.050000 67.190000 71.200000 ;
        RECT 65.890000 70.900000 67.340000 71.050000 ;
        RECT 66.040000 70.750000 67.490000 70.900000 ;
        RECT 66.190000 70.600000 67.640000 70.750000 ;
        RECT 66.340000 70.450000 67.790000 70.600000 ;
        RECT 66.490000 70.300000 67.940000 70.450000 ;
        RECT 66.640000 70.150000 68.090000 70.300000 ;
        RECT 66.790000 70.000000 68.240000 70.150000 ;
        RECT 66.940000 69.850000 68.390000 70.000000 ;
        RECT 67.090000 69.700000 68.540000 69.850000 ;
        RECT 67.240000 69.550000 68.690000 69.700000 ;
        RECT 67.390000 69.400000 68.840000 69.550000 ;
        RECT 67.540000 69.250000 68.990000 69.400000 ;
        RECT 67.690000 69.100000 69.140000 69.250000 ;
        RECT 67.840000 68.950000 69.290000 69.100000 ;
        RECT 67.990000 68.800000 69.440000 68.950000 ;
        RECT 68.140000 68.650000 69.590000 68.800000 ;
        RECT 68.290000 68.500000 69.740000 68.650000 ;
        RECT 68.440000 68.350000 69.890000 68.500000 ;
        RECT 68.590000 68.200000 70.040000 68.350000 ;
        RECT 68.740000 68.050000 70.190000 68.200000 ;
        RECT 68.890000 67.900000 70.340000 68.050000 ;
        RECT 69.040000 67.750000 70.490000 67.900000 ;
        RECT 69.190000 67.600000 70.640000 67.750000 ;
        RECT 69.340000 67.450000 70.790000 67.600000 ;
        RECT 69.490000 67.300000 70.940000 67.450000 ;
        RECT 69.640000 67.150000 71.090000 67.300000 ;
        RECT 69.790000 67.000000 71.240000 67.150000 ;
        RECT 69.940000 66.850000 71.390000 67.000000 ;
        RECT 70.090000 66.700000 71.540000 66.850000 ;
        RECT 70.240000 66.550000 71.690000 66.700000 ;
        RECT 70.390000 66.400000 71.840000 66.550000 ;
        RECT 70.540000 66.250000 71.990000 66.400000 ;
        RECT 70.690000 66.100000 72.140000 66.250000 ;
        RECT 70.840000 65.950000 72.290000 66.100000 ;
        RECT 70.990000 65.800000 72.440000 65.950000 ;
        RECT 71.140000 65.650000 72.590000 65.800000 ;
        RECT 71.290000 65.500000 72.740000 65.650000 ;
        RECT 71.440000 65.350000 72.890000 65.500000 ;
        RECT 71.590000 65.200000 73.040000 65.350000 ;
        RECT 71.740000 65.050000 73.190000 65.200000 ;
        RECT 71.890000 64.900000 73.340000 65.050000 ;
        RECT 72.040000 64.750000 73.490000 64.900000 ;
        RECT 72.190000  0.000000 73.260000 49.320000 ;
        RECT 72.190000 49.320000 73.260000 49.470000 ;
        RECT 72.190000 49.470000 73.410000 49.620000 ;
        RECT 72.190000 49.620000 73.560000 49.770000 ;
        RECT 72.190000 49.770000 73.710000 49.920000 ;
        RECT 72.190000 49.920000 73.860000 49.985000 ;
        RECT 72.190000 49.985000 73.925000 64.465000 ;
        RECT 72.190000 64.465000 73.860000 64.530000 ;
        RECT 72.190000 64.530000 73.795000 64.595000 ;
        RECT 72.190000 64.595000 73.790000 64.600000 ;
        RECT 72.190000 64.600000 73.640000 64.750000 ;
    END
  END TIE_WEAK_HI_H
  PIN XRES_H_N
    ANTENNAPARTIALCUTAREA  0.240000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.915000 0.000000 29.685000 0.335000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.170000 10.610000 29.050000 10.760000 ;
        RECT 28.170000 10.760000 28.900000 10.910000 ;
        RECT 28.170000 10.910000 28.900000 14.770000 ;
        RECT 28.185000 10.595000 29.200000 10.610000 ;
        RECT 28.335000 10.445000 29.215000 10.595000 ;
        RECT 28.485000 10.295000 29.365000 10.445000 ;
        RECT 28.635000 10.145000 29.515000 10.295000 ;
        RECT 28.785000  9.995000 29.665000 10.145000 ;
        RECT 28.935000  0.000000 29.665000  9.845000 ;
        RECT 28.935000  9.845000 29.665000  9.995000 ;
    END
  END XRES_H_N
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 1.270000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 8.885000 75.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 1.270000 13.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 2.035000 75.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 1.270000 7.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 14.935000 75.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 0.965000 18.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 1.270000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 19.785000 75.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 70.035000 75.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 1.270000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 1.270000 94.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 19.885000 75.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 1.270000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 64.085000 75.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 1.270000 68.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 1.270000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 1.270000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 36.735000 75.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 47.735000 75.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.645000 75.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.405000 75.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.840000 1.270000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 1.270000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 36.840000 75.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 1.270000 41.655000 ;
        RECT 0.000000 41.655000 3.720000 46.170000 ;
        RECT 0.000000 46.170000 1.270000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.655000 41.630000 75.000000 46.190000 ;
        RECT 73.730000 41.585000 75.000000 41.630000 ;
        RECT 73.730000 46.190000 75.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 1.270000 46.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 1.270000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 25.835000 75.000000 30.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 1.270000 30.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 1.270000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 58.235000 75.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 1.270000 62.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 31.885000 75.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 1.270000 35.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT -0.265000 125.265000 75.000000 129.185000 ;
      RECT -0.265000 129.185000 41.620000 130.225000 ;
      RECT -0.160000 140.815000 75.160000 144.435000 ;
      RECT  0.000000  96.860000 58.340000  96.865000 ;
      RECT  0.000000  96.865000 75.000000  97.865000 ;
      RECT  0.000000  97.865000 58.340000  99.360000 ;
      RECT  0.000000  99.360000 75.000000 101.740000 ;
      RECT  0.000000 101.740000 58.340000 101.780000 ;
      RECT  0.000000 101.780000  0.165000 102.385000 ;
      RECT  0.000000 102.385000  0.455000 102.395000 ;
      RECT  0.000000 102.395000  0.595000 125.265000 ;
      RECT  0.000000 130.995000 38.355000 131.325000 ;
      RECT  0.000000 131.325000 13.200000 134.390000 ;
      RECT  0.000000 134.390000 75.000000 134.950000 ;
      RECT  0.000000 134.950000 52.445000 136.970000 ;
      RECT  0.000000 136.970000  1.045000 138.600000 ;
      RECT  0.000000 138.600000 75.000000 140.050000 ;
      RECT  0.700000 130.425000 42.015000 130.795000 ;
      RECT  0.700000 130.795000 38.355000 130.995000 ;
      RECT  0.985000   0.185000 33.890000   0.645000 ;
      RECT  0.985000   0.645000  4.525000   3.740000 ;
      RECT  0.985000   3.740000  7.065000   4.105000 ;
      RECT  0.985000 101.780000  2.645000 102.395000 ;
      RECT  1.015000   4.105000  7.065000   8.600000 ;
      RECT  1.015000   8.600000  5.625000  12.860000 ;
      RECT  1.015000  12.860000  6.055000  13.870000 ;
      RECT  1.015000  13.870000  5.625000  17.770000 ;
      RECT  1.015000  17.770000 14.130000  18.870000 ;
      RECT  1.015000  18.870000  5.605000  37.435000 ;
      RECT  1.015000  37.435000 14.270000  38.625000 ;
      RECT  1.015000  38.625000  4.525000  71.780000 ;
      RECT  1.015000  71.780000 31.450000  84.665000 ;
      RECT  1.100000  85.320000  2.790000  96.860000 ;
      RECT  1.145000  84.665000 31.450000  85.320000 ;
      RECT 11.005000  17.765000 11.270000  17.770000 ;
      RECT 11.270000  18.870000 14.130000  25.580000 ;
      RECT 13.095000   3.770000 16.800000   6.465000 ;
      RECT 13.095000   6.465000 32.410000   6.520000 ;
      RECT 13.095000   6.520000 32.395000   8.665000 ;
      RECT 13.460000  25.580000 14.130000  27.375000 ;
      RECT 13.460000  27.375000 20.685000  27.545000 ;
      RECT 13.460000  27.545000 14.130000  34.045000 ;
      RECT 14.130000 136.970000 52.445000 137.930000 ;
      RECT 14.130000 137.930000 75.000000 138.600000 ;
      RECT 14.165000  13.360000 14.435000  13.735000 ;
      RECT 14.185000   8.665000 14.385000  12.750000 ;
      RECT 14.480000  13.050000 24.760000  15.670000 ;
      RECT 16.115000  10.105000 16.285000  10.160000 ;
      RECT 16.115000  10.160000 16.800000  10.330000 ;
      RECT 16.115000  10.330000 16.285000  10.635000 ;
      RECT 16.130000  11.590000 16.800000  11.760000 ;
      RECT 16.630000  11.480000 16.800000  11.590000 ;
      RECT 16.630000  11.760000 16.800000  12.010000 ;
      RECT 16.950000  15.670000 24.760000  15.930000 ;
      RECT 16.950000  15.930000 32.350000  16.600000 ;
      RECT 16.950000  16.600000 26.460000  18.815000 ;
      RECT 17.885000   0.645000 33.890000   3.235000 ;
      RECT 18.700000  18.815000 26.460000  20.255000 ;
      RECT 18.885000  24.405000 20.685000  27.375000 ;
      RECT 19.155000  39.220000 26.270000  41.890000 ;
      RECT 19.155000  41.890000 32.495000  42.120000 ;
      RECT 19.155000  42.120000 32.435000  43.020000 ;
      RECT 20.685000  20.255000 26.460000  20.490000 ;
      RECT 20.855000  20.490000 26.460000  21.035000 ;
      RECT 20.855000  24.480000 26.460000  25.800000 ;
      RECT 21.135000  37.530000 26.270000  39.220000 ;
      RECT 23.730000  21.035000 26.460000  24.480000 ;
      RECT 24.035000 131.325000 25.835000 134.390000 ;
      RECT 24.435000  11.465000 25.140000  11.995000 ;
      RECT 24.470000   9.975000 25.105000  10.160000 ;
      RECT 24.470000  10.160000 25.140000  10.330000 ;
      RECT 24.470000  10.330000 25.105000  10.505000 ;
      RECT 25.070000  25.800000 26.460000  26.780000 ;
      RECT 25.070000  26.780000 32.625000  27.950000 ;
      RECT 25.070000  27.950000 27.385000  33.830000 ;
      RECT 25.070000  33.830000 32.435000  33.940000 ;
      RECT 25.070000  33.940000 32.495000  34.170000 ;
      RECT 25.070000  34.170000 26.270000  37.530000 ;
      RECT 25.140000  47.770000 31.450000  71.780000 ;
      RECT 26.480000  14.880000 26.650000  15.410000 ;
      RECT 26.975000  34.730000 31.525000  34.960000 ;
      RECT 26.975000  34.960000 27.205000  40.965000 ;
      RECT 26.975000  40.965000 31.525000  41.195000 ;
      RECT 27.370000  17.445000 27.540000  25.820000 ;
      RECT 27.760000  14.880000 27.930000  15.410000 ;
      RECT 27.850000  35.215000 30.690000  35.385000 ;
      RECT 28.665000  30.760000 28.835000  31.290000 ;
      RECT 28.665000  31.845000 28.835000  32.375000 ;
      RECT 29.035000  28.960000 29.205000  29.490000 ;
      RECT 29.035000  30.070000 29.205000  30.600000 ;
      RECT 29.065000  31.460000 29.595000  31.630000 ;
      RECT 29.150000  18.365000 29.680000  18.535000 ;
      RECT 29.150000  20.125000 29.680000  20.295000 ;
      RECT 29.330000  24.890000 30.490000  25.220000 ;
      RECT 29.455000   3.235000 32.410000   6.465000 ;
      RECT 30.105000  25.405000 30.635000  25.575000 ;
      RECT 30.115000  29.700000 30.645000  29.870000 ;
      RECT 30.215000  14.720000 30.385000  15.250000 ;
      RECT 30.415000  19.390000 30.585000  19.920000 ;
      RECT 30.415000  20.510000 30.585000  21.040000 ;
      RECT 30.835000  17.635000 31.005000  18.165000 ;
      RECT 30.835000  18.755000 31.005000  19.285000 ;
      RECT 30.960000  46.750000 31.490000  46.920000 ;
      RECT 31.130000  46.485000 31.490000  46.750000 ;
      RECT 31.130000  46.920000 31.490000  47.155000 ;
      RECT 31.295000  34.960000 31.525000  40.965000 ;
      RECT 31.495000  14.720000 31.665000  15.250000 ;
      RECT 32.155000  28.780000 32.325000  32.550000 ;
      RECT 32.265000  34.170000 32.495000  41.890000 ;
      RECT 33.420000  73.960000 33.870000  81.465000 ;
      RECT 33.445000  82.260000 34.600000  83.340000 ;
      RECT 33.535000  81.905000 34.065000  82.075000 ;
      RECT 34.850000  83.100000 35.380000  83.270000 ;
      RECT 35.090000   0.900000 38.860000   1.070000 ;
      RECT 35.160000   1.070000 38.860000   1.080000 ;
      RECT 36.555000 131.325000 38.355000 134.390000 ;
      RECT 38.970000 133.145000 40.600000 133.825000 ;
      RECT 40.040000   0.195000 74.560000   5.755000 ;
      RECT 40.335000   5.755000 74.560000   5.960000 ;
      RECT 40.495000 130.795000 42.015000 130.995000 ;
      RECT 40.495000 130.995000 75.000000 132.595000 ;
      RECT 42.840000 129.770000 43.730000 130.440000 ;
      RECT 43.350000  60.495000 43.720000  78.760000 ;
      RECT 48.290000 129.770000 50.440000 130.440000 ;
      RECT 51.880000 133.145000 52.770000 133.815000 ;
      RECT 53.575000 135.430000 55.095000 137.450000 ;
      RECT 53.970000   5.960000 74.560000   6.580000 ;
      RECT 55.000000 129.770000 56.460000 130.440000 ;
      RECT 58.340000 102.310000 72.060000 102.395000 ;
      RECT 60.770000 133.145000 61.800000 133.815000 ;
      RECT 60.855000 129.760000 61.780000 130.430000 ;
      RECT 62.040000 129.185000 75.000000 130.225000 ;
      RECT 62.065000 132.595000 75.000000 134.390000 ;
      RECT 62.730000   6.580000 63.170000  59.670000 ;
      RECT 63.130000  60.940000 63.180000  85.005000 ;
      RECT 67.105000 134.950000 75.000000 137.930000 ;
      RECT 68.960000  85.895000 71.490000  86.125000 ;
      RECT 68.960000  86.125000 74.315000  94.410000 ;
      RECT 69.260000  94.410000 74.315000  96.865000 ;
      RECT 72.060000  97.865000 75.000000  99.360000 ;
      RECT 72.060000 101.740000 75.000000 101.780000 ;
      RECT 73.265000   6.580000 74.560000  84.995000 ;
      RECT 73.265000  84.995000 73.855000  85.020000 ;
      RECT 74.355000 101.780000 75.000000 125.265000 ;
    LAYER met1 ;
      RECT -0.145000  95.895000  2.680000  95.965000 ;
      RECT -0.145000  95.965000  2.750000  96.035000 ;
      RECT -0.145000  96.035000  2.820000  96.105000 ;
      RECT -0.145000  96.105000  2.890000  96.175000 ;
      RECT -0.145000  96.175000  2.960000  96.245000 ;
      RECT -0.145000  96.245000  3.030000  96.315000 ;
      RECT -0.145000  96.315000  3.100000  96.385000 ;
      RECT -0.145000  96.385000  3.170000  96.455000 ;
      RECT -0.145000  96.455000  3.240000  96.525000 ;
      RECT -0.145000  96.525000  3.310000  96.595000 ;
      RECT -0.145000  96.545000  3.325000  96.610000 ;
      RECT -0.145000  96.545000  3.325000  96.610000 ;
      RECT -0.145000  96.595000  3.380000  96.665000 ;
      RECT -0.145000  96.610000  3.395000  96.680000 ;
      RECT -0.145000  96.610000  3.395000  96.680000 ;
      RECT -0.145000  96.665000  3.450000  96.735000 ;
      RECT -0.145000  96.680000  3.465000  96.750000 ;
      RECT -0.145000  96.680000  3.465000  96.750000 ;
      RECT -0.145000  96.735000  3.520000  96.805000 ;
      RECT -0.145000  96.750000  3.535000  96.820000 ;
      RECT -0.145000  96.750000  3.535000  96.820000 ;
      RECT -0.145000  96.805000  3.590000  96.875000 ;
      RECT -0.145000  96.820000  3.605000  96.890000 ;
      RECT -0.145000  96.820000  3.605000  96.890000 ;
      RECT -0.145000  96.875000  3.660000  96.945000 ;
      RECT -0.145000  96.890000  3.675000  96.960000 ;
      RECT -0.145000  96.890000  3.675000  96.960000 ;
      RECT -0.145000  96.945000  3.730000  97.015000 ;
      RECT -0.145000  96.960000  3.745000  97.030000 ;
      RECT -0.145000  96.960000  3.745000  97.030000 ;
      RECT -0.145000  97.015000  3.800000  97.085000 ;
      RECT -0.145000  97.030000  3.815000  97.100000 ;
      RECT -0.145000  97.030000  3.815000  97.100000 ;
      RECT -0.145000  97.085000  3.870000  97.155000 ;
      RECT -0.145000  97.100000  3.885000  97.170000 ;
      RECT -0.145000  97.100000  3.885000  97.170000 ;
      RECT -0.145000  97.155000  3.940000  97.225000 ;
      RECT -0.145000  97.170000  3.955000  97.240000 ;
      RECT -0.145000  97.170000  3.955000  97.240000 ;
      RECT -0.145000  97.225000  4.010000  97.295000 ;
      RECT -0.145000  97.240000  4.025000  97.310000 ;
      RECT -0.145000  97.240000  4.025000  97.310000 ;
      RECT -0.145000  97.295000  4.080000  97.365000 ;
      RECT -0.145000  97.310000  4.095000  97.380000 ;
      RECT -0.145000  97.310000  4.095000  97.380000 ;
      RECT -0.145000  97.365000  4.150000  97.435000 ;
      RECT -0.145000  97.380000  4.165000  97.450000 ;
      RECT -0.145000  97.380000  4.165000  97.450000 ;
      RECT -0.145000  97.435000  4.220000  97.505000 ;
      RECT -0.145000  97.450000  4.235000  97.520000 ;
      RECT -0.145000  97.450000  4.235000  97.520000 ;
      RECT -0.145000  97.505000  4.290000  97.530000 ;
      RECT -0.145000  97.520000  4.305000  97.530000 ;
      RECT -0.145000  97.520000  4.305000  97.530000 ;
      RECT -0.145000  97.530000 56.545000 100.330000 ;
      RECT -0.145000 100.330000 56.545000 101.420000 ;
      RECT -0.145000 125.440000 14.680000 125.510000 ;
      RECT -0.145000 125.440000 14.680000 125.510000 ;
      RECT -0.145000 125.510000 14.610000 125.580000 ;
      RECT -0.145000 125.510000 14.610000 125.580000 ;
      RECT -0.145000 125.580000 14.540000 125.650000 ;
      RECT -0.145000 125.580000 14.540000 125.650000 ;
      RECT -0.145000 125.650000 14.470000 125.720000 ;
      RECT -0.145000 125.650000 14.470000 125.720000 ;
      RECT -0.145000 125.720000 14.400000 125.790000 ;
      RECT -0.145000 125.720000 14.400000 125.790000 ;
      RECT -0.145000 125.790000 14.330000 125.860000 ;
      RECT -0.145000 125.790000 14.330000 125.860000 ;
      RECT -0.145000 125.860000 14.260000 125.930000 ;
      RECT -0.145000 125.860000 14.260000 125.930000 ;
      RECT -0.145000 125.930000 14.190000 126.000000 ;
      RECT -0.145000 125.930000 14.190000 126.000000 ;
      RECT -0.145000 126.000000 14.120000 126.070000 ;
      RECT -0.145000 126.000000 14.120000 126.070000 ;
      RECT -0.145000 126.070000 14.050000 126.140000 ;
      RECT -0.145000 126.070000 14.050000 126.140000 ;
      RECT -0.145000 126.140000 13.980000 126.210000 ;
      RECT -0.145000 126.140000 13.980000 126.210000 ;
      RECT -0.145000 126.210000 13.910000 126.280000 ;
      RECT -0.145000 126.210000 13.910000 126.280000 ;
      RECT -0.145000 126.280000 13.840000 126.350000 ;
      RECT -0.145000 126.280000 13.840000 126.350000 ;
      RECT -0.145000 126.350000 13.770000 126.420000 ;
      RECT -0.145000 126.350000 13.770000 126.420000 ;
      RECT -0.145000 126.420000 13.700000 126.490000 ;
      RECT -0.145000 126.420000 13.700000 126.490000 ;
      RECT -0.145000 126.490000 13.630000 126.560000 ;
      RECT -0.145000 126.490000 13.630000 126.560000 ;
      RECT -0.145000 126.560000 13.560000 126.630000 ;
      RECT -0.145000 126.560000 13.560000 126.630000 ;
      RECT -0.145000 126.630000 13.490000 126.700000 ;
      RECT -0.145000 126.630000 13.490000 126.700000 ;
      RECT -0.145000 126.700000 13.420000 126.770000 ;
      RECT -0.145000 126.700000 13.420000 126.770000 ;
      RECT -0.145000 126.770000 13.350000 126.840000 ;
      RECT -0.145000 126.770000 13.350000 126.840000 ;
      RECT -0.145000 126.840000 13.280000 126.910000 ;
      RECT -0.145000 126.840000 13.280000 126.910000 ;
      RECT -0.145000 126.910000 13.210000 126.980000 ;
      RECT -0.145000 126.910000 13.210000 126.980000 ;
      RECT -0.145000 126.980000 13.140000 127.050000 ;
      RECT -0.145000 126.980000 13.140000 127.050000 ;
      RECT -0.145000 127.050000 13.070000 127.120000 ;
      RECT -0.145000 127.050000 13.070000 127.120000 ;
      RECT -0.145000 127.120000 13.000000 127.190000 ;
      RECT -0.145000 127.120000 13.000000 127.190000 ;
      RECT -0.145000 127.190000 12.930000 127.260000 ;
      RECT -0.145000 127.190000 12.930000 127.260000 ;
      RECT -0.145000 127.260000 12.860000 127.330000 ;
      RECT -0.145000 127.260000 12.860000 127.330000 ;
      RECT -0.145000 127.330000 12.790000 127.400000 ;
      RECT -0.145000 127.330000 12.790000 127.400000 ;
      RECT -0.145000 127.400000 12.720000 127.470000 ;
      RECT -0.145000 127.400000 12.720000 127.470000 ;
      RECT -0.145000 127.470000 12.650000 127.540000 ;
      RECT -0.145000 127.470000 12.650000 127.540000 ;
      RECT -0.145000 127.540000 12.580000 127.610000 ;
      RECT -0.145000 127.540000 12.580000 127.610000 ;
      RECT -0.145000 127.610000 12.510000 127.680000 ;
      RECT -0.145000 127.610000 12.510000 127.680000 ;
      RECT -0.145000 127.680000 12.440000 127.750000 ;
      RECT -0.145000 127.680000 12.440000 127.750000 ;
      RECT -0.145000 127.750000 12.370000 127.820000 ;
      RECT -0.145000 127.750000 12.370000 127.820000 ;
      RECT -0.145000 127.820000 12.300000 127.890000 ;
      RECT -0.145000 127.820000 12.300000 127.890000 ;
      RECT -0.145000 127.890000 12.230000 127.960000 ;
      RECT -0.145000 127.890000 12.230000 127.960000 ;
      RECT -0.145000 127.960000 12.160000 128.030000 ;
      RECT -0.145000 127.960000 12.160000 128.030000 ;
      RECT -0.145000 128.030000 12.090000 128.100000 ;
      RECT -0.145000 128.030000 12.090000 128.100000 ;
      RECT -0.145000 128.100000 12.020000 128.170000 ;
      RECT -0.145000 128.100000 12.020000 128.170000 ;
      RECT -0.145000 128.170000 11.950000 128.240000 ;
      RECT -0.145000 128.170000 11.950000 128.240000 ;
      RECT -0.145000 128.240000 11.930000 128.260000 ;
      RECT -0.145000 128.240000 11.930000 128.260000 ;
      RECT -0.145000 128.260000 11.860000 128.330000 ;
      RECT -0.145000 128.260000 11.860000 128.330000 ;
      RECT -0.145000 128.330000 11.790000 128.400000 ;
      RECT -0.145000 128.330000 11.790000 128.400000 ;
      RECT -0.145000 128.400000 11.720000 128.470000 ;
      RECT -0.145000 128.400000 11.720000 128.470000 ;
      RECT -0.145000 128.470000 11.650000 128.540000 ;
      RECT -0.145000 128.470000 11.650000 128.540000 ;
      RECT -0.145000 128.540000 11.580000 128.610000 ;
      RECT -0.145000 128.540000 11.580000 128.610000 ;
      RECT -0.145000 128.610000 11.510000 128.680000 ;
      RECT -0.145000 128.610000 11.510000 128.680000 ;
      RECT -0.145000 128.680000 11.440000 128.750000 ;
      RECT -0.145000 128.680000 11.440000 128.750000 ;
      RECT -0.145000 128.750000 11.370000 128.820000 ;
      RECT -0.145000 128.750000 11.370000 128.820000 ;
      RECT -0.145000 128.820000 11.300000 128.890000 ;
      RECT -0.145000 128.820000 11.300000 128.890000 ;
      RECT -0.145000 128.890000 11.230000 128.960000 ;
      RECT -0.145000 128.890000 11.230000 128.960000 ;
      RECT -0.145000 128.960000 11.160000 129.030000 ;
      RECT -0.145000 128.960000 11.160000 129.030000 ;
      RECT -0.145000 129.030000 11.090000 129.100000 ;
      RECT -0.145000 129.030000 11.090000 129.100000 ;
      RECT -0.145000 129.100000 11.020000 129.170000 ;
      RECT -0.145000 129.100000 11.020000 129.170000 ;
      RECT -0.145000 129.170000 10.950000 129.240000 ;
      RECT -0.145000 129.170000 10.950000 129.240000 ;
      RECT -0.145000 129.240000 10.880000 129.310000 ;
      RECT -0.145000 129.240000 10.880000 129.310000 ;
      RECT -0.145000 129.310000 10.810000 129.380000 ;
      RECT -0.145000 129.310000 10.810000 129.380000 ;
      RECT -0.145000 129.380000 10.740000 129.450000 ;
      RECT -0.145000 129.380000 10.740000 129.450000 ;
      RECT -0.145000 129.450000 10.670000 129.520000 ;
      RECT -0.145000 129.450000 10.670000 129.520000 ;
      RECT -0.145000 129.520000 10.600000 129.590000 ;
      RECT -0.145000 129.520000 10.600000 129.590000 ;
      RECT -0.145000 129.590000 10.530000 129.660000 ;
      RECT -0.145000 129.590000 10.530000 129.660000 ;
      RECT -0.145000 129.660000 10.460000 129.730000 ;
      RECT -0.145000 129.660000 10.460000 129.730000 ;
      RECT -0.145000 129.730000 10.390000 129.800000 ;
      RECT -0.145000 129.730000 10.390000 129.800000 ;
      RECT -0.145000 129.800000 10.320000 129.870000 ;
      RECT -0.145000 129.800000 10.320000 129.870000 ;
      RECT -0.145000 129.870000 10.250000 129.940000 ;
      RECT -0.145000 129.870000 10.250000 129.940000 ;
      RECT -0.145000 129.940000 10.180000 130.010000 ;
      RECT -0.145000 129.940000 10.180000 130.010000 ;
      RECT -0.145000 130.010000 10.110000 130.080000 ;
      RECT -0.145000 130.010000 10.110000 130.080000 ;
      RECT -0.145000 130.080000 10.040000 130.150000 ;
      RECT -0.145000 130.080000 10.040000 130.150000 ;
      RECT -0.145000 130.150000  9.970000 130.220000 ;
      RECT -0.145000 130.150000  9.970000 130.220000 ;
      RECT -0.145000 131.275000  0.940000 131.345000 ;
      RECT -0.145000 131.275000  0.940000 131.345000 ;
      RECT -0.145000 131.345000  1.010000 131.415000 ;
      RECT -0.145000 131.345000  1.010000 131.415000 ;
      RECT -0.145000 131.415000  1.080000 131.485000 ;
      RECT -0.145000 131.415000  1.080000 131.485000 ;
      RECT -0.145000 131.485000  1.150000 131.555000 ;
      RECT -0.145000 131.485000  1.150000 131.555000 ;
      RECT -0.145000 131.555000  1.220000 131.625000 ;
      RECT -0.145000 131.555000  1.220000 131.625000 ;
      RECT -0.145000 131.625000  1.290000 131.695000 ;
      RECT -0.145000 131.625000  1.290000 131.695000 ;
      RECT -0.145000 131.695000  1.360000 131.765000 ;
      RECT -0.145000 131.695000  1.360000 131.765000 ;
      RECT -0.145000 131.765000  1.430000 131.835000 ;
      RECT -0.145000 131.765000  1.430000 131.835000 ;
      RECT -0.145000 131.835000  1.500000 131.905000 ;
      RECT -0.145000 131.835000  1.500000 131.905000 ;
      RECT -0.145000 131.905000  1.570000 131.975000 ;
      RECT -0.145000 131.905000  1.570000 131.975000 ;
      RECT -0.145000 131.975000  1.640000 132.045000 ;
      RECT -0.145000 131.975000  1.640000 132.045000 ;
      RECT -0.145000 132.045000  1.710000 132.115000 ;
      RECT -0.145000 132.045000  1.710000 132.115000 ;
      RECT -0.145000 132.115000  1.780000 132.185000 ;
      RECT -0.145000 132.115000  1.780000 132.185000 ;
      RECT -0.145000 132.185000  1.850000 132.255000 ;
      RECT -0.145000 132.185000  1.850000 132.255000 ;
      RECT -0.145000 132.255000  1.920000 132.325000 ;
      RECT -0.145000 132.255000  1.920000 132.325000 ;
      RECT -0.145000 132.325000  1.990000 132.395000 ;
      RECT -0.145000 132.325000  1.990000 132.395000 ;
      RECT -0.145000 132.395000  2.060000 132.465000 ;
      RECT -0.145000 132.395000  2.060000 132.465000 ;
      RECT -0.145000 132.465000  2.130000 132.535000 ;
      RECT -0.145000 132.465000  2.130000 132.535000 ;
      RECT -0.145000 132.535000  2.200000 132.605000 ;
      RECT -0.145000 132.535000  2.200000 132.605000 ;
      RECT -0.145000 132.605000  2.270000 132.675000 ;
      RECT -0.145000 132.605000  2.270000 132.675000 ;
      RECT -0.145000 132.675000  2.340000 132.740000 ;
      RECT -0.145000 132.675000  2.340000 132.740000 ;
      RECT -0.145000 132.740000  2.405000 132.810000 ;
      RECT -0.145000 132.740000  2.405000 132.810000 ;
      RECT -0.145000 132.810000  2.475000 132.880000 ;
      RECT -0.145000 132.810000  2.475000 132.880000 ;
      RECT -0.145000 132.880000  2.545000 132.950000 ;
      RECT -0.145000 132.880000  2.545000 132.950000 ;
      RECT -0.145000 132.950000  2.615000 133.020000 ;
      RECT -0.145000 132.950000  2.615000 133.020000 ;
      RECT -0.145000 133.020000  2.685000 133.090000 ;
      RECT -0.145000 133.020000  2.685000 133.090000 ;
      RECT -0.145000 133.090000  2.755000 133.160000 ;
      RECT -0.145000 133.090000  2.755000 133.160000 ;
      RECT -0.145000 133.160000  2.825000 133.230000 ;
      RECT -0.145000 133.160000  2.825000 133.230000 ;
      RECT -0.145000 133.230000  2.895000 133.300000 ;
      RECT -0.145000 133.230000  2.895000 133.300000 ;
      RECT -0.145000 133.300000  2.965000 133.370000 ;
      RECT -0.145000 133.300000  2.965000 133.370000 ;
      RECT -0.145000 133.370000  3.035000 133.440000 ;
      RECT -0.145000 133.370000  3.035000 133.440000 ;
      RECT -0.145000 133.440000  3.105000 133.510000 ;
      RECT -0.145000 133.440000  3.105000 133.510000 ;
      RECT -0.145000 133.510000  3.175000 133.580000 ;
      RECT -0.145000 133.510000  3.175000 133.580000 ;
      RECT -0.145000 133.580000  3.245000 133.650000 ;
      RECT -0.145000 133.580000  3.245000 133.650000 ;
      RECT -0.145000 133.650000  3.315000 133.720000 ;
      RECT -0.145000 133.650000  3.315000 133.720000 ;
      RECT -0.145000 133.720000  3.385000 133.790000 ;
      RECT -0.145000 133.720000  3.385000 133.790000 ;
      RECT -0.145000 133.790000  3.455000 133.860000 ;
      RECT -0.145000 133.790000  3.455000 133.860000 ;
      RECT -0.145000 133.860000  3.525000 133.930000 ;
      RECT -0.145000 133.860000  3.525000 133.930000 ;
      RECT -0.145000 133.930000  3.595000 134.000000 ;
      RECT -0.145000 133.930000  3.595000 134.000000 ;
      RECT -0.145000 134.000000  3.665000 134.070000 ;
      RECT -0.145000 134.000000  3.665000 134.070000 ;
      RECT -0.145000 134.070000  3.735000 134.140000 ;
      RECT -0.145000 134.070000  3.735000 134.140000 ;
      RECT -0.145000 134.140000  3.805000 134.180000 ;
      RECT -0.145000 134.140000  3.805000 134.180000 ;
      RECT -0.145000 134.180000  3.775000 134.250000 ;
      RECT -0.145000 134.180000  3.775000 134.250000 ;
      RECT -0.145000 134.250000  3.700000 134.320000 ;
      RECT -0.145000 134.250000  3.700000 134.320000 ;
      RECT -0.145000 134.320000  3.635000 134.390000 ;
      RECT -0.145000 134.320000  3.635000 134.390000 ;
      RECT -0.145000 134.390000  3.560000 134.460000 ;
      RECT -0.145000 134.390000  3.560000 134.460000 ;
      RECT -0.145000 134.460000  3.490000 134.530000 ;
      RECT -0.145000 134.460000  3.490000 134.530000 ;
      RECT -0.145000 134.530000  3.420000 134.600000 ;
      RECT -0.145000 134.530000  3.420000 134.600000 ;
      RECT -0.145000 134.600000  3.350000 134.670000 ;
      RECT -0.145000 134.600000  3.350000 134.670000 ;
      RECT -0.145000 134.670000  3.280000 134.740000 ;
      RECT -0.145000 134.670000  3.280000 134.740000 ;
      RECT -0.145000 134.740000  3.210000 134.810000 ;
      RECT -0.145000 134.740000  3.210000 134.810000 ;
      RECT -0.145000 134.810000  3.140000 134.880000 ;
      RECT -0.145000 134.810000  3.140000 134.880000 ;
      RECT -0.145000 134.880000  3.070000 134.950000 ;
      RECT -0.145000 134.880000  3.070000 134.950000 ;
      RECT -0.145000 134.950000  3.000000 135.020000 ;
      RECT -0.145000 134.950000  3.000000 135.020000 ;
      RECT -0.145000 135.020000  2.930000 135.090000 ;
      RECT -0.145000 135.020000  2.930000 135.090000 ;
      RECT -0.145000 135.090000  2.860000 135.160000 ;
      RECT -0.145000 135.090000  2.860000 135.160000 ;
      RECT -0.145000 135.160000  2.790000 135.230000 ;
      RECT -0.145000 135.160000  2.790000 135.230000 ;
      RECT -0.145000 135.230000  2.720000 135.300000 ;
      RECT -0.145000 135.230000  2.720000 135.300000 ;
      RECT -0.145000 135.300000  2.650000 135.370000 ;
      RECT -0.145000 135.300000  2.650000 135.370000 ;
      RECT -0.145000 135.370000  2.580000 135.440000 ;
      RECT -0.145000 135.370000  2.580000 135.440000 ;
      RECT -0.145000 135.440000  2.550000 135.470000 ;
      RECT -0.145000 135.440000  2.550000 135.470000 ;
      RECT -0.145000 135.470000  2.480000 135.540000 ;
      RECT -0.145000 135.470000  2.480000 135.540000 ;
      RECT -0.145000 135.540000  2.410000 135.610000 ;
      RECT -0.145000 135.540000  2.410000 135.610000 ;
      RECT -0.145000 135.610000  2.340000 135.680000 ;
      RECT -0.145000 135.610000  2.340000 135.680000 ;
      RECT -0.145000 135.680000  2.270000 135.750000 ;
      RECT -0.145000 135.680000  2.270000 135.750000 ;
      RECT -0.145000 135.750000  2.200000 135.820000 ;
      RECT -0.145000 135.750000  2.200000 135.820000 ;
      RECT -0.145000 135.820000  2.130000 135.890000 ;
      RECT -0.145000 135.820000  2.130000 135.890000 ;
      RECT -0.145000 135.890000  2.060000 135.960000 ;
      RECT -0.145000 135.890000  2.060000 135.960000 ;
      RECT -0.145000 135.960000  1.990000 136.030000 ;
      RECT -0.145000 135.960000  1.990000 136.030000 ;
      RECT -0.145000 136.030000  1.920000 136.100000 ;
      RECT -0.145000 136.030000  1.920000 136.100000 ;
      RECT -0.145000 136.100000  1.850000 136.170000 ;
      RECT -0.145000 136.100000  1.850000 136.170000 ;
      RECT -0.145000 136.170000  1.780000 136.240000 ;
      RECT -0.145000 136.170000  1.780000 136.240000 ;
      RECT -0.145000 136.240000  1.710000 136.310000 ;
      RECT -0.145000 136.240000  1.710000 136.310000 ;
      RECT -0.145000 136.310000  1.640000 136.380000 ;
      RECT -0.145000 136.310000  1.640000 136.380000 ;
      RECT -0.145000 136.380000  1.570000 136.450000 ;
      RECT -0.145000 136.380000  1.570000 136.450000 ;
      RECT -0.145000 136.450000  1.495000 136.520000 ;
      RECT -0.145000 136.450000  1.495000 136.520000 ;
      RECT -0.145000 136.520000  1.425000 136.590000 ;
      RECT -0.145000 136.520000  1.425000 136.590000 ;
      RECT -0.145000 136.590000  1.355000 136.660000 ;
      RECT -0.145000 136.590000  1.355000 136.660000 ;
      RECT -0.145000 136.660000  1.285000 136.730000 ;
      RECT -0.145000 136.660000  1.285000 136.730000 ;
      RECT -0.145000 136.730000  1.215000 136.800000 ;
      RECT -0.145000 136.730000  1.215000 136.800000 ;
      RECT -0.145000 136.800000  1.145000 136.870000 ;
      RECT -0.145000 136.800000  1.145000 136.870000 ;
      RECT -0.145000 136.870000  1.075000 136.940000 ;
      RECT -0.145000 136.870000  1.075000 136.940000 ;
      RECT -0.145000 136.940000  1.005000 137.010000 ;
      RECT -0.145000 136.940000  1.005000 137.010000 ;
      RECT -0.145000 137.010000  0.935000 137.080000 ;
      RECT -0.145000 137.010000  0.935000 137.080000 ;
      RECT -0.145000 137.080000  0.865000 137.150000 ;
      RECT -0.145000 137.080000  0.865000 137.150000 ;
      RECT -0.145000 137.150000  0.795000 137.220000 ;
      RECT -0.145000 137.150000  0.795000 137.220000 ;
      RECT -0.145000 137.220000  0.725000 137.290000 ;
      RECT -0.145000 137.220000  0.725000 137.290000 ;
      RECT -0.145000 137.290000  0.655000 137.360000 ;
      RECT -0.145000 137.290000  0.655000 137.360000 ;
      RECT -0.145000 137.360000  0.585000 137.430000 ;
      RECT -0.145000 137.360000  0.585000 137.430000 ;
      RECT -0.145000 137.430000  0.515000 137.500000 ;
      RECT -0.145000 137.430000  0.515000 137.500000 ;
      RECT -0.145000 137.500000  0.445000 137.570000 ;
      RECT -0.145000 137.500000  0.445000 137.570000 ;
      RECT -0.145000 137.570000  0.375000 137.640000 ;
      RECT -0.145000 137.570000  0.375000 137.640000 ;
      RECT -0.145000 137.640000  0.305000 137.710000 ;
      RECT -0.145000 137.640000  0.305000 137.710000 ;
      RECT -0.145000 137.710000  0.235000 137.780000 ;
      RECT -0.145000 137.710000  0.235000 137.780000 ;
      RECT -0.145000 137.780000  0.165000 137.850000 ;
      RECT -0.145000 137.780000  0.165000 137.850000 ;
      RECT -0.145000 137.850000  0.095000 137.920000 ;
      RECT -0.145000 137.850000  0.095000 137.920000 ;
      RECT -0.145000 137.920000  0.025000 137.990000 ;
      RECT -0.145000 137.920000  0.025000 137.990000 ;
      RECT -0.145000 137.990000 -0.045000 138.060000 ;
      RECT -0.145000 137.990000 -0.045000 138.060000 ;
      RECT -0.145000 138.060000 -0.115000 138.130000 ;
      RECT -0.145000 138.060000 -0.115000 138.130000 ;
      RECT -0.145000 138.160000  0.940000 139.015000 ;
      RECT -0.145000 139.015000  0.940000 139.085000 ;
      RECT -0.145000 139.085000  1.010000 139.155000 ;
      RECT -0.145000 139.155000  1.080000 139.225000 ;
      RECT -0.145000 139.225000  1.150000 139.295000 ;
      RECT -0.145000 139.295000  1.220000 139.365000 ;
      RECT -0.145000 139.365000  1.290000 139.435000 ;
      RECT -0.145000 139.435000  1.360000 139.505000 ;
      RECT -0.145000 139.505000 11.105000 139.540000 ;
      RECT -0.145000 139.540000 11.140000 139.575000 ;
      RECT -0.145000 139.575000 69.715000 139.645000 ;
      RECT -0.145000 139.645000 69.785000 139.715000 ;
      RECT -0.145000 139.715000 69.855000 139.785000 ;
      RECT -0.145000 139.785000 69.925000 139.850000 ;
      RECT -0.145000 139.850000  1.385000 139.920000 ;
      RECT -0.145000 139.920000  1.315000 139.990000 ;
      RECT -0.145000 139.990000  1.245000 140.060000 ;
      RECT -0.145000 140.060000  1.175000 140.130000 ;
      RECT -0.145000 140.130000  1.105000 140.200000 ;
      RECT -0.145000 140.200000  1.035000 140.270000 ;
      RECT -0.145000 140.270000  0.965000 140.340000 ;
      RECT -0.145000 140.340000  0.940000 140.365000 ;
      RECT -0.145000 140.365000  0.940000 143.640000 ;
      RECT -0.145000 143.640000  0.940000 143.710000 ;
      RECT -0.145000 143.710000  1.010000 143.780000 ;
      RECT -0.145000 143.780000  1.080000 143.850000 ;
      RECT -0.145000 143.850000  1.150000 143.920000 ;
      RECT -0.145000 143.920000  1.220000 143.990000 ;
      RECT -0.145000 143.990000  1.290000 144.060000 ;
      RECT -0.145000 144.060000  1.360000 144.130000 ;
      RECT -0.145000 144.130000  1.430000 144.200000 ;
      RECT -0.145000 144.200000  1.500000 144.270000 ;
      RECT -0.145000 144.270000  1.570000 144.340000 ;
      RECT -0.145000 144.340000  1.640000 144.410000 ;
      RECT -0.145000 144.410000  1.710000 144.480000 ;
      RECT -0.145000 144.480000  1.780000 144.550000 ;
      RECT -0.145000 144.550000  1.850000 144.620000 ;
      RECT -0.145000 144.620000  1.920000 144.690000 ;
      RECT -0.145000 144.690000  1.990000 144.760000 ;
      RECT -0.145000 144.760000  2.060000 144.830000 ;
      RECT -0.145000 144.830000  2.130000 144.900000 ;
      RECT -0.145000 144.900000  2.200000 144.970000 ;
      RECT -0.145000 144.970000  2.270000 145.040000 ;
      RECT -0.145000 145.040000  2.340000 145.110000 ;
      RECT -0.145000 145.110000  2.410000 145.130000 ;
      RECT -0.125000  96.525000  3.310000  96.545000 ;
      RECT -0.125000  96.525000  3.310000  96.545000 ;
      RECT -0.115000 138.130000  0.940000 138.160000 ;
      RECT -0.055000  96.455000  3.240000  96.525000 ;
      RECT -0.055000  96.455000  3.240000  96.525000 ;
      RECT -0.045000 138.060000  0.940000 138.130000 ;
      RECT  0.000000   0.000000  0.705000  84.590000 ;
      RECT  0.000000   0.000000 12.145000   6.435000 ;
      RECT  0.000000   6.435000 11.775000   6.805000 ;
      RECT  0.000000   6.805000 12.230000   6.980000 ;
      RECT  0.000000   6.980000 12.555000   7.310000 ;
      RECT  0.000000   7.310000 12.555000  10.370000 ;
      RECT  0.000000  10.370000 12.660000  10.445000 ;
      RECT  0.000000  10.445000 14.415000  12.400000 ;
      RECT  0.000000  12.400000 18.075000  16.060000 ;
      RECT  0.000000  16.060000 24.085000  18.665000 ;
      RECT  0.000000  18.665000 24.085000  25.415000 ;
      RECT  0.000000  25.415000 24.675000  26.005000 ;
      RECT  0.000000  26.005000 24.675000  42.680000 ;
      RECT  0.000000  42.680000 24.210000  43.145000 ;
      RECT  0.000000  43.145000  5.925000  43.685000 ;
      RECT  0.000000  43.685000 75.000000 200.000000 ;
      RECT  0.000000  84.590000  0.705000  84.660000 ;
      RECT  0.000000  84.660000  0.775000  84.730000 ;
      RECT  0.000000  84.730000  0.845000  84.800000 ;
      RECT  0.000000  84.800000  0.915000  84.825000 ;
      RECT  0.000000  84.825000  0.940000  95.065000 ;
      RECT  0.000000  95.065000  0.870000  95.135000 ;
      RECT  0.000000  95.135000  0.800000  95.205000 ;
      RECT  0.000000  95.205000  0.730000  95.275000 ;
      RECT  0.000000  95.275000  0.660000  95.345000 ;
      RECT  0.000000  95.345000  0.590000  95.415000 ;
      RECT  0.000000  95.415000  0.520000  95.485000 ;
      RECT  0.000000  95.485000  0.450000  95.555000 ;
      RECT  0.000000  95.555000  0.390000  95.615000 ;
      RECT  0.000000 101.700000 73.490000 104.845000 ;
      RECT  0.000000 104.845000 74.035000 125.160000 ;
      RECT  0.000000 130.500000 10.015000 130.570000 ;
      RECT  0.000000 130.570000  9.945000 130.640000 ;
      RECT  0.000000 130.640000  9.875000 130.710000 ;
      RECT  0.000000 130.710000  9.805000 130.780000 ;
      RECT  0.000000 130.780000  9.735000 130.850000 ;
      RECT  0.000000 130.850000  9.665000 130.920000 ;
      RECT  0.000000 130.920000  9.595000 130.990000 ;
      RECT  0.000000 130.990000  9.590000 130.995000 ;
      RECT  0.000000 145.410000  2.595000 146.420000 ;
      RECT  0.000000 146.420000 59.500000 199.490000 ;
      RECT  0.000000 146.420000 70.525000 146.425000 ;
      RECT  0.000000 146.420000 70.525000 195.970000 ;
      RECT  0.000000 146.425000 73.405000 195.970000 ;
      RECT  0.000000 146.425000 75.000000 174.220000 ;
      RECT  0.000000 174.220000 73.405000 175.420000 ;
      RECT  0.000000 175.420000 75.000000 195.970000 ;
      RECT  0.000000 195.970000 59.500000 199.490000 ;
      RECT  0.000000 199.490000 59.500000 200.000000 ;
      RECT  0.015000  96.385000  3.170000  96.455000 ;
      RECT  0.015000  96.385000  3.170000  96.455000 ;
      RECT  0.025000 137.990000  0.940000 138.060000 ;
      RECT  0.085000  96.315000  3.100000  96.385000 ;
      RECT  0.085000  96.315000  3.100000  96.385000 ;
      RECT  0.095000 137.920000  0.940000 137.990000 ;
      RECT  0.155000  96.245000  3.030000  96.315000 ;
      RECT  0.155000  96.245000  3.030000  96.315000 ;
      RECT  0.165000 137.850000  0.940000 137.920000 ;
      RECT  0.225000  96.175000  2.960000  96.245000 ;
      RECT  0.225000  96.175000  2.960000  96.245000 ;
      RECT  0.235000 137.780000  0.940000 137.850000 ;
      RECT  0.295000  96.105000  2.890000  96.175000 ;
      RECT  0.295000  96.105000  2.890000  96.175000 ;
      RECT  0.305000 137.710000  0.940000 137.780000 ;
      RECT  0.365000  96.035000  2.820000  96.105000 ;
      RECT  0.365000  96.035000  2.820000  96.105000 ;
      RECT  0.375000 137.640000  0.940000 137.710000 ;
      RECT  0.435000  95.965000  2.750000  96.035000 ;
      RECT  0.435000  95.965000  2.750000  96.035000 ;
      RECT  0.445000 137.570000  0.940000 137.640000 ;
      RECT  0.505000  95.895000  2.680000  95.965000 ;
      RECT  0.505000  95.895000  2.680000  95.965000 ;
      RECT  0.515000 137.500000  0.940000 137.570000 ;
      RECT  0.520000  95.880000  2.665000  95.895000 ;
      RECT  0.520000  95.880000  2.665000  95.895000 ;
      RECT  0.520000  95.880000  2.665000  95.895000 ;
      RECT  0.535000  95.865000  2.650000  95.880000 ;
      RECT  0.535000  95.865000  2.650000  95.880000 ;
      RECT  0.535000  95.865000  2.650000  95.880000 ;
      RECT  0.585000 137.430000  0.940000 137.500000 ;
      RECT  0.590000  95.810000  2.595000  95.865000 ;
      RECT  0.590000  95.810000  2.595000  95.865000 ;
      RECT  0.590000  95.810000  2.650000  95.865000 ;
      RECT  0.655000 137.360000  0.940000 137.430000 ;
      RECT  0.660000  95.740000  2.525000  95.810000 ;
      RECT  0.660000  95.740000  2.525000  95.810000 ;
      RECT  0.660000  95.740000  2.650000  95.810000 ;
      RECT  0.725000 137.290000  0.940000 137.360000 ;
      RECT  0.730000  95.670000  2.455000  95.740000 ;
      RECT  0.730000  95.670000  2.455000  95.740000 ;
      RECT  0.730000  95.670000  2.650000  95.740000 ;
      RECT  0.795000 137.220000  0.940000 137.290000 ;
      RECT  0.800000  95.600000  2.385000  95.670000 ;
      RECT  0.800000  95.600000  2.385000  95.670000 ;
      RECT  0.800000  95.600000  2.650000  95.670000 ;
      RECT  0.865000 137.150000  0.940000 137.220000 ;
      RECT  0.870000  95.530000  2.315000  95.600000 ;
      RECT  0.870000  95.530000  2.315000  95.600000 ;
      RECT  0.870000  95.530000  2.650000  95.600000 ;
      RECT  0.935000 137.080000  0.940000 137.150000 ;
      RECT  0.940000  95.460000  2.650000  95.530000 ;
      RECT  0.945000  95.460000  2.245000  95.530000 ;
      RECT  0.945000  95.460000  2.245000  95.530000 ;
      RECT  0.985000   0.240000 11.975000   0.590000 ;
      RECT  0.985000   0.590000  3.300000   0.660000 ;
      RECT  0.985000   0.660000  3.230000   0.730000 ;
      RECT  0.985000   0.730000  3.160000   0.800000 ;
      RECT  0.985000   0.800000  3.090000   0.870000 ;
      RECT  0.985000   0.870000  3.020000   0.940000 ;
      RECT  0.985000   0.940000  2.950000   1.010000 ;
      RECT  0.985000   1.010000  2.880000   1.080000 ;
      RECT  0.985000   1.080000  2.810000   1.150000 ;
      RECT  0.985000   1.150000  2.740000   1.220000 ;
      RECT  0.985000   1.220000  2.670000   1.290000 ;
      RECT  0.985000   1.290000  2.600000   1.360000 ;
      RECT  0.985000   1.360000  2.530000   1.430000 ;
      RECT  0.985000   1.430000  2.460000   1.500000 ;
      RECT  0.985000   1.500000  2.415000   1.545000 ;
      RECT  0.985000   1.545000  2.415000   3.150000 ;
      RECT  0.985000   3.150000  2.415000   3.220000 ;
      RECT  0.985000   3.220000  2.485000   3.290000 ;
      RECT  0.985000   3.290000  2.555000   3.360000 ;
      RECT  0.985000   3.360000  2.625000   3.430000 ;
      RECT  0.985000   3.430000  2.695000   3.500000 ;
      RECT  0.985000   3.500000  2.765000   3.570000 ;
      RECT  0.985000   3.570000  2.835000   3.640000 ;
      RECT  0.985000   3.640000  2.905000   3.710000 ;
      RECT  0.985000   3.710000  2.975000   3.780000 ;
      RECT  0.985000   3.780000  3.045000   3.850000 ;
      RECT  0.985000   3.850000  3.115000   3.920000 ;
      RECT  0.985000   3.920000  3.185000   3.990000 ;
      RECT  0.985000   3.990000  3.255000   4.060000 ;
      RECT  0.985000   4.060000  3.325000   4.105000 ;
      RECT  0.985000   4.105000  4.515000  71.340000 ;
      RECT  0.985000  71.910000 19.260000  79.760000 ;
      RECT  0.985000  80.435000 30.155000  84.475000 ;
      RECT  1.010000  95.390000  2.175000  95.460000 ;
      RECT  1.010000  95.390000  2.175000  95.460000 ;
      RECT  1.010000  95.390000  2.650000  95.460000 ;
      RECT  1.055000  84.475000  3.865000  84.545000 ;
      RECT  1.055000  84.475000  3.865000  84.545000 ;
      RECT  1.080000  95.320000  2.650000  95.390000 ;
      RECT  1.085000  95.320000  2.105000  95.390000 ;
      RECT  1.085000  95.320000  2.105000  95.390000 ;
      RECT  1.125000  84.545000  3.795000  84.615000 ;
      RECT  1.125000  84.545000  3.795000  84.615000 ;
      RECT  1.125000 130.995000 72.380000 131.065000 ;
      RECT  1.150000  95.250000  2.650000  95.320000 ;
      RECT  1.155000  95.250000  2.035000  95.320000 ;
      RECT  1.155000  95.250000  2.035000  95.320000 ;
      RECT  1.195000  84.615000  3.725000  84.685000 ;
      RECT  1.195000  84.615000  3.725000  84.685000 ;
      RECT  1.195000 131.065000 72.380000 131.135000 ;
      RECT  1.220000  81.705000  2.650000  85.760000 ;
      RECT  1.220000  84.685000  3.700000  84.710000 ;
      RECT  1.220000  84.685000  3.700000  84.710000 ;
      RECT  1.220000  84.710000  3.630000  84.780000 ;
      RECT  1.220000  84.780000  3.560000  84.850000 ;
      RECT  1.220000  84.850000  3.490000  84.920000 ;
      RECT  1.220000  84.920000  3.420000  84.990000 ;
      RECT  1.220000  84.990000  3.350000  85.060000 ;
      RECT  1.220000  85.060000  3.280000  85.130000 ;
      RECT  1.220000  85.130000  3.210000  85.200000 ;
      RECT  1.220000  85.200000  3.140000  85.270000 ;
      RECT  1.220000  85.270000  3.070000  85.340000 ;
      RECT  1.220000  85.340000  3.000000  85.410000 ;
      RECT  1.220000  85.410000  2.930000  85.480000 ;
      RECT  1.220000  85.480000  2.860000  85.550000 ;
      RECT  1.220000  85.550000  2.790000  85.620000 ;
      RECT  1.220000  85.620000  2.720000  85.690000 ;
      RECT  1.220000  85.690000  2.650000  85.760000 ;
      RECT  1.220000  85.760000  2.580000  85.830000 ;
      RECT  1.220000  85.760000  2.580000  85.830000 ;
      RECT  1.220000  85.830000  2.510000  85.900000 ;
      RECT  1.220000  85.830000  2.510000  85.900000 ;
      RECT  1.220000  85.900000  2.440000  85.970000 ;
      RECT  1.220000  85.900000  2.440000  85.970000 ;
      RECT  1.220000  85.970000  2.370000  86.040000 ;
      RECT  1.220000  85.970000  2.370000  86.040000 ;
      RECT  1.220000  86.040000  2.300000  86.110000 ;
      RECT  1.220000  86.040000  2.300000  86.110000 ;
      RECT  1.220000  86.110000  2.230000  86.180000 ;
      RECT  1.220000  86.110000  2.230000  86.180000 ;
      RECT  1.220000  86.180000  2.160000  86.250000 ;
      RECT  1.220000  86.180000  2.160000  86.250000 ;
      RECT  1.220000  86.250000  2.090000  86.320000 ;
      RECT  1.220000  86.250000  2.090000  86.320000 ;
      RECT  1.220000  86.320000  2.020000  86.390000 ;
      RECT  1.220000  86.320000  2.020000  86.390000 ;
      RECT  1.220000  86.390000  1.950000  86.460000 ;
      RECT  1.220000  86.390000  1.950000  86.460000 ;
      RECT  1.220000  86.460000  1.880000  86.530000 ;
      RECT  1.220000  86.460000  1.880000  86.530000 ;
      RECT  1.220000  86.530000  1.810000  86.600000 ;
      RECT  1.220000  86.530000  1.810000  86.600000 ;
      RECT  1.220000  86.600000  1.740000  86.670000 ;
      RECT  1.220000  86.600000  1.740000  86.670000 ;
      RECT  1.220000  86.670000  1.670000  86.740000 ;
      RECT  1.220000  86.670000  1.670000  86.740000 ;
      RECT  1.220000  86.740000  1.600000  86.810000 ;
      RECT  1.220000  86.740000  1.600000  86.810000 ;
      RECT  1.220000  86.810000  1.530000  86.880000 ;
      RECT  1.220000  86.810000  1.530000  86.880000 ;
      RECT  1.220000  86.880000  1.460000  86.950000 ;
      RECT  1.220000  86.880000  1.460000  86.950000 ;
      RECT  1.220000  86.950000  1.390000  87.020000 ;
      RECT  1.220000  86.950000  1.390000  87.020000 ;
      RECT  1.220000  87.020000  1.320000  87.090000 ;
      RECT  1.220000  87.020000  1.320000  87.090000 ;
      RECT  1.220000  87.090000  1.250000  87.160000 ;
      RECT  1.220000  87.090000  1.250000  87.160000 ;
      RECT  1.220000  87.190000  2.650000  94.810000 ;
      RECT  1.220000  94.810000  1.525000  94.880000 ;
      RECT  1.220000  94.880000  1.455000  94.950000 ;
      RECT  1.220000  94.950000  1.385000  95.020000 ;
      RECT  1.220000  95.020000  1.315000  95.090000 ;
      RECT  1.220000  95.090000  1.245000  95.160000 ;
      RECT  1.220000  95.160000  1.225000  95.180000 ;
      RECT  1.220000  95.180000  2.650000  95.250000 ;
      RECT  1.220000 135.750000 14.920000 139.225000 ;
      RECT  1.220000 137.195000 70.400000 137.265000 ;
      RECT  1.220000 137.195000 70.400000 137.265000 ;
      RECT  1.220000 137.265000 70.330000 137.335000 ;
      RECT  1.220000 137.265000 70.330000 137.335000 ;
      RECT  1.220000 137.335000 70.260000 137.405000 ;
      RECT  1.220000 137.335000 70.260000 137.405000 ;
      RECT  1.220000 137.405000 70.190000 137.475000 ;
      RECT  1.220000 137.405000 70.190000 137.475000 ;
      RECT  1.220000 137.475000 70.120000 137.545000 ;
      RECT  1.220000 137.475000 70.120000 137.545000 ;
      RECT  1.220000 137.545000 70.050000 137.615000 ;
      RECT  1.220000 137.545000 70.050000 137.615000 ;
      RECT  1.220000 137.615000 69.980000 137.685000 ;
      RECT  1.220000 137.615000 69.980000 137.685000 ;
      RECT  1.220000 137.685000 69.910000 137.755000 ;
      RECT  1.220000 137.685000 69.910000 137.755000 ;
      RECT  1.220000 137.755000 69.840000 137.825000 ;
      RECT  1.220000 137.755000 69.840000 137.825000 ;
      RECT  1.220000 137.825000 69.770000 137.895000 ;
      RECT  1.220000 137.825000 69.770000 137.895000 ;
      RECT  1.220000 137.895000 69.700000 137.965000 ;
      RECT  1.220000 137.895000 69.700000 137.965000 ;
      RECT  1.220000 137.965000 69.630000 138.035000 ;
      RECT  1.220000 137.965000 69.630000 138.035000 ;
      RECT  1.220000 138.035000 69.560000 138.105000 ;
      RECT  1.220000 138.035000 69.560000 138.105000 ;
      RECT  1.220000 138.105000 69.490000 138.175000 ;
      RECT  1.220000 138.105000 69.490000 138.175000 ;
      RECT  1.220000 138.175000 69.420000 138.245000 ;
      RECT  1.220000 138.175000 69.420000 138.245000 ;
      RECT  1.220000 138.245000 69.350000 138.315000 ;
      RECT  1.220000 138.245000 69.350000 138.315000 ;
      RECT  1.220000 138.315000 69.280000 138.385000 ;
      RECT  1.220000 138.315000 69.280000 138.385000 ;
      RECT  1.220000 138.385000 69.210000 138.455000 ;
      RECT  1.220000 138.385000 69.210000 138.455000 ;
      RECT  1.220000 138.455000 69.140000 138.525000 ;
      RECT  1.220000 138.455000 69.140000 138.525000 ;
      RECT  1.220000 138.525000 69.070000 138.595000 ;
      RECT  1.220000 138.525000 69.070000 138.595000 ;
      RECT  1.220000 138.595000 69.000000 138.665000 ;
      RECT  1.220000 138.595000 69.000000 138.665000 ;
      RECT  1.220000 138.665000 16.790000 138.685000 ;
      RECT  1.220000 138.665000 16.790000 138.685000 ;
      RECT  1.220000 138.685000 16.770000 138.705000 ;
      RECT  1.220000 138.685000 16.770000 138.705000 ;
      RECT  1.220000 138.705000 16.765000 138.710000 ;
      RECT  1.220000 138.705000 16.765000 138.710000 ;
      RECT  1.220000 138.710000 14.920000 138.900000 ;
      RECT  1.220000 140.480000 70.225000 140.550000 ;
      RECT  1.220000 140.550000 70.295000 140.620000 ;
      RECT  1.220000 140.620000 70.365000 140.690000 ;
      RECT  1.220000 140.690000 70.435000 140.760000 ;
      RECT  1.220000 140.760000 70.505000 140.780000 ;
      RECT  1.220000 140.780000 70.525000 141.095000 ;
      RECT  1.225000  95.180000  1.965000  95.250000 ;
      RECT  1.225000  95.180000  1.965000  95.250000 ;
      RECT  1.245000  95.160000  1.945000  95.180000 ;
      RECT  1.245000  95.160000  1.945000  95.180000 ;
      RECT  1.265000 131.135000 72.380000 131.205000 ;
      RECT  1.265000 137.150000 70.470000 137.195000 ;
      RECT  1.265000 137.150000 70.470000 137.195000 ;
      RECT  1.290000 138.900000 14.920000 138.970000 ;
      RECT  1.290000 138.900000 14.920000 138.970000 ;
      RECT  1.290000 140.410000 70.155000 140.480000 ;
      RECT  1.315000  95.090000  1.875000  95.160000 ;
      RECT  1.315000  95.090000  1.875000  95.160000 ;
      RECT  1.335000 131.205000 72.380000 131.275000 ;
      RECT  1.335000 137.080000 70.515000 137.150000 ;
      RECT  1.335000 137.080000 70.515000 137.150000 ;
      RECT  1.340000 141.375000 69.645000 143.595000 ;
      RECT  1.360000 138.970000 14.920000 139.040000 ;
      RECT  1.360000 138.970000 14.920000 139.040000 ;
      RECT  1.360000 140.340000 70.085000 140.410000 ;
      RECT  1.385000  95.020000  1.805000  95.090000 ;
      RECT  1.385000  95.020000  1.805000  95.090000 ;
      RECT  1.405000 131.275000 72.380000 131.345000 ;
      RECT  1.405000 137.010000 70.585000 137.080000 ;
      RECT  1.405000 137.010000 70.585000 137.080000 ;
      RECT  1.430000 139.040000 14.920000 139.110000 ;
      RECT  1.430000 139.040000 14.920000 139.110000 ;
      RECT  1.430000 140.270000 70.015000 140.340000 ;
      RECT  1.455000  94.950000  1.735000  95.020000 ;
      RECT  1.455000  94.950000  1.735000  95.020000 ;
      RECT  1.475000 131.345000 72.380000 131.415000 ;
      RECT  1.475000 136.940000 70.655000 137.010000 ;
      RECT  1.475000 136.940000 70.655000 137.010000 ;
      RECT  1.500000 139.110000 14.920000 139.180000 ;
      RECT  1.500000 139.110000 14.920000 139.180000 ;
      RECT  1.500000 140.200000 69.945000 140.270000 ;
      RECT  1.525000  94.880000  1.665000  94.950000 ;
      RECT  1.525000  94.880000  1.665000  94.950000 ;
      RECT  1.545000 131.415000 72.380000 131.485000 ;
      RECT  1.545000 136.870000 70.725000 136.940000 ;
      RECT  1.545000 136.870000 70.725000 136.940000 ;
      RECT  1.545000 139.180000 14.920000 139.225000 ;
      RECT  1.545000 139.180000 14.920000 139.225000 ;
      RECT  1.570000 140.130000 69.875000 140.200000 ;
      RECT  1.615000 131.485000 72.380000 131.555000 ;
      RECT  1.615000 136.800000 70.795000 136.870000 ;
      RECT  1.615000 136.800000 70.795000 136.870000 ;
      RECT  1.640000 143.875000 70.525000 143.945000 ;
      RECT  1.665000  94.810000  2.650000  94.880000 ;
      RECT  1.685000 131.555000 72.380000 131.625000 ;
      RECT  1.685000 136.730000 70.865000 136.800000 ;
      RECT  1.685000 136.730000 70.865000 136.800000 ;
      RECT  1.710000 143.945000 70.525000 144.015000 ;
      RECT  1.735000  94.880000  2.650000  94.950000 ;
      RECT  1.755000 131.625000 72.380000 131.695000 ;
      RECT  1.755000 136.660000 70.935000 136.730000 ;
      RECT  1.755000 136.660000 70.935000 136.730000 ;
      RECT  1.780000 144.015000 70.525000 144.085000 ;
      RECT  1.805000  94.950000  2.650000  95.020000 ;
      RECT  1.825000 131.695000 72.380000 131.765000 ;
      RECT  1.825000 136.590000 71.005000 136.660000 ;
      RECT  1.825000 136.590000 71.005000 136.660000 ;
      RECT  1.850000 144.085000 70.525000 144.155000 ;
      RECT  1.875000  95.020000  2.650000  95.090000 ;
      RECT  1.895000 131.765000 72.380000 131.835000 ;
      RECT  1.895000 136.520000 71.075000 136.590000 ;
      RECT  1.895000 136.520000 71.075000 136.590000 ;
      RECT  1.920000 144.155000 70.525000 144.225000 ;
      RECT  1.945000  95.090000  2.650000  95.160000 ;
      RECT  1.965000  95.160000  2.650000  95.180000 ;
      RECT  1.965000 131.835000 72.380000 131.905000 ;
      RECT  1.965000 136.450000 71.145000 136.520000 ;
      RECT  1.965000 136.450000 71.145000 136.520000 ;
      RECT  1.980000 144.225000 70.525000 144.285000 ;
      RECT  2.035000 131.905000 72.380000 131.975000 ;
      RECT  2.035000 136.380000 71.215000 136.450000 ;
      RECT  2.035000 136.380000 71.215000 136.450000 ;
      RECT  2.050000 144.285000 70.455000 144.355000 ;
      RECT  2.105000 131.975000 72.380000 132.045000 ;
      RECT  2.105000 136.310000 71.285000 136.380000 ;
      RECT  2.105000 136.310000 71.285000 136.380000 ;
      RECT  2.120000 144.355000 70.385000 144.425000 ;
      RECT  2.175000 132.045000 72.380000 132.115000 ;
      RECT  2.175000 136.240000 71.355000 136.310000 ;
      RECT  2.175000 136.240000 71.355000 136.310000 ;
      RECT  2.190000 144.425000 70.315000 144.495000 ;
      RECT  2.245000 132.115000 72.380000 132.185000 ;
      RECT  2.245000 136.170000 71.425000 136.240000 ;
      RECT  2.245000 136.170000 71.425000 136.240000 ;
      RECT  2.260000 144.495000 70.245000 144.565000 ;
      RECT  2.315000 132.185000 72.380000 132.255000 ;
      RECT  2.315000 136.100000 71.495000 136.170000 ;
      RECT  2.315000 136.100000 71.495000 136.170000 ;
      RECT  2.330000 144.565000 70.175000 144.635000 ;
      RECT  2.385000 132.255000 72.380000 132.325000 ;
      RECT  2.385000 136.030000 71.565000 136.100000 ;
      RECT  2.385000 136.030000 71.565000 136.100000 ;
      RECT  2.400000 144.635000 70.105000 144.705000 ;
      RECT  2.455000 132.325000 72.380000 132.395000 ;
      RECT  2.455000 135.960000 71.635000 136.030000 ;
      RECT  2.455000 135.960000 71.635000 136.030000 ;
      RECT  2.470000 144.705000 70.035000 144.775000 ;
      RECT  2.475000 132.740000 13.110000 132.810000 ;
      RECT  2.520000 132.395000 72.380000 132.460000 ;
      RECT  2.525000 135.890000 71.705000 135.960000 ;
      RECT  2.525000 135.890000 71.705000 135.960000 ;
      RECT  2.540000 144.775000 69.965000 144.845000 ;
      RECT  2.545000 132.810000 13.110000 132.880000 ;
      RECT  2.545000 144.845000 69.960000 144.850000 ;
      RECT  2.580000 135.440000 13.110000 135.470000 ;
      RECT  2.595000 135.820000 71.775000 135.890000 ;
      RECT  2.595000 135.820000 71.775000 135.890000 ;
      RECT  2.615000 132.880000 13.110000 132.950000 ;
      RECT  2.650000 135.370000 13.110000 135.440000 ;
      RECT  2.665000 135.750000 71.845000 135.820000 ;
      RECT  2.665000 135.750000 71.845000 135.820000 ;
      RECT  2.685000 132.950000 13.110000 133.020000 ;
      RECT  2.695000   1.660000  3.625000   3.035000 ;
      RECT  2.715000   1.640000  3.625000   1.660000 ;
      RECT  2.720000 135.300000 13.110000 135.370000 ;
      RECT  2.755000 133.020000 13.110000 133.090000 ;
      RECT  2.765000   3.035000  3.625000   3.105000 ;
      RECT  2.785000   1.570000  3.625000   1.640000 ;
      RECT  2.790000 135.230000 13.110000 135.300000 ;
      RECT  2.825000 133.090000 13.110000 133.160000 ;
      RECT  2.835000   3.105000  3.625000   3.175000 ;
      RECT  2.855000   1.500000  3.625000   1.570000 ;
      RECT  2.860000 135.160000 13.110000 135.230000 ;
      RECT  2.875000 145.130000  5.945000 146.140000 ;
      RECT  2.895000 133.160000 13.110000 133.230000 ;
      RECT  2.905000   3.175000  3.625000   3.245000 ;
      RECT  2.925000   1.430000  3.625000   1.500000 ;
      RECT  2.930000  85.875000 71.475000  94.750000 ;
      RECT  2.930000  94.750000 75.000000  95.615000 ;
      RECT  2.930000  95.615000 73.545000  95.680000 ;
      RECT  2.930000  95.680000 73.480000  95.745000 ;
      RECT  2.930000  95.745000 73.475000  95.750000 ;
      RECT  2.930000 135.090000 13.110000 135.160000 ;
      RECT  2.965000 133.230000 13.110000 133.300000 ;
      RECT  2.970000  85.835000 71.475000  85.875000 ;
      RECT  2.970000  85.835000 71.475000  85.875000 ;
      RECT  2.975000   3.245000  3.625000   3.315000 ;
      RECT  2.995000   1.360000  3.625000   1.430000 ;
      RECT  3.000000  95.750000 71.475000  95.820000 ;
      RECT  3.000000  95.750000 71.475000  95.820000 ;
      RECT  3.000000  95.750000 73.405000  95.820000 ;
      RECT  3.000000 135.020000 13.110000 135.090000 ;
      RECT  3.035000 133.300000 13.110000 133.370000 ;
      RECT  3.040000  85.765000 71.475000  85.835000 ;
      RECT  3.040000  85.765000 71.475000  85.835000 ;
      RECT  3.045000   3.315000  3.625000   3.385000 ;
      RECT  3.065000   1.290000  3.625000   1.360000 ;
      RECT  3.070000  95.820000 71.475000  95.890000 ;
      RECT  3.070000  95.820000 71.475000  95.890000 ;
      RECT  3.070000  95.820000 73.335000  95.890000 ;
      RECT  3.070000 134.950000 13.110000 135.020000 ;
      RECT  3.090000   3.385000  3.625000   3.430000 ;
      RECT  3.105000 133.370000 13.110000 133.440000 ;
      RECT  3.110000  85.695000 71.475000  85.765000 ;
      RECT  3.110000  85.695000 71.475000  85.765000 ;
      RECT  3.135000   1.220000  3.625000   1.290000 ;
      RECT  3.140000  95.890000 71.475000  95.960000 ;
      RECT  3.140000  95.890000 71.475000  95.960000 ;
      RECT  3.140000  95.890000 73.265000  95.960000 ;
      RECT  3.140000 134.880000 13.110000 134.950000 ;
      RECT  3.160000   3.430000 12.005000   3.500000 ;
      RECT  3.175000 133.440000 13.110000 133.510000 ;
      RECT  3.180000  85.625000 71.475000  85.695000 ;
      RECT  3.180000  85.625000 71.475000  85.695000 ;
      RECT  3.205000   1.150000  3.625000   1.220000 ;
      RECT  3.210000  95.960000 71.475000  96.030000 ;
      RECT  3.210000  95.960000 71.475000  96.030000 ;
      RECT  3.210000  95.960000 73.195000  96.030000 ;
      RECT  3.210000 134.810000 13.110000 134.880000 ;
      RECT  3.230000   3.500000 12.005000   3.570000 ;
      RECT  3.245000 133.510000 13.110000 133.580000 ;
      RECT  3.250000  85.555000 71.475000  85.625000 ;
      RECT  3.250000  85.555000 71.475000  85.625000 ;
      RECT  3.260000  85.545000 71.475000  85.555000 ;
      RECT  3.260000  85.545000 71.475000  85.555000 ;
      RECT  3.260000  85.545000 75.000000  85.555000 ;
      RECT  3.275000   1.080000  3.625000   1.150000 ;
      RECT  3.280000  96.030000 71.475000  96.100000 ;
      RECT  3.280000  96.030000 71.475000  96.100000 ;
      RECT  3.280000  96.030000 73.125000  96.100000 ;
      RECT  3.280000 134.740000 13.110000 134.810000 ;
      RECT  3.300000   3.570000 12.005000   3.640000 ;
      RECT  3.315000 133.580000 13.110000 133.650000 ;
      RECT  3.330000  85.475000 71.475000  85.545000 ;
      RECT  3.330000  85.475000 71.475000  85.545000 ;
      RECT  3.330000  85.475000 75.000000  85.545000 ;
      RECT  3.345000   1.010000  3.625000   1.080000 ;
      RECT  3.350000  96.100000 71.475000  96.170000 ;
      RECT  3.350000  96.100000 71.475000  96.170000 ;
      RECT  3.350000  96.100000 73.055000  96.170000 ;
      RECT  3.350000 134.670000 13.110000 134.740000 ;
      RECT  3.370000   3.640000 12.005000   3.710000 ;
      RECT  3.385000 133.650000 13.110000 133.720000 ;
      RECT  3.400000  85.405000 71.475000  85.475000 ;
      RECT  3.400000  85.405000 71.475000  85.475000 ;
      RECT  3.400000  85.405000 75.000000  85.475000 ;
      RECT  3.415000   0.940000  3.625000   1.010000 ;
      RECT  3.420000  96.170000 71.475000  96.240000 ;
      RECT  3.420000  96.170000 71.475000  96.240000 ;
      RECT  3.420000  96.170000 72.985000  96.240000 ;
      RECT  3.420000 134.600000 13.110000 134.670000 ;
      RECT  3.440000   3.710000 12.005000   3.780000 ;
      RECT  3.455000 133.720000 13.110000 133.790000 ;
      RECT  3.470000  85.335000 71.475000  85.405000 ;
      RECT  3.470000  85.335000 71.475000  85.405000 ;
      RECT  3.470000  85.335000 75.000000  85.405000 ;
      RECT  3.485000   0.870000  3.625000   0.940000 ;
      RECT  3.485000   3.780000 12.005000   3.825000 ;
      RECT  3.490000  85.315000 33.105000  85.335000 ;
      RECT  3.490000  85.315000 33.105000  85.335000 ;
      RECT  3.490000  96.240000 71.475000  96.310000 ;
      RECT  3.490000  96.240000 71.475000  96.310000 ;
      RECT  3.490000  96.240000 72.915000  96.310000 ;
      RECT  3.490000 134.530000 13.110000 134.600000 ;
      RECT  3.525000 133.790000 13.110000 133.860000 ;
      RECT  3.560000  85.245000 33.105000  85.315000 ;
      RECT  3.560000  85.245000 33.105000  85.315000 ;
      RECT  3.560000  96.310000 71.475000  96.380000 ;
      RECT  3.560000  96.310000 71.475000  96.380000 ;
      RECT  3.560000  96.310000 72.845000  96.380000 ;
      RECT  3.560000 134.460000 13.110000 134.530000 ;
      RECT  3.595000 133.860000 13.110000 133.930000 ;
      RECT  3.630000  85.175000 33.105000  85.245000 ;
      RECT  3.630000  85.175000 33.105000  85.245000 ;
      RECT  3.630000  96.380000 71.475000  96.450000 ;
      RECT  3.630000  96.380000 71.475000  96.450000 ;
      RECT  3.630000  96.380000 72.775000  96.450000 ;
      RECT  3.635000 134.390000 13.110000 134.460000 ;
      RECT  3.665000 133.930000 13.110000 134.000000 ;
      RECT  3.700000  85.105000 33.105000  85.175000 ;
      RECT  3.700000  85.105000 33.105000  85.175000 ;
      RECT  3.700000  96.450000 71.475000  96.520000 ;
      RECT  3.700000  96.450000 71.475000  96.520000 ;
      RECT  3.700000  96.450000 72.705000  96.520000 ;
      RECT  3.700000 134.320000 13.110000 134.390000 ;
      RECT  3.735000 134.000000 13.110000 134.070000 ;
      RECT  3.770000  85.035000 33.105000  85.105000 ;
      RECT  3.770000  85.035000 33.105000  85.105000 ;
      RECT  3.770000  96.520000 71.475000  96.590000 ;
      RECT  3.770000  96.520000 71.475000  96.590000 ;
      RECT  3.770000  96.520000 72.635000  96.590000 ;
      RECT  3.775000 134.250000 13.110000 134.320000 ;
      RECT  3.805000 134.070000 13.110000 134.140000 ;
      RECT  3.840000  84.965000 33.105000  85.035000 ;
      RECT  3.840000  84.965000 33.105000  85.035000 ;
      RECT  3.840000  96.590000 71.475000  96.660000 ;
      RECT  3.840000  96.590000 71.475000  96.660000 ;
      RECT  3.840000  96.590000 72.565000  96.660000 ;
      RECT  3.845000 134.140000 13.110000 134.180000 ;
      RECT  3.845000 134.180000 13.110000 134.250000 ;
      RECT  3.905000   1.140000  5.710000   3.150000 ;
      RECT  3.910000  84.895000 33.105000  84.965000 ;
      RECT  3.910000  84.895000 33.105000  84.965000 ;
      RECT  3.910000  96.660000 71.475000  96.730000 ;
      RECT  3.910000  96.660000 71.475000  96.730000 ;
      RECT  3.910000  96.660000 72.495000  96.730000 ;
      RECT  3.980000  84.825000 33.105000  84.895000 ;
      RECT  3.980000  84.825000 33.105000  84.895000 ;
      RECT  3.980000  96.730000 71.475000  96.800000 ;
      RECT  3.980000  96.730000 71.475000  96.800000 ;
      RECT  3.980000  96.730000 72.425000  96.800000 ;
      RECT  4.050000  84.755000 33.105000  84.825000 ;
      RECT  4.050000  84.755000 33.105000  84.825000 ;
      RECT  4.050000  96.800000 71.475000  96.870000 ;
      RECT  4.050000  96.800000 71.475000  96.870000 ;
      RECT  4.050000  96.800000 72.355000  96.870000 ;
      RECT  4.120000  96.870000 71.475000  96.940000 ;
      RECT  4.120000  96.870000 71.475000  96.940000 ;
      RECT  4.120000  96.870000 72.285000  96.940000 ;
      RECT  4.190000  96.940000 71.475000  97.010000 ;
      RECT  4.190000  96.940000 71.475000  97.010000 ;
      RECT  4.190000  96.940000 72.215000  97.010000 ;
      RECT  4.260000  97.010000 71.475000  97.080000 ;
      RECT  4.260000  97.010000 71.475000  97.080000 ;
      RECT  4.260000  97.010000 72.145000  97.080000 ;
      RECT  4.330000  97.080000 71.475000  97.150000 ;
      RECT  4.330000  97.080000 71.475000  97.150000 ;
      RECT  4.330000  97.080000 72.075000  97.150000 ;
      RECT  4.400000  97.150000 71.475000  97.220000 ;
      RECT  4.400000  97.150000 71.475000  97.220000 ;
      RECT  4.400000  97.150000 72.005000  97.220000 ;
      RECT  4.430000  97.220000 71.475000  97.250000 ;
      RECT  4.430000  97.220000 71.475000  97.250000 ;
      RECT  4.430000  97.220000 71.975000  97.250000 ;
      RECT  4.795000   3.430000 12.005000   3.825000 ;
      RECT  4.795000   3.825000 12.005000   6.380000 ;
      RECT  4.795000   6.380000 11.935000   6.450000 ;
      RECT  4.795000   6.380000 11.935000   6.450000 ;
      RECT  4.795000   6.450000 11.865000   6.520000 ;
      RECT  4.795000   6.450000 11.865000   6.520000 ;
      RECT  4.795000   6.520000 11.795000   6.590000 ;
      RECT  4.795000   6.520000 11.795000   6.590000 ;
      RECT  4.795000   6.590000 11.725000   6.660000 ;
      RECT  4.795000   6.590000 11.725000   6.660000 ;
      RECT  4.795000   6.660000 11.655000   6.730000 ;
      RECT  4.795000   6.660000 11.655000   6.730000 ;
      RECT  4.795000   6.730000 11.585000   6.800000 ;
      RECT  4.795000   6.730000 11.585000   6.800000 ;
      RECT  4.795000   6.800000 11.515000   6.870000 ;
      RECT  4.795000   6.800000 11.515000   6.870000 ;
      RECT  4.795000   6.870000 11.445000   6.940000 ;
      RECT  4.795000   6.870000 11.445000   6.940000 ;
      RECT  4.795000   6.940000 11.440000   6.945000 ;
      RECT  4.795000   6.940000 11.440000   6.945000 ;
      RECT  4.795000   6.945000 12.090000   7.040000 ;
      RECT  4.795000   7.040000 12.090000   7.110000 ;
      RECT  4.795000   7.040000 12.090000   7.110000 ;
      RECT  4.795000   7.110000 12.160000   7.180000 ;
      RECT  4.795000   7.110000 12.160000   7.180000 ;
      RECT  4.795000   7.180000 12.230000   7.250000 ;
      RECT  4.795000   7.180000 12.230000   7.250000 ;
      RECT  4.795000   7.250000 12.300000   7.320000 ;
      RECT  4.795000   7.250000 12.300000   7.320000 ;
      RECT  4.795000   7.320000 12.370000   7.365000 ;
      RECT  4.795000   7.320000 12.370000   7.365000 ;
      RECT  4.795000   7.365000 12.415000  10.510000 ;
      RECT  4.795000   7.365000 12.415000  12.455000 ;
      RECT  4.795000   7.365000 12.415000  12.455000 ;
      RECT  4.795000  10.510000 12.520000  10.585000 ;
      RECT  4.795000  10.585000 14.275000  12.455000 ;
      RECT  4.795000  10.585000 14.275000  16.200000 ;
      RECT  4.795000  12.455000 14.275000  12.525000 ;
      RECT  4.795000  12.455000 14.275000  12.525000 ;
      RECT  4.795000  12.525000 14.345000  12.595000 ;
      RECT  4.795000  12.525000 14.345000  12.595000 ;
      RECT  4.795000  12.595000 14.415000  12.665000 ;
      RECT  4.795000  12.595000 14.415000  12.665000 ;
      RECT  4.795000  12.665000 14.485000  12.735000 ;
      RECT  4.795000  12.665000 14.485000  12.735000 ;
      RECT  4.795000  12.735000 14.555000  12.805000 ;
      RECT  4.795000  12.735000 14.555000  12.805000 ;
      RECT  4.795000  12.805000 14.625000  12.875000 ;
      RECT  4.795000  12.805000 14.625000  12.875000 ;
      RECT  4.795000  12.875000 14.695000  12.945000 ;
      RECT  4.795000  12.875000 14.695000  12.945000 ;
      RECT  4.795000  12.945000 14.765000  13.015000 ;
      RECT  4.795000  12.945000 14.765000  13.015000 ;
      RECT  4.795000  13.015000 14.835000  13.085000 ;
      RECT  4.795000  13.015000 14.835000  13.085000 ;
      RECT  4.795000  13.085000 14.905000  13.155000 ;
      RECT  4.795000  13.085000 14.905000  13.155000 ;
      RECT  4.795000  13.155000 14.975000  13.225000 ;
      RECT  4.795000  13.155000 14.975000  13.225000 ;
      RECT  4.795000  13.225000 15.045000  13.295000 ;
      RECT  4.795000  13.225000 15.045000  13.295000 ;
      RECT  4.795000  13.295000 15.115000  13.365000 ;
      RECT  4.795000  13.295000 15.115000  13.365000 ;
      RECT  4.795000  13.365000 15.185000  13.435000 ;
      RECT  4.795000  13.365000 15.185000  13.435000 ;
      RECT  4.795000  13.435000 15.255000  13.505000 ;
      RECT  4.795000  13.435000 15.255000  13.505000 ;
      RECT  4.795000  13.505000 15.325000  13.575000 ;
      RECT  4.795000  13.505000 15.325000  13.575000 ;
      RECT  4.795000  13.575000 15.395000  13.645000 ;
      RECT  4.795000  13.575000 15.395000  13.645000 ;
      RECT  4.795000  13.645000 15.465000  13.715000 ;
      RECT  4.795000  13.645000 15.465000  13.715000 ;
      RECT  4.795000  13.715000 15.535000  13.785000 ;
      RECT  4.795000  13.715000 15.535000  13.785000 ;
      RECT  4.795000  13.785000 15.605000  13.855000 ;
      RECT  4.795000  13.785000 15.605000  13.855000 ;
      RECT  4.795000  13.855000 15.675000  13.925000 ;
      RECT  4.795000  13.855000 15.675000  13.925000 ;
      RECT  4.795000  13.925000 15.745000  13.995000 ;
      RECT  4.795000  13.925000 15.745000  13.995000 ;
      RECT  4.795000  13.995000 15.815000  14.065000 ;
      RECT  4.795000  13.995000 15.815000  14.065000 ;
      RECT  4.795000  14.065000 15.885000  14.135000 ;
      RECT  4.795000  14.065000 15.885000  14.135000 ;
      RECT  4.795000  14.135000 15.955000  14.205000 ;
      RECT  4.795000  14.135000 15.955000  14.205000 ;
      RECT  4.795000  14.205000 16.025000  14.275000 ;
      RECT  4.795000  14.205000 16.025000  14.275000 ;
      RECT  4.795000  14.275000 16.095000  14.345000 ;
      RECT  4.795000  14.275000 16.095000  14.345000 ;
      RECT  4.795000  14.345000 16.165000  14.415000 ;
      RECT  4.795000  14.345000 16.165000  14.415000 ;
      RECT  4.795000  14.415000 16.235000  14.485000 ;
      RECT  4.795000  14.415000 16.235000  14.485000 ;
      RECT  4.795000  14.485000 16.305000  14.555000 ;
      RECT  4.795000  14.485000 16.305000  14.555000 ;
      RECT  4.795000  14.555000 16.375000  14.625000 ;
      RECT  4.795000  14.555000 16.375000  14.625000 ;
      RECT  4.795000  14.625000 16.445000  14.695000 ;
      RECT  4.795000  14.625000 16.445000  14.695000 ;
      RECT  4.795000  14.695000 16.515000  14.765000 ;
      RECT  4.795000  14.695000 16.515000  14.765000 ;
      RECT  4.795000  14.765000 16.585000  14.835000 ;
      RECT  4.795000  14.765000 16.585000  14.835000 ;
      RECT  4.795000  14.835000 16.655000  14.905000 ;
      RECT  4.795000  14.835000 16.655000  14.905000 ;
      RECT  4.795000  14.905000 16.725000  14.975000 ;
      RECT  4.795000  14.905000 16.725000  14.975000 ;
      RECT  4.795000  14.975000 16.795000  15.045000 ;
      RECT  4.795000  14.975000 16.795000  15.045000 ;
      RECT  4.795000  15.045000 16.865000  15.115000 ;
      RECT  4.795000  15.045000 16.865000  15.115000 ;
      RECT  4.795000  15.115000 16.935000  15.185000 ;
      RECT  4.795000  15.115000 16.935000  15.185000 ;
      RECT  4.795000  15.185000 17.005000  15.255000 ;
      RECT  4.795000  15.185000 17.005000  15.255000 ;
      RECT  4.795000  15.255000 17.075000  15.325000 ;
      RECT  4.795000  15.255000 17.075000  15.325000 ;
      RECT  4.795000  15.325000 17.145000  15.395000 ;
      RECT  4.795000  15.325000 17.145000  15.395000 ;
      RECT  4.795000  15.395000 17.215000  15.465000 ;
      RECT  4.795000  15.395000 17.215000  15.465000 ;
      RECT  4.795000  15.465000 17.285000  15.535000 ;
      RECT  4.795000  15.465000 17.285000  15.535000 ;
      RECT  4.795000  15.535000 17.355000  15.605000 ;
      RECT  4.795000  15.535000 17.355000  15.605000 ;
      RECT  4.795000  15.605000 17.425000  15.675000 ;
      RECT  4.795000  15.605000 17.425000  15.675000 ;
      RECT  4.795000  15.675000 17.495000  15.745000 ;
      RECT  4.795000  15.675000 17.495000  15.745000 ;
      RECT  4.795000  15.745000 17.565000  15.815000 ;
      RECT  4.795000  15.745000 17.565000  15.815000 ;
      RECT  4.795000  15.815000 17.635000  15.885000 ;
      RECT  4.795000  15.815000 17.635000  15.885000 ;
      RECT  4.795000  15.885000 17.705000  15.955000 ;
      RECT  4.795000  15.885000 17.705000  15.955000 ;
      RECT  4.795000  15.955000 17.775000  16.025000 ;
      RECT  4.795000  15.955000 17.775000  16.025000 ;
      RECT  4.795000  16.025000 17.845000  16.095000 ;
      RECT  4.795000  16.025000 17.845000  16.095000 ;
      RECT  4.795000  16.095000 17.915000  16.165000 ;
      RECT  4.795000  16.095000 17.915000  16.165000 ;
      RECT  4.795000  16.165000 17.985000  16.200000 ;
      RECT  4.795000  16.165000 17.985000  16.200000 ;
      RECT  4.795000  16.200000 21.420000  16.270000 ;
      RECT  4.795000  16.200000 21.420000  16.270000 ;
      RECT  4.795000  16.270000 21.490000  16.340000 ;
      RECT  4.795000  16.270000 21.490000  16.340000 ;
      RECT  4.795000  16.340000 21.560000  16.410000 ;
      RECT  4.795000  16.340000 21.560000  16.410000 ;
      RECT  4.795000  16.410000 21.630000  16.480000 ;
      RECT  4.795000  16.410000 21.630000  16.480000 ;
      RECT  4.795000  16.480000 21.700000  16.550000 ;
      RECT  4.795000  16.480000 21.700000  16.550000 ;
      RECT  4.795000  16.550000 21.770000  16.620000 ;
      RECT  4.795000  16.550000 21.770000  16.620000 ;
      RECT  4.795000  16.620000 21.840000  16.690000 ;
      RECT  4.795000  16.620000 21.840000  16.690000 ;
      RECT  4.795000  16.690000 21.910000  16.760000 ;
      RECT  4.795000  16.690000 21.910000  16.760000 ;
      RECT  4.795000  16.760000 21.980000  16.830000 ;
      RECT  4.795000  16.760000 21.980000  16.830000 ;
      RECT  4.795000  16.830000 22.050000  16.900000 ;
      RECT  4.795000  16.830000 22.050000  16.900000 ;
      RECT  4.795000  16.900000 22.120000  16.970000 ;
      RECT  4.795000  16.900000 22.120000  16.970000 ;
      RECT  4.795000  16.970000 22.190000  17.040000 ;
      RECT  4.795000  16.970000 22.190000  17.040000 ;
      RECT  4.795000  17.040000 22.260000  17.110000 ;
      RECT  4.795000  17.040000 22.260000  17.110000 ;
      RECT  4.795000  17.110000 22.330000  17.180000 ;
      RECT  4.795000  17.110000 22.330000  17.180000 ;
      RECT  4.795000  17.180000 22.400000  17.250000 ;
      RECT  4.795000  17.180000 22.400000  17.250000 ;
      RECT  4.795000  17.250000 22.470000  17.320000 ;
      RECT  4.795000  17.250000 22.470000  17.320000 ;
      RECT  4.795000  17.320000 22.540000  17.390000 ;
      RECT  4.795000  17.320000 22.540000  17.390000 ;
      RECT  4.795000  17.390000 22.610000  17.460000 ;
      RECT  4.795000  17.390000 22.610000  17.460000 ;
      RECT  4.795000  17.460000 22.680000  17.530000 ;
      RECT  4.795000  17.460000 22.680000  17.530000 ;
      RECT  4.795000  17.530000 22.750000  17.600000 ;
      RECT  4.795000  17.530000 22.750000  17.600000 ;
      RECT  4.795000  17.600000 22.820000  17.670000 ;
      RECT  4.795000  17.600000 22.820000  17.670000 ;
      RECT  4.795000  17.670000 22.890000  17.740000 ;
      RECT  4.795000  17.670000 22.890000  17.740000 ;
      RECT  4.795000  17.740000 22.960000  17.810000 ;
      RECT  4.795000  17.740000 22.960000  17.810000 ;
      RECT  4.795000  17.810000 23.030000  17.880000 ;
      RECT  4.795000  17.810000 23.030000  17.880000 ;
      RECT  4.795000  17.880000 23.100000  17.950000 ;
      RECT  4.795000  17.880000 23.100000  17.950000 ;
      RECT  4.795000  17.950000 23.170000  18.020000 ;
      RECT  4.795000  17.950000 23.170000  18.020000 ;
      RECT  4.795000  18.020000 23.240000  18.090000 ;
      RECT  4.795000  18.020000 23.240000  18.090000 ;
      RECT  4.795000  18.090000 23.310000  18.160000 ;
      RECT  4.795000  18.090000 23.310000  18.160000 ;
      RECT  4.795000  18.160000 23.380000  18.230000 ;
      RECT  4.795000  18.160000 23.380000  18.230000 ;
      RECT  4.795000  18.230000 23.450000  18.300000 ;
      RECT  4.795000  18.230000 23.450000  18.300000 ;
      RECT  4.795000  18.300000 23.520000  18.370000 ;
      RECT  4.795000  18.300000 23.520000  18.370000 ;
      RECT  4.795000  18.370000 23.590000  18.440000 ;
      RECT  4.795000  18.370000 23.590000  18.440000 ;
      RECT  4.795000  18.440000 23.660000  18.510000 ;
      RECT  4.795000  18.440000 23.660000  18.510000 ;
      RECT  4.795000  18.510000 23.730000  18.580000 ;
      RECT  4.795000  18.510000 23.730000  18.580000 ;
      RECT  4.795000  18.580000 23.800000  18.650000 ;
      RECT  4.795000  18.580000 23.800000  18.650000 ;
      RECT  4.795000  18.650000 23.870000  18.720000 ;
      RECT  4.795000  18.650000 23.870000  18.720000 ;
      RECT  4.795000  18.720000 23.940000  18.725000 ;
      RECT  4.795000  18.720000 23.940000  18.725000 ;
      RECT  4.795000  18.725000 23.945000  25.470000 ;
      RECT  4.795000  18.725000 23.945000  26.060000 ;
      RECT  4.795000  25.470000 23.945000  25.540000 ;
      RECT  4.795000  25.470000 23.945000  25.540000 ;
      RECT  4.795000  25.540000 24.015000  25.610000 ;
      RECT  4.795000  25.540000 24.015000  25.610000 ;
      RECT  4.795000  25.610000 24.085000  25.680000 ;
      RECT  4.795000  25.610000 24.085000  25.680000 ;
      RECT  4.795000  25.680000 24.155000  25.750000 ;
      RECT  4.795000  25.680000 24.155000  25.750000 ;
      RECT  4.795000  25.750000 24.225000  25.820000 ;
      RECT  4.795000  25.750000 24.225000  25.820000 ;
      RECT  4.795000  25.820000 24.295000  25.890000 ;
      RECT  4.795000  25.820000 24.295000  25.890000 ;
      RECT  4.795000  25.890000 24.365000  25.960000 ;
      RECT  4.795000  25.890000 24.365000  25.960000 ;
      RECT  4.795000  25.960000 24.435000  26.030000 ;
      RECT  4.795000  25.960000 24.435000  26.030000 ;
      RECT  4.795000  26.030000 24.505000  26.060000 ;
      RECT  4.795000  26.030000 24.505000  26.060000 ;
      RECT  4.795000  26.060000 24.535000  42.625000 ;
      RECT  4.795000  42.625000 24.465000  42.695000 ;
      RECT  4.795000  42.625000 24.465000  42.695000 ;
      RECT  4.795000  42.695000 24.395000  42.765000 ;
      RECT  4.795000  42.695000 24.395000  42.765000 ;
      RECT  4.795000  42.765000 24.325000  42.835000 ;
      RECT  4.795000  42.765000 24.325000  42.835000 ;
      RECT  4.795000  42.835000 24.255000  42.905000 ;
      RECT  4.795000  42.835000 24.255000  42.905000 ;
      RECT  4.795000  42.905000 24.185000  42.975000 ;
      RECT  4.795000  42.905000 24.185000  42.975000 ;
      RECT  4.795000  42.975000 24.155000  43.005000 ;
      RECT  4.795000  42.975000 24.155000  43.005000 ;
      RECT  4.795000  43.005000  5.785000  43.825000 ;
      RECT  4.795000  43.825000 73.380000  71.630000 ;
      RECT  5.990000   0.870000 12.005000   3.430000 ;
      RECT  6.225000 143.875000 70.525000 144.285000 ;
      RECT  6.225000 144.285000 70.455000 144.355000 ;
      RECT  6.225000 144.285000 70.455000 144.355000 ;
      RECT  6.225000 144.355000 70.385000 144.425000 ;
      RECT  6.225000 144.355000 70.385000 144.425000 ;
      RECT  6.225000 144.425000 70.315000 144.495000 ;
      RECT  6.225000 144.425000 70.315000 144.495000 ;
      RECT  6.225000 144.495000 70.245000 144.565000 ;
      RECT  6.225000 144.495000 70.245000 144.565000 ;
      RECT  6.225000 144.565000 70.175000 144.635000 ;
      RECT  6.225000 144.565000 70.175000 144.635000 ;
      RECT  6.225000 144.635000 70.105000 144.705000 ;
      RECT  6.225000 144.635000 70.105000 144.705000 ;
      RECT  6.225000 144.705000 70.035000 144.775000 ;
      RECT  6.225000 144.705000 70.035000 144.775000 ;
      RECT  6.225000 144.775000 69.965000 144.845000 ;
      RECT  6.225000 144.775000 69.965000 144.845000 ;
      RECT  6.225000 144.845000 69.960000 144.850000 ;
      RECT  6.225000 144.845000 69.960000 144.850000 ;
      RECT  6.225000 144.850000 69.890000 144.920000 ;
      RECT  6.225000 144.850000 69.890000 144.920000 ;
      RECT  6.225000 144.920000 69.820000 144.990000 ;
      RECT  6.225000 144.920000 69.820000 144.990000 ;
      RECT  6.225000 144.990000 69.750000 145.060000 ;
      RECT  6.225000 144.990000 69.750000 145.060000 ;
      RECT  6.225000 145.060000 69.680000 145.130000 ;
      RECT  6.225000 145.060000 69.680000 145.130000 ;
      RECT  6.225000 145.130000 69.610000 145.200000 ;
      RECT  6.225000 145.130000 69.610000 145.200000 ;
      RECT  6.225000 145.200000 69.540000 145.270000 ;
      RECT  6.225000 145.200000 69.540000 145.270000 ;
      RECT  6.225000 145.270000 69.470000 145.340000 ;
      RECT  6.225000 145.270000 69.470000 145.340000 ;
      RECT  6.225000 145.340000 69.400000 145.410000 ;
      RECT  6.225000 145.340000 69.400000 145.410000 ;
      RECT  6.225000 145.410000 70.525000 146.420000 ;
      RECT  6.225000 145.410000 70.525000 195.970000 ;
      RECT  8.190000 132.395000 72.380000 132.460000 ;
      RECT  8.190000 132.395000 72.380000 132.460000 ;
      RECT  8.260000 132.325000 72.380000 132.395000 ;
      RECT  8.260000 132.325000 72.380000 132.395000 ;
      RECT  8.330000 132.255000 72.380000 132.325000 ;
      RECT  8.330000 132.255000 72.380000 132.325000 ;
      RECT  8.400000 132.185000 72.380000 132.255000 ;
      RECT  8.400000 132.185000 72.380000 132.255000 ;
      RECT  8.470000 132.115000 72.380000 132.185000 ;
      RECT  8.470000 132.115000 72.380000 132.185000 ;
      RECT  8.540000 132.045000 72.380000 132.115000 ;
      RECT  8.540000 132.045000 72.380000 132.115000 ;
      RECT  8.610000 131.975000 72.380000 132.045000 ;
      RECT  8.610000 131.975000 72.380000 132.045000 ;
      RECT  8.680000 131.905000 72.380000 131.975000 ;
      RECT  8.680000 131.905000 72.380000 131.975000 ;
      RECT  8.750000 131.835000 72.380000 131.905000 ;
      RECT  8.750000 131.835000 72.380000 131.905000 ;
      RECT  8.820000 131.765000 72.380000 131.835000 ;
      RECT  8.820000 131.765000 72.380000 131.835000 ;
      RECT  8.890000 131.695000 72.380000 131.765000 ;
      RECT  8.890000 131.695000 72.380000 131.765000 ;
      RECT  8.960000 131.625000 72.380000 131.695000 ;
      RECT  8.960000 131.625000 72.380000 131.695000 ;
      RECT  9.030000 131.555000 72.380000 131.625000 ;
      RECT  9.030000 131.555000 72.380000 131.625000 ;
      RECT  9.100000 131.485000 72.380000 131.555000 ;
      RECT  9.100000 131.485000 72.380000 131.555000 ;
      RECT  9.170000 131.415000 72.380000 131.485000 ;
      RECT  9.170000 131.415000 72.380000 131.485000 ;
      RECT  9.240000 131.345000 72.380000 131.415000 ;
      RECT  9.240000 131.345000 72.380000 131.415000 ;
      RECT  9.310000 131.275000 72.380000 131.345000 ;
      RECT  9.310000 131.275000 72.380000 131.345000 ;
      RECT  9.380000 131.205000 72.380000 131.275000 ;
      RECT  9.380000 131.205000 72.380000 131.275000 ;
      RECT  9.450000 131.135000 72.380000 131.205000 ;
      RECT  9.450000 131.135000 72.380000 131.205000 ;
      RECT  9.520000 131.065000 72.380000 131.135000 ;
      RECT  9.520000 131.065000 72.380000 131.135000 ;
      RECT  9.590000 130.995000 72.380000 131.065000 ;
      RECT  9.590000 130.995000 72.380000 131.065000 ;
      RECT  9.595000 130.990000 72.380000 130.995000 ;
      RECT  9.595000 130.990000 72.380000 130.995000 ;
      RECT  9.665000 130.920000 72.380000 130.990000 ;
      RECT  9.665000 130.920000 72.380000 130.990000 ;
      RECT  9.735000 130.850000 72.380000 130.920000 ;
      RECT  9.735000 130.850000 72.380000 130.920000 ;
      RECT  9.805000 130.780000 72.380000 130.850000 ;
      RECT  9.805000 130.780000 72.380000 130.850000 ;
      RECT  9.875000 130.710000 72.380000 130.780000 ;
      RECT  9.875000 130.710000 72.380000 130.780000 ;
      RECT  9.945000 130.640000 72.380000 130.710000 ;
      RECT  9.945000 130.640000 72.380000 130.710000 ;
      RECT 10.015000 130.570000 72.380000 130.640000 ;
      RECT 10.015000 130.570000 72.380000 130.640000 ;
      RECT 10.085000 130.500000 72.380000 130.570000 ;
      RECT 10.085000 130.500000 72.380000 130.570000 ;
      RECT 10.155000 130.430000 64.845000 130.500000 ;
      RECT 10.155000 130.430000 64.845000 130.500000 ;
      RECT 10.225000 130.360000 64.775000 130.430000 ;
      RECT 10.225000 130.360000 64.775000 130.430000 ;
      RECT 10.295000 130.290000 64.705000 130.360000 ;
      RECT 10.295000 130.290000 64.705000 130.360000 ;
      RECT 10.365000 130.220000 64.635000 130.290000 ;
      RECT 10.365000 130.220000 64.635000 130.290000 ;
      RECT 10.435000 130.150000 64.565000 130.220000 ;
      RECT 10.435000 130.150000 64.565000 130.220000 ;
      RECT 10.505000 130.080000 64.495000 130.150000 ;
      RECT 10.505000 130.080000 64.495000 130.150000 ;
      RECT 10.575000 130.010000 64.425000 130.080000 ;
      RECT 10.575000 130.010000 64.425000 130.080000 ;
      RECT 10.645000 129.940000 64.355000 130.010000 ;
      RECT 10.645000 129.940000 64.355000 130.010000 ;
      RECT 10.715000 129.870000 64.285000 129.940000 ;
      RECT 10.715000 129.870000 64.285000 129.940000 ;
      RECT 10.785000 129.800000 64.215000 129.870000 ;
      RECT 10.785000 129.800000 64.215000 129.870000 ;
      RECT 10.855000 129.730000 64.145000 129.800000 ;
      RECT 10.855000 129.730000 64.145000 129.800000 ;
      RECT 10.925000 129.660000 64.075000 129.730000 ;
      RECT 10.925000 129.660000 64.075000 129.730000 ;
      RECT 10.995000 129.590000 64.005000 129.660000 ;
      RECT 10.995000 129.590000 64.005000 129.660000 ;
      RECT 11.065000 129.520000 63.935000 129.590000 ;
      RECT 11.065000 129.520000 63.935000 129.590000 ;
      RECT 11.135000 129.450000 63.865000 129.520000 ;
      RECT 11.135000 129.450000 63.865000 129.520000 ;
      RECT 11.205000 129.380000 63.795000 129.450000 ;
      RECT 11.205000 129.380000 63.795000 129.450000 ;
      RECT 11.255000 139.225000 14.920000 139.260000 ;
      RECT 11.255000 139.225000 14.920000 139.260000 ;
      RECT 11.275000 129.310000 63.725000 129.380000 ;
      RECT 11.275000 129.310000 63.725000 129.380000 ;
      RECT 11.290000 139.260000 14.920000 139.295000 ;
      RECT 11.290000 139.260000 14.920000 139.295000 ;
      RECT 11.345000 129.240000 63.655000 129.310000 ;
      RECT 11.345000 129.240000 63.655000 129.310000 ;
      RECT 11.415000 129.170000 63.585000 129.240000 ;
      RECT 11.415000 129.170000 63.585000 129.240000 ;
      RECT 11.485000 129.100000 63.515000 129.170000 ;
      RECT 11.485000 129.100000 63.515000 129.170000 ;
      RECT 11.555000 129.030000 63.445000 129.100000 ;
      RECT 11.555000 129.030000 63.445000 129.100000 ;
      RECT 11.625000 128.960000 63.375000 129.030000 ;
      RECT 11.625000 128.960000 63.375000 129.030000 ;
      RECT 11.695000 128.890000 63.305000 128.960000 ;
      RECT 11.695000 128.890000 63.305000 128.960000 ;
      RECT 11.765000 128.820000 63.235000 128.890000 ;
      RECT 11.765000 128.820000 63.235000 128.890000 ;
      RECT 11.835000 128.750000 63.165000 128.820000 ;
      RECT 11.835000 128.750000 63.165000 128.820000 ;
      RECT 11.905000 128.680000 63.095000 128.750000 ;
      RECT 11.905000 128.680000 63.095000 128.750000 ;
      RECT 11.950000 128.240000 63.050000 128.260000 ;
      RECT 11.975000 128.610000 63.025000 128.680000 ;
      RECT 11.975000 128.610000 63.025000 128.680000 ;
      RECT 12.020000 128.170000 62.980000 128.240000 ;
      RECT 12.045000 128.540000 62.955000 128.610000 ;
      RECT 12.045000 128.540000 62.955000 128.610000 ;
      RECT 12.090000 128.100000 62.910000 128.170000 ;
      RECT 12.160000 128.030000 62.840000 128.100000 ;
      RECT 12.230000 127.960000 62.770000 128.030000 ;
      RECT 12.300000 127.890000 62.700000 127.960000 ;
      RECT 12.370000 127.820000 62.630000 127.890000 ;
      RECT 12.440000 127.750000 62.560000 127.820000 ;
      RECT 12.510000 127.680000 62.490000 127.750000 ;
      RECT 12.580000 127.610000 62.420000 127.680000 ;
      RECT 12.650000 127.540000 62.350000 127.610000 ;
      RECT 12.685000   0.000000 14.415000   6.715000 ;
      RECT 12.685000   6.715000 14.415000   7.070000 ;
      RECT 12.720000 127.470000 62.280000 127.540000 ;
      RECT 12.790000 127.400000 62.210000 127.470000 ;
      RECT 12.825000   3.550000 14.275000   6.660000 ;
      RECT 12.860000 127.330000 62.140000 127.400000 ;
      RECT 12.895000   6.660000 14.275000   6.730000 ;
      RECT 12.920000   0.240000 13.915000   3.270000 ;
      RECT 12.930000 127.260000 62.070000 127.330000 ;
      RECT 12.965000   6.730000 14.275000   6.800000 ;
      RECT 12.970000  10.555000 14.275000  10.585000 ;
      RECT 13.000000 127.190000 62.000000 127.260000 ;
      RECT 13.035000   6.800000 14.275000   6.870000 ;
      RECT 13.040000   7.070000 14.415000  10.290000 ;
      RECT 13.040000  10.290000 14.415000  10.445000 ;
      RECT 13.040000  10.485000 14.275000  10.555000 ;
      RECT 13.070000 127.120000 61.930000 127.190000 ;
      RECT 13.105000   6.870000 14.275000   6.940000 ;
      RECT 13.110000  10.415000 14.275000  10.485000 ;
      RECT 13.140000 127.050000 61.860000 127.120000 ;
      RECT 13.175000   6.940000 14.275000   7.010000 ;
      RECT 13.180000   7.010000 14.275000   7.015000 ;
      RECT 13.180000   7.015000 14.275000  10.345000 ;
      RECT 13.180000  10.345000 14.275000  10.415000 ;
      RECT 13.210000 126.980000 61.790000 127.050000 ;
      RECT 13.280000 126.910000 61.720000 126.980000 ;
      RECT 13.350000 126.840000 61.650000 126.910000 ;
      RECT 13.390000 130.500000 72.380000 135.750000 ;
      RECT 13.390000 132.460000 72.380000 135.285000 ;
      RECT 13.390000 135.285000 72.310000 135.355000 ;
      RECT 13.390000 135.285000 72.310000 135.355000 ;
      RECT 13.390000 135.355000 72.240000 135.425000 ;
      RECT 13.390000 135.355000 72.240000 135.425000 ;
      RECT 13.390000 135.425000 72.170000 135.495000 ;
      RECT 13.390000 135.425000 72.170000 135.495000 ;
      RECT 13.390000 135.495000 72.100000 135.565000 ;
      RECT 13.390000 135.495000 72.100000 135.565000 ;
      RECT 13.390000 135.565000 72.030000 135.635000 ;
      RECT 13.390000 135.565000 72.030000 135.635000 ;
      RECT 13.390000 135.635000 71.960000 135.705000 ;
      RECT 13.390000 135.635000 71.960000 135.705000 ;
      RECT 13.390000 135.705000 71.915000 135.750000 ;
      RECT 13.390000 135.705000 71.915000 135.750000 ;
      RECT 13.420000 126.770000 61.580000 126.840000 ;
      RECT 13.490000 126.700000 61.510000 126.770000 ;
      RECT 13.560000 126.630000 61.440000 126.700000 ;
      RECT 13.630000 126.560000 61.370000 126.630000 ;
      RECT 13.700000 126.490000 61.300000 126.560000 ;
      RECT 13.770000 126.420000 61.230000 126.490000 ;
      RECT 13.840000 126.350000 61.160000 126.420000 ;
      RECT 13.910000 126.280000 61.090000 126.350000 ;
      RECT 13.980000 126.210000 61.020000 126.280000 ;
      RECT 14.050000 126.140000 60.950000 126.210000 ;
      RECT 14.120000 126.070000 60.880000 126.140000 ;
      RECT 14.190000 126.000000 60.810000 126.070000 ;
      RECT 14.260000 125.930000 60.740000 126.000000 ;
      RECT 14.330000 125.860000 60.670000 125.930000 ;
      RECT 14.400000 125.790000 60.600000 125.860000 ;
      RECT 14.470000 125.720000 60.530000 125.790000 ;
      RECT 14.540000 125.650000 60.460000 125.720000 ;
      RECT 14.610000 125.580000 60.390000 125.650000 ;
      RECT 14.680000 125.510000 60.320000 125.580000 ;
      RECT 14.750000 125.440000 60.250000 125.510000 ;
      RECT 15.200000 138.990000 69.130000 139.060000 ;
      RECT 15.200000 139.060000 69.200000 139.130000 ;
      RECT 15.200000 139.130000 69.270000 139.200000 ;
      RECT 15.200000 139.200000 69.340000 139.270000 ;
      RECT 15.200000 139.270000 69.410000 139.340000 ;
      RECT 15.200000 139.340000 69.480000 139.410000 ;
      RECT 15.200000 139.410000 69.550000 139.480000 ;
      RECT 15.200000 139.480000 69.620000 139.550000 ;
      RECT 15.200000 139.550000 69.690000 139.575000 ;
      RECT 15.275000   0.000000 22.220000   1.345000 ;
      RECT 15.275000   1.345000 24.765000  11.280000 ;
      RECT 15.275000  11.280000 16.460000  12.150000 ;
      RECT 15.275000  12.150000 16.460000  12.470000 ;
      RECT 15.415000   0.830000 16.780000   3.430000 ;
      RECT 15.415000   3.430000 24.625000  11.140000 ;
      RECT 15.415000  11.140000 16.320000  12.095000 ;
      RECT 15.485000  12.095000 16.320000  12.165000 ;
      RECT 15.525000   0.200000 21.315000   0.550000 ;
      RECT 15.555000  12.165000 16.320000  12.235000 ;
      RECT 15.590000  12.470000 16.995000  13.005000 ;
      RECT 15.625000  12.235000 16.320000  12.305000 ;
      RECT 15.695000  12.305000 16.320000  12.375000 ;
      RECT 15.765000  12.375000 16.320000  12.445000 ;
      RECT 15.835000  12.445000 16.320000  12.515000 ;
      RECT 15.845000  12.515000 16.320000  12.525000 ;
      RECT 15.915000  12.525000 16.320000  12.595000 ;
      RECT 15.985000  12.595000 16.390000  12.665000 ;
      RECT 16.055000  12.665000 16.460000  12.735000 ;
      RECT 16.125000  12.735000 16.530000  12.805000 ;
      RECT 16.125000  13.005000 25.015000  13.175000 ;
      RECT 16.195000  12.805000 16.600000  12.875000 ;
      RECT 16.265000  12.875000 16.670000  12.945000 ;
      RECT 16.295000  13.175000 25.015000  15.195000 ;
      RECT 16.335000  12.945000 16.740000  13.015000 ;
      RECT 16.405000  13.015000 16.810000  13.085000 ;
      RECT 16.465000  13.085000 16.880000  13.145000 ;
      RECT 16.510000  13.145000 24.790000  13.190000 ;
      RECT 16.550000  13.190000 24.835000  13.230000 ;
      RECT 16.620000  13.230000 24.875000  13.300000 ;
      RECT 16.690000  13.300000 24.875000  13.370000 ;
      RECT 16.760000  13.370000 24.875000  13.440000 ;
      RECT 16.830000  13.440000 24.875000  13.510000 ;
      RECT 16.885000 138.985000 75.145000 138.990000 ;
      RECT 16.900000  13.510000 24.875000  13.580000 ;
      RECT 16.905000 138.965000 75.145000 138.985000 ;
      RECT 16.925000 138.945000 75.145000 138.965000 ;
      RECT 16.970000  11.280000 24.765000  12.250000 ;
      RECT 16.970000  12.250000 24.765000  12.290000 ;
      RECT 16.970000  13.580000 24.875000  13.650000 ;
      RECT 17.010000  12.290000 24.560000  12.495000 ;
      RECT 17.040000  13.650000 24.875000  13.720000 ;
      RECT 17.060000   1.140000 18.910000   3.150000 ;
      RECT 17.110000   3.430000 24.625000  12.195000 ;
      RECT 17.110000  11.140000 24.625000  12.195000 ;
      RECT 17.110000  13.720000 24.875000  13.790000 ;
      RECT 17.130000  12.195000 24.625000  12.215000 ;
      RECT 17.130000  12.195000 24.625000  12.215000 ;
      RECT 17.150000  12.215000 24.625000  12.235000 ;
      RECT 17.150000  12.215000 24.625000  12.235000 ;
      RECT 17.180000  13.790000 24.875000  13.860000 ;
      RECT 17.210000  12.235000 24.565000  12.295000 ;
      RECT 17.210000  12.235000 24.565000  12.295000 ;
      RECT 17.250000  13.860000 24.875000  13.930000 ;
      RECT 17.270000  12.295000 24.505000  12.355000 ;
      RECT 17.270000  12.295000 24.505000  12.355000 ;
      RECT 17.320000  13.930000 24.875000  14.000000 ;
      RECT 17.390000  14.000000 24.875000  14.070000 ;
      RECT 17.460000  14.070000 24.875000  14.140000 ;
      RECT 17.530000  14.140000 24.875000  14.210000 ;
      RECT 17.600000  14.210000 24.875000  14.280000 ;
      RECT 17.670000  14.280000 24.875000  14.350000 ;
      RECT 17.740000  14.350000 24.875000  14.420000 ;
      RECT 17.810000  14.420000 24.875000  14.490000 ;
      RECT 17.880000  14.490000 24.875000  14.560000 ;
      RECT 17.950000  14.560000 24.875000  14.630000 ;
      RECT 18.020000  14.630000 24.875000  14.700000 ;
      RECT 18.090000  14.700000 24.875000  14.770000 ;
      RECT 18.160000  14.770000 24.875000  14.840000 ;
      RECT 18.230000  14.840000 24.875000  14.910000 ;
      RECT 18.300000  14.910000 24.875000  14.980000 ;
      RECT 18.315000  15.195000 25.100000  15.280000 ;
      RECT 18.370000  14.980000 24.875000  15.050000 ;
      RECT 18.440000  15.050000 24.875000  15.120000 ;
      RECT 18.460000  15.120000 24.875000  15.140000 ;
      RECT 18.985000   0.550000 21.315000   0.620000 ;
      RECT 19.055000   0.620000 21.315000   0.690000 ;
      RECT 19.125000   0.690000 21.315000   0.760000 ;
      RECT 19.190000   2.785000 22.900000   2.855000 ;
      RECT 19.190000   2.785000 22.900000   2.855000 ;
      RECT 19.190000   2.855000 22.970000   2.925000 ;
      RECT 19.190000   2.855000 22.970000   2.925000 ;
      RECT 19.190000   2.925000 23.040000   2.995000 ;
      RECT 19.190000   2.925000 23.040000   2.995000 ;
      RECT 19.190000   2.995000 23.110000   3.065000 ;
      RECT 19.190000   2.995000 23.110000   3.065000 ;
      RECT 19.190000   3.065000 23.180000   3.135000 ;
      RECT 19.190000   3.065000 23.180000   3.135000 ;
      RECT 19.190000   3.135000 23.250000   3.205000 ;
      RECT 19.190000   3.135000 23.250000   3.205000 ;
      RECT 19.190000   3.205000 23.320000   3.275000 ;
      RECT 19.190000   3.205000 23.320000   3.275000 ;
      RECT 19.190000   3.275000 23.390000   3.280000 ;
      RECT 19.190000   3.275000 23.390000   3.280000 ;
      RECT 19.190000   3.280000 24.625000   3.430000 ;
      RECT 19.190000   3.280000 24.625000  11.140000 ;
      RECT 19.190000   3.280000 24.625000  11.140000 ;
      RECT 19.195000   0.760000 21.315000   0.830000 ;
      RECT 19.265000   0.830000 21.385000   0.900000 ;
      RECT 19.335000   0.900000 21.455000   0.970000 ;
      RECT 19.405000   0.970000 21.525000   1.040000 ;
      RECT 19.475000   1.040000 21.595000   1.110000 ;
      RECT 19.540000  71.630000 73.380000  80.155000 ;
      RECT 19.545000   1.110000 21.665000   1.180000 ;
      RECT 19.580000   1.180000 21.735000   1.215000 ;
      RECT 19.580000   1.215000 21.770000   1.285000 ;
      RECT 19.580000   1.285000 21.840000   1.355000 ;
      RECT 19.580000   1.355000 21.910000   1.425000 ;
      RECT 19.580000   1.425000 21.980000   1.495000 ;
      RECT 19.580000   1.495000 22.050000   1.565000 ;
      RECT 19.580000   1.565000 22.120000   1.585000 ;
      RECT 19.580000   1.585000 24.585000   2.505000 ;
      RECT 21.595000   0.000000 22.080000   0.645000 ;
      RECT 21.665000   0.645000 22.080000   0.715000 ;
      RECT 21.735000   0.715000 22.080000   0.785000 ;
      RECT 21.805000   0.785000 22.080000   0.855000 ;
      RECT 21.805000  15.280000 25.805000  15.985000 ;
      RECT 21.875000   0.855000 22.080000   0.925000 ;
      RECT 21.915000  15.140000 24.875000  15.195000 ;
      RECT 21.945000   0.925000 22.080000   0.995000 ;
      RECT 21.970000  15.195000 24.875000  15.250000 ;
      RECT 22.015000   0.995000 22.080000   1.065000 ;
      RECT 22.040000  15.250000 24.875000  15.320000 ;
      RECT 22.110000  15.320000 24.945000  15.390000 ;
      RECT 22.180000  15.390000 25.015000  15.460000 ;
      RECT 22.250000  15.460000 25.085000  15.530000 ;
      RECT 22.320000  15.530000 25.155000  15.600000 ;
      RECT 22.390000  15.600000 25.225000  15.670000 ;
      RECT 22.460000  15.670000 25.295000  15.740000 ;
      RECT 22.505000  15.985000 30.665000  16.845000 ;
      RECT 22.530000  15.740000 25.365000  15.810000 ;
      RECT 22.600000  15.810000 25.435000  15.880000 ;
      RECT 22.670000  15.880000 25.505000  15.950000 ;
      RECT 22.740000  15.950000 25.575000  16.020000 ;
      RECT 22.790000   1.560000 24.585000   1.585000 ;
      RECT 22.800000   0.000000 24.765000   1.345000 ;
      RECT 22.810000  16.020000 25.645000  16.090000 ;
      RECT 22.845000  16.090000 25.715000  16.125000 ;
      RECT 22.860000   1.490000 24.585000   1.560000 ;
      RECT 22.915000  16.125000 29.750000  16.195000 ;
      RECT 22.915000  16.125000 29.750000  16.195000 ;
      RECT 22.930000   1.420000 24.585000   1.490000 ;
      RECT 22.940000   0.000000 24.625000   0.390000 ;
      RECT 22.940000   0.390000 23.210000   0.745000 ;
      RECT 22.940000   0.745000 23.140000   0.815000 ;
      RECT 22.940000   0.815000 23.070000   0.885000 ;
      RECT 22.940000   0.885000 23.000000   0.955000 ;
      RECT 22.985000  16.195000 29.820000  16.265000 ;
      RECT 22.985000  16.195000 29.820000  16.265000 ;
      RECT 23.000000   1.350000 24.585000   1.420000 ;
      RECT 23.055000  16.265000 29.890000  16.335000 ;
      RECT 23.055000  16.265000 29.890000  16.335000 ;
      RECT 23.070000   1.280000 24.585000   1.350000 ;
      RECT 23.085000   2.505000 24.585000   2.575000 ;
      RECT 23.125000  16.335000 29.960000  16.405000 ;
      RECT 23.125000  16.335000 29.960000  16.405000 ;
      RECT 23.140000   1.210000 24.585000   1.280000 ;
      RECT 23.155000   2.575000 24.585000   2.645000 ;
      RECT 23.195000  16.405000 30.030000  16.475000 ;
      RECT 23.195000  16.405000 30.030000  16.475000 ;
      RECT 23.210000   1.140000 24.585000   1.210000 ;
      RECT 23.225000   2.645000 24.585000   2.715000 ;
      RECT 23.265000  16.475000 30.100000  16.545000 ;
      RECT 23.265000  16.475000 30.100000  16.545000 ;
      RECT 23.280000   1.070000 24.585000   1.140000 ;
      RECT 23.295000   2.715000 24.585000   2.785000 ;
      RECT 23.335000  16.545000 30.170000  16.615000 ;
      RECT 23.335000  16.545000 30.170000  16.615000 ;
      RECT 23.350000   1.000000 24.585000   1.070000 ;
      RECT 23.365000   2.785000 24.585000   2.855000 ;
      RECT 23.365000  16.845000 30.665000  18.340000 ;
      RECT 23.405000  16.615000 30.240000  16.685000 ;
      RECT 23.405000  16.615000 30.240000  16.685000 ;
      RECT 23.420000   0.930000 24.585000   1.000000 ;
      RECT 23.435000   2.855000 24.585000   2.925000 ;
      RECT 23.475000  16.685000 30.310000  16.755000 ;
      RECT 23.475000  16.685000 30.310000  16.755000 ;
      RECT 23.490000   0.670000 24.585000   0.860000 ;
      RECT 23.490000   0.860000 24.585000   0.930000 ;
      RECT 23.505000   2.925000 24.585000   2.995000 ;
      RECT 23.510000   2.995000 24.585000   3.000000 ;
      RECT 23.545000  16.755000 30.380000  16.825000 ;
      RECT 23.545000  16.755000 30.380000  16.825000 ;
      RECT 23.615000  16.825000 30.450000  16.895000 ;
      RECT 23.615000  16.825000 30.450000  16.895000 ;
      RECT 23.620000  16.895000 30.520000  16.900000 ;
      RECT 23.620000  16.895000 30.520000  16.900000 ;
      RECT 23.690000  16.900000 30.525000  16.970000 ;
      RECT 23.690000  16.900000 30.525000  16.970000 ;
      RECT 23.760000  16.970000 30.525000  17.040000 ;
      RECT 23.760000  16.970000 30.525000  17.040000 ;
      RECT 23.830000  17.040000 30.525000  17.110000 ;
      RECT 23.830000  17.040000 30.525000  17.110000 ;
      RECT 23.900000  17.110000 30.525000  17.180000 ;
      RECT 23.900000  17.110000 30.525000  17.180000 ;
      RECT 23.970000  17.180000 30.525000  17.250000 ;
      RECT 23.970000  17.180000 30.525000  17.250000 ;
      RECT 24.040000  17.250000 30.525000  17.320000 ;
      RECT 24.040000  17.250000 30.525000  17.320000 ;
      RECT 24.110000  17.320000 30.525000  17.390000 ;
      RECT 24.110000  17.320000 30.525000  17.390000 ;
      RECT 24.180000  17.390000 30.525000  17.460000 ;
      RECT 24.180000  17.390000 30.525000  17.460000 ;
      RECT 24.250000  17.460000 30.525000  17.530000 ;
      RECT 24.250000  17.460000 30.525000  17.530000 ;
      RECT 24.320000  17.530000 30.525000  17.600000 ;
      RECT 24.320000  17.530000 30.525000  17.600000 ;
      RECT 24.390000  17.600000 30.525000  17.670000 ;
      RECT 24.390000  17.600000 30.525000  17.670000 ;
      RECT 24.460000  17.670000 30.525000  17.740000 ;
      RECT 24.460000  17.670000 30.525000  17.740000 ;
      RECT 24.530000  17.740000 30.525000  17.810000 ;
      RECT 24.530000  17.740000 30.525000  17.810000 ;
      RECT 24.545000  43.775000 73.380000  43.825000 ;
      RECT 24.545000  43.775000 73.380000  43.825000 ;
      RECT 24.600000  17.810000 30.525000  17.880000 ;
      RECT 24.600000  17.810000 30.525000  17.880000 ;
      RECT 24.615000  43.705000 73.380000  43.775000 ;
      RECT 24.615000  43.705000 73.380000  43.775000 ;
      RECT 24.670000  17.880000 30.525000  17.950000 ;
      RECT 24.670000  17.880000 30.525000  17.950000 ;
      RECT 24.685000  43.635000 73.380000  43.705000 ;
      RECT 24.685000  43.635000 73.380000  43.705000 ;
      RECT 24.740000  17.950000 30.525000  18.020000 ;
      RECT 24.740000  17.950000 30.525000  18.020000 ;
      RECT 24.755000  43.565000 73.380000  43.635000 ;
      RECT 24.755000  43.565000 73.380000  43.635000 ;
      RECT 24.810000  18.020000 30.525000  18.090000 ;
      RECT 24.810000  18.020000 30.525000  18.090000 ;
      RECT 24.825000  43.495000 73.380000  43.565000 ;
      RECT 24.825000  43.495000 73.380000  43.565000 ;
      RECT 24.865000  18.340000 30.665000  19.485000 ;
      RECT 24.865000  19.485000 32.625000  25.085000 ;
      RECT 24.865000  25.085000 32.625000  25.675000 ;
      RECT 24.880000  18.090000 30.525000  18.160000 ;
      RECT 24.880000  18.090000 30.525000  18.160000 ;
      RECT 24.895000  43.425000 73.380000  43.495000 ;
      RECT 24.895000  43.425000 73.380000  43.495000 ;
      RECT 24.950000  18.160000 30.525000  18.230000 ;
      RECT 24.950000  18.160000 30.525000  18.230000 ;
      RECT 24.965000  43.355000 73.380000  43.425000 ;
      RECT 24.965000  43.355000 73.380000  43.425000 ;
      RECT 25.005000  16.900000 30.525000  25.030000 ;
      RECT 25.005000  18.230000 30.525000  18.285000 ;
      RECT 25.005000  18.230000 30.525000  18.285000 ;
      RECT 25.005000  18.285000 30.525000  19.625000 ;
      RECT 25.005000  19.625000 32.485000  25.030000 ;
      RECT 25.035000  43.285000 73.380000  43.355000 ;
      RECT 25.035000  43.285000 73.380000  43.355000 ;
      RECT 25.075000  25.030000 32.485000  25.100000 ;
      RECT 25.075000  25.030000 32.485000  25.100000 ;
      RECT 25.105000  43.215000 73.380000  43.285000 ;
      RECT 25.105000  43.215000 73.380000  43.285000 ;
      RECT 25.145000  25.100000 32.485000  25.170000 ;
      RECT 25.145000  25.100000 32.485000  25.170000 ;
      RECT 25.175000  43.145000 73.380000  43.215000 ;
      RECT 25.175000  43.145000 73.380000  43.215000 ;
      RECT 25.215000  25.170000 32.485000  25.240000 ;
      RECT 25.215000  25.170000 32.485000  25.240000 ;
      RECT 25.245000  43.075000 73.380000  43.145000 ;
      RECT 25.245000  43.075000 73.380000  43.145000 ;
      RECT 25.275000   0.000000 27.440000   3.180000 ;
      RECT 25.275000   3.180000 28.045000   3.785000 ;
      RECT 25.275000   3.785000 28.045000   4.245000 ;
      RECT 25.275000   4.245000 29.310000   4.755000 ;
      RECT 25.275000   4.755000 28.045000   5.685000 ;
      RECT 25.275000   5.685000 32.620000   8.890000 ;
      RECT 25.275000   8.890000 32.625000   8.895000 ;
      RECT 25.275000   8.895000 32.625000  12.415000 ;
      RECT 25.275000  12.415000 32.625000  12.665000 ;
      RECT 25.285000  25.240000 32.485000  25.310000 ;
      RECT 25.285000  25.240000 32.485000  25.310000 ;
      RECT 25.315000  43.005000 73.380000  43.075000 ;
      RECT 25.315000  43.005000 73.380000  43.075000 ;
      RECT 25.355000  25.310000 32.485000  25.380000 ;
      RECT 25.355000  25.310000 32.485000  25.380000 ;
      RECT 25.385000  42.935000 73.380000  43.005000 ;
      RECT 25.385000  42.935000 73.380000  43.005000 ;
      RECT 25.415000   3.515000 27.575000   3.585000 ;
      RECT 25.415000   3.585000 27.645000   3.655000 ;
      RECT 25.415000   3.655000 27.715000   3.725000 ;
      RECT 25.415000   3.725000 27.785000   3.795000 ;
      RECT 25.415000   3.795000 27.855000   3.845000 ;
      RECT 25.415000   3.845000 27.905000   4.385000 ;
      RECT 25.415000   4.385000 29.415000   4.455000 ;
      RECT 25.415000   4.455000 29.345000   4.525000 ;
      RECT 25.415000   4.525000 29.275000   4.595000 ;
      RECT 25.415000   4.595000 29.255000   4.615000 ;
      RECT 25.415000   4.615000 27.905000   5.825000 ;
      RECT 25.415000   5.825000 31.165000   6.800000 ;
      RECT 25.415000   5.825000 31.165000   8.950000 ;
      RECT 25.415000   5.825000 31.165000   8.950000 ;
      RECT 25.415000   5.825000 31.165000   8.950000 ;
      RECT 25.415000   6.800000 32.480000   8.945000 ;
      RECT 25.415000   8.945000 32.480000   8.950000 ;
      RECT 25.415000   8.945000 32.480000   8.950000 ;
      RECT 25.415000   8.950000 32.485000  12.360000 ;
      RECT 25.425000  25.380000 32.485000  25.450000 ;
      RECT 25.425000  25.380000 32.485000  25.450000 ;
      RECT 25.455000  25.675000 32.625000  28.070000 ;
      RECT 25.455000  28.070000 32.485000  28.210000 ;
      RECT 25.455000  28.210000 28.495000  28.480000 ;
      RECT 25.455000  28.480000 28.495000  32.575000 ;
      RECT 25.455000  32.575000 75.000000  42.670000 ;
      RECT 25.455000  42.670000 75.000000  43.685000 ;
      RECT 25.455000  42.865000 73.380000  42.935000 ;
      RECT 25.455000  42.865000 73.380000  42.935000 ;
      RECT 25.485000  12.360000 32.485000  12.430000 ;
      RECT 25.485000  12.360000 32.485000  12.430000 ;
      RECT 25.495000  25.450000 32.485000  25.520000 ;
      RECT 25.495000  25.450000 32.485000  25.520000 ;
      RECT 25.525000  12.665000 32.625000  14.975000 ;
      RECT 25.525000  14.975000 32.625000  15.475000 ;
      RECT 25.525000  42.795000 73.380000  42.865000 ;
      RECT 25.525000  42.795000 73.380000  42.865000 ;
      RECT 25.555000  12.430000 32.485000  12.500000 ;
      RECT 25.555000  12.430000 32.485000  12.500000 ;
      RECT 25.560000   0.185000 27.265000   3.235000 ;
      RECT 25.565000  25.520000 32.485000  25.590000 ;
      RECT 25.565000  25.520000 32.485000  25.590000 ;
      RECT 25.595000  25.590000 32.485000  25.620000 ;
      RECT 25.595000  25.590000 32.485000  25.620000 ;
      RECT 25.595000  25.620000 32.485000  28.015000 ;
      RECT 25.595000  28.015000 32.460000  28.040000 ;
      RECT 25.595000  28.015000 32.460000  28.040000 ;
      RECT 25.595000  28.040000 32.430000  28.070000 ;
      RECT 25.595000  28.040000 32.430000  28.070000 ;
      RECT 25.595000  28.070000 28.640000  28.140000 ;
      RECT 25.595000  28.070000 28.640000  28.140000 ;
      RECT 25.595000  28.140000 28.570000  28.210000 ;
      RECT 25.595000  28.140000 28.570000  28.210000 ;
      RECT 25.595000  28.210000 28.500000  28.280000 ;
      RECT 25.595000  28.210000 28.500000  28.280000 ;
      RECT 25.595000  28.280000 28.430000  28.350000 ;
      RECT 25.595000  28.280000 28.430000  28.350000 ;
      RECT 25.595000  28.350000 28.360000  28.420000 ;
      RECT 25.595000  28.350000 28.360000  28.420000 ;
      RECT 25.595000  28.420000 28.355000  28.425000 ;
      RECT 25.595000  28.420000 28.355000  28.425000 ;
      RECT 25.595000  28.425000 28.355000  32.715000 ;
      RECT 25.595000  32.715000 73.380000  42.725000 ;
      RECT 25.595000  42.725000 73.380000  42.795000 ;
      RECT 25.595000  42.725000 73.380000  42.795000 ;
      RECT 25.625000  12.500000 32.485000  12.570000 ;
      RECT 25.625000  12.500000 32.485000  12.570000 ;
      RECT 25.665000  12.570000 32.485000  12.610000 ;
      RECT 25.665000  12.570000 32.485000  12.610000 ;
      RECT 25.665000  12.610000 32.485000  14.920000 ;
      RECT 25.735000  14.920000 32.485000  14.990000 ;
      RECT 25.735000  14.920000 32.485000  14.990000 ;
      RECT 25.805000  14.990000 32.485000  15.060000 ;
      RECT 25.805000  14.990000 32.485000  15.060000 ;
      RECT 25.875000  15.060000 32.485000  15.130000 ;
      RECT 25.875000  15.060000 32.485000  15.130000 ;
      RECT 25.945000  15.130000 32.485000  15.200000 ;
      RECT 25.945000  15.130000 32.485000  15.200000 ;
      RECT 26.015000  15.200000 32.485000  15.270000 ;
      RECT 26.015000  15.200000 32.485000  15.270000 ;
      RECT 26.080000  15.270000 32.485000  15.335000 ;
      RECT 26.080000  15.270000 32.485000  15.335000 ;
      RECT 28.370000   0.000000 30.365000   2.795000 ;
      RECT 28.370000   2.795000 30.365000   3.400000 ;
      RECT 28.500000   0.185000 30.205000   2.395000 ;
      RECT 28.515000   2.675000 30.225000   2.745000 ;
      RECT 28.585000   2.745000 30.225000   2.815000 ;
      RECT 28.655000   2.815000 30.225000   2.885000 ;
      RECT 28.725000   2.885000 30.225000   2.955000 ;
      RECT 28.795000   2.955000 30.225000   3.025000 ;
      RECT 28.865000   3.025000 30.225000   3.095000 ;
      RECT 28.935000   3.095000 30.225000   3.165000 ;
      RECT 28.975000   3.400000 30.365000   3.700000 ;
      RECT 28.975000   3.700000 29.820000   4.245000 ;
      RECT 29.005000   3.165000 30.225000   3.235000 ;
      RECT 29.005000  28.790000 75.000000  32.575000 ;
      RECT 29.075000   3.235000 30.225000   3.305000 ;
      RECT 29.080000  28.720000 75.000000  28.790000 ;
      RECT 29.115000   3.305000 30.225000   3.345000 ;
      RECT 29.115000   3.345000 30.225000   3.645000 ;
      RECT 29.115000   3.645000 30.155000   3.715000 ;
      RECT 29.115000   3.715000 30.085000   3.785000 ;
      RECT 29.115000   3.785000 30.015000   3.855000 ;
      RECT 29.115000   3.855000 29.945000   3.925000 ;
      RECT 29.115000   3.925000 29.875000   3.995000 ;
      RECT 29.115000   3.995000 29.805000   4.065000 ;
      RECT 29.115000   4.065000 29.735000   4.135000 ;
      RECT 29.115000   4.135000 29.665000   4.205000 ;
      RECT 29.115000   4.205000 29.595000   4.275000 ;
      RECT 29.115000   4.275000 29.525000   4.345000 ;
      RECT 29.115000   4.345000 29.485000   4.385000 ;
      RECT 29.145000  28.860000 73.380000  32.715000 ;
      RECT 29.765000   5.815000 31.165000   5.825000 ;
      RECT 29.835000   5.745000 31.165000   5.815000 ;
      RECT 29.905000   5.675000 31.165000   5.745000 ;
      RECT 29.975000   5.605000 31.165000   5.675000 ;
      RECT 30.025000  15.475000 32.625000  16.625000 ;
      RECT 30.045000   5.535000 31.165000   5.605000 ;
      RECT 30.115000   5.465000 31.165000   5.535000 ;
      RECT 30.150000  15.335000 32.485000  15.405000 ;
      RECT 30.150000  15.335000 32.485000  15.405000 ;
      RECT 30.185000   5.395000 31.165000   5.465000 ;
      RECT 30.220000  15.405000 32.485000  15.475000 ;
      RECT 30.220000  15.405000 32.485000  15.475000 ;
      RECT 30.255000   5.325000 31.165000   5.395000 ;
      RECT 30.290000  15.475000 32.485000  15.545000 ;
      RECT 30.290000  15.475000 32.485000  15.545000 ;
      RECT 30.325000   5.255000 31.165000   5.325000 ;
      RECT 30.360000  15.545000 32.485000  15.615000 ;
      RECT 30.360000  15.545000 32.485000  15.615000 ;
      RECT 30.395000   5.185000 31.165000   5.255000 ;
      RECT 30.430000  15.615000 32.485000  15.685000 ;
      RECT 30.430000  15.615000 32.485000  15.685000 ;
      RECT 30.435000  80.155000 73.380000  84.520000 ;
      RECT 30.435000  84.520000 33.105000  84.755000 ;
      RECT 30.465000   5.115000 31.165000   5.185000 ;
      RECT 30.500000  15.685000 32.485000  15.755000 ;
      RECT 30.500000  15.685000 32.485000  15.755000 ;
      RECT 30.535000   5.045000 31.165000   5.115000 ;
      RECT 30.570000  15.755000 32.485000  15.825000 ;
      RECT 30.570000  15.755000 32.485000  15.825000 ;
      RECT 30.605000   4.975000 31.165000   5.045000 ;
      RECT 30.640000  15.825000 32.485000  15.895000 ;
      RECT 30.640000  15.825000 32.485000  15.895000 ;
      RECT 30.675000   4.905000 31.165000   4.975000 ;
      RECT 30.710000  15.895000 32.485000  15.965000 ;
      RECT 30.710000  15.895000 32.485000  15.965000 ;
      RECT 30.745000   4.835000 31.165000   4.905000 ;
      RECT 30.780000  15.965000 32.485000  16.035000 ;
      RECT 30.780000  15.965000 32.485000  16.035000 ;
      RECT 30.815000   4.765000 31.165000   4.835000 ;
      RECT 30.850000  16.035000 32.485000  16.105000 ;
      RECT 30.850000  16.035000 32.485000  16.105000 ;
      RECT 30.885000   4.695000 31.165000   4.765000 ;
      RECT 30.920000  16.105000 32.485000  16.175000 ;
      RECT 30.920000  16.105000 32.485000  16.175000 ;
      RECT 30.955000   4.625000 31.165000   4.695000 ;
      RECT 30.990000  16.175000 32.485000  16.245000 ;
      RECT 30.990000  16.175000 32.485000  16.245000 ;
      RECT 31.025000   4.555000 31.165000   4.625000 ;
      RECT 31.060000  16.245000 32.485000  16.315000 ;
      RECT 31.060000  16.245000 32.485000  16.315000 ;
      RECT 31.095000   4.485000 31.165000   4.555000 ;
      RECT 31.130000  16.315000 32.485000  16.385000 ;
      RECT 31.130000  16.315000 32.485000  16.385000 ;
      RECT 31.175000  16.625000 32.625000  19.485000 ;
      RECT 31.200000  16.385000 32.485000  16.455000 ;
      RECT 31.200000  16.385000 32.485000  16.455000 ;
      RECT 31.270000  16.455000 32.485000  16.525000 ;
      RECT 31.270000  16.455000 32.485000  16.525000 ;
      RECT 31.295000   0.000000 32.620000   4.090000 ;
      RECT 31.295000   4.090000 32.620000   5.685000 ;
      RECT 31.315000  16.525000 32.485000  16.570000 ;
      RECT 31.315000  16.525000 32.485000  16.570000 ;
      RECT 31.315000  16.570000 32.485000  19.625000 ;
      RECT 31.435000   0.000000 32.480000   0.390000 ;
      RECT 31.445000   0.670000 32.410000   6.520000 ;
      RECT 33.160000   0.000000 75.000000   8.660000 ;
      RECT 33.160000   8.660000 75.000000   8.665000 ;
      RECT 33.165000   8.665000 75.000000  28.720000 ;
      RECT 33.300000   0.000000 75.000000   0.600000 ;
      RECT 33.300000   0.600000 34.820000   0.620000 ;
      RECT 33.300000   0.620000 34.615000   2.160000 ;
      RECT 33.300000   2.160000 39.940000   6.270000 ;
      RECT 33.300000   6.270000 73.110000   6.340000 ;
      RECT 33.300000   6.270000 73.110000   6.340000 ;
      RECT 33.300000   6.340000 73.180000   6.410000 ;
      RECT 33.300000   6.340000 73.180000   6.410000 ;
      RECT 33.300000   6.410000 73.250000   6.480000 ;
      RECT 33.300000   6.410000 73.250000   6.480000 ;
      RECT 33.300000   6.480000 73.320000   6.540000 ;
      RECT 33.300000   6.480000 73.320000   6.540000 ;
      RECT 33.300000   6.540000 73.380000   8.605000 ;
      RECT 33.305000   8.605000 73.380000   8.610000 ;
      RECT 33.305000   8.605000 73.380000   8.610000 ;
      RECT 33.305000   8.610000 73.380000  28.860000 ;
      RECT 33.305000   8.610000 73.380000  32.715000 ;
      RECT 33.385000  84.800000 74.700000  85.055000 ;
      RECT 34.895000   0.900000 38.965000   1.880000 ;
      RECT 35.100000   0.880000 38.920000   0.900000 ;
      RECT 39.200000   0.600000 75.000000   0.620000 ;
      RECT 39.245000   0.620000 75.000000   0.740000 ;
      RECT 39.245000   0.740000 39.940000   2.160000 ;
      RECT 40.220000   1.020000 74.590000   5.990000 ;
      RECT 56.545000 100.330000 72.090000 101.420000 ;
      RECT 56.725000  97.530000 72.090000  97.760000 ;
      RECT 56.825000  98.040000 71.245000  98.110000 ;
      RECT 56.825000  98.110000 71.315000  98.180000 ;
      RECT 56.825000  98.180000 71.385000  98.250000 ;
      RECT 56.825000  98.250000 71.455000  98.320000 ;
      RECT 56.825000  98.320000 71.525000  98.390000 ;
      RECT 56.825000  98.390000 71.595000  98.460000 ;
      RECT 56.825000  98.460000 71.665000  98.530000 ;
      RECT 56.825000  98.530000 71.735000  98.600000 ;
      RECT 56.825000  98.600000 71.805000  98.605000 ;
      RECT 56.825000  98.605000 71.810000  99.405000 ;
      RECT 56.825000  99.405000 71.740000  99.475000 ;
      RECT 56.825000  99.475000 71.670000  99.545000 ;
      RECT 56.825000  99.545000 71.600000  99.615000 ;
      RECT 56.825000  99.615000 71.530000  99.685000 ;
      RECT 56.825000  99.685000 71.460000  99.755000 ;
      RECT 56.825000  99.755000 71.390000  99.825000 ;
      RECT 56.825000  99.825000 71.320000  99.895000 ;
      RECT 56.825000  99.895000 71.250000  99.965000 ;
      RECT 56.825000  99.965000 71.180000 100.035000 ;
      RECT 56.825000 100.035000 71.165000 100.050000 ;
      RECT 59.500000 199.490000 64.600000 200.000000 ;
      RECT 59.780000 196.250000 64.320000 199.210000 ;
      RECT 60.320000 125.440000 75.145000 125.510000 ;
      RECT 60.320000 125.440000 75.145000 125.510000 ;
      RECT 60.390000 125.510000 75.145000 125.580000 ;
      RECT 60.390000 125.510000 75.145000 125.580000 ;
      RECT 60.460000 125.580000 75.145000 125.650000 ;
      RECT 60.460000 125.580000 75.145000 125.650000 ;
      RECT 60.530000 125.650000 75.145000 125.720000 ;
      RECT 60.530000 125.650000 75.145000 125.720000 ;
      RECT 60.600000 125.720000 75.145000 125.790000 ;
      RECT 60.600000 125.720000 75.145000 125.790000 ;
      RECT 60.670000 125.790000 75.145000 125.860000 ;
      RECT 60.670000 125.790000 75.145000 125.860000 ;
      RECT 60.740000 125.860000 75.145000 125.930000 ;
      RECT 60.740000 125.860000 75.145000 125.930000 ;
      RECT 60.810000 125.930000 75.145000 126.000000 ;
      RECT 60.810000 125.930000 75.145000 126.000000 ;
      RECT 60.880000 126.000000 75.145000 126.070000 ;
      RECT 60.880000 126.000000 75.145000 126.070000 ;
      RECT 60.950000 126.070000 75.145000 126.140000 ;
      RECT 60.950000 126.070000 75.145000 126.140000 ;
      RECT 61.020000 126.140000 75.145000 126.210000 ;
      RECT 61.020000 126.140000 75.145000 126.210000 ;
      RECT 61.090000 126.210000 75.145000 126.280000 ;
      RECT 61.090000 126.210000 75.145000 126.280000 ;
      RECT 61.160000 126.280000 75.145000 126.350000 ;
      RECT 61.160000 126.280000 75.145000 126.350000 ;
      RECT 61.230000 126.350000 75.145000 126.420000 ;
      RECT 61.230000 126.350000 75.145000 126.420000 ;
      RECT 61.300000 126.420000 75.145000 126.490000 ;
      RECT 61.300000 126.420000 75.145000 126.490000 ;
      RECT 61.370000 126.490000 75.145000 126.560000 ;
      RECT 61.370000 126.490000 75.145000 126.560000 ;
      RECT 61.440000 126.560000 75.145000 126.630000 ;
      RECT 61.440000 126.560000 75.145000 126.630000 ;
      RECT 61.510000 126.630000 75.145000 126.700000 ;
      RECT 61.510000 126.630000 75.145000 126.700000 ;
      RECT 61.580000 126.700000 75.145000 126.770000 ;
      RECT 61.580000 126.700000 75.145000 126.770000 ;
      RECT 61.650000 126.770000 75.145000 126.840000 ;
      RECT 61.650000 126.770000 75.145000 126.840000 ;
      RECT 61.720000 126.840000 75.145000 126.910000 ;
      RECT 61.720000 126.840000 75.145000 126.910000 ;
      RECT 61.790000 126.910000 75.145000 126.980000 ;
      RECT 61.790000 126.910000 75.145000 126.980000 ;
      RECT 61.860000 126.980000 75.145000 127.050000 ;
      RECT 61.860000 126.980000 75.145000 127.050000 ;
      RECT 61.930000 127.050000 75.145000 127.120000 ;
      RECT 61.930000 127.050000 75.145000 127.120000 ;
      RECT 62.000000 127.120000 75.145000 127.190000 ;
      RECT 62.000000 127.120000 75.145000 127.190000 ;
      RECT 62.070000 127.190000 75.145000 127.260000 ;
      RECT 62.070000 127.190000 75.145000 127.260000 ;
      RECT 62.140000 127.260000 75.145000 127.330000 ;
      RECT 62.140000 127.260000 75.145000 127.330000 ;
      RECT 62.210000 127.330000 75.145000 127.400000 ;
      RECT 62.210000 127.330000 75.145000 127.400000 ;
      RECT 62.280000 127.400000 75.145000 127.470000 ;
      RECT 62.280000 127.400000 75.145000 127.470000 ;
      RECT 62.350000 127.470000 75.145000 127.540000 ;
      RECT 62.350000 127.470000 75.145000 127.540000 ;
      RECT 62.420000 127.540000 75.145000 127.610000 ;
      RECT 62.420000 127.540000 75.145000 127.610000 ;
      RECT 62.490000 127.610000 75.145000 127.680000 ;
      RECT 62.490000 127.610000 75.145000 127.680000 ;
      RECT 62.560000 127.680000 75.145000 127.750000 ;
      RECT 62.560000 127.680000 75.145000 127.750000 ;
      RECT 62.630000 127.750000 75.145000 127.820000 ;
      RECT 62.630000 127.750000 75.145000 127.820000 ;
      RECT 62.700000 127.820000 75.145000 127.890000 ;
      RECT 62.700000 127.820000 75.145000 127.890000 ;
      RECT 62.770000 127.890000 75.145000 127.960000 ;
      RECT 62.770000 127.890000 75.145000 127.960000 ;
      RECT 62.840000 127.960000 75.145000 128.030000 ;
      RECT 62.840000 127.960000 75.145000 128.030000 ;
      RECT 62.910000 128.030000 75.145000 128.100000 ;
      RECT 62.910000 128.030000 75.145000 128.100000 ;
      RECT 62.980000 128.100000 75.145000 128.170000 ;
      RECT 62.980000 128.100000 75.145000 128.170000 ;
      RECT 63.050000 128.170000 75.145000 128.240000 ;
      RECT 63.050000 128.170000 75.145000 128.240000 ;
      RECT 63.070000 128.240000 75.145000 128.260000 ;
      RECT 63.070000 128.240000 75.145000 128.260000 ;
      RECT 63.140000 128.260000 75.145000 128.330000 ;
      RECT 63.140000 128.260000 75.145000 128.330000 ;
      RECT 63.210000 128.330000 75.145000 128.400000 ;
      RECT 63.210000 128.330000 75.145000 128.400000 ;
      RECT 63.280000 128.400000 75.145000 128.470000 ;
      RECT 63.280000 128.400000 75.145000 128.470000 ;
      RECT 63.350000 128.470000 75.145000 128.540000 ;
      RECT 63.350000 128.470000 75.145000 128.540000 ;
      RECT 63.420000 128.540000 75.145000 128.610000 ;
      RECT 63.420000 128.540000 75.145000 128.610000 ;
      RECT 63.490000 128.610000 75.145000 128.680000 ;
      RECT 63.490000 128.610000 75.145000 128.680000 ;
      RECT 63.560000 128.680000 75.145000 128.750000 ;
      RECT 63.560000 128.680000 75.145000 128.750000 ;
      RECT 63.630000 128.750000 75.145000 128.820000 ;
      RECT 63.630000 128.750000 75.145000 128.820000 ;
      RECT 63.700000 128.820000 75.145000 128.890000 ;
      RECT 63.700000 128.820000 75.145000 128.890000 ;
      RECT 63.770000 128.890000 75.145000 128.960000 ;
      RECT 63.770000 128.890000 75.145000 128.960000 ;
      RECT 63.840000 128.960000 75.145000 129.030000 ;
      RECT 63.840000 128.960000 75.145000 129.030000 ;
      RECT 63.910000 129.030000 75.145000 129.100000 ;
      RECT 63.910000 129.030000 75.145000 129.100000 ;
      RECT 63.980000 129.100000 75.145000 129.170000 ;
      RECT 63.980000 129.100000 75.145000 129.170000 ;
      RECT 64.050000 129.170000 75.145000 129.240000 ;
      RECT 64.050000 129.170000 75.145000 129.240000 ;
      RECT 64.120000 129.240000 75.145000 129.310000 ;
      RECT 64.120000 129.240000 75.145000 129.310000 ;
      RECT 64.190000 129.310000 75.145000 129.380000 ;
      RECT 64.190000 129.310000 75.145000 129.380000 ;
      RECT 64.260000 129.380000 75.145000 129.450000 ;
      RECT 64.260000 129.380000 75.145000 129.450000 ;
      RECT 64.330000 129.450000 75.145000 129.520000 ;
      RECT 64.330000 129.450000 75.145000 129.520000 ;
      RECT 64.400000 129.520000 75.145000 129.590000 ;
      RECT 64.400000 129.520000 75.145000 129.590000 ;
      RECT 64.470000 129.590000 75.145000 129.660000 ;
      RECT 64.470000 129.590000 75.145000 129.660000 ;
      RECT 64.540000 129.660000 75.145000 129.730000 ;
      RECT 64.540000 129.660000 75.145000 129.730000 ;
      RECT 64.600000 175.420000 75.000000 200.000000 ;
      RECT 64.600000 195.970000 75.000000 199.490000 ;
      RECT 64.600000 199.490000 75.000000 200.000000 ;
      RECT 64.610000 129.730000 75.145000 129.800000 ;
      RECT 64.610000 129.730000 75.145000 129.800000 ;
      RECT 64.680000 129.800000 75.145000 129.870000 ;
      RECT 64.680000 129.800000 75.145000 129.870000 ;
      RECT 64.750000 129.870000 75.145000 129.940000 ;
      RECT 64.750000 129.870000 75.145000 129.940000 ;
      RECT 64.820000 129.940000 75.145000 130.010000 ;
      RECT 64.820000 129.940000 75.145000 130.010000 ;
      RECT 64.890000 130.010000 75.145000 130.080000 ;
      RECT 64.890000 130.010000 75.145000 130.080000 ;
      RECT 64.960000 130.080000 75.145000 130.150000 ;
      RECT 64.960000 130.080000 75.145000 130.150000 ;
      RECT 65.030000 130.150000 75.145000 130.220000 ;
      RECT 65.030000 130.150000 75.145000 130.220000 ;
      RECT 69.105000 138.955000 75.145000 138.960000 ;
      RECT 69.105000 138.955000 75.145000 138.960000 ;
      RECT 69.110000 138.950000 75.145000 138.955000 ;
      RECT 69.110000 138.950000 75.145000 138.955000 ;
      RECT 69.115000 138.945000 75.145000 138.950000 ;
      RECT 69.115000 138.945000 75.145000 138.950000 ;
      RECT 69.115000 138.960000 75.145000 138.975000 ;
      RECT 69.115000 138.960000 75.145000 138.975000 ;
      RECT 69.130000 138.975000 75.145000 138.990000 ;
      RECT 69.130000 138.975000 75.145000 138.990000 ;
      RECT 69.160000 138.900000 75.145000 138.945000 ;
      RECT 69.160000 138.900000 75.145000 138.945000 ;
      RECT 69.200000 138.990000 75.145000 139.060000 ;
      RECT 69.200000 138.990000 75.145000 139.060000 ;
      RECT 69.230000 138.830000 75.145000 138.900000 ;
      RECT 69.230000 138.830000 75.145000 138.900000 ;
      RECT 69.270000 139.060000 75.145000 139.130000 ;
      RECT 69.270000 139.060000 75.145000 139.130000 ;
      RECT 69.300000 138.760000 75.145000 138.830000 ;
      RECT 69.300000 138.760000 75.145000 138.830000 ;
      RECT 69.340000 139.130000 75.145000 139.200000 ;
      RECT 69.340000 139.130000 75.145000 139.200000 ;
      RECT 69.370000 138.690000 75.145000 138.760000 ;
      RECT 69.370000 138.690000 75.145000 138.760000 ;
      RECT 69.410000 139.200000 75.145000 139.270000 ;
      RECT 69.410000 139.200000 75.145000 139.270000 ;
      RECT 69.440000 138.620000 75.145000 138.690000 ;
      RECT 69.440000 138.620000 75.145000 138.690000 ;
      RECT 69.480000 139.270000 75.145000 139.340000 ;
      RECT 69.480000 139.270000 75.145000 139.340000 ;
      RECT 69.510000 138.550000 75.145000 138.620000 ;
      RECT 69.510000 138.550000 75.145000 138.620000 ;
      RECT 69.550000 139.340000 75.145000 139.410000 ;
      RECT 69.550000 139.340000 75.145000 139.410000 ;
      RECT 69.580000 138.480000 75.145000 138.550000 ;
      RECT 69.580000 138.480000 75.145000 138.550000 ;
      RECT 69.620000 139.410000 75.145000 139.480000 ;
      RECT 69.620000 139.410000 75.145000 139.480000 ;
      RECT 69.650000 138.410000 75.145000 138.480000 ;
      RECT 69.650000 138.410000 75.145000 138.480000 ;
      RECT 69.690000 139.480000 75.145000 139.550000 ;
      RECT 69.690000 139.480000 75.145000 139.550000 ;
      RECT 69.715000 139.550000 75.145000 139.575000 ;
      RECT 69.715000 139.550000 75.145000 139.575000 ;
      RECT 69.720000 138.340000 75.145000 138.410000 ;
      RECT 69.720000 138.340000 75.145000 138.410000 ;
      RECT 69.785000 139.575000 75.145000 139.645000 ;
      RECT 69.785000 139.575000 75.145000 139.645000 ;
      RECT 69.790000 138.270000 75.145000 138.340000 ;
      RECT 69.790000 138.270000 75.145000 138.340000 ;
      RECT 69.855000 139.645000 75.145000 139.715000 ;
      RECT 69.855000 139.645000 75.145000 139.715000 ;
      RECT 69.860000 138.200000 75.145000 138.270000 ;
      RECT 69.860000 138.200000 75.145000 138.270000 ;
      RECT 69.925000 139.715000 75.145000 139.785000 ;
      RECT 69.925000 139.715000 75.145000 139.785000 ;
      RECT 69.925000 141.095000 70.525000 143.875000 ;
      RECT 69.930000 138.130000 75.145000 138.200000 ;
      RECT 69.930000 138.130000 75.145000 138.200000 ;
      RECT 69.990000 139.785000 75.145000 139.850000 ;
      RECT 69.990000 139.785000 75.145000 139.850000 ;
      RECT 70.000000 138.060000 75.145000 138.130000 ;
      RECT 70.000000 138.060000 75.145000 138.130000 ;
      RECT 70.060000 139.850000 75.145000 139.920000 ;
      RECT 70.060000 139.850000 75.145000 139.920000 ;
      RECT 70.070000 137.990000 75.145000 138.060000 ;
      RECT 70.070000 137.990000 75.145000 138.060000 ;
      RECT 70.105000 145.100000 75.145000 145.130000 ;
      RECT 70.130000 139.920000 75.145000 139.990000 ;
      RECT 70.130000 139.920000 75.145000 139.990000 ;
      RECT 70.140000 137.920000 75.145000 137.990000 ;
      RECT 70.140000 137.920000 75.145000 137.990000 ;
      RECT 70.175000 145.030000 75.145000 145.100000 ;
      RECT 70.200000 139.990000 75.145000 140.060000 ;
      RECT 70.200000 139.990000 75.145000 140.060000 ;
      RECT 70.210000 137.850000 75.145000 137.920000 ;
      RECT 70.210000 137.850000 75.145000 137.920000 ;
      RECT 70.245000 144.960000 75.145000 145.030000 ;
      RECT 70.270000 140.060000 75.145000 140.130000 ;
      RECT 70.270000 140.060000 75.145000 140.130000 ;
      RECT 70.280000 137.780000 75.145000 137.850000 ;
      RECT 70.280000 137.780000 75.145000 137.850000 ;
      RECT 70.315000 144.890000 75.145000 144.960000 ;
      RECT 70.340000 140.130000 75.145000 140.200000 ;
      RECT 70.340000 140.130000 75.145000 140.200000 ;
      RECT 70.350000 137.710000 75.145000 137.780000 ;
      RECT 70.350000 137.710000 75.145000 137.780000 ;
      RECT 70.385000 144.820000 75.145000 144.890000 ;
      RECT 70.410000 140.200000 75.145000 140.270000 ;
      RECT 70.410000 140.200000 75.145000 140.270000 ;
      RECT 70.420000 137.640000 75.145000 137.710000 ;
      RECT 70.420000 137.640000 75.145000 137.710000 ;
      RECT 70.455000 144.750000 75.145000 144.820000 ;
      RECT 70.480000 140.270000 75.145000 140.340000 ;
      RECT 70.480000 140.270000 75.145000 140.340000 ;
      RECT 70.490000 137.570000 75.145000 137.640000 ;
      RECT 70.490000 137.570000 75.145000 137.640000 ;
      RECT 70.525000 144.680000 75.145000 144.750000 ;
      RECT 70.550000 140.340000 75.145000 140.410000 ;
      RECT 70.550000 140.340000 75.145000 140.410000 ;
      RECT 70.560000 137.500000 75.145000 137.570000 ;
      RECT 70.560000 137.500000 75.145000 137.570000 ;
      RECT 70.595000 144.610000 75.145000 144.680000 ;
      RECT 70.620000 140.410000 75.145000 140.480000 ;
      RECT 70.620000 140.410000 75.145000 140.480000 ;
      RECT 70.630000 137.430000 75.145000 137.500000 ;
      RECT 70.630000 137.430000 75.145000 137.500000 ;
      RECT 70.665000 144.540000 75.145000 144.610000 ;
      RECT 70.690000 140.480000 75.145000 140.550000 ;
      RECT 70.690000 140.480000 75.145000 140.550000 ;
      RECT 70.700000 137.360000 75.145000 137.430000 ;
      RECT 70.700000 137.360000 75.145000 137.430000 ;
      RECT 70.735000 144.470000 75.145000 144.540000 ;
      RECT 70.760000 140.550000 75.145000 140.620000 ;
      RECT 70.760000 140.550000 75.145000 140.620000 ;
      RECT 70.770000 137.290000 75.145000 137.360000 ;
      RECT 70.770000 137.290000 75.145000 137.360000 ;
      RECT 70.805000 139.850000 75.145000 145.130000 ;
      RECT 70.805000 140.620000 75.145000 140.665000 ;
      RECT 70.805000 140.620000 75.145000 140.665000 ;
      RECT 70.805000 140.665000 75.145000 144.400000 ;
      RECT 70.805000 144.400000 75.145000 144.470000 ;
      RECT 70.805000 144.400000 75.145000 145.130000 ;
      RECT 70.805000 145.130000 73.195000 146.145000 ;
      RECT 70.840000 137.220000 75.145000 137.290000 ;
      RECT 70.840000 137.220000 75.145000 137.290000 ;
      RECT 70.910000 137.150000 75.145000 137.220000 ;
      RECT 70.910000 137.150000 75.145000 137.220000 ;
      RECT 70.980000 137.080000 75.145000 137.150000 ;
      RECT 70.980000 137.080000 75.145000 137.150000 ;
      RECT 71.050000 137.010000 75.145000 137.080000 ;
      RECT 71.050000 137.010000 75.145000 137.080000 ;
      RECT 71.120000 136.940000 75.145000 137.010000 ;
      RECT 71.120000 136.940000 75.145000 137.010000 ;
      RECT 71.190000 136.870000 75.145000 136.940000 ;
      RECT 71.190000 136.870000 75.145000 136.940000 ;
      RECT 71.260000 136.800000 75.145000 136.870000 ;
      RECT 71.260000 136.800000 75.145000 136.870000 ;
      RECT 71.320000 100.290000 75.145000 100.330000 ;
      RECT 71.330000 136.730000 75.145000 136.800000 ;
      RECT 71.330000 136.730000 75.145000 136.800000 ;
      RECT 71.390000 100.220000 75.145000 100.290000 ;
      RECT 71.400000 136.660000 75.145000 136.730000 ;
      RECT 71.400000 136.660000 75.145000 136.730000 ;
      RECT 71.430000  97.760000 75.145000  97.830000 ;
      RECT 71.460000 100.150000 75.145000 100.220000 ;
      RECT 71.470000 136.590000 75.145000 136.660000 ;
      RECT 71.470000 136.590000 75.145000 136.660000 ;
      RECT 71.500000  97.830000 75.145000  97.900000 ;
      RECT 71.530000 100.080000 75.145000 100.150000 ;
      RECT 71.540000 136.520000 75.145000 136.590000 ;
      RECT 71.540000 136.520000 75.145000 136.590000 ;
      RECT 71.570000  97.900000 75.145000  97.970000 ;
      RECT 71.600000 100.010000 75.145000 100.080000 ;
      RECT 71.610000 136.450000 75.145000 136.520000 ;
      RECT 71.610000 136.450000 75.145000 136.520000 ;
      RECT 71.640000  97.970000 75.145000  98.040000 ;
      RECT 71.670000  99.940000 75.145000 100.010000 ;
      RECT 71.680000 136.380000 75.145000 136.450000 ;
      RECT 71.680000 136.380000 75.145000 136.450000 ;
      RECT 71.710000  98.040000 75.145000  98.110000 ;
      RECT 71.740000  99.870000 75.145000  99.940000 ;
      RECT 71.750000 136.310000 75.145000 136.380000 ;
      RECT 71.750000 136.310000 75.145000 136.380000 ;
      RECT 71.755000  85.835000 74.700000  94.470000 ;
      RECT 71.780000  98.110000 75.145000  98.180000 ;
      RECT 71.810000  99.800000 75.145000  99.870000 ;
      RECT 71.820000 136.240000 75.145000 136.310000 ;
      RECT 71.820000 136.240000 75.145000 136.310000 ;
      RECT 71.850000  98.180000 75.145000  98.250000 ;
      RECT 71.880000  99.730000 75.145000  99.800000 ;
      RECT 71.890000 136.170000 75.145000 136.240000 ;
      RECT 71.890000 136.170000 75.145000 136.240000 ;
      RECT 71.920000  98.250000 75.145000  98.320000 ;
      RECT 71.950000  99.660000 75.145000  99.730000 ;
      RECT 71.960000 136.100000 75.145000 136.170000 ;
      RECT 71.960000 136.100000 75.145000 136.170000 ;
      RECT 71.990000  98.320000 75.145000  98.390000 ;
      RECT 72.020000  99.590000 75.145000  99.660000 ;
      RECT 72.030000 136.030000 75.145000 136.100000 ;
      RECT 72.030000 136.030000 75.145000 136.100000 ;
      RECT 72.060000  98.390000 75.145000  98.460000 ;
      RECT 72.090000  97.530000 75.145000 100.765000 ;
      RECT 72.090000  97.760000 75.145000  98.490000 ;
      RECT 72.090000  98.460000 75.145000  98.490000 ;
      RECT 72.090000  98.490000 75.145000  99.520000 ;
      RECT 72.090000  99.520000 75.145000  99.590000 ;
      RECT 72.090000  99.520000 75.145000 100.330000 ;
      RECT 72.090000 100.330000 75.145000 101.420000 ;
      RECT 72.100000 135.960000 75.145000 136.030000 ;
      RECT 72.100000 135.960000 75.145000 136.030000 ;
      RECT 72.115000  97.505000 75.145000  97.530000 ;
      RECT 72.170000 135.890000 75.145000 135.960000 ;
      RECT 72.170000 135.890000 75.145000 135.960000 ;
      RECT 72.185000  97.435000 75.145000  97.505000 ;
      RECT 72.240000 135.820000 75.145000 135.890000 ;
      RECT 72.240000 135.820000 75.145000 135.890000 ;
      RECT 72.255000  97.365000 75.145000  97.435000 ;
      RECT 72.310000 135.750000 75.145000 135.820000 ;
      RECT 72.310000 135.750000 75.145000 135.820000 ;
      RECT 72.325000  97.295000 75.145000  97.365000 ;
      RECT 72.380000 130.500000 75.000000 130.995000 ;
      RECT 72.380000 135.680000 75.145000 135.750000 ;
      RECT 72.380000 135.680000 75.145000 135.750000 ;
      RECT 72.395000  97.225000 75.145000  97.295000 ;
      RECT 72.450000 135.610000 75.145000 135.680000 ;
      RECT 72.450000 135.610000 75.145000 135.680000 ;
      RECT 72.465000  97.155000 75.145000  97.225000 ;
      RECT 72.520000 135.540000 75.145000 135.610000 ;
      RECT 72.520000 135.540000 75.145000 135.610000 ;
      RECT 72.535000  97.085000 75.145000  97.155000 ;
      RECT 72.590000 135.470000 75.145000 135.540000 ;
      RECT 72.590000 135.470000 75.145000 135.540000 ;
      RECT 72.605000  97.015000 75.145000  97.085000 ;
      RECT 72.660000 131.275000 75.145000 132.915000 ;
      RECT 72.660000 135.400000 75.145000 135.470000 ;
      RECT 72.660000 135.400000 75.145000 135.470000 ;
      RECT 72.675000  96.945000 75.145000  97.015000 ;
      RECT 72.695000 135.365000 75.145000 135.400000 ;
      RECT 72.695000 135.365000 75.145000 135.400000 ;
      RECT 72.745000  96.875000 75.145000  96.945000 ;
      RECT 72.765000 135.295000 75.145000 135.365000 ;
      RECT 72.765000 135.295000 75.145000 135.365000 ;
      RECT 72.815000  96.805000 75.145000  96.875000 ;
      RECT 72.835000 135.225000 75.145000 135.295000 ;
      RECT 72.835000 135.225000 75.145000 135.295000 ;
      RECT 72.885000  96.735000 75.145000  96.805000 ;
      RECT 72.905000 135.155000 75.145000 135.225000 ;
      RECT 72.905000 135.155000 75.145000 135.225000 ;
      RECT 72.955000  96.665000 75.145000  96.735000 ;
      RECT 72.975000 135.085000 75.145000 135.155000 ;
      RECT 72.975000 135.085000 75.145000 135.155000 ;
      RECT 73.025000  96.595000 75.145000  96.665000 ;
      RECT 73.045000 135.015000 75.145000 135.085000 ;
      RECT 73.045000 135.015000 75.145000 135.085000 ;
      RECT 73.095000  96.525000 75.145000  96.595000 ;
      RECT 73.115000 134.945000 75.145000 135.015000 ;
      RECT 73.115000 134.945000 75.145000 135.015000 ;
      RECT 73.165000  96.455000 75.145000  96.525000 ;
      RECT 73.185000 134.875000 75.145000 134.945000 ;
      RECT 73.185000 134.875000 75.145000 134.945000 ;
      RECT 73.235000  96.385000 75.145000  96.455000 ;
      RECT 73.255000 134.805000 75.145000 134.875000 ;
      RECT 73.255000 134.805000 75.145000 134.875000 ;
      RECT 73.295000   5.990000 74.590000   6.060000 ;
      RECT 73.305000  96.315000 75.145000  96.385000 ;
      RECT 73.325000 134.735000 75.145000 134.805000 ;
      RECT 73.325000 134.735000 75.145000 134.805000 ;
      RECT 73.365000   6.060000 74.590000   6.130000 ;
      RECT 73.375000  96.245000 75.145000  96.315000 ;
      RECT 73.395000 134.665000 75.145000 134.735000 ;
      RECT 73.395000 134.665000 75.145000 134.735000 ;
      RECT 73.435000   6.130000 74.590000   6.200000 ;
      RECT 73.445000  96.175000 75.145000  96.245000 ;
      RECT 73.465000 134.595000 75.145000 134.665000 ;
      RECT 73.465000 134.595000 75.145000 134.665000 ;
      RECT 73.475000 145.410000 75.000000 146.425000 ;
      RECT 73.505000   6.200000 74.590000   6.270000 ;
      RECT 73.515000  96.105000 75.145000  96.175000 ;
      RECT 73.535000 134.525000 75.145000 134.595000 ;
      RECT 73.535000 134.525000 75.145000 134.595000 ;
      RECT 73.575000   6.270000 74.590000   6.340000 ;
      RECT 73.585000  96.035000 75.145000  96.105000 ;
      RECT 73.605000 134.455000 75.145000 134.525000 ;
      RECT 73.605000 134.455000 75.145000 134.525000 ;
      RECT 73.645000   6.340000 74.590000   6.410000 ;
      RECT 73.655000  95.965000 75.145000  96.035000 ;
      RECT 73.660000   6.410000 74.590000   6.425000 ;
      RECT 73.660000   6.425000 74.590000  79.620000 ;
      RECT 73.660000  79.620000 74.590000  79.675000 ;
      RECT 73.660000  79.675000 74.645000  79.730000 ;
      RECT 73.660000  79.730000 74.700000  84.800000 ;
      RECT 73.675000 134.385000 75.145000 134.455000 ;
      RECT 73.675000 134.385000 75.145000 134.455000 ;
      RECT 73.685000 174.500000 74.745000 175.140000 ;
      RECT 73.725000  95.895000 75.145000  95.965000 ;
      RECT 73.725000  95.895000 75.145000 100.535000 ;
      RECT 73.745000 134.315000 75.145000 134.385000 ;
      RECT 73.745000 134.315000 75.145000 134.385000 ;
      RECT 73.770000 101.420000 74.700000 104.565000 ;
      RECT 73.815000 134.245000 75.145000 134.315000 ;
      RECT 73.815000 134.245000 75.145000 134.315000 ;
      RECT 73.885000 134.175000 75.145000 134.245000 ;
      RECT 73.885000 134.175000 75.145000 134.245000 ;
      RECT 73.955000 134.105000 75.145000 134.175000 ;
      RECT 73.955000 134.105000 75.145000 134.175000 ;
      RECT 74.025000 134.035000 75.145000 134.105000 ;
      RECT 74.025000 134.035000 75.145000 134.105000 ;
      RECT 74.035000 104.845000 75.000000 105.150000 ;
      RECT 74.095000 133.965000 75.145000 134.035000 ;
      RECT 74.095000 133.965000 75.145000 134.035000 ;
      RECT 74.165000 133.895000 75.145000 133.965000 ;
      RECT 74.165000 133.895000 75.145000 133.965000 ;
      RECT 74.235000 133.825000 75.145000 133.895000 ;
      RECT 74.235000 133.825000 75.145000 133.895000 ;
      RECT 74.305000 133.755000 75.145000 133.825000 ;
      RECT 74.305000 133.755000 75.145000 133.825000 ;
      RECT 74.315000 105.430000 74.915000 125.440000 ;
      RECT 74.375000 133.685000 75.145000 133.755000 ;
      RECT 74.375000 133.685000 75.145000 133.755000 ;
      RECT 74.445000 133.615000 75.145000 133.685000 ;
      RECT 74.445000 133.615000 75.145000 133.685000 ;
      RECT 74.515000 133.545000 75.145000 133.615000 ;
      RECT 74.515000 133.545000 75.145000 133.615000 ;
      RECT 74.585000 133.475000 75.145000 133.545000 ;
      RECT 74.585000 133.475000 75.145000 133.545000 ;
      RECT 74.655000 133.405000 75.145000 133.475000 ;
      RECT 74.655000 133.405000 75.145000 133.475000 ;
      RECT 74.725000 133.335000 75.145000 133.405000 ;
      RECT 74.725000 133.335000 75.145000 133.405000 ;
      RECT 74.795000 133.265000 75.145000 133.335000 ;
      RECT 74.795000 133.265000 75.145000 133.335000 ;
      RECT 74.855000 102.200000 74.925000 102.270000 ;
      RECT 74.855000 102.270000 74.995000 102.340000 ;
      RECT 74.855000 102.340000 75.065000 102.410000 ;
      RECT 74.855000 102.410000 75.135000 102.420000 ;
      RECT 74.865000 133.195000 75.145000 133.265000 ;
      RECT 74.865000 133.195000 75.145000 133.265000 ;
      RECT 74.935000 133.125000 75.145000 133.195000 ;
      RECT 74.935000 133.125000 75.145000 133.195000 ;
      RECT 75.005000 133.055000 75.145000 133.125000 ;
      RECT 75.005000 133.055000 75.145000 133.125000 ;
      RECT 75.075000 132.985000 75.145000 133.055000 ;
      RECT 75.075000 132.985000 75.145000 133.055000 ;
    LAYER met2 ;
      RECT  0.000000   0.000000  8.145000   4.405000 ;
      RECT  0.000000   0.000000  8.285000   1.320000 ;
      RECT  0.000000   1.320000 12.145000   1.610000 ;
      RECT  0.000000   1.610000 17.105000   3.275000 ;
      RECT  0.000000   3.155000 10.635000   3.225000 ;
      RECT  0.000000   3.225000 10.565000   3.295000 ;
      RECT  0.000000   3.275000 19.935000   3.295000 ;
      RECT  0.000000   3.295000  9.595000   4.460000 ;
      RECT  0.000000   3.295000 10.495000   3.365000 ;
      RECT  0.000000   3.365000 10.425000   3.435000 ;
      RECT  0.000000   3.435000 10.355000   3.505000 ;
      RECT  0.000000   3.505000 10.285000   3.575000 ;
      RECT  0.000000   3.575000 10.215000   3.645000 ;
      RECT  0.000000   3.645000 10.145000   3.715000 ;
      RECT  0.000000   3.715000 10.075000   3.785000 ;
      RECT  0.000000   3.785000 10.005000   3.855000 ;
      RECT  0.000000   3.855000  9.935000   3.925000 ;
      RECT  0.000000   3.925000  9.865000   3.995000 ;
      RECT  0.000000   3.995000  9.795000   4.065000 ;
      RECT  0.000000   4.065000  9.725000   4.135000 ;
      RECT  0.000000   4.135000  9.655000   4.205000 ;
      RECT  0.000000   4.205000  9.585000   4.275000 ;
      RECT  0.000000   4.275000  9.515000   4.345000 ;
      RECT  0.000000   4.345000  9.455000   4.405000 ;
      RECT  0.000000   4.405000  3.005000  26.495000 ;
      RECT  0.000000   4.460000  9.595000   9.030000 ;
      RECT  0.000000   9.030000 10.725000  10.160000 ;
      RECT  0.000000   9.085000  9.455000   9.155000 ;
      RECT  0.000000   9.155000  9.525000   9.225000 ;
      RECT  0.000000   9.225000  9.595000   9.295000 ;
      RECT  0.000000   9.295000  9.665000   9.365000 ;
      RECT  0.000000   9.365000  9.735000   9.435000 ;
      RECT  0.000000   9.435000  9.805000   9.505000 ;
      RECT  0.000000   9.505000  9.875000   9.575000 ;
      RECT  0.000000   9.575000  9.945000   9.645000 ;
      RECT  0.000000   9.645000 10.015000   9.715000 ;
      RECT  0.000000   9.715000 10.085000   9.785000 ;
      RECT  0.000000   9.785000 10.155000   9.855000 ;
      RECT  0.000000   9.855000 10.225000   9.925000 ;
      RECT  0.000000   9.925000 10.295000   9.995000 ;
      RECT  0.000000   9.995000 10.365000  10.065000 ;
      RECT  0.000000  10.065000 10.435000  10.135000 ;
      RECT  0.000000  10.135000 10.505000  10.205000 ;
      RECT  0.000000  10.160000 10.725000  26.550000 ;
      RECT  0.000000  10.205000 10.575000  10.215000 ;
      RECT  0.000000  26.495000 10.515000  26.565000 ;
      RECT  0.000000  26.550000 10.510000  26.765000 ;
      RECT  0.000000  26.565000 10.445000  26.635000 ;
      RECT  0.000000  26.635000 10.375000  26.705000 ;
      RECT  0.000000  26.705000 10.370000  26.710000 ;
      RECT  0.000000  26.710000  3.005000 196.995000 ;
      RECT  0.000000  26.765000 10.510000  28.470000 ;
      RECT  0.000000  28.470000 10.725000  28.685000 ;
      RECT  0.000000  28.525000 10.370000  28.595000 ;
      RECT  0.000000  28.595000 10.440000  28.665000 ;
      RECT  0.000000  28.665000 10.510000  28.735000 ;
      RECT  0.000000  28.685000 10.725000  31.255000 ;
      RECT  0.000000  28.735000 10.580000  28.740000 ;
      RECT  0.000000  31.255000 11.120000  31.650000 ;
      RECT  0.000000  31.310000 10.585000  31.380000 ;
      RECT  0.000000  31.380000 10.655000  31.450000 ;
      RECT  0.000000  31.450000 10.725000  31.520000 ;
      RECT  0.000000  31.520000 10.795000  31.590000 ;
      RECT  0.000000  31.590000 10.865000  31.660000 ;
      RECT  0.000000  31.650000 11.120000  36.420000 ;
      RECT  0.000000  31.660000 10.935000  31.705000 ;
      RECT  0.000000  36.420000 75.000000 200.000000 ;
      RECT  0.000000 196.995000 75.000000 200.000000 ;
      RECT  3.000000   3.002000  5.145000   4.460000 ;
      RECT  3.000000   4.460000  6.455000  10.330000 ;
      RECT  3.000000  10.330000  6.455000  10.400000 ;
      RECT  3.000000  10.330000  6.455000  10.400000 ;
      RECT  3.000000  10.400000  6.520000  10.470000 ;
      RECT  3.000000  10.400000  6.520000  10.470000 ;
      RECT  3.000000  10.470000  6.595000  10.540000 ;
      RECT  3.000000  10.470000  6.595000  10.540000 ;
      RECT  3.000000  10.540000  6.665000  10.610000 ;
      RECT  3.000000  10.540000  6.665000  10.610000 ;
      RECT  3.000000  10.610000  6.730000  10.680000 ;
      RECT  3.000000  10.610000  6.730000  10.680000 ;
      RECT  3.000000  10.680000  6.805000  10.750000 ;
      RECT  3.000000  10.680000  6.805000  10.750000 ;
      RECT  3.000000  10.750000  6.875000  10.820000 ;
      RECT  3.000000  10.750000  6.875000  10.820000 ;
      RECT  3.000000  10.820000  6.940000  10.890000 ;
      RECT  3.000000  10.820000  6.940000  10.890000 ;
      RECT  3.000000  10.890000  7.015000  10.960000 ;
      RECT  3.000000  10.890000  7.015000  10.960000 ;
      RECT  3.000000  10.960000  7.085000  11.030000 ;
      RECT  3.000000  10.960000  7.085000  11.030000 ;
      RECT  3.000000  11.030000  7.150000  11.100000 ;
      RECT  3.000000  11.030000  7.150000  11.100000 ;
      RECT  3.000000  11.100000  7.225000  11.170000 ;
      RECT  3.000000  11.100000  7.225000  11.170000 ;
      RECT  3.000000  11.170000  7.295000  11.240000 ;
      RECT  3.000000  11.170000  7.295000  11.240000 ;
      RECT  3.000000  11.240000  7.365000  11.310000 ;
      RECT  3.000000  11.240000  7.365000  11.310000 ;
      RECT  3.000000  11.310000  7.435000  11.380000 ;
      RECT  3.000000  11.310000  7.435000  11.380000 ;
      RECT  3.000000  11.380000  7.505000  11.450000 ;
      RECT  3.000000  11.380000  7.505000  11.450000 ;
      RECT  3.000000  11.450000  7.575000  11.460000 ;
      RECT  3.000000  11.450000  7.575000  11.460000 ;
      RECT  3.000000  11.460000  7.585000  25.250000 ;
      RECT  3.000000  25.250000  7.515000  25.320000 ;
      RECT  3.000000  25.250000  7.515000  25.320000 ;
      RECT  3.000000  25.320000  7.440000  25.390000 ;
      RECT  3.000000  25.320000  7.440000  25.390000 ;
      RECT  3.000000  25.390000  7.375000  25.460000 ;
      RECT  3.000000  25.390000  7.375000  25.460000 ;
      RECT  3.000000  25.460000  7.370000  25.465000 ;
      RECT  3.000000  25.460000  7.370000  25.465000 ;
      RECT  3.000000  25.465000  7.370000  29.770000 ;
      RECT  3.000000  29.770000  7.370000  29.840000 ;
      RECT  3.000000  29.770000  7.370000  29.840000 ;
      RECT  3.000000  29.840000  7.435000  29.910000 ;
      RECT  3.000000  29.840000  7.435000  29.910000 ;
      RECT  3.000000  29.910000  7.510000  29.980000 ;
      RECT  3.000000  29.910000  7.510000  29.980000 ;
      RECT  3.000000  29.980000  7.580000  29.985000 ;
      RECT  3.000000  29.980000  7.580000  29.985000 ;
      RECT  3.000000  29.985000  7.585000  32.555000 ;
      RECT  3.000000  32.555000  7.585000  32.625000 ;
      RECT  3.000000  32.555000  7.585000  32.625000 ;
      RECT  3.000000  32.625000  7.650000  32.695000 ;
      RECT  3.000000  32.625000  7.650000  32.695000 ;
      RECT  3.000000  32.695000  7.725000  32.765000 ;
      RECT  3.000000  32.695000  7.725000  32.765000 ;
      RECT  3.000000  32.765000  7.795000  32.835000 ;
      RECT  3.000000  32.765000  7.795000  32.835000 ;
      RECT  3.000000  32.835000  7.865000  32.905000 ;
      RECT  3.000000  32.835000  7.865000  32.905000 ;
      RECT  3.000000  32.905000  7.935000  32.950000 ;
      RECT  3.000000  32.905000  7.935000  32.950000 ;
      RECT  3.000000  32.950000  7.975000  39.560000 ;
      RECT  3.000000  39.560000 72.000000 197.000000 ;
      RECT  5.145000   4.405000  9.455000   7.410000 ;
      RECT  6.450000   1.750000 16.965000   3.155000 ;
      RECT  6.450000   3.155000  9.455000   4.405000 ;
      RECT  6.450000   7.410000  9.455000  10.215000 ;
      RECT  6.455000  10.215000 10.585000  13.220000 ;
      RECT  7.365000  26.710000 10.370000  28.740000 ;
      RECT  7.365000  28.740000 10.585000  31.310000 ;
      RECT  7.370000  23.490000 10.585000  26.495000 ;
      RECT  7.370000  31.310000 10.585000  31.705000 ;
      RECT  7.370000  31.705000 10.980000  31.745000 ;
      RECT  7.580000  13.220000 10.585000  23.490000 ;
      RECT  7.580000  31.745000 10.980000  36.560000 ;
      RECT  7.975000  36.560000 15.435000  39.560000 ;
      RECT  7.975000  39.560000 15.430000  39.565000 ;
      RECT  8.145000   1.460000 12.005000   1.750000 ;
      RECT  9.035000   0.000000 12.145000   1.320000 ;
      RECT  9.175000   0.000000 12.005000   1.460000 ;
      RECT 10.135000   4.685000 15.825000   4.945000 ;
      RECT 10.135000   4.945000 29.180000   5.525000 ;
      RECT 10.135000   5.525000 29.180000   8.800000 ;
      RECT 10.135000   8.800000 29.180000   9.930000 ;
      RECT 10.275000   4.745000 15.430000   4.815000 ;
      RECT 10.275000   4.815000 15.500000   4.885000 ;
      RECT 10.275000   4.885000 15.570000   4.955000 ;
      RECT 10.275000   4.955000 15.640000   5.025000 ;
      RECT 10.275000   5.025000 15.710000   5.085000 ;
      RECT 10.275000   5.085000 28.540000   5.155000 ;
      RECT 10.275000   5.155000 28.610000   5.225000 ;
      RECT 10.275000   5.225000 28.680000   5.295000 ;
      RECT 10.275000   5.295000 28.750000   5.365000 ;
      RECT 10.275000   5.365000 28.820000   5.435000 ;
      RECT 10.275000   5.435000 28.890000   5.505000 ;
      RECT 10.275000   5.505000 28.960000   5.575000 ;
      RECT 10.275000   5.575000 29.030000   5.585000 ;
      RECT 10.275000   5.585000 29.040000   8.590000 ;
      RECT 10.275000   8.590000 14.405000   8.745000 ;
      RECT 10.345000   4.675000 15.360000   4.745000 ;
      RECT 10.345000   8.745000 29.040000   8.815000 ;
      RECT 10.415000   4.605000 15.290000   4.675000 ;
      RECT 10.415000   8.815000 29.040000   8.885000 ;
      RECT 10.485000   4.535000 15.220000   4.605000 ;
      RECT 10.485000   8.885000 29.040000   8.955000 ;
      RECT 10.555000   4.465000 15.150000   4.535000 ;
      RECT 10.555000   8.955000 29.040000   9.025000 ;
      RECT 10.625000   4.395000 15.080000   4.465000 ;
      RECT 10.625000   9.025000 29.040000   9.095000 ;
      RECT 10.695000   4.325000 15.010000   4.395000 ;
      RECT 10.695000   9.095000 29.040000   9.165000 ;
      RECT 10.765000   4.255000 14.940000   4.325000 ;
      RECT 10.765000   9.165000 29.040000   9.235000 ;
      RECT 10.835000   4.185000 14.870000   4.255000 ;
      RECT 10.835000   9.235000 29.040000   9.305000 ;
      RECT 10.905000   4.115000 14.800000   4.185000 ;
      RECT 10.905000   9.305000 29.040000   9.375000 ;
      RECT 10.975000   4.045000 14.730000   4.115000 ;
      RECT 10.975000   9.375000 29.040000   9.445000 ;
      RECT 10.990000   3.835000 15.570000   4.685000 ;
      RECT 11.045000   3.975000 14.660000   4.045000 ;
      RECT 11.045000   9.445000 29.040000   9.515000 ;
      RECT 11.050000  27.360000 75.000000  27.875000 ;
      RECT 11.050000  27.875000 75.000000  28.090000 ;
      RECT 11.115000   9.515000 29.040000   9.585000 ;
      RECT 11.185000   9.585000 29.040000   9.655000 ;
      RECT 11.190000  27.415000 14.805000  27.820000 ;
      RECT 11.195000  27.410000 75.000000  27.415000 ;
      RECT 11.255000   9.655000 29.040000   9.725000 ;
      RECT 11.260000  27.820000 75.000000  27.890000 ;
      RECT 11.265000   9.930000 29.180000  11.145000 ;
      RECT 11.265000  11.145000 29.630000  11.595000 ;
      RECT 11.265000  11.595000 29.630000  15.815000 ;
      RECT 11.265000  15.815000 30.225000  16.410000 ;
      RECT 11.265000  16.410000 30.225000  20.635000 ;
      RECT 11.265000  20.635000 75.000000  27.145000 ;
      RECT 11.265000  27.145000 75.000000  27.360000 ;
      RECT 11.265000  27.340000 75.000000  27.410000 ;
      RECT 11.265000  28.090000 75.000000  31.025000 ;
      RECT 11.265000  31.025000 75.000000  31.420000 ;
      RECT 11.325000   9.725000 29.040000   9.795000 ;
      RECT 11.330000  27.890000 75.000000  27.960000 ;
      RECT 11.335000  27.270000 75.000000  27.340000 ;
      RECT 11.395000   9.795000 29.040000   9.865000 ;
      RECT 11.400000  27.960000 75.000000  28.030000 ;
      RECT 11.405000   9.865000 29.040000   9.875000 ;
      RECT 11.405000   9.875000 14.405000  11.200000 ;
      RECT 11.405000  11.200000 29.040000  11.270000 ;
      RECT 11.405000  11.270000 29.110000  11.340000 ;
      RECT 11.405000  11.340000 29.180000  11.410000 ;
      RECT 11.405000  11.410000 29.250000  11.480000 ;
      RECT 11.405000  11.480000 29.320000  11.550000 ;
      RECT 11.405000  11.550000 29.390000  11.620000 ;
      RECT 11.405000  11.620000 29.460000  11.650000 ;
      RECT 11.405000  11.650000 14.410000  15.870000 ;
      RECT 11.405000  15.870000 29.490000  15.940000 ;
      RECT 11.405000  15.940000 29.560000  16.010000 ;
      RECT 11.405000  16.010000 29.630000  16.080000 ;
      RECT 11.405000  16.080000 29.700000  16.150000 ;
      RECT 11.405000  16.150000 29.770000  16.220000 ;
      RECT 11.405000  16.220000 29.840000  16.290000 ;
      RECT 11.405000  16.290000 29.910000  16.360000 ;
      RECT 11.405000  16.360000 29.980000  16.430000 ;
      RECT 11.405000  16.430000 30.050000  16.465000 ;
      RECT 11.405000  16.465000 14.410000  20.775000 ;
      RECT 11.405000  20.775000 14.805000  27.415000 ;
      RECT 11.405000  27.200000 75.000000  27.270000 ;
      RECT 11.405000  27.820000 14.805000  30.970000 ;
      RECT 11.405000  28.030000 75.000000  28.035000 ;
      RECT 11.475000  30.970000 75.000000  31.040000 ;
      RECT 11.545000  31.040000 75.000000  31.110000 ;
      RECT 11.615000  31.110000 75.000000  31.180000 ;
      RECT 11.660000  31.420000 75.000000  35.880000 ;
      RECT 11.685000  31.180000 75.000000  31.250000 ;
      RECT 11.755000  31.250000 75.000000  31.320000 ;
      RECT 11.800000  30.970000 14.805000  35.740000 ;
      RECT 11.800000  31.320000 75.000000  31.365000 ;
      RECT 12.290000  35.880000 75.000000  36.420000 ;
      RECT 12.430000  20.775000 75.000000  36.560000 ;
      RECT 12.685000   0.000000 14.415000   1.125000 ;
      RECT 12.685000   1.125000 17.105000   1.610000 ;
      RECT 12.795000   1.745000 16.965000   1.750000 ;
      RECT 12.810000   1.730000 16.965000   1.745000 ;
      RECT 12.825000   0.000000 14.275000   1.265000 ;
      RECT 12.825000   1.265000 16.965000   1.715000 ;
      RECT 12.825000   1.715000 16.965000   1.730000 ;
      RECT 13.275000   6.975000 13.415000   7.045000 ;
      RECT 13.275000   6.975000 13.415000   7.045000 ;
      RECT 13.275000   7.045000 13.485000   7.115000 ;
      RECT 13.275000   7.045000 13.485000   7.115000 ;
      RECT 13.275000   7.115000 13.555000   7.185000 ;
      RECT 13.275000   7.115000 13.555000   7.185000 ;
      RECT 13.275000   7.185000 13.625000   7.255000 ;
      RECT 13.275000   7.185000 13.625000   7.255000 ;
      RECT 13.275000   7.255000 13.695000   7.325000 ;
      RECT 13.275000   7.255000 13.695000   7.325000 ;
      RECT 13.275000   7.325000 13.765000   7.395000 ;
      RECT 13.275000   7.325000 13.765000   7.395000 ;
      RECT 13.275000   7.395000 13.835000   7.465000 ;
      RECT 13.275000   7.395000 13.835000   7.465000 ;
      RECT 13.275000   7.465000 13.905000   7.500000 ;
      RECT 13.275000   7.465000 13.905000   7.500000 ;
      RECT 13.345000   7.500000 13.940000   7.570000 ;
      RECT 13.345000   7.500000 13.940000   7.570000 ;
      RECT 13.415000   7.570000 14.010000   7.640000 ;
      RECT 13.415000   7.570000 14.010000   7.640000 ;
      RECT 13.485000   7.640000 14.080000   7.710000 ;
      RECT 13.485000   7.640000 14.080000   7.710000 ;
      RECT 13.555000   7.710000 14.150000   7.780000 ;
      RECT 13.555000   7.710000 14.150000   7.780000 ;
      RECT 13.625000   7.780000 14.220000   7.850000 ;
      RECT 13.625000   7.780000 14.220000   7.850000 ;
      RECT 13.695000   7.850000 14.290000   7.920000 ;
      RECT 13.695000   7.850000 14.290000   7.920000 ;
      RECT 13.765000   7.920000 14.360000   7.990000 ;
      RECT 13.765000   7.920000 14.360000   7.990000 ;
      RECT 13.835000   7.990000 14.430000   8.060000 ;
      RECT 13.835000   7.990000 14.430000   8.060000 ;
      RECT 13.860000   8.060000 14.500000   8.085000 ;
      RECT 13.860000   8.060000 14.500000   8.085000 ;
      RECT 13.930000   8.085000 26.040000   8.155000 ;
      RECT 13.930000   8.085000 26.040000   8.155000 ;
      RECT 14.000000   8.155000 26.040000   8.225000 ;
      RECT 14.000000   8.155000 26.040000   8.225000 ;
      RECT 14.070000   8.225000 26.040000   8.295000 ;
      RECT 14.070000   8.225000 26.040000   8.295000 ;
      RECT 14.140000   8.295000 26.040000   8.365000 ;
      RECT 14.140000   8.295000 26.040000   8.365000 ;
      RECT 14.210000   8.365000 26.040000   8.435000 ;
      RECT 14.210000   8.365000 26.040000   8.435000 ;
      RECT 14.280000   8.435000 26.040000   8.505000 ;
      RECT 14.280000   8.435000 26.040000   8.505000 ;
      RECT 14.350000   8.505000 26.040000   8.575000 ;
      RECT 14.350000   8.505000 26.040000   8.575000 ;
      RECT 14.405000   8.575000 26.040000   8.630000 ;
      RECT 14.405000   8.575000 26.040000   8.630000 ;
      RECT 14.405000   8.630000 26.040000  12.445000 ;
      RECT 14.405000  12.445000 26.040000  12.515000 ;
      RECT 14.405000  12.445000 26.040000  12.515000 ;
      RECT 14.405000  12.515000 26.110000  12.585000 ;
      RECT 14.405000  12.515000 26.110000  12.585000 ;
      RECT 14.405000  12.585000 26.180000  12.655000 ;
      RECT 14.405000  12.585000 26.180000  12.655000 ;
      RECT 14.405000  12.655000 26.250000  12.725000 ;
      RECT 14.405000  12.655000 26.250000  12.725000 ;
      RECT 14.405000  12.725000 26.320000  12.795000 ;
      RECT 14.405000  12.725000 26.320000  12.795000 ;
      RECT 14.405000  12.795000 26.390000  12.865000 ;
      RECT 14.405000  12.795000 26.390000  12.865000 ;
      RECT 14.405000  12.865000 26.455000  12.895000 ;
      RECT 14.405000  12.865000 26.455000  12.895000 ;
      RECT 14.405000  12.895000 26.490000  17.115000 ;
      RECT 14.405000  17.115000 26.490000  17.185000 ;
      RECT 14.405000  17.115000 26.490000  17.185000 ;
      RECT 14.405000  17.185000 26.560000  17.255000 ;
      RECT 14.405000  17.185000 26.560000  17.255000 ;
      RECT 14.405000  17.255000 26.630000  17.325000 ;
      RECT 14.405000  17.255000 26.630000  17.325000 ;
      RECT 14.405000  17.325000 26.700000  17.395000 ;
      RECT 14.405000  17.325000 26.700000  17.395000 ;
      RECT 14.405000  17.395000 26.770000  17.465000 ;
      RECT 14.405000  17.395000 26.770000  17.465000 ;
      RECT 14.405000  17.465000 26.840000  17.535000 ;
      RECT 14.405000  17.465000 26.840000  17.535000 ;
      RECT 14.405000  17.535000 26.910000  17.605000 ;
      RECT 14.405000  17.535000 26.910000  17.605000 ;
      RECT 14.405000  17.605000 26.980000  17.675000 ;
      RECT 14.405000  17.605000 26.980000  17.675000 ;
      RECT 14.405000  17.675000 27.045000  17.710000 ;
      RECT 14.405000  17.675000 27.045000  17.710000 ;
      RECT 14.405000  17.710000 27.080000  23.775000 ;
      RECT 14.405000  23.775000 72.000000  29.725000 ;
      RECT 14.475000  29.725000 72.000000  29.795000 ;
      RECT 14.475000  29.725000 72.000000  29.795000 ;
      RECT 14.545000  29.795000 72.000000  29.865000 ;
      RECT 14.545000  29.795000 72.000000  29.865000 ;
      RECT 14.615000  29.865000 72.000000  29.935000 ;
      RECT 14.615000  29.865000 72.000000  29.935000 ;
      RECT 14.685000  29.935000 72.000000  30.005000 ;
      RECT 14.685000  29.935000 72.000000  30.005000 ;
      RECT 14.755000  30.005000 72.000000  30.075000 ;
      RECT 14.755000  30.005000 72.000000  30.075000 ;
      RECT 14.800000  30.075000 72.000000  30.120000 ;
      RECT 14.800000  30.075000 72.000000  30.120000 ;
      RECT 14.800000  30.120000 72.000000  32.740000 ;
      RECT 14.945000   3.295000 19.935000   3.595000 ;
      RECT 15.070000   3.155000 16.965000   3.225000 ;
      RECT 15.140000   3.225000 16.965000   3.295000 ;
      RECT 15.210000   3.295000 16.965000   3.365000 ;
      RECT 15.245000   3.595000 22.220000   4.185000 ;
      RECT 15.260000   3.365000 16.965000   3.415000 ;
      RECT 15.275000   0.000000 17.105000   1.125000 ;
      RECT 15.330000   3.415000 19.795000   3.485000 ;
      RECT 15.400000   3.485000 19.795000   3.555000 ;
      RECT 15.415000   0.000000 16.965000   1.265000 ;
      RECT 15.430000  32.740000 72.000000  39.560000 ;
      RECT 15.470000   3.555000 19.795000   3.625000 ;
      RECT 15.540000   3.625000 19.795000   3.695000 ;
      RECT 15.580000   3.695000 19.795000   3.735000 ;
      RECT 15.650000   3.735000 22.080000   3.805000 ;
      RECT 15.720000   3.805000 22.080000   3.875000 ;
      RECT 15.790000   3.875000 22.080000   3.945000 ;
      RECT 15.835000   4.185000 22.000000   4.405000 ;
      RECT 15.860000   3.945000 22.080000   4.015000 ;
      RECT 15.930000   4.015000 22.080000   4.085000 ;
      RECT 15.975000   4.085000 22.080000   4.130000 ;
      RECT 16.040000   4.130000 22.015000   4.195000 ;
      RECT 16.110000   4.195000 21.945000   4.265000 ;
      RECT 19.050000   0.000000 19.935000   3.275000 ;
      RECT 19.190000   0.000000 19.795000   3.415000 ;
      RECT 21.365000   0.000000 22.220000   3.595000 ;
      RECT 21.505000   0.000000 22.080000   3.735000 ;
      RECT 22.800000   0.000000 27.440000   0.470000 ;
      RECT 22.800000   0.470000 28.775000   0.475000 ;
      RECT 22.800000   0.475000 32.620000   0.780000 ;
      RECT 22.800000   0.780000 72.075000   0.910000 ;
      RECT 22.800000   0.910000 75.000000   4.200000 ;
      RECT 22.800000   4.200000 75.000000   4.405000 ;
      RECT 22.940000   0.000000 27.300000   0.610000 ;
      RECT 22.940000   0.610000 28.635000   0.615000 ;
      RECT 22.940000   0.615000 32.480000   0.920000 ;
      RECT 22.940000   0.920000 33.300000   3.925000 ;
      RECT 22.940000   3.925000 29.860000   4.145000 ;
      RECT 23.000000   4.145000 75.000000   4.205000 ;
      RECT 23.060000   4.205000 75.000000   4.265000 ;
      RECT 26.035000   8.590000 29.040000   8.745000 ;
      RECT 26.040000   9.875000 29.040000  11.200000 ;
      RECT 26.040000  11.650000 29.490000  14.655000 ;
      RECT 26.485000  14.655000 29.490000  15.870000 ;
      RECT 26.490000  16.465000 30.085000  19.470000 ;
      RECT 27.080000  19.470000 30.085000  20.775000 ;
      RECT 28.370000   0.000000 28.775000   0.470000 ;
      RECT 28.825000   4.405000 75.000000   5.300000 ;
      RECT 28.950000   4.265000 75.000000   4.335000 ;
      RECT 29.020000   4.335000 75.000000   4.405000 ;
      RECT 29.090000   4.405000 75.000000   4.475000 ;
      RECT 29.160000   4.475000 75.000000   4.545000 ;
      RECT 29.230000   4.545000 75.000000   4.615000 ;
      RECT 29.300000   4.615000 75.000000   4.685000 ;
      RECT 29.370000   4.685000 75.000000   4.755000 ;
      RECT 29.440000   4.755000 75.000000   4.825000 ;
      RECT 29.510000   4.825000 75.000000   4.895000 ;
      RECT 29.580000   4.895000 75.000000   4.965000 ;
      RECT 29.650000   4.965000 75.000000   5.035000 ;
      RECT 29.720000   5.035000 75.000000   5.105000 ;
      RECT 29.720000   5.300000 75.000000  10.915000 ;
      RECT 29.720000  10.915000 75.000000  11.365000 ;
      RECT 29.790000   5.105000 75.000000   5.175000 ;
      RECT 29.825000   0.000000 30.365000   0.470000 ;
      RECT 29.825000   0.470000 32.620000   0.475000 ;
      RECT 29.860000   1.050000 75.000000  10.860000 ;
      RECT 29.860000   1.050000 75.000000  10.860000 ;
      RECT 29.860000   5.175000 75.000000   5.245000 ;
      RECT 29.930000  10.860000 75.000000  10.930000 ;
      RECT 29.965000   0.000000 30.225000   0.610000 ;
      RECT 29.965000   0.610000 32.480000   0.615000 ;
      RECT 30.000000  10.930000 75.000000  11.000000 ;
      RECT 30.070000  11.000000 75.000000  11.070000 ;
      RECT 30.140000  11.070000 75.000000  11.140000 ;
      RECT 30.170000  11.365000 75.000000  15.585000 ;
      RECT 30.170000  15.585000 75.000000  16.180000 ;
      RECT 30.210000  11.140000 75.000000  11.210000 ;
      RECT 30.280000  11.210000 75.000000  11.280000 ;
      RECT 30.310000  10.860000 33.315000  12.525000 ;
      RECT 30.310000  11.280000 75.000000  11.310000 ;
      RECT 30.310000  12.525000 33.905000  15.530000 ;
      RECT 30.380000  15.530000 75.000000  15.600000 ;
      RECT 30.450000  15.600000 75.000000  15.670000 ;
      RECT 30.520000  15.670000 75.000000  15.740000 ;
      RECT 30.590000  15.740000 75.000000  15.810000 ;
      RECT 30.660000  15.810000 75.000000  15.880000 ;
      RECT 30.730000  15.880000 75.000000  15.950000 ;
      RECT 30.765000  16.180000 75.000000  20.635000 ;
      RECT 30.800000  15.950000 75.000000  16.020000 ;
      RECT 30.870000  16.020000 75.000000  16.090000 ;
      RECT 30.905000  16.090000 75.000000  16.125000 ;
      RECT 30.905000  16.125000 33.910000  20.775000 ;
      RECT 31.295000   0.000000 32.620000   0.470000 ;
      RECT 31.435000   0.000000 32.480000   0.610000 ;
      RECT 32.820000   3.920000 68.935000   3.960000 ;
      RECT 32.820000   3.920000 68.935000   3.960000 ;
      RECT 32.860000   3.960000 68.935000   4.000000 ;
      RECT 32.860000   3.960000 68.935000   4.000000 ;
      RECT 32.860000   4.000000 68.935000   4.050000 ;
      RECT 32.860000   4.050000 72.000000   9.615000 ;
      RECT 32.930000   9.615000 72.000000   9.685000 ;
      RECT 32.930000   9.615000 72.000000   9.685000 ;
      RECT 33.000000   9.685000 72.000000   9.755000 ;
      RECT 33.000000   9.685000 72.000000   9.755000 ;
      RECT 33.070000   9.755000 72.000000   9.825000 ;
      RECT 33.070000   9.755000 72.000000   9.825000 ;
      RECT 33.140000   9.825000 72.000000   9.895000 ;
      RECT 33.140000   9.825000 72.000000   9.895000 ;
      RECT 33.160000   0.000000 72.075000   0.780000 ;
      RECT 33.210000   9.895000 72.000000   9.965000 ;
      RECT 33.210000   9.895000 72.000000   9.965000 ;
      RECT 33.280000   9.965000 72.000000  10.035000 ;
      RECT 33.280000   9.965000 72.000000  10.035000 ;
      RECT 33.300000   0.000000 71.935000  10.860000 ;
      RECT 33.300000   0.000000 71.935000  10.860000 ;
      RECT 33.310000  10.035000 72.000000  10.065000 ;
      RECT 33.310000  10.035000 72.000000  10.065000 ;
      RECT 33.310000  10.065000 72.000000  14.285000 ;
      RECT 33.380000  14.285000 72.000000  14.355000 ;
      RECT 33.380000  14.285000 72.000000  14.355000 ;
      RECT 33.450000  14.355000 72.000000  14.425000 ;
      RECT 33.450000  14.355000 72.000000  14.425000 ;
      RECT 33.520000  14.425000 72.000000  14.495000 ;
      RECT 33.520000  14.425000 72.000000  14.495000 ;
      RECT 33.590000  14.495000 72.000000  14.565000 ;
      RECT 33.590000  14.495000 72.000000  14.565000 ;
      RECT 33.660000  14.565000 72.000000  14.635000 ;
      RECT 33.660000  14.565000 72.000000  14.635000 ;
      RECT 33.730000  14.635000 72.000000  14.705000 ;
      RECT 33.730000  14.635000 72.000000  14.705000 ;
      RECT 33.800000  14.705000 72.000000  14.775000 ;
      RECT 33.800000  14.705000 72.000000  14.775000 ;
      RECT 33.870000  14.775000 72.000000  14.845000 ;
      RECT 33.870000  14.775000 72.000000  14.845000 ;
      RECT 33.905000  14.845000 72.000000  14.880000 ;
      RECT 33.905000  14.845000 72.000000  14.880000 ;
      RECT 33.905000  14.880000 72.000000  23.775000 ;
      RECT 36.300000   3.000000 68.935000   3.920000 ;
      RECT 71.995000  10.860000 75.000000  15.530000 ;
      RECT 71.995000  16.125000 75.000000  20.775000 ;
      RECT 71.995000  36.560000 75.000000 196.995000 ;
      RECT 73.130000   1.020000 75.000000   1.050000 ;
      RECT 73.375000   0.000000 75.000000   0.910000 ;
      RECT 73.515000   0.000000 75.000000   1.020000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000  8.000000   3.005000 ;
      RECT  0.000000   0.000000  8.100000  15.660000 ;
      RECT  0.000000   3.005000  3.005000  17.245000 ;
      RECT  0.000000  15.620000  7.850000  15.770000 ;
      RECT  0.000000  15.660000  6.475000  17.285000 ;
      RECT  0.000000  15.770000  7.700000  15.920000 ;
      RECT  0.000000  15.920000  7.550000  16.070000 ;
      RECT  0.000000  16.070000  7.400000  16.220000 ;
      RECT  0.000000  16.220000  7.250000  16.370000 ;
      RECT  0.000000  16.370000  7.100000  16.520000 ;
      RECT  0.000000  16.520000  6.950000  16.670000 ;
      RECT  0.000000  16.670000  6.800000  16.820000 ;
      RECT  0.000000  16.820000  6.650000  16.970000 ;
      RECT  0.000000  16.970000  6.500000  17.120000 ;
      RECT  0.000000  17.120000  6.375000  17.245000 ;
      RECT  0.000000  17.245000  6.375000  64.435000 ;
      RECT  0.000000  17.285000  6.475000  31.630000 ;
      RECT  0.000000  31.630000  9.270000  34.425000 ;
      RECT  0.000000  31.670000  6.375000  31.820000 ;
      RECT  0.000000  31.820000  6.525000  31.970000 ;
      RECT  0.000000  31.970000  6.675000  32.120000 ;
      RECT  0.000000  32.120000  6.825000  32.270000 ;
      RECT  0.000000  32.270000  6.975000  32.420000 ;
      RECT  0.000000  32.420000  7.125000  32.570000 ;
      RECT  0.000000  32.570000  7.275000  32.720000 ;
      RECT  0.000000  32.720000  7.425000  32.870000 ;
      RECT  0.000000  32.870000  7.575000  33.020000 ;
      RECT  0.000000  33.020000  7.725000  33.170000 ;
      RECT  0.000000  33.170000  7.875000  33.320000 ;
      RECT  0.000000  33.320000  8.025000  33.470000 ;
      RECT  0.000000  33.470000  8.175000  33.620000 ;
      RECT  0.000000  33.620000  8.325000  33.770000 ;
      RECT  0.000000  33.770000  8.475000  33.920000 ;
      RECT  0.000000  33.920000  8.625000  34.070000 ;
      RECT  0.000000  34.070000  8.775000  34.220000 ;
      RECT  0.000000  34.220000  8.925000  34.370000 ;
      RECT  0.000000  34.370000  9.075000  34.520000 ;
      RECT  0.000000  34.425000 71.890000  64.475000 ;
      RECT  0.000000  34.520000  9.225000  34.525000 ;
      RECT  0.000000  64.435000 71.640000  64.585000 ;
      RECT  0.000000  64.475000 64.560000  71.805000 ;
      RECT  0.000000  64.585000 71.490000  64.735000 ;
      RECT  0.000000  64.735000 71.340000  64.885000 ;
      RECT  0.000000  64.885000 71.190000  65.035000 ;
      RECT  0.000000  65.035000 71.040000  65.185000 ;
      RECT  0.000000  65.185000 70.890000  65.335000 ;
      RECT  0.000000  65.335000 70.740000  65.485000 ;
      RECT  0.000000  65.485000 70.590000  65.635000 ;
      RECT  0.000000  65.635000 70.440000  65.785000 ;
      RECT  0.000000  65.785000 70.290000  65.935000 ;
      RECT  0.000000  65.935000 70.140000  66.085000 ;
      RECT  0.000000  66.085000 69.990000  66.235000 ;
      RECT  0.000000  66.235000 69.840000  66.385000 ;
      RECT  0.000000  66.385000 69.690000  66.535000 ;
      RECT  0.000000  66.535000 69.540000  66.685000 ;
      RECT  0.000000  66.685000 69.390000  66.835000 ;
      RECT  0.000000  66.835000 69.240000  66.985000 ;
      RECT  0.000000  66.985000 69.090000  67.135000 ;
      RECT  0.000000  67.135000 68.940000  67.285000 ;
      RECT  0.000000  67.285000 68.790000  67.435000 ;
      RECT  0.000000  67.435000 68.640000  67.585000 ;
      RECT  0.000000  67.585000 68.490000  67.735000 ;
      RECT  0.000000  67.735000 68.340000  67.885000 ;
      RECT  0.000000  67.885000 68.190000  68.035000 ;
      RECT  0.000000  68.035000 68.040000  68.185000 ;
      RECT  0.000000  68.185000 67.890000  68.335000 ;
      RECT  0.000000  68.335000 67.740000  68.485000 ;
      RECT  0.000000  68.485000 67.590000  68.635000 ;
      RECT  0.000000  68.635000 67.440000  68.785000 ;
      RECT  0.000000  68.785000 67.290000  68.935000 ;
      RECT  0.000000  68.935000 67.140000  69.085000 ;
      RECT  0.000000  69.085000 66.990000  69.235000 ;
      RECT  0.000000  69.235000 66.840000  69.385000 ;
      RECT  0.000000  69.385000 66.690000  69.535000 ;
      RECT  0.000000  69.535000 66.540000  69.685000 ;
      RECT  0.000000  69.685000 66.390000  69.835000 ;
      RECT  0.000000  69.835000 66.240000  69.985000 ;
      RECT  0.000000  69.985000 66.090000  70.135000 ;
      RECT  0.000000  70.135000 65.940000  70.285000 ;
      RECT  0.000000  70.285000 65.790000  70.435000 ;
      RECT  0.000000  70.435000 65.640000  70.585000 ;
      RECT  0.000000  70.585000 65.490000  70.735000 ;
      RECT  0.000000  70.735000 65.340000  70.885000 ;
      RECT  0.000000  70.885000 65.190000  71.035000 ;
      RECT  0.000000  71.035000 65.040000  71.185000 ;
      RECT  0.000000  71.185000 64.890000  71.335000 ;
      RECT  0.000000  71.335000 64.740000  71.485000 ;
      RECT  0.000000  71.485000 64.590000  71.635000 ;
      RECT  0.000000  71.635000 64.460000  71.765000 ;
      RECT  0.000000  71.765000  3.005000 196.995000 ;
      RECT  0.000000  71.805000 64.560000  94.945000 ;
      RECT  0.000000  94.945000 75.000000 200.000000 ;
      RECT  0.000000 196.995000 75.000000 200.000000 ;
      RECT  3.000000   3.002000  5.000000  14.375000 ;
      RECT  3.000000  14.375000  4.850000  14.525000 ;
      RECT  3.000000  14.375000  4.850000  14.525000 ;
      RECT  3.000000  14.525000  4.700000  14.675000 ;
      RECT  3.000000  14.525000  4.700000  14.675000 ;
      RECT  3.000000  14.675000  4.550000  14.825000 ;
      RECT  3.000000  14.675000  4.550000  14.825000 ;
      RECT  3.000000  14.825000  4.395000  14.975000 ;
      RECT  3.000000  14.825000  4.395000  14.975000 ;
      RECT  3.000000  14.975000  4.250000  15.125000 ;
      RECT  3.000000  14.975000  4.250000  15.125000 ;
      RECT  3.000000  15.125000  4.100000  15.275000 ;
      RECT  3.000000  15.125000  4.100000  15.275000 ;
      RECT  3.000000  15.275000  3.945000  15.425000 ;
      RECT  3.000000  15.275000  3.945000  15.425000 ;
      RECT  3.000000  15.425000  3.800000  15.575000 ;
      RECT  3.000000  15.425000  3.800000  15.575000 ;
      RECT  3.000000  15.575000  3.650000  15.725000 ;
      RECT  3.000000  15.575000  3.650000  15.725000 ;
      RECT  3.000000  15.725000  3.500000  15.875000 ;
      RECT  3.000000  15.725000  3.500000  15.875000 ;
      RECT  3.000000  15.875000  3.375000  16.000000 ;
      RECT  3.000000  15.875000  3.375000  16.000000 ;
      RECT  3.000000  16.000000  3.375000  32.915000 ;
      RECT  3.000000  32.915000  3.375000  33.065000 ;
      RECT  3.000000  32.915000  3.375000  33.065000 ;
      RECT  3.000000  33.065000  3.525000  33.215000 ;
      RECT  3.000000  33.065000  3.525000  33.215000 ;
      RECT  3.000000  33.215000  3.675000  33.365000 ;
      RECT  3.000000  33.215000  3.675000  33.365000 ;
      RECT  3.000000  33.365000  3.820000  33.515000 ;
      RECT  3.000000  33.365000  3.820000  33.515000 ;
      RECT  3.000000  33.515000  3.970000  33.665000 ;
      RECT  3.000000  33.515000  3.970000  33.665000 ;
      RECT  3.000000  33.665000  4.125000  33.815000 ;
      RECT  3.000000  33.665000  4.125000  33.815000 ;
      RECT  3.000000  33.815000  4.270000  33.965000 ;
      RECT  3.000000  33.815000  4.270000  33.965000 ;
      RECT  3.000000  33.965000  4.425000  34.115000 ;
      RECT  3.000000  33.965000  4.425000  34.115000 ;
      RECT  3.000000  34.115000  4.575000  34.265000 ;
      RECT  3.000000  34.115000  4.575000  34.265000 ;
      RECT  3.000000  34.265000  4.725000  34.415000 ;
      RECT  3.000000  34.265000  4.725000  34.415000 ;
      RECT  3.000000  34.415000  4.875000  34.565000 ;
      RECT  3.000000  34.415000  4.875000  34.565000 ;
      RECT  3.000000  34.565000  5.020000  34.715000 ;
      RECT  3.000000  34.565000  5.020000  34.715000 ;
      RECT  3.000000  34.715000  5.175000  34.865000 ;
      RECT  3.000000  34.715000  5.175000  34.865000 ;
      RECT  3.000000  34.865000  5.325000  35.015000 ;
      RECT  3.000000  34.865000  5.325000  35.015000 ;
      RECT  3.000000  35.015000  5.475000  35.165000 ;
      RECT  3.000000  35.015000  5.475000  35.165000 ;
      RECT  3.000000  35.165000  5.625000  35.315000 ;
      RECT  3.000000  35.165000  5.625000  35.315000 ;
      RECT  3.000000  35.315000  5.770000  35.465000 ;
      RECT  3.000000  35.315000  5.770000  35.465000 ;
      RECT  3.000000  35.465000  5.925000  35.615000 ;
      RECT  3.000000  35.465000  5.925000  35.615000 ;
      RECT  3.000000  35.615000  6.075000  35.765000 ;
      RECT  3.000000  35.615000  6.075000  35.765000 ;
      RECT  3.000000  35.765000  6.225000  35.915000 ;
      RECT  3.000000  35.765000  6.225000  35.915000 ;
      RECT  3.000000  35.915000  6.375000  36.065000 ;
      RECT  3.000000  35.915000  6.375000  36.065000 ;
      RECT  3.000000  36.065000  6.520000  36.215000 ;
      RECT  3.000000  36.065000  6.520000  36.215000 ;
      RECT  3.000000  36.215000  6.675000  36.365000 ;
      RECT  3.000000  36.215000  6.675000  36.365000 ;
      RECT  3.000000  36.365000  6.825000  36.515000 ;
      RECT  3.000000  36.365000  6.825000  36.515000 ;
      RECT  3.000000  36.515000  6.975000  36.665000 ;
      RECT  3.000000  36.515000  6.975000  36.665000 ;
      RECT  3.000000  36.665000  7.125000  36.815000 ;
      RECT  3.000000  36.665000  7.125000  36.815000 ;
      RECT  3.000000  36.815000  7.270000  36.965000 ;
      RECT  3.000000  36.815000  7.270000  36.965000 ;
      RECT  3.000000  36.965000  7.425000  37.115000 ;
      RECT  3.000000  36.965000  7.425000  37.115000 ;
      RECT  3.000000  37.115000  7.575000  37.265000 ;
      RECT  3.000000  37.115000  7.575000  37.265000 ;
      RECT  3.000000  37.265000  7.725000  37.415000 ;
      RECT  3.000000  37.265000  7.725000  37.415000 ;
      RECT  3.000000  37.415000  7.875000  37.525000 ;
      RECT  3.000000  37.415000  7.875000  37.525000 ;
      RECT  3.000000  37.525000 68.785000  63.190000 ;
      RECT  3.000000  63.190000 68.640000  63.340000 ;
      RECT  3.000000  63.190000 68.640000  63.340000 ;
      RECT  3.000000  63.340000 68.490000  63.490000 ;
      RECT  3.000000  63.340000 68.490000  63.490000 ;
      RECT  3.000000  63.490000 68.335000  63.640000 ;
      RECT  3.000000  63.490000 68.335000  63.640000 ;
      RECT  3.000000  63.640000 68.190000  63.790000 ;
      RECT  3.000000  63.640000 68.190000  63.790000 ;
      RECT  3.000000  63.790000 68.035000  63.940000 ;
      RECT  3.000000  63.790000 68.035000  63.940000 ;
      RECT  3.000000  63.940000 67.890000  64.090000 ;
      RECT  3.000000  63.940000 67.890000  64.090000 ;
      RECT  3.000000  64.090000 67.740000  64.240000 ;
      RECT  3.000000  64.090000 67.740000  64.240000 ;
      RECT  3.000000  64.240000 67.585000  64.390000 ;
      RECT  3.000000  64.240000 67.585000  64.390000 ;
      RECT  3.000000  64.390000 67.440000  64.540000 ;
      RECT  3.000000  64.390000 67.440000  64.540000 ;
      RECT  3.000000  64.540000 67.285000  64.690000 ;
      RECT  3.000000  64.540000 67.285000  64.690000 ;
      RECT  3.000000  64.690000 67.140000  64.840000 ;
      RECT  3.000000  64.690000 67.140000  64.840000 ;
      RECT  3.000000  64.840000 66.990000  64.990000 ;
      RECT  3.000000  64.840000 66.990000  64.990000 ;
      RECT  3.000000  64.990000 66.835000  65.140000 ;
      RECT  3.000000  64.990000 66.835000  65.140000 ;
      RECT  3.000000  65.140000 66.690000  65.290000 ;
      RECT  3.000000  65.140000 66.690000  65.290000 ;
      RECT  3.000000  65.290000 66.535000  65.440000 ;
      RECT  3.000000  65.290000 66.535000  65.440000 ;
      RECT  3.000000  65.440000 66.390000  65.590000 ;
      RECT  3.000000  65.440000 66.390000  65.590000 ;
      RECT  3.000000  65.590000 66.240000  65.740000 ;
      RECT  3.000000  65.590000 66.240000  65.740000 ;
      RECT  3.000000  65.740000 66.085000  65.890000 ;
      RECT  3.000000  65.740000 66.085000  65.890000 ;
      RECT  3.000000  65.890000 65.940000  66.040000 ;
      RECT  3.000000  65.890000 65.940000  66.040000 ;
      RECT  3.000000  66.040000 65.785000  66.190000 ;
      RECT  3.000000  66.040000 65.785000  66.190000 ;
      RECT  3.000000  66.190000 65.640000  66.340000 ;
      RECT  3.000000  66.190000 65.640000  66.340000 ;
      RECT  3.000000  66.340000 65.485000  66.490000 ;
      RECT  3.000000  66.340000 65.485000  66.490000 ;
      RECT  3.000000  66.490000 65.335000  66.640000 ;
      RECT  3.000000  66.490000 65.335000  66.640000 ;
      RECT  3.000000  66.640000 65.190000  66.790000 ;
      RECT  3.000000  66.640000 65.190000  66.790000 ;
      RECT  3.000000  66.790000 65.035000  66.940000 ;
      RECT  3.000000  66.790000 65.035000  66.940000 ;
      RECT  3.000000  66.940000 64.890000  67.090000 ;
      RECT  3.000000  66.940000 64.890000  67.090000 ;
      RECT  3.000000  67.090000 64.735000  67.240000 ;
      RECT  3.000000  67.090000 64.735000  67.240000 ;
      RECT  3.000000  67.240000 64.585000  67.390000 ;
      RECT  3.000000  67.240000 64.585000  67.390000 ;
      RECT  3.000000  67.390000 64.440000  67.540000 ;
      RECT  3.000000  67.390000 64.440000  67.540000 ;
      RECT  3.000000  67.540000 64.285000  67.690000 ;
      RECT  3.000000  67.540000 64.285000  67.690000 ;
      RECT  3.000000  67.690000 64.140000  67.840000 ;
      RECT  3.000000  67.690000 64.140000  67.840000 ;
      RECT  3.000000  67.840000 63.990000  67.990000 ;
      RECT  3.000000  67.840000 63.990000  67.990000 ;
      RECT  3.000000  67.990000 63.840000  68.140000 ;
      RECT  3.000000  67.990000 63.840000  68.140000 ;
      RECT  3.000000  68.140000 63.690000  68.290000 ;
      RECT  3.000000  68.140000 63.690000  68.290000 ;
      RECT  3.000000  68.290000 63.540000  68.440000 ;
      RECT  3.000000  68.290000 63.540000  68.440000 ;
      RECT  3.000000  68.440000 63.390000  68.590000 ;
      RECT  3.000000  68.440000 63.390000  68.590000 ;
      RECT  3.000000  68.590000 63.240000  68.740000 ;
      RECT  3.000000  68.590000 63.240000  68.740000 ;
      RECT  3.000000  68.740000 63.090000  68.890000 ;
      RECT  3.000000  68.740000 63.090000  68.890000 ;
      RECT  3.000000  68.890000 62.940000  69.040000 ;
      RECT  3.000000  68.890000 62.940000  69.040000 ;
      RECT  3.000000  69.040000 62.790000  69.190000 ;
      RECT  3.000000  69.040000 62.790000  69.190000 ;
      RECT  3.000000  69.190000 62.640000  69.340000 ;
      RECT  3.000000  69.190000 62.640000  69.340000 ;
      RECT  3.000000  69.340000 62.490000  69.490000 ;
      RECT  3.000000  69.340000 62.490000  69.490000 ;
      RECT  3.000000  69.490000 62.340000  69.640000 ;
      RECT  3.000000  69.490000 62.340000  69.640000 ;
      RECT  3.000000  69.640000 62.190000  69.790000 ;
      RECT  3.000000  69.640000 62.190000  69.790000 ;
      RECT  3.000000  69.790000 62.040000  69.940000 ;
      RECT  3.000000  69.790000 62.040000  69.940000 ;
      RECT  3.000000  69.940000 61.890000  70.090000 ;
      RECT  3.000000  69.940000 61.890000  70.090000 ;
      RECT  3.000000  70.090000 61.740000  70.240000 ;
      RECT  3.000000  70.090000 61.740000  70.240000 ;
      RECT  3.000000  70.240000 61.590000  70.390000 ;
      RECT  3.000000  70.240000 61.590000  70.390000 ;
      RECT  3.000000  70.390000 61.460000  70.520000 ;
      RECT  3.000000  70.390000 61.460000  70.520000 ;
      RECT  3.000000  70.520000 61.460000  98.045000 ;
      RECT  3.000000  98.045000 72.000000 197.000000 ;
      RECT  3.370000   3.005000  8.000000  15.620000 ;
      RECT  3.370000  15.620000  6.375000  17.245000 ;
      RECT  6.375000  34.525000 25.680000  37.525000 ;
      RECT  6.375000  37.525000 25.675000  37.530000 ;
      RECT  7.595000  17.745000 71.890000  31.170000 ;
      RECT  7.595000  31.170000 71.890000  33.095000 ;
      RECT  7.695000  17.785000 12.325000  28.125000 ;
      RECT  7.695000  28.125000 25.675000  29.990000 ;
      RECT  7.695000  29.990000 25.680000  31.130000 ;
      RECT  7.820000  17.660000 71.790000  17.785000 ;
      RECT  7.845000  31.130000 71.790000  31.280000 ;
      RECT  7.970000  17.510000 71.790000  17.660000 ;
      RECT  7.995000  31.280000 71.790000  31.430000 ;
      RECT  8.120000  17.360000 71.790000  17.510000 ;
      RECT  8.145000  31.430000 71.790000  31.580000 ;
      RECT  8.270000  17.210000 71.790000  17.360000 ;
      RECT  8.295000  31.580000 71.790000  31.730000 ;
      RECT  8.420000  17.060000 71.790000  17.210000 ;
      RECT  8.445000  31.730000 71.790000  31.880000 ;
      RECT  8.570000  16.910000 71.790000  17.060000 ;
      RECT  8.595000  31.880000 71.790000  32.030000 ;
      RECT  8.720000  16.760000 71.790000  16.910000 ;
      RECT  8.745000  32.030000 71.790000  32.180000 ;
      RECT  8.870000  16.610000 71.790000  16.760000 ;
      RECT  8.895000  32.180000 71.790000  32.330000 ;
      RECT  9.020000  16.460000 71.790000  16.610000 ;
      RECT  9.045000  32.330000 71.790000  32.480000 ;
      RECT  9.170000  16.310000 71.790000  16.460000 ;
      RECT  9.195000  32.480000 71.790000  32.630000 ;
      RECT  9.220000   0.000000 16.945000   3.435000 ;
      RECT  9.220000   3.435000 19.775000   7.275000 ;
      RECT  9.220000   7.275000 22.605000  10.105000 ;
      RECT  9.220000  10.105000 22.605000  12.565000 ;
      RECT  9.220000  12.565000 27.870000  15.070000 ;
      RECT  9.220000  15.070000 71.890000  16.120000 ;
      RECT  9.220000  16.120000 71.890000  17.745000 ;
      RECT  9.320000   0.000000 16.845000   7.315000 ;
      RECT  9.320000   0.000000 16.845000  10.145000 ;
      RECT  9.320000   3.535000 19.675000  12.665000 ;
      RECT  9.320000   7.315000 19.675000   7.465000 ;
      RECT  9.320000   7.465000 19.825000   7.615000 ;
      RECT  9.320000   7.615000 19.975000   7.765000 ;
      RECT  9.320000   7.765000 20.125000   7.915000 ;
      RECT  9.320000   7.915000 20.275000   8.065000 ;
      RECT  9.320000   8.065000 20.425000   8.215000 ;
      RECT  9.320000   8.215000 20.575000   8.365000 ;
      RECT  9.320000   8.365000 20.725000   8.515000 ;
      RECT  9.320000   8.515000 20.875000   8.665000 ;
      RECT  9.320000   8.665000 21.025000   8.815000 ;
      RECT  9.320000   8.815000 21.175000   8.965000 ;
      RECT  9.320000   8.965000 21.325000   9.115000 ;
      RECT  9.320000   9.115000 21.475000   9.265000 ;
      RECT  9.320000   9.265000 21.625000   9.415000 ;
      RECT  9.320000   9.415000 21.775000   9.565000 ;
      RECT  9.320000   9.565000 21.925000   9.715000 ;
      RECT  9.320000   9.715000 22.075000   9.865000 ;
      RECT  9.320000   9.865000 22.225000  10.015000 ;
      RECT  9.320000  10.015000 22.375000  10.145000 ;
      RECT  9.320000  12.665000 12.325000  17.785000 ;
      RECT  9.320000  16.160000 71.790000  16.310000 ;
      RECT  9.345000  32.630000 71.790000  32.780000 ;
      RECT  9.495000  32.780000 71.790000  32.930000 ;
      RECT  9.560000  32.930000 71.790000  32.995000 ;
      RECT 10.695000  19.030000 68.785000  29.885000 ;
      RECT 10.750000  29.885000 68.785000  29.940000 ;
      RECT 10.750000  29.885000 68.785000  29.940000 ;
      RECT 10.805000  18.920000 68.785000  19.030000 ;
      RECT 10.805000  18.920000 68.785000  19.030000 ;
      RECT 10.805000  29.940000 68.785000  29.995000 ;
      RECT 10.805000  29.940000 68.785000  29.995000 ;
      RECT 10.955000  18.770000 68.785000  18.920000 ;
      RECT 10.955000  18.770000 68.785000  18.920000 ;
      RECT 11.105000  18.620000 68.785000  18.770000 ;
      RECT 11.105000  18.620000 68.785000  18.770000 ;
      RECT 11.255000  18.470000 68.785000  18.620000 ;
      RECT 11.255000  18.470000 68.785000  18.620000 ;
      RECT 11.405000  18.320000 68.785000  18.470000 ;
      RECT 11.405000  18.320000 68.785000  18.470000 ;
      RECT 11.555000  18.170000 68.785000  18.320000 ;
      RECT 11.555000  18.170000 68.785000  18.320000 ;
      RECT 11.570000  18.155000 24.770000  18.170000 ;
      RECT 11.570000  18.155000 24.770000  18.170000 ;
      RECT 11.720000  18.005000 24.770000  18.155000 ;
      RECT 11.720000  18.005000 24.770000  18.155000 ;
      RECT 11.870000  17.855000 24.770000  18.005000 ;
      RECT 11.870000  17.855000 24.770000  18.005000 ;
      RECT 12.020000  17.705000 24.770000  17.855000 ;
      RECT 12.020000  17.705000 24.770000  17.855000 ;
      RECT 12.170000  17.555000 24.770000  17.705000 ;
      RECT 12.170000  17.555000 24.770000  17.705000 ;
      RECT 12.320000   3.000000 13.845000   6.535000 ;
      RECT 12.320000   6.535000 16.670000   8.560000 ;
      RECT 12.320000   8.560000 16.670000   8.710000 ;
      RECT 12.320000   8.560000 16.670000   8.710000 ;
      RECT 12.320000   8.710000 16.825000   8.860000 ;
      RECT 12.320000   8.710000 16.825000   8.860000 ;
      RECT 12.320000   8.860000 16.970000   9.010000 ;
      RECT 12.320000   8.860000 16.970000   9.010000 ;
      RECT 12.320000   9.010000 17.125000   9.160000 ;
      RECT 12.320000   9.010000 17.125000   9.160000 ;
      RECT 12.320000   9.160000 17.275000   9.310000 ;
      RECT 12.320000   9.160000 17.275000   9.310000 ;
      RECT 12.320000   9.310000 17.420000   9.460000 ;
      RECT 12.320000   9.310000 17.420000   9.460000 ;
      RECT 12.320000   9.460000 17.575000   9.610000 ;
      RECT 12.320000   9.460000 17.575000   9.610000 ;
      RECT 12.320000   9.610000 17.720000   9.760000 ;
      RECT 12.320000   9.610000 17.720000   9.760000 ;
      RECT 12.320000   9.760000 17.875000   9.910000 ;
      RECT 12.320000   9.760000 17.875000   9.910000 ;
      RECT 12.320000   9.910000 18.025000  10.060000 ;
      RECT 12.320000   9.910000 18.025000  10.060000 ;
      RECT 12.320000  10.060000 18.170000  10.210000 ;
      RECT 12.320000  10.060000 18.170000  10.210000 ;
      RECT 12.320000  10.210000 18.325000  10.360000 ;
      RECT 12.320000  10.210000 18.325000  10.360000 ;
      RECT 12.320000  10.360000 18.470000  10.510000 ;
      RECT 12.320000  10.360000 18.470000  10.510000 ;
      RECT 12.320000  10.510000 18.625000  10.660000 ;
      RECT 12.320000  10.510000 18.625000  10.660000 ;
      RECT 12.320000  10.660000 18.775000  10.810000 ;
      RECT 12.320000  10.660000 18.775000  10.810000 ;
      RECT 12.320000  10.810000 18.920000  10.960000 ;
      RECT 12.320000  10.810000 18.920000  10.960000 ;
      RECT 12.320000  10.960000 19.075000  11.110000 ;
      RECT 12.320000  10.960000 19.075000  11.110000 ;
      RECT 12.320000  11.110000 19.220000  11.260000 ;
      RECT 12.320000  11.110000 19.220000  11.260000 ;
      RECT 12.320000  11.260000 19.375000  11.390000 ;
      RECT 12.320000  11.260000 19.375000  11.390000 ;
      RECT 12.320000  11.390000 19.505000  15.665000 ;
      RECT 12.320000  15.665000 24.770000  17.405000 ;
      RECT 12.320000  17.405000 24.770000  17.555000 ;
      RECT 12.320000  17.405000 24.770000  17.555000 ;
      RECT 19.210000   0.000000 19.775000   3.435000 ;
      RECT 19.310000   0.000000 19.675000   3.535000 ;
      RECT 19.500000  10.145000 22.505000  12.665000 ;
      RECT 19.500000  12.665000 27.770000  15.170000 ;
      RECT 19.505000  15.170000 32.305000  18.170000 ;
      RECT 19.505000  18.170000 32.300000  18.175000 ;
      RECT 21.525000   0.000000 28.635000   6.545000 ;
      RECT 21.525000   6.545000 28.635000   9.370000 ;
      RECT 21.625000   0.000000 28.535000   3.005000 ;
      RECT 21.625000   3.005000 24.630000   3.500000 ;
      RECT 21.625000   3.500000 28.535000   6.505000 ;
      RECT 21.775000   6.505000 28.535000   6.655000 ;
      RECT 21.925000   6.655000 28.535000   6.805000 ;
      RECT 22.075000   6.805000 28.535000   6.955000 ;
      RECT 22.225000   6.955000 28.535000   7.105000 ;
      RECT 22.375000   7.105000 28.535000   7.255000 ;
      RECT 22.525000   7.255000 28.535000   7.405000 ;
      RECT 22.575000  33.095000 71.890000  34.425000 ;
      RECT 22.675000   7.405000 28.535000   7.555000 ;
      RECT 22.675000  31.130000 25.680000  34.525000 ;
      RECT 22.825000   7.555000 28.535000   7.705000 ;
      RECT 22.975000   7.705000 28.535000   7.855000 ;
      RECT 23.125000   7.855000 28.535000   8.005000 ;
      RECT 23.275000   8.005000 28.535000   8.155000 ;
      RECT 23.425000   8.155000 28.535000   8.305000 ;
      RECT 23.575000   8.305000 28.535000   8.455000 ;
      RECT 23.725000   8.455000 28.535000   8.605000 ;
      RECT 23.875000   8.605000 28.535000   8.755000 ;
      RECT 24.025000   8.755000 28.535000   8.905000 ;
      RECT 24.175000   8.905000 28.535000   9.055000 ;
      RECT 24.325000   9.055000 28.535000   9.205000 ;
      RECT 24.350000   9.370000 28.635000   9.720000 ;
      RECT 24.350000   9.720000 27.870000  10.485000 ;
      RECT 24.350000  10.485000 27.870000  12.565000 ;
      RECT 24.450000   9.205000 28.535000   9.330000 ;
      RECT 24.450000   9.330000 28.535000   9.680000 ;
      RECT 24.450000   9.680000 27.770000  12.665000 ;
      RECT 24.450000   9.680000 28.385000   9.830000 ;
      RECT 24.450000   9.830000 28.235000   9.980000 ;
      RECT 24.450000   9.980000 28.085000  10.130000 ;
      RECT 24.450000  10.130000 27.935000  10.280000 ;
      RECT 24.450000  10.280000 27.785000  10.430000 ;
      RECT 24.450000  10.430000 27.770000  10.445000 ;
      RECT 24.625000   3.000000 25.535000   5.260000 ;
      RECT 24.625000   3.000000 25.535000   5.260000 ;
      RECT 24.770000  18.175000 32.300000  20.790000 ;
      RECT 25.530000   3.005000 28.535000   3.500000 ;
      RECT 25.675000  29.990000 68.785000  37.525000 ;
      RECT 29.200000  11.035000 71.890000  15.070000 ;
      RECT 29.300000  11.075000 33.065000  14.080000 ;
      RECT 29.300000  14.080000 32.305000  15.170000 ;
      RECT 29.315000  11.060000 71.790000  11.075000 ;
      RECT 29.465000  10.910000 71.790000  11.060000 ;
      RECT 29.615000  10.760000 71.790000  10.910000 ;
      RECT 29.765000  10.610000 71.790000  10.760000 ;
      RECT 29.915000  10.460000 71.790000  10.610000 ;
      RECT 29.965000   0.000000 71.890000  10.270000 ;
      RECT 29.965000  10.270000 71.890000  11.035000 ;
      RECT 30.065000   0.000000 71.790000   3.005000 ;
      RECT 30.065000   3.005000 33.070000  11.075000 ;
      RECT 30.065000  10.310000 71.790000  10.460000 ;
      RECT 32.300000  12.320000 68.785000  18.170000 ;
      RECT 32.315000  12.305000 68.785000  12.320000 ;
      RECT 32.315000  12.305000 68.785000  12.320000 ;
      RECT 32.465000  12.155000 68.785000  12.305000 ;
      RECT 32.465000  12.155000 68.785000  12.305000 ;
      RECT 32.615000  12.005000 68.785000  12.155000 ;
      RECT 32.615000  12.005000 68.785000  12.155000 ;
      RECT 32.765000  11.855000 68.785000  12.005000 ;
      RECT 32.765000  11.855000 68.785000  12.005000 ;
      RECT 32.915000  11.705000 68.785000  11.855000 ;
      RECT 32.915000  11.705000 68.785000  11.855000 ;
      RECT 33.065000   3.000000 68.785000  11.555000 ;
      RECT 33.065000  11.555000 68.785000  11.705000 ;
      RECT 33.065000  11.555000 68.785000  11.705000 ;
      RECT 61.455000  71.765000 64.460000  95.045000 ;
      RECT 61.460000  95.045000 69.390000  98.050000 ;
      RECT 66.290000  72.525000 75.000000  94.945000 ;
      RECT 66.390000  72.565000 70.635000  75.570000 ;
      RECT 66.390000  75.570000 69.395000  95.045000 ;
      RECT 66.525000  72.430000 75.000000  72.565000 ;
      RECT 66.675000  72.280000 75.000000  72.430000 ;
      RECT 66.825000  72.130000 75.000000  72.280000 ;
      RECT 66.975000  71.980000 75.000000  72.130000 ;
      RECT 67.125000  71.830000 75.000000  71.980000 ;
      RECT 67.275000  71.680000 75.000000  71.830000 ;
      RECT 67.425000  71.530000 75.000000  71.680000 ;
      RECT 67.545000  61.430000 71.790000  64.435000 ;
      RECT 67.575000  71.380000 75.000000  71.530000 ;
      RECT 67.725000  71.230000 75.000000  71.380000 ;
      RECT 67.875000  71.080000 75.000000  71.230000 ;
      RECT 68.025000  70.930000 75.000000  71.080000 ;
      RECT 68.175000  70.780000 75.000000  70.930000 ;
      RECT 68.325000  70.630000 75.000000  70.780000 ;
      RECT 68.475000  70.480000 75.000000  70.630000 ;
      RECT 68.625000  70.330000 75.000000  70.480000 ;
      RECT 68.775000  70.180000 75.000000  70.330000 ;
      RECT 68.785000   3.005000 71.790000  61.430000 ;
      RECT 68.925000  70.030000 75.000000  70.180000 ;
      RECT 69.075000  69.880000 75.000000  70.030000 ;
      RECT 69.225000  69.730000 75.000000  69.880000 ;
      RECT 69.375000  69.580000 75.000000  69.730000 ;
      RECT 69.390000  73.810000 72.000000  98.045000 ;
      RECT 69.445000  73.755000 72.000000  73.810000 ;
      RECT 69.445000  73.755000 72.000000  73.810000 ;
      RECT 69.525000  69.430000 75.000000  69.580000 ;
      RECT 69.595000  73.605000 72.000000  73.755000 ;
      RECT 69.595000  73.605000 72.000000  73.755000 ;
      RECT 69.675000  69.280000 75.000000  69.430000 ;
      RECT 69.745000  73.455000 72.000000  73.605000 ;
      RECT 69.745000  73.455000 72.000000  73.605000 ;
      RECT 69.825000  69.130000 75.000000  69.280000 ;
      RECT 69.895000  73.305000 72.000000  73.455000 ;
      RECT 69.895000  73.305000 72.000000  73.455000 ;
      RECT 69.975000  68.980000 75.000000  69.130000 ;
      RECT 70.045000  73.155000 72.000000  73.305000 ;
      RECT 70.045000  73.155000 72.000000  73.305000 ;
      RECT 70.125000  68.830000 75.000000  68.980000 ;
      RECT 70.195000  73.005000 72.000000  73.155000 ;
      RECT 70.195000  73.005000 72.000000  73.155000 ;
      RECT 70.275000  68.680000 75.000000  68.830000 ;
      RECT 70.345000  72.855000 72.000000  73.005000 ;
      RECT 70.345000  72.855000 72.000000  73.005000 ;
      RECT 70.425000  68.530000 75.000000  68.680000 ;
      RECT 70.495000  72.705000 72.000000  72.855000 ;
      RECT 70.495000  72.705000 72.000000  72.855000 ;
      RECT 70.575000  68.380000 75.000000  68.530000 ;
      RECT 70.645000  72.555000 72.000000  72.705000 ;
      RECT 70.645000  72.555000 72.000000  72.705000 ;
      RECT 70.725000  68.230000 75.000000  68.380000 ;
      RECT 70.795000  72.405000 72.000000  72.555000 ;
      RECT 70.795000  72.405000 72.000000  72.555000 ;
      RECT 70.875000  68.080000 75.000000  68.230000 ;
      RECT 70.945000  72.255000 72.000000  72.405000 ;
      RECT 70.945000  72.255000 72.000000  72.405000 ;
      RECT 71.025000  67.930000 75.000000  68.080000 ;
      RECT 71.095000  72.105000 72.000000  72.255000 ;
      RECT 71.095000  72.105000 72.000000  72.255000 ;
      RECT 71.175000  67.780000 75.000000  67.930000 ;
      RECT 71.245000  71.955000 72.000000  72.105000 ;
      RECT 71.245000  71.955000 72.000000  72.105000 ;
      RECT 71.325000  67.630000 75.000000  67.780000 ;
      RECT 71.395000  71.805000 72.000000  71.955000 ;
      RECT 71.395000  71.805000 72.000000  71.955000 ;
      RECT 71.475000  67.480000 75.000000  67.630000 ;
      RECT 71.545000  71.655000 72.000000  71.805000 ;
      RECT 71.545000  71.655000 72.000000  71.805000 ;
      RECT 71.625000  67.330000 75.000000  67.480000 ;
      RECT 71.695000  71.505000 72.000000  71.655000 ;
      RECT 71.695000  71.505000 72.000000  71.655000 ;
      RECT 71.775000  67.180000 75.000000  67.330000 ;
      RECT 71.845000  71.355000 72.000000  71.505000 ;
      RECT 71.845000  71.355000 72.000000  71.505000 ;
      RECT 71.925000  67.030000 75.000000  67.180000 ;
      RECT 71.995000  72.565000 75.000000 196.995000 ;
      RECT 72.075000  66.880000 75.000000  67.030000 ;
      RECT 72.225000  66.730000 75.000000  66.880000 ;
      RECT 72.375000  66.580000 75.000000  66.730000 ;
      RECT 72.525000  66.430000 75.000000  66.580000 ;
      RECT 72.675000  66.280000 75.000000  66.430000 ;
      RECT 72.825000  66.130000 75.000000  66.280000 ;
      RECT 72.975000  65.980000 75.000000  66.130000 ;
      RECT 73.125000  65.830000 75.000000  65.980000 ;
      RECT 73.275000  65.680000 75.000000  65.830000 ;
      RECT 73.425000  65.530000 75.000000  65.680000 ;
      RECT 73.560000   0.000000 75.000000  49.195000 ;
      RECT 73.560000  49.195000 75.000000  49.860000 ;
      RECT 73.575000  65.380000 75.000000  65.530000 ;
      RECT 73.660000   0.000000 75.000000  49.155000 ;
      RECT 73.725000  65.230000 75.000000  65.380000 ;
      RECT 73.810000  49.155000 75.000000  49.305000 ;
      RECT 73.875000  65.080000 75.000000  65.230000 ;
      RECT 73.960000  49.305000 75.000000  49.455000 ;
      RECT 74.025000  64.930000 75.000000  65.080000 ;
      RECT 74.110000  49.455000 75.000000  49.605000 ;
      RECT 74.175000  64.780000 75.000000  64.930000 ;
      RECT 74.225000  49.860000 75.000000  64.590000 ;
      RECT 74.225000  64.590000 75.000000  72.525000 ;
      RECT 74.260000  49.605000 75.000000  49.755000 ;
      RECT 74.325000  49.755000 75.000000  49.820000 ;
      RECT 74.325000  49.820000 75.000000  64.630000 ;
      RECT 74.325000  64.630000 75.000000  64.780000 ;
    LAYER met4 ;
      RECT  0.000000   0.000000  1.670000   1.635000 ;
      RECT  0.000000   0.000000 75.000000   1.635000 ;
      RECT  0.000000   7.885000  1.670000   8.485000 ;
      RECT  0.000000   7.885000 75.000000   8.485000 ;
      RECT  0.000000  13.935000  1.365000  14.535000 ;
      RECT  0.000000  13.935000 75.000000  14.535000 ;
      RECT  0.000000  18.785000  1.365000  19.385000 ;
      RECT  0.000000  18.785000 75.000000  19.385000 ;
      RECT  0.000000  24.835000  1.670000  25.435000 ;
      RECT  0.000000  24.835000 75.000000  25.435000 ;
      RECT  0.000000  30.885000  1.670000  31.485000 ;
      RECT  0.000000  30.885000 75.000000  31.485000 ;
      RECT  0.000000  35.735000  1.670000  36.335000 ;
      RECT  0.000000  35.735000 75.000000  36.335000 ;
      RECT  0.000000  40.585000  1.670000  41.185000 ;
      RECT  0.000000  40.585000 75.000000  41.185000 ;
      RECT  0.000000  46.635000  1.670000  47.335000 ;
      RECT  0.000000  46.635000 75.000000  47.435000 ;
      RECT  0.000000  57.035000 75.000000  57.835000 ;
      RECT  0.000000  57.135000  1.670000  57.835000 ;
      RECT  0.000000  63.085000  1.670000  63.685000 ;
      RECT  0.000000  63.085000 75.000000  63.685000 ;
      RECT  0.000000  68.935000  1.670000  69.635000 ;
      RECT  0.000000  68.935000 75.000000  69.635000 ;
      RECT  0.000000  95.400000 75.000000 175.385000 ;
      RECT  1.365000  13.935000 73.635000  19.385000 ;
      RECT  1.570000  47.435000 73.430000  57.035000 ;
      RECT  1.670000   0.000000 73.330000  13.935000 ;
      RECT  1.670000  19.385000 73.330000  41.230000 ;
      RECT  1.670000  36.335000 73.330000  41.230000 ;
      RECT  1.670000  36.335000 73.330000  41.230000 ;
      RECT  1.670000  41.185000 75.000000  41.255000 ;
      RECT  1.670000  41.230000 73.255000  41.255000 ;
      RECT  1.670000  46.570000 73.255000  46.590000 ;
      RECT  1.670000  46.570000 73.255000  57.135000 ;
      RECT  1.670000  46.570000 75.000000  46.635000 ;
      RECT  1.670000  46.590000 73.330000  57.135000 ;
      RECT  1.670000  46.590000 73.330000  57.135000 ;
      RECT  1.670000  46.590000 73.330000  95.400000 ;
      RECT  1.670000 175.385000 73.330000 200.000000 ;
      RECT  4.120000  41.230000 73.255000  46.570000 ;
      RECT  4.120000  41.255000 73.255000  46.570000 ;
      RECT  4.120000  41.255000 73.255000  57.135000 ;
      RECT  4.120000  41.255000 75.000000  41.285000 ;
      RECT  4.120000  41.285000 73.430000  41.330000 ;
      RECT  4.120000  41.330000 73.355000  46.490000 ;
      RECT  4.120000  46.490000 73.430000  46.535000 ;
      RECT  4.120000  46.535000 75.000000  46.570000 ;
      RECT 73.330000   0.000000 75.000000   1.635000 ;
      RECT 73.330000   7.885000 75.000000   8.485000 ;
      RECT 73.330000  24.835000 75.000000  25.435000 ;
      RECT 73.330000  30.885000 75.000000  31.485000 ;
      RECT 73.330000  35.735000 75.000000  36.335000 ;
      RECT 73.330000  40.585000 75.000000  41.185000 ;
      RECT 73.330000  46.635000 75.000000  47.335000 ;
      RECT 73.330000  57.135000 75.000000  57.835000 ;
      RECT 73.330000  63.085000 75.000000  63.685000 ;
      RECT 73.330000  68.935000 75.000000  69.635000 ;
      RECT 73.635000  13.935000 75.000000  14.535000 ;
      RECT 73.635000  18.785000 75.000000  19.385000 ;
    LAYER met5 ;
      RECT  0.000000   0.000000 75.000000   1.335000 ;
      RECT  0.000000  36.035000 75.000000  36.040000 ;
      RECT  0.000000  95.785000 75.000000 126.315000 ;
      RECT  0.000000 126.315000 28.895000 146.425000 ;
      RECT  0.000000 146.425000 75.000000 174.985000 ;
      RECT  1.765000  14.235000 73.235000  19.085000 ;
      RECT  2.070000   1.335000 72.930000  14.235000 ;
      RECT  2.070000  19.085000 72.930000  95.785000 ;
      RECT  2.070000 174.985000 72.930000 200.000000 ;
      RECT 42.790000 126.315000 75.000000 146.425000 ;
  END
END sky130_fd_io__top_xres4v2
END LIBRARY
