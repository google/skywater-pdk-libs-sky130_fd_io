# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__overlay_vssd_lvc
  CLASS BLOCK ;
  FOREIGN sky130_fd_io__overlay_vssd_lvc ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  75.00000 BY  198.0000 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.530000 39.600000 0.850000 39.920000 ;
      LAYER met4 ;
        RECT 0.530000 39.600000 0.850000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 40.030000 0.850000 40.350000 ;
      LAYER met4 ;
        RECT 0.530000 40.030000 0.850000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 40.460000 0.850000 40.780000 ;
      LAYER met4 ;
        RECT 0.530000 40.460000 0.850000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 40.890000 0.850000 41.210000 ;
      LAYER met4 ;
        RECT 0.530000 40.890000 0.850000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 41.320000 0.850000 41.640000 ;
      LAYER met4 ;
        RECT 0.530000 41.320000 0.850000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 41.750000 0.850000 42.070000 ;
      LAYER met4 ;
        RECT 0.530000 41.750000 0.850000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 42.180000 0.850000 42.500000 ;
      LAYER met4 ;
        RECT 0.530000 42.180000 0.850000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 42.610000 0.850000 42.930000 ;
      LAYER met4 ;
        RECT 0.530000 42.610000 0.850000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 43.040000 0.850000 43.360000 ;
      LAYER met4 ;
        RECT 0.530000 43.040000 0.850000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 43.470000 0.850000 43.790000 ;
      LAYER met4 ;
        RECT 0.530000 43.470000 0.850000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 43.900000 0.850000 44.220000 ;
      LAYER met4 ;
        RECT 0.530000 43.900000 0.850000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 39.600000 1.255000 39.920000 ;
      LAYER met4 ;
        RECT 0.935000 39.600000 1.255000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 40.030000 1.255000 40.350000 ;
      LAYER met4 ;
        RECT 0.935000 40.030000 1.255000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 40.460000 1.255000 40.780000 ;
      LAYER met4 ;
        RECT 0.935000 40.460000 1.255000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 40.890000 1.255000 41.210000 ;
      LAYER met4 ;
        RECT 0.935000 40.890000 1.255000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 41.320000 1.255000 41.640000 ;
      LAYER met4 ;
        RECT 0.935000 41.320000 1.255000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 41.750000 1.255000 42.070000 ;
      LAYER met4 ;
        RECT 0.935000 41.750000 1.255000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 42.180000 1.255000 42.500000 ;
      LAYER met4 ;
        RECT 0.935000 42.180000 1.255000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 42.610000 1.255000 42.930000 ;
      LAYER met4 ;
        RECT 0.935000 42.610000 1.255000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 43.040000 1.255000 43.360000 ;
      LAYER met4 ;
        RECT 0.935000 43.040000 1.255000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 43.470000 1.255000 43.790000 ;
      LAYER met4 ;
        RECT 0.935000 43.470000 1.255000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 43.900000 1.255000 44.220000 ;
      LAYER met4 ;
        RECT 0.935000 43.900000 1.255000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.340000 39.600000 1.660000 39.920000 ;
      LAYER met4 ;
        RECT 1.340000 39.600000 1.660000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.340000 40.030000 1.660000 40.350000 ;
      LAYER met4 ;
        RECT 1.340000 40.030000 1.660000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.340000 40.460000 1.660000 40.780000 ;
      LAYER met4 ;
        RECT 1.340000 40.460000 1.660000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.340000 40.890000 1.660000 41.210000 ;
      LAYER met4 ;
        RECT 1.340000 40.890000 1.660000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.340000 41.320000 1.660000 41.640000 ;
      LAYER met4 ;
        RECT 1.340000 41.320000 1.660000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.340000 41.750000 1.660000 42.070000 ;
      LAYER met4 ;
        RECT 1.340000 41.750000 1.660000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.340000 42.180000 1.660000 42.500000 ;
      LAYER met4 ;
        RECT 1.340000 42.180000 1.660000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.340000 42.610000 1.660000 42.930000 ;
      LAYER met4 ;
        RECT 1.340000 42.610000 1.660000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.340000 43.040000 1.660000 43.360000 ;
      LAYER met4 ;
        RECT 1.340000 43.040000 1.660000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.340000 43.470000 1.660000 43.790000 ;
      LAYER met4 ;
        RECT 1.340000 43.470000 1.660000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.340000 43.900000 1.660000 44.220000 ;
      LAYER met4 ;
        RECT 1.340000 43.900000 1.660000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.745000 39.600000 2.065000 39.920000 ;
      LAYER met4 ;
        RECT 1.745000 39.600000 2.065000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.745000 40.030000 2.065000 40.350000 ;
      LAYER met4 ;
        RECT 1.745000 40.030000 2.065000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.745000 40.460000 2.065000 40.780000 ;
      LAYER met4 ;
        RECT 1.745000 40.460000 2.065000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.745000 40.890000 2.065000 41.210000 ;
      LAYER met4 ;
        RECT 1.745000 40.890000 2.065000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.745000 41.320000 2.065000 41.640000 ;
      LAYER met4 ;
        RECT 1.745000 41.320000 2.065000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.745000 41.750000 2.065000 42.070000 ;
      LAYER met4 ;
        RECT 1.745000 41.750000 2.065000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.745000 42.180000 2.065000 42.500000 ;
      LAYER met4 ;
        RECT 1.745000 42.180000 2.065000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.745000 42.610000 2.065000 42.930000 ;
      LAYER met4 ;
        RECT 1.745000 42.610000 2.065000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.745000 43.040000 2.065000 43.360000 ;
      LAYER met4 ;
        RECT 1.745000 43.040000 2.065000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.745000 43.470000 2.065000 43.790000 ;
      LAYER met4 ;
        RECT 1.745000 43.470000 2.065000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.745000 43.900000 2.065000 44.220000 ;
      LAYER met4 ;
        RECT 1.745000 43.900000 2.065000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.150000 39.600000 10.470000 39.920000 ;
      LAYER met4 ;
        RECT 10.150000 39.600000 10.470000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.150000 40.030000 10.470000 40.350000 ;
      LAYER met4 ;
        RECT 10.150000 40.030000 10.470000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.150000 40.460000 10.470000 40.780000 ;
      LAYER met4 ;
        RECT 10.150000 40.460000 10.470000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.150000 40.890000 10.470000 41.210000 ;
      LAYER met4 ;
        RECT 10.150000 40.890000 10.470000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.150000 41.320000 10.470000 41.640000 ;
      LAYER met4 ;
        RECT 10.150000 41.320000 10.470000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.150000 41.750000 10.470000 42.070000 ;
      LAYER met4 ;
        RECT 10.150000 41.750000 10.470000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.150000 42.180000 10.470000 42.500000 ;
      LAYER met4 ;
        RECT 10.150000 42.180000 10.470000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.150000 42.610000 10.470000 42.930000 ;
      LAYER met4 ;
        RECT 10.150000 42.610000 10.470000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.150000 43.040000 10.470000 43.360000 ;
      LAYER met4 ;
        RECT 10.150000 43.040000 10.470000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.150000 43.470000 10.470000 43.790000 ;
      LAYER met4 ;
        RECT 10.150000 43.470000 10.470000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.150000 43.900000 10.470000 44.220000 ;
      LAYER met4 ;
        RECT 10.150000 43.900000 10.470000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550000 39.600000 10.870000 39.920000 ;
      LAYER met4 ;
        RECT 10.550000 39.600000 10.870000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550000 40.030000 10.870000 40.350000 ;
      LAYER met4 ;
        RECT 10.550000 40.030000 10.870000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550000 40.460000 10.870000 40.780000 ;
      LAYER met4 ;
        RECT 10.550000 40.460000 10.870000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550000 40.890000 10.870000 41.210000 ;
      LAYER met4 ;
        RECT 10.550000 40.890000 10.870000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550000 41.320000 10.870000 41.640000 ;
      LAYER met4 ;
        RECT 10.550000 41.320000 10.870000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550000 41.750000 10.870000 42.070000 ;
      LAYER met4 ;
        RECT 10.550000 41.750000 10.870000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550000 42.180000 10.870000 42.500000 ;
      LAYER met4 ;
        RECT 10.550000 42.180000 10.870000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550000 42.610000 10.870000 42.930000 ;
      LAYER met4 ;
        RECT 10.550000 42.610000 10.870000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550000 43.040000 10.870000 43.360000 ;
      LAYER met4 ;
        RECT 10.550000 43.040000 10.870000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550000 43.470000 10.870000 43.790000 ;
      LAYER met4 ;
        RECT 10.550000 43.470000 10.870000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550000 43.900000 10.870000 44.220000 ;
      LAYER met4 ;
        RECT 10.550000 43.900000 10.870000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950000 39.600000 11.270000 39.920000 ;
      LAYER met4 ;
        RECT 10.950000 39.600000 11.270000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950000 40.030000 11.270000 40.350000 ;
      LAYER met4 ;
        RECT 10.950000 40.030000 11.270000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950000 40.460000 11.270000 40.780000 ;
      LAYER met4 ;
        RECT 10.950000 40.460000 11.270000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950000 40.890000 11.270000 41.210000 ;
      LAYER met4 ;
        RECT 10.950000 40.890000 11.270000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950000 41.320000 11.270000 41.640000 ;
      LAYER met4 ;
        RECT 10.950000 41.320000 11.270000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950000 41.750000 11.270000 42.070000 ;
      LAYER met4 ;
        RECT 10.950000 41.750000 11.270000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950000 42.180000 11.270000 42.500000 ;
      LAYER met4 ;
        RECT 10.950000 42.180000 11.270000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950000 42.610000 11.270000 42.930000 ;
      LAYER met4 ;
        RECT 10.950000 42.610000 11.270000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950000 43.040000 11.270000 43.360000 ;
      LAYER met4 ;
        RECT 10.950000 43.040000 11.270000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950000 43.470000 11.270000 43.790000 ;
      LAYER met4 ;
        RECT 10.950000 43.470000 11.270000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950000 43.900000 11.270000 44.220000 ;
      LAYER met4 ;
        RECT 10.950000 43.900000 11.270000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.350000 39.600000 11.670000 39.920000 ;
      LAYER met4 ;
        RECT 11.350000 39.600000 11.670000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.350000 40.030000 11.670000 40.350000 ;
      LAYER met4 ;
        RECT 11.350000 40.030000 11.670000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.350000 40.460000 11.670000 40.780000 ;
      LAYER met4 ;
        RECT 11.350000 40.460000 11.670000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.350000 40.890000 11.670000 41.210000 ;
      LAYER met4 ;
        RECT 11.350000 40.890000 11.670000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.350000 41.320000 11.670000 41.640000 ;
      LAYER met4 ;
        RECT 11.350000 41.320000 11.670000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.350000 41.750000 11.670000 42.070000 ;
      LAYER met4 ;
        RECT 11.350000 41.750000 11.670000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.350000 42.180000 11.670000 42.500000 ;
      LAYER met4 ;
        RECT 11.350000 42.180000 11.670000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.350000 42.610000 11.670000 42.930000 ;
      LAYER met4 ;
        RECT 11.350000 42.610000 11.670000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.350000 43.040000 11.670000 43.360000 ;
      LAYER met4 ;
        RECT 11.350000 43.040000 11.670000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.350000 43.470000 11.670000 43.790000 ;
      LAYER met4 ;
        RECT 11.350000 43.470000 11.670000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.350000 43.900000 11.670000 44.220000 ;
      LAYER met4 ;
        RECT 11.350000 43.900000 11.670000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.750000 39.600000 12.070000 39.920000 ;
      LAYER met4 ;
        RECT 11.750000 39.600000 12.070000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.750000 40.030000 12.070000 40.350000 ;
      LAYER met4 ;
        RECT 11.750000 40.030000 12.070000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.750000 40.460000 12.070000 40.780000 ;
      LAYER met4 ;
        RECT 11.750000 40.460000 12.070000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.750000 40.890000 12.070000 41.210000 ;
      LAYER met4 ;
        RECT 11.750000 40.890000 12.070000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.750000 41.320000 12.070000 41.640000 ;
      LAYER met4 ;
        RECT 11.750000 41.320000 12.070000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.750000 41.750000 12.070000 42.070000 ;
      LAYER met4 ;
        RECT 11.750000 41.750000 12.070000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.750000 42.180000 12.070000 42.500000 ;
      LAYER met4 ;
        RECT 11.750000 42.180000 12.070000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.750000 42.610000 12.070000 42.930000 ;
      LAYER met4 ;
        RECT 11.750000 42.610000 12.070000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.750000 43.040000 12.070000 43.360000 ;
      LAYER met4 ;
        RECT 11.750000 43.040000 12.070000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.750000 43.470000 12.070000 43.790000 ;
      LAYER met4 ;
        RECT 11.750000 43.470000 12.070000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.750000 43.900000 12.070000 44.220000 ;
      LAYER met4 ;
        RECT 11.750000 43.900000 12.070000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.150000 39.600000 12.470000 39.920000 ;
      LAYER met4 ;
        RECT 12.150000 39.600000 12.470000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.150000 40.030000 12.470000 40.350000 ;
      LAYER met4 ;
        RECT 12.150000 40.030000 12.470000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.150000 40.460000 12.470000 40.780000 ;
      LAYER met4 ;
        RECT 12.150000 40.460000 12.470000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.150000 40.890000 12.470000 41.210000 ;
      LAYER met4 ;
        RECT 12.150000 40.890000 12.470000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.150000 41.320000 12.470000 41.640000 ;
      LAYER met4 ;
        RECT 12.150000 41.320000 12.470000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.150000 41.750000 12.470000 42.070000 ;
      LAYER met4 ;
        RECT 12.150000 41.750000 12.470000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.150000 42.180000 12.470000 42.500000 ;
      LAYER met4 ;
        RECT 12.150000 42.180000 12.470000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.150000 42.610000 12.470000 42.930000 ;
      LAYER met4 ;
        RECT 12.150000 42.610000 12.470000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.150000 43.040000 12.470000 43.360000 ;
      LAYER met4 ;
        RECT 12.150000 43.040000 12.470000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.150000 43.470000 12.470000 43.790000 ;
      LAYER met4 ;
        RECT 12.150000 43.470000 12.470000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.150000 43.900000 12.470000 44.220000 ;
      LAYER met4 ;
        RECT 12.150000 43.900000 12.470000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.550000 39.600000 12.870000 39.920000 ;
      LAYER met4 ;
        RECT 12.550000 39.600000 12.870000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.550000 40.030000 12.870000 40.350000 ;
      LAYER met4 ;
        RECT 12.550000 40.030000 12.870000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.550000 40.460000 12.870000 40.780000 ;
      LAYER met4 ;
        RECT 12.550000 40.460000 12.870000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.550000 40.890000 12.870000 41.210000 ;
      LAYER met4 ;
        RECT 12.550000 40.890000 12.870000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.550000 41.320000 12.870000 41.640000 ;
      LAYER met4 ;
        RECT 12.550000 41.320000 12.870000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.550000 41.750000 12.870000 42.070000 ;
      LAYER met4 ;
        RECT 12.550000 41.750000 12.870000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.550000 42.180000 12.870000 42.500000 ;
      LAYER met4 ;
        RECT 12.550000 42.180000 12.870000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.550000 42.610000 12.870000 42.930000 ;
      LAYER met4 ;
        RECT 12.550000 42.610000 12.870000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.550000 43.040000 12.870000 43.360000 ;
      LAYER met4 ;
        RECT 12.550000 43.040000 12.870000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.550000 43.470000 12.870000 43.790000 ;
      LAYER met4 ;
        RECT 12.550000 43.470000 12.870000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.550000 43.900000 12.870000 44.220000 ;
      LAYER met4 ;
        RECT 12.550000 43.900000 12.870000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.950000 39.600000 13.270000 39.920000 ;
      LAYER met4 ;
        RECT 12.950000 39.600000 13.270000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.950000 40.030000 13.270000 40.350000 ;
      LAYER met4 ;
        RECT 12.950000 40.030000 13.270000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.950000 40.460000 13.270000 40.780000 ;
      LAYER met4 ;
        RECT 12.950000 40.460000 13.270000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.950000 40.890000 13.270000 41.210000 ;
      LAYER met4 ;
        RECT 12.950000 40.890000 13.270000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.950000 41.320000 13.270000 41.640000 ;
      LAYER met4 ;
        RECT 12.950000 41.320000 13.270000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.950000 41.750000 13.270000 42.070000 ;
      LAYER met4 ;
        RECT 12.950000 41.750000 13.270000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.950000 42.180000 13.270000 42.500000 ;
      LAYER met4 ;
        RECT 12.950000 42.180000 13.270000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.950000 42.610000 13.270000 42.930000 ;
      LAYER met4 ;
        RECT 12.950000 42.610000 13.270000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.950000 43.040000 13.270000 43.360000 ;
      LAYER met4 ;
        RECT 12.950000 43.040000 13.270000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.950000 43.470000 13.270000 43.790000 ;
      LAYER met4 ;
        RECT 12.950000 43.470000 13.270000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.950000 43.900000 13.270000 44.220000 ;
      LAYER met4 ;
        RECT 12.950000 43.900000 13.270000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.350000 39.600000 13.670000 39.920000 ;
      LAYER met4 ;
        RECT 13.350000 39.600000 13.670000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.350000 40.030000 13.670000 40.350000 ;
      LAYER met4 ;
        RECT 13.350000 40.030000 13.670000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.350000 40.460000 13.670000 40.780000 ;
      LAYER met4 ;
        RECT 13.350000 40.460000 13.670000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.350000 40.890000 13.670000 41.210000 ;
      LAYER met4 ;
        RECT 13.350000 40.890000 13.670000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.350000 41.320000 13.670000 41.640000 ;
      LAYER met4 ;
        RECT 13.350000 41.320000 13.670000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.350000 41.750000 13.670000 42.070000 ;
      LAYER met4 ;
        RECT 13.350000 41.750000 13.670000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.350000 42.180000 13.670000 42.500000 ;
      LAYER met4 ;
        RECT 13.350000 42.180000 13.670000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.350000 42.610000 13.670000 42.930000 ;
      LAYER met4 ;
        RECT 13.350000 42.610000 13.670000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.350000 43.040000 13.670000 43.360000 ;
      LAYER met4 ;
        RECT 13.350000 43.040000 13.670000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.350000 43.470000 13.670000 43.790000 ;
      LAYER met4 ;
        RECT 13.350000 43.470000 13.670000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.350000 43.900000 13.670000 44.220000 ;
      LAYER met4 ;
        RECT 13.350000 43.900000 13.670000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.750000 39.600000 14.070000 39.920000 ;
      LAYER met4 ;
        RECT 13.750000 39.600000 14.070000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.750000 40.030000 14.070000 40.350000 ;
      LAYER met4 ;
        RECT 13.750000 40.030000 14.070000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.750000 40.460000 14.070000 40.780000 ;
      LAYER met4 ;
        RECT 13.750000 40.460000 14.070000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.750000 40.890000 14.070000 41.210000 ;
      LAYER met4 ;
        RECT 13.750000 40.890000 14.070000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.750000 41.320000 14.070000 41.640000 ;
      LAYER met4 ;
        RECT 13.750000 41.320000 14.070000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.750000 41.750000 14.070000 42.070000 ;
      LAYER met4 ;
        RECT 13.750000 41.750000 14.070000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.750000 42.180000 14.070000 42.500000 ;
      LAYER met4 ;
        RECT 13.750000 42.180000 14.070000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.750000 42.610000 14.070000 42.930000 ;
      LAYER met4 ;
        RECT 13.750000 42.610000 14.070000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.750000 43.040000 14.070000 43.360000 ;
      LAYER met4 ;
        RECT 13.750000 43.040000 14.070000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.750000 43.470000 14.070000 43.790000 ;
      LAYER met4 ;
        RECT 13.750000 43.470000 14.070000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.750000 43.900000 14.070000 44.220000 ;
      LAYER met4 ;
        RECT 13.750000 43.900000 14.070000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.150000 39.600000 14.470000 39.920000 ;
      LAYER met4 ;
        RECT 14.150000 39.600000 14.470000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.150000 40.030000 14.470000 40.350000 ;
      LAYER met4 ;
        RECT 14.150000 40.030000 14.470000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.150000 40.460000 14.470000 40.780000 ;
      LAYER met4 ;
        RECT 14.150000 40.460000 14.470000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.150000 40.890000 14.470000 41.210000 ;
      LAYER met4 ;
        RECT 14.150000 40.890000 14.470000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.150000 41.320000 14.470000 41.640000 ;
      LAYER met4 ;
        RECT 14.150000 41.320000 14.470000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.150000 41.750000 14.470000 42.070000 ;
      LAYER met4 ;
        RECT 14.150000 41.750000 14.470000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.150000 42.180000 14.470000 42.500000 ;
      LAYER met4 ;
        RECT 14.150000 42.180000 14.470000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.150000 42.610000 14.470000 42.930000 ;
      LAYER met4 ;
        RECT 14.150000 42.610000 14.470000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.150000 43.040000 14.470000 43.360000 ;
      LAYER met4 ;
        RECT 14.150000 43.040000 14.470000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.150000 43.470000 14.470000 43.790000 ;
      LAYER met4 ;
        RECT 14.150000 43.470000 14.470000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.150000 43.900000 14.470000 44.220000 ;
      LAYER met4 ;
        RECT 14.150000 43.900000 14.470000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.550000 39.600000 14.870000 39.920000 ;
      LAYER met4 ;
        RECT 14.550000 39.600000 14.870000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.550000 40.030000 14.870000 40.350000 ;
      LAYER met4 ;
        RECT 14.550000 40.030000 14.870000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.550000 40.460000 14.870000 40.780000 ;
      LAYER met4 ;
        RECT 14.550000 40.460000 14.870000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.550000 40.890000 14.870000 41.210000 ;
      LAYER met4 ;
        RECT 14.550000 40.890000 14.870000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.550000 41.320000 14.870000 41.640000 ;
      LAYER met4 ;
        RECT 14.550000 41.320000 14.870000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.550000 41.750000 14.870000 42.070000 ;
      LAYER met4 ;
        RECT 14.550000 41.750000 14.870000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.550000 42.180000 14.870000 42.500000 ;
      LAYER met4 ;
        RECT 14.550000 42.180000 14.870000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.550000 42.610000 14.870000 42.930000 ;
      LAYER met4 ;
        RECT 14.550000 42.610000 14.870000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.550000 43.040000 14.870000 43.360000 ;
      LAYER met4 ;
        RECT 14.550000 43.040000 14.870000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.550000 43.470000 14.870000 43.790000 ;
      LAYER met4 ;
        RECT 14.550000 43.470000 14.870000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.550000 43.900000 14.870000 44.220000 ;
      LAYER met4 ;
        RECT 14.550000 43.900000 14.870000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.950000 39.600000 15.270000 39.920000 ;
      LAYER met4 ;
        RECT 14.950000 39.600000 15.270000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.950000 40.030000 15.270000 40.350000 ;
      LAYER met4 ;
        RECT 14.950000 40.030000 15.270000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.950000 40.460000 15.270000 40.780000 ;
      LAYER met4 ;
        RECT 14.950000 40.460000 15.270000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.950000 40.890000 15.270000 41.210000 ;
      LAYER met4 ;
        RECT 14.950000 40.890000 15.270000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.950000 41.320000 15.270000 41.640000 ;
      LAYER met4 ;
        RECT 14.950000 41.320000 15.270000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.950000 41.750000 15.270000 42.070000 ;
      LAYER met4 ;
        RECT 14.950000 41.750000 15.270000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.950000 42.180000 15.270000 42.500000 ;
      LAYER met4 ;
        RECT 14.950000 42.180000 15.270000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.950000 42.610000 15.270000 42.930000 ;
      LAYER met4 ;
        RECT 14.950000 42.610000 15.270000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.950000 43.040000 15.270000 43.360000 ;
      LAYER met4 ;
        RECT 14.950000 43.040000 15.270000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.950000 43.470000 15.270000 43.790000 ;
      LAYER met4 ;
        RECT 14.950000 43.470000 15.270000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.950000 43.900000 15.270000 44.220000 ;
      LAYER met4 ;
        RECT 14.950000 43.900000 15.270000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.350000 39.600000 15.670000 39.920000 ;
      LAYER met4 ;
        RECT 15.350000 39.600000 15.670000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.350000 40.030000 15.670000 40.350000 ;
      LAYER met4 ;
        RECT 15.350000 40.030000 15.670000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.350000 40.460000 15.670000 40.780000 ;
      LAYER met4 ;
        RECT 15.350000 40.460000 15.670000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.350000 40.890000 15.670000 41.210000 ;
      LAYER met4 ;
        RECT 15.350000 40.890000 15.670000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.350000 41.320000 15.670000 41.640000 ;
      LAYER met4 ;
        RECT 15.350000 41.320000 15.670000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.350000 41.750000 15.670000 42.070000 ;
      LAYER met4 ;
        RECT 15.350000 41.750000 15.670000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.350000 42.180000 15.670000 42.500000 ;
      LAYER met4 ;
        RECT 15.350000 42.180000 15.670000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.350000 42.610000 15.670000 42.930000 ;
      LAYER met4 ;
        RECT 15.350000 42.610000 15.670000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.350000 43.040000 15.670000 43.360000 ;
      LAYER met4 ;
        RECT 15.350000 43.040000 15.670000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.350000 43.470000 15.670000 43.790000 ;
      LAYER met4 ;
        RECT 15.350000 43.470000 15.670000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.350000 43.900000 15.670000 44.220000 ;
      LAYER met4 ;
        RECT 15.350000 43.900000 15.670000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.750000 39.600000 16.070000 39.920000 ;
      LAYER met4 ;
        RECT 15.750000 39.600000 16.070000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.750000 40.030000 16.070000 40.350000 ;
      LAYER met4 ;
        RECT 15.750000 40.030000 16.070000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.750000 40.460000 16.070000 40.780000 ;
      LAYER met4 ;
        RECT 15.750000 40.460000 16.070000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.750000 40.890000 16.070000 41.210000 ;
      LAYER met4 ;
        RECT 15.750000 40.890000 16.070000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.750000 41.320000 16.070000 41.640000 ;
      LAYER met4 ;
        RECT 15.750000 41.320000 16.070000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.750000 41.750000 16.070000 42.070000 ;
      LAYER met4 ;
        RECT 15.750000 41.750000 16.070000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.750000 42.180000 16.070000 42.500000 ;
      LAYER met4 ;
        RECT 15.750000 42.180000 16.070000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.750000 42.610000 16.070000 42.930000 ;
      LAYER met4 ;
        RECT 15.750000 42.610000 16.070000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.750000 43.040000 16.070000 43.360000 ;
      LAYER met4 ;
        RECT 15.750000 43.040000 16.070000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.750000 43.470000 16.070000 43.790000 ;
      LAYER met4 ;
        RECT 15.750000 43.470000 16.070000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.750000 43.900000 16.070000 44.220000 ;
      LAYER met4 ;
        RECT 15.750000 43.900000 16.070000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.150000 39.600000 16.470000 39.920000 ;
      LAYER met4 ;
        RECT 16.150000 39.600000 16.470000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.150000 40.030000 16.470000 40.350000 ;
      LAYER met4 ;
        RECT 16.150000 40.030000 16.470000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.150000 40.460000 16.470000 40.780000 ;
      LAYER met4 ;
        RECT 16.150000 40.460000 16.470000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.150000 40.890000 16.470000 41.210000 ;
      LAYER met4 ;
        RECT 16.150000 40.890000 16.470000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.150000 41.320000 16.470000 41.640000 ;
      LAYER met4 ;
        RECT 16.150000 41.320000 16.470000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.150000 41.750000 16.470000 42.070000 ;
      LAYER met4 ;
        RECT 16.150000 41.750000 16.470000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.150000 42.180000 16.470000 42.500000 ;
      LAYER met4 ;
        RECT 16.150000 42.180000 16.470000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.150000 42.610000 16.470000 42.930000 ;
      LAYER met4 ;
        RECT 16.150000 42.610000 16.470000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.150000 43.040000 16.470000 43.360000 ;
      LAYER met4 ;
        RECT 16.150000 43.040000 16.470000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.150000 43.470000 16.470000 43.790000 ;
      LAYER met4 ;
        RECT 16.150000 43.470000 16.470000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.150000 43.900000 16.470000 44.220000 ;
      LAYER met4 ;
        RECT 16.150000 43.900000 16.470000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.550000 39.600000 16.870000 39.920000 ;
      LAYER met4 ;
        RECT 16.550000 39.600000 16.870000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.550000 40.030000 16.870000 40.350000 ;
      LAYER met4 ;
        RECT 16.550000 40.030000 16.870000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.550000 40.460000 16.870000 40.780000 ;
      LAYER met4 ;
        RECT 16.550000 40.460000 16.870000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.550000 40.890000 16.870000 41.210000 ;
      LAYER met4 ;
        RECT 16.550000 40.890000 16.870000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.550000 41.320000 16.870000 41.640000 ;
      LAYER met4 ;
        RECT 16.550000 41.320000 16.870000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.550000 41.750000 16.870000 42.070000 ;
      LAYER met4 ;
        RECT 16.550000 41.750000 16.870000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.550000 42.180000 16.870000 42.500000 ;
      LAYER met4 ;
        RECT 16.550000 42.180000 16.870000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.550000 42.610000 16.870000 42.930000 ;
      LAYER met4 ;
        RECT 16.550000 42.610000 16.870000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.550000 43.040000 16.870000 43.360000 ;
      LAYER met4 ;
        RECT 16.550000 43.040000 16.870000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.550000 43.470000 16.870000 43.790000 ;
      LAYER met4 ;
        RECT 16.550000 43.470000 16.870000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.550000 43.900000 16.870000 44.220000 ;
      LAYER met4 ;
        RECT 16.550000 43.900000 16.870000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.950000 39.600000 17.270000 39.920000 ;
      LAYER met4 ;
        RECT 16.950000 39.600000 17.270000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.950000 40.030000 17.270000 40.350000 ;
      LAYER met4 ;
        RECT 16.950000 40.030000 17.270000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.950000 40.460000 17.270000 40.780000 ;
      LAYER met4 ;
        RECT 16.950000 40.460000 17.270000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.950000 40.890000 17.270000 41.210000 ;
      LAYER met4 ;
        RECT 16.950000 40.890000 17.270000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.950000 41.320000 17.270000 41.640000 ;
      LAYER met4 ;
        RECT 16.950000 41.320000 17.270000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.950000 41.750000 17.270000 42.070000 ;
      LAYER met4 ;
        RECT 16.950000 41.750000 17.270000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.950000 42.180000 17.270000 42.500000 ;
      LAYER met4 ;
        RECT 16.950000 42.180000 17.270000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.950000 42.610000 17.270000 42.930000 ;
      LAYER met4 ;
        RECT 16.950000 42.610000 17.270000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.950000 43.040000 17.270000 43.360000 ;
      LAYER met4 ;
        RECT 16.950000 43.040000 17.270000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.950000 43.470000 17.270000 43.790000 ;
      LAYER met4 ;
        RECT 16.950000 43.470000 17.270000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.950000 43.900000 17.270000 44.220000 ;
      LAYER met4 ;
        RECT 16.950000 43.900000 17.270000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.350000 39.600000 17.670000 39.920000 ;
      LAYER met4 ;
        RECT 17.350000 39.600000 17.670000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.350000 40.030000 17.670000 40.350000 ;
      LAYER met4 ;
        RECT 17.350000 40.030000 17.670000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.350000 40.460000 17.670000 40.780000 ;
      LAYER met4 ;
        RECT 17.350000 40.460000 17.670000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.350000 40.890000 17.670000 41.210000 ;
      LAYER met4 ;
        RECT 17.350000 40.890000 17.670000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.350000 41.320000 17.670000 41.640000 ;
      LAYER met4 ;
        RECT 17.350000 41.320000 17.670000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.350000 41.750000 17.670000 42.070000 ;
      LAYER met4 ;
        RECT 17.350000 41.750000 17.670000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.350000 42.180000 17.670000 42.500000 ;
      LAYER met4 ;
        RECT 17.350000 42.180000 17.670000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.350000 42.610000 17.670000 42.930000 ;
      LAYER met4 ;
        RECT 17.350000 42.610000 17.670000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.350000 43.040000 17.670000 43.360000 ;
      LAYER met4 ;
        RECT 17.350000 43.040000 17.670000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.350000 43.470000 17.670000 43.790000 ;
      LAYER met4 ;
        RECT 17.350000 43.470000 17.670000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.350000 43.900000 17.670000 44.220000 ;
      LAYER met4 ;
        RECT 17.350000 43.900000 17.670000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.750000 39.600000 18.070000 39.920000 ;
      LAYER met4 ;
        RECT 17.750000 39.600000 18.070000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.750000 40.030000 18.070000 40.350000 ;
      LAYER met4 ;
        RECT 17.750000 40.030000 18.070000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.750000 40.460000 18.070000 40.780000 ;
      LAYER met4 ;
        RECT 17.750000 40.460000 18.070000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.750000 40.890000 18.070000 41.210000 ;
      LAYER met4 ;
        RECT 17.750000 40.890000 18.070000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.750000 41.320000 18.070000 41.640000 ;
      LAYER met4 ;
        RECT 17.750000 41.320000 18.070000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.750000 41.750000 18.070000 42.070000 ;
      LAYER met4 ;
        RECT 17.750000 41.750000 18.070000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.750000 42.180000 18.070000 42.500000 ;
      LAYER met4 ;
        RECT 17.750000 42.180000 18.070000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.750000 42.610000 18.070000 42.930000 ;
      LAYER met4 ;
        RECT 17.750000 42.610000 18.070000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.750000 43.040000 18.070000 43.360000 ;
      LAYER met4 ;
        RECT 17.750000 43.040000 18.070000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.750000 43.470000 18.070000 43.790000 ;
      LAYER met4 ;
        RECT 17.750000 43.470000 18.070000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.750000 43.900000 18.070000 44.220000 ;
      LAYER met4 ;
        RECT 17.750000 43.900000 18.070000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.150000 39.600000 18.470000 39.920000 ;
      LAYER met4 ;
        RECT 18.150000 39.600000 18.470000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.150000 40.030000 18.470000 40.350000 ;
      LAYER met4 ;
        RECT 18.150000 40.030000 18.470000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.150000 40.460000 18.470000 40.780000 ;
      LAYER met4 ;
        RECT 18.150000 40.460000 18.470000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.150000 40.890000 18.470000 41.210000 ;
      LAYER met4 ;
        RECT 18.150000 40.890000 18.470000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.150000 41.320000 18.470000 41.640000 ;
      LAYER met4 ;
        RECT 18.150000 41.320000 18.470000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.150000 41.750000 18.470000 42.070000 ;
      LAYER met4 ;
        RECT 18.150000 41.750000 18.470000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.150000 42.180000 18.470000 42.500000 ;
      LAYER met4 ;
        RECT 18.150000 42.180000 18.470000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.150000 42.610000 18.470000 42.930000 ;
      LAYER met4 ;
        RECT 18.150000 42.610000 18.470000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.150000 43.040000 18.470000 43.360000 ;
      LAYER met4 ;
        RECT 18.150000 43.040000 18.470000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.150000 43.470000 18.470000 43.790000 ;
      LAYER met4 ;
        RECT 18.150000 43.470000 18.470000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.150000 43.900000 18.470000 44.220000 ;
      LAYER met4 ;
        RECT 18.150000 43.900000 18.470000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.550000 39.600000 18.870000 39.920000 ;
      LAYER met4 ;
        RECT 18.550000 39.600000 18.870000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.550000 40.030000 18.870000 40.350000 ;
      LAYER met4 ;
        RECT 18.550000 40.030000 18.870000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.550000 40.460000 18.870000 40.780000 ;
      LAYER met4 ;
        RECT 18.550000 40.460000 18.870000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.550000 40.890000 18.870000 41.210000 ;
      LAYER met4 ;
        RECT 18.550000 40.890000 18.870000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.550000 41.320000 18.870000 41.640000 ;
      LAYER met4 ;
        RECT 18.550000 41.320000 18.870000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.550000 41.750000 18.870000 42.070000 ;
      LAYER met4 ;
        RECT 18.550000 41.750000 18.870000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.550000 42.180000 18.870000 42.500000 ;
      LAYER met4 ;
        RECT 18.550000 42.180000 18.870000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.550000 42.610000 18.870000 42.930000 ;
      LAYER met4 ;
        RECT 18.550000 42.610000 18.870000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.550000 43.040000 18.870000 43.360000 ;
      LAYER met4 ;
        RECT 18.550000 43.040000 18.870000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.550000 43.470000 18.870000 43.790000 ;
      LAYER met4 ;
        RECT 18.550000 43.470000 18.870000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.550000 43.900000 18.870000 44.220000 ;
      LAYER met4 ;
        RECT 18.550000 43.900000 18.870000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.950000 39.600000 19.270000 39.920000 ;
      LAYER met4 ;
        RECT 18.950000 39.600000 19.270000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.950000 40.030000 19.270000 40.350000 ;
      LAYER met4 ;
        RECT 18.950000 40.030000 19.270000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.950000 40.460000 19.270000 40.780000 ;
      LAYER met4 ;
        RECT 18.950000 40.460000 19.270000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.950000 40.890000 19.270000 41.210000 ;
      LAYER met4 ;
        RECT 18.950000 40.890000 19.270000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.950000 41.320000 19.270000 41.640000 ;
      LAYER met4 ;
        RECT 18.950000 41.320000 19.270000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.950000 41.750000 19.270000 42.070000 ;
      LAYER met4 ;
        RECT 18.950000 41.750000 19.270000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.950000 42.180000 19.270000 42.500000 ;
      LAYER met4 ;
        RECT 18.950000 42.180000 19.270000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.950000 42.610000 19.270000 42.930000 ;
      LAYER met4 ;
        RECT 18.950000 42.610000 19.270000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.950000 43.040000 19.270000 43.360000 ;
      LAYER met4 ;
        RECT 18.950000 43.040000 19.270000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.950000 43.470000 19.270000 43.790000 ;
      LAYER met4 ;
        RECT 18.950000 43.470000 19.270000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.950000 43.900000 19.270000 44.220000 ;
      LAYER met4 ;
        RECT 18.950000 43.900000 19.270000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.350000 39.600000 19.670000 39.920000 ;
      LAYER met4 ;
        RECT 19.350000 39.600000 19.670000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.350000 40.030000 19.670000 40.350000 ;
      LAYER met4 ;
        RECT 19.350000 40.030000 19.670000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.350000 40.460000 19.670000 40.780000 ;
      LAYER met4 ;
        RECT 19.350000 40.460000 19.670000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.350000 40.890000 19.670000 41.210000 ;
      LAYER met4 ;
        RECT 19.350000 40.890000 19.670000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.350000 41.320000 19.670000 41.640000 ;
      LAYER met4 ;
        RECT 19.350000 41.320000 19.670000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.350000 41.750000 19.670000 42.070000 ;
      LAYER met4 ;
        RECT 19.350000 41.750000 19.670000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.350000 42.180000 19.670000 42.500000 ;
      LAYER met4 ;
        RECT 19.350000 42.180000 19.670000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.350000 42.610000 19.670000 42.930000 ;
      LAYER met4 ;
        RECT 19.350000 42.610000 19.670000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.350000 43.040000 19.670000 43.360000 ;
      LAYER met4 ;
        RECT 19.350000 43.040000 19.670000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.350000 43.470000 19.670000 43.790000 ;
      LAYER met4 ;
        RECT 19.350000 43.470000 19.670000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.350000 43.900000 19.670000 44.220000 ;
      LAYER met4 ;
        RECT 19.350000 43.900000 19.670000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.750000 39.600000 20.070000 39.920000 ;
      LAYER met4 ;
        RECT 19.750000 39.600000 20.070000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.750000 40.030000 20.070000 40.350000 ;
      LAYER met4 ;
        RECT 19.750000 40.030000 20.070000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.750000 40.460000 20.070000 40.780000 ;
      LAYER met4 ;
        RECT 19.750000 40.460000 20.070000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.750000 40.890000 20.070000 41.210000 ;
      LAYER met4 ;
        RECT 19.750000 40.890000 20.070000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.750000 41.320000 20.070000 41.640000 ;
      LAYER met4 ;
        RECT 19.750000 41.320000 20.070000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.750000 41.750000 20.070000 42.070000 ;
      LAYER met4 ;
        RECT 19.750000 41.750000 20.070000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.750000 42.180000 20.070000 42.500000 ;
      LAYER met4 ;
        RECT 19.750000 42.180000 20.070000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.750000 42.610000 20.070000 42.930000 ;
      LAYER met4 ;
        RECT 19.750000 42.610000 20.070000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.750000 43.040000 20.070000 43.360000 ;
      LAYER met4 ;
        RECT 19.750000 43.040000 20.070000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.750000 43.470000 20.070000 43.790000 ;
      LAYER met4 ;
        RECT 19.750000 43.470000 20.070000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.750000 43.900000 20.070000 44.220000 ;
      LAYER met4 ;
        RECT 19.750000 43.900000 20.070000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.150000 39.600000 2.470000 39.920000 ;
      LAYER met4 ;
        RECT 2.150000 39.600000 2.470000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.150000 40.030000 2.470000 40.350000 ;
      LAYER met4 ;
        RECT 2.150000 40.030000 2.470000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.150000 40.460000 2.470000 40.780000 ;
      LAYER met4 ;
        RECT 2.150000 40.460000 2.470000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.150000 40.890000 2.470000 41.210000 ;
      LAYER met4 ;
        RECT 2.150000 40.890000 2.470000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.150000 41.320000 2.470000 41.640000 ;
      LAYER met4 ;
        RECT 2.150000 41.320000 2.470000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.150000 41.750000 2.470000 42.070000 ;
      LAYER met4 ;
        RECT 2.150000 41.750000 2.470000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.150000 42.180000 2.470000 42.500000 ;
      LAYER met4 ;
        RECT 2.150000 42.180000 2.470000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.150000 42.610000 2.470000 42.930000 ;
      LAYER met4 ;
        RECT 2.150000 42.610000 2.470000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.150000 43.040000 2.470000 43.360000 ;
      LAYER met4 ;
        RECT 2.150000 43.040000 2.470000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.150000 43.470000 2.470000 43.790000 ;
      LAYER met4 ;
        RECT 2.150000 43.470000 2.470000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.150000 43.900000 2.470000 44.220000 ;
      LAYER met4 ;
        RECT 2.150000 43.900000 2.470000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.550000 39.600000 2.870000 39.920000 ;
      LAYER met4 ;
        RECT 2.550000 39.600000 2.870000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.550000 40.030000 2.870000 40.350000 ;
      LAYER met4 ;
        RECT 2.550000 40.030000 2.870000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.550000 40.460000 2.870000 40.780000 ;
      LAYER met4 ;
        RECT 2.550000 40.460000 2.870000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.550000 40.890000 2.870000 41.210000 ;
      LAYER met4 ;
        RECT 2.550000 40.890000 2.870000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.550000 41.320000 2.870000 41.640000 ;
      LAYER met4 ;
        RECT 2.550000 41.320000 2.870000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.550000 41.750000 2.870000 42.070000 ;
      LAYER met4 ;
        RECT 2.550000 41.750000 2.870000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.550000 42.180000 2.870000 42.500000 ;
      LAYER met4 ;
        RECT 2.550000 42.180000 2.870000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.550000 42.610000 2.870000 42.930000 ;
      LAYER met4 ;
        RECT 2.550000 42.610000 2.870000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.550000 43.040000 2.870000 43.360000 ;
      LAYER met4 ;
        RECT 2.550000 43.040000 2.870000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.550000 43.470000 2.870000 43.790000 ;
      LAYER met4 ;
        RECT 2.550000 43.470000 2.870000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.550000 43.900000 2.870000 44.220000 ;
      LAYER met4 ;
        RECT 2.550000 43.900000 2.870000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.950000 39.600000 3.270000 39.920000 ;
      LAYER met4 ;
        RECT 2.950000 39.600000 3.270000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.950000 40.030000 3.270000 40.350000 ;
      LAYER met4 ;
        RECT 2.950000 40.030000 3.270000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.950000 40.460000 3.270000 40.780000 ;
      LAYER met4 ;
        RECT 2.950000 40.460000 3.270000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.950000 40.890000 3.270000 41.210000 ;
      LAYER met4 ;
        RECT 2.950000 40.890000 3.270000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.950000 41.320000 3.270000 41.640000 ;
      LAYER met4 ;
        RECT 2.950000 41.320000 3.270000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.950000 41.750000 3.270000 42.070000 ;
      LAYER met4 ;
        RECT 2.950000 41.750000 3.270000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.950000 42.180000 3.270000 42.500000 ;
      LAYER met4 ;
        RECT 2.950000 42.180000 3.270000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.950000 42.610000 3.270000 42.930000 ;
      LAYER met4 ;
        RECT 2.950000 42.610000 3.270000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.950000 43.040000 3.270000 43.360000 ;
      LAYER met4 ;
        RECT 2.950000 43.040000 3.270000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.950000 43.470000 3.270000 43.790000 ;
      LAYER met4 ;
        RECT 2.950000 43.470000 3.270000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.950000 43.900000 3.270000 44.220000 ;
      LAYER met4 ;
        RECT 2.950000 43.900000 3.270000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150000 39.600000 20.470000 39.920000 ;
      LAYER met4 ;
        RECT 20.150000 39.600000 20.470000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150000 40.030000 20.470000 40.350000 ;
      LAYER met4 ;
        RECT 20.150000 40.030000 20.470000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150000 40.460000 20.470000 40.780000 ;
      LAYER met4 ;
        RECT 20.150000 40.460000 20.470000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150000 40.890000 20.470000 41.210000 ;
      LAYER met4 ;
        RECT 20.150000 40.890000 20.470000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150000 41.320000 20.470000 41.640000 ;
      LAYER met4 ;
        RECT 20.150000 41.320000 20.470000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150000 41.750000 20.470000 42.070000 ;
      LAYER met4 ;
        RECT 20.150000 41.750000 20.470000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150000 42.180000 20.470000 42.500000 ;
      LAYER met4 ;
        RECT 20.150000 42.180000 20.470000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150000 42.610000 20.470000 42.930000 ;
      LAYER met4 ;
        RECT 20.150000 42.610000 20.470000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150000 43.040000 20.470000 43.360000 ;
      LAYER met4 ;
        RECT 20.150000 43.040000 20.470000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150000 43.470000 20.470000 43.790000 ;
      LAYER met4 ;
        RECT 20.150000 43.470000 20.470000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150000 43.900000 20.470000 44.220000 ;
      LAYER met4 ;
        RECT 20.150000 43.900000 20.470000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.550000 39.600000 20.870000 39.920000 ;
      LAYER met4 ;
        RECT 20.550000 39.600000 20.870000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.550000 40.030000 20.870000 40.350000 ;
      LAYER met4 ;
        RECT 20.550000 40.030000 20.870000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.550000 40.460000 20.870000 40.780000 ;
      LAYER met4 ;
        RECT 20.550000 40.460000 20.870000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.550000 40.890000 20.870000 41.210000 ;
      LAYER met4 ;
        RECT 20.550000 40.890000 20.870000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.550000 41.320000 20.870000 41.640000 ;
      LAYER met4 ;
        RECT 20.550000 41.320000 20.870000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.550000 41.750000 20.870000 42.070000 ;
      LAYER met4 ;
        RECT 20.550000 41.750000 20.870000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.550000 42.180000 20.870000 42.500000 ;
      LAYER met4 ;
        RECT 20.550000 42.180000 20.870000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.550000 42.610000 20.870000 42.930000 ;
      LAYER met4 ;
        RECT 20.550000 42.610000 20.870000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.550000 43.040000 20.870000 43.360000 ;
      LAYER met4 ;
        RECT 20.550000 43.040000 20.870000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.550000 43.470000 20.870000 43.790000 ;
      LAYER met4 ;
        RECT 20.550000 43.470000 20.870000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.550000 43.900000 20.870000 44.220000 ;
      LAYER met4 ;
        RECT 20.550000 43.900000 20.870000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.950000 39.600000 21.270000 39.920000 ;
      LAYER met4 ;
        RECT 20.950000 39.600000 21.270000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.950000 40.030000 21.270000 40.350000 ;
      LAYER met4 ;
        RECT 20.950000 40.030000 21.270000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.950000 40.460000 21.270000 40.780000 ;
      LAYER met4 ;
        RECT 20.950000 40.460000 21.270000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.950000 40.890000 21.270000 41.210000 ;
      LAYER met4 ;
        RECT 20.950000 40.890000 21.270000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.950000 41.320000 21.270000 41.640000 ;
      LAYER met4 ;
        RECT 20.950000 41.320000 21.270000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.950000 41.750000 21.270000 42.070000 ;
      LAYER met4 ;
        RECT 20.950000 41.750000 21.270000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.950000 42.180000 21.270000 42.500000 ;
      LAYER met4 ;
        RECT 20.950000 42.180000 21.270000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.950000 42.610000 21.270000 42.930000 ;
      LAYER met4 ;
        RECT 20.950000 42.610000 21.270000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.950000 43.040000 21.270000 43.360000 ;
      LAYER met4 ;
        RECT 20.950000 43.040000 21.270000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.950000 43.470000 21.270000 43.790000 ;
      LAYER met4 ;
        RECT 20.950000 43.470000 21.270000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.950000 43.900000 21.270000 44.220000 ;
      LAYER met4 ;
        RECT 20.950000 43.900000 21.270000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.350000 39.600000 21.670000 39.920000 ;
      LAYER met4 ;
        RECT 21.350000 39.600000 21.670000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.350000 40.030000 21.670000 40.350000 ;
      LAYER met4 ;
        RECT 21.350000 40.030000 21.670000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.350000 40.460000 21.670000 40.780000 ;
      LAYER met4 ;
        RECT 21.350000 40.460000 21.670000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.350000 40.890000 21.670000 41.210000 ;
      LAYER met4 ;
        RECT 21.350000 40.890000 21.670000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.350000 41.320000 21.670000 41.640000 ;
      LAYER met4 ;
        RECT 21.350000 41.320000 21.670000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.350000 41.750000 21.670000 42.070000 ;
      LAYER met4 ;
        RECT 21.350000 41.750000 21.670000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.350000 42.180000 21.670000 42.500000 ;
      LAYER met4 ;
        RECT 21.350000 42.180000 21.670000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.350000 42.610000 21.670000 42.930000 ;
      LAYER met4 ;
        RECT 21.350000 42.610000 21.670000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.350000 43.040000 21.670000 43.360000 ;
      LAYER met4 ;
        RECT 21.350000 43.040000 21.670000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.350000 43.470000 21.670000 43.790000 ;
      LAYER met4 ;
        RECT 21.350000 43.470000 21.670000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.350000 43.900000 21.670000 44.220000 ;
      LAYER met4 ;
        RECT 21.350000 43.900000 21.670000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750000 39.600000 22.070000 39.920000 ;
      LAYER met4 ;
        RECT 21.750000 39.600000 22.070000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750000 40.030000 22.070000 40.350000 ;
      LAYER met4 ;
        RECT 21.750000 40.030000 22.070000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750000 40.460000 22.070000 40.780000 ;
      LAYER met4 ;
        RECT 21.750000 40.460000 22.070000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750000 40.890000 22.070000 41.210000 ;
      LAYER met4 ;
        RECT 21.750000 40.890000 22.070000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750000 41.320000 22.070000 41.640000 ;
      LAYER met4 ;
        RECT 21.750000 41.320000 22.070000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750000 41.750000 22.070000 42.070000 ;
      LAYER met4 ;
        RECT 21.750000 41.750000 22.070000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750000 42.180000 22.070000 42.500000 ;
      LAYER met4 ;
        RECT 21.750000 42.180000 22.070000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750000 42.610000 22.070000 42.930000 ;
      LAYER met4 ;
        RECT 21.750000 42.610000 22.070000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750000 43.040000 22.070000 43.360000 ;
      LAYER met4 ;
        RECT 21.750000 43.040000 22.070000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750000 43.470000 22.070000 43.790000 ;
      LAYER met4 ;
        RECT 21.750000 43.470000 22.070000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750000 43.900000 22.070000 44.220000 ;
      LAYER met4 ;
        RECT 21.750000 43.900000 22.070000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.150000 39.600000 22.470000 39.920000 ;
      LAYER met4 ;
        RECT 22.150000 39.600000 22.470000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.150000 40.030000 22.470000 40.350000 ;
      LAYER met4 ;
        RECT 22.150000 40.030000 22.470000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.150000 40.460000 22.470000 40.780000 ;
      LAYER met4 ;
        RECT 22.150000 40.460000 22.470000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.150000 40.890000 22.470000 41.210000 ;
      LAYER met4 ;
        RECT 22.150000 40.890000 22.470000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.150000 41.320000 22.470000 41.640000 ;
      LAYER met4 ;
        RECT 22.150000 41.320000 22.470000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.150000 41.750000 22.470000 42.070000 ;
      LAYER met4 ;
        RECT 22.150000 41.750000 22.470000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.150000 42.180000 22.470000 42.500000 ;
      LAYER met4 ;
        RECT 22.150000 42.180000 22.470000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.150000 42.610000 22.470000 42.930000 ;
      LAYER met4 ;
        RECT 22.150000 42.610000 22.470000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.150000 43.040000 22.470000 43.360000 ;
      LAYER met4 ;
        RECT 22.150000 43.040000 22.470000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.150000 43.470000 22.470000 43.790000 ;
      LAYER met4 ;
        RECT 22.150000 43.470000 22.470000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.150000 43.900000 22.470000 44.220000 ;
      LAYER met4 ;
        RECT 22.150000 43.900000 22.470000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.550000 39.600000 22.870000 39.920000 ;
      LAYER met4 ;
        RECT 22.550000 39.600000 22.870000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.550000 40.030000 22.870000 40.350000 ;
      LAYER met4 ;
        RECT 22.550000 40.030000 22.870000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.550000 40.460000 22.870000 40.780000 ;
      LAYER met4 ;
        RECT 22.550000 40.460000 22.870000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.550000 40.890000 22.870000 41.210000 ;
      LAYER met4 ;
        RECT 22.550000 40.890000 22.870000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.550000 41.320000 22.870000 41.640000 ;
      LAYER met4 ;
        RECT 22.550000 41.320000 22.870000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.550000 41.750000 22.870000 42.070000 ;
      LAYER met4 ;
        RECT 22.550000 41.750000 22.870000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.550000 42.180000 22.870000 42.500000 ;
      LAYER met4 ;
        RECT 22.550000 42.180000 22.870000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.550000 42.610000 22.870000 42.930000 ;
      LAYER met4 ;
        RECT 22.550000 42.610000 22.870000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.550000 43.040000 22.870000 43.360000 ;
      LAYER met4 ;
        RECT 22.550000 43.040000 22.870000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.550000 43.470000 22.870000 43.790000 ;
      LAYER met4 ;
        RECT 22.550000 43.470000 22.870000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.550000 43.900000 22.870000 44.220000 ;
      LAYER met4 ;
        RECT 22.550000 43.900000 22.870000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950000 39.600000 23.270000 39.920000 ;
      LAYER met4 ;
        RECT 22.950000 39.600000 23.270000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950000 40.030000 23.270000 40.350000 ;
      LAYER met4 ;
        RECT 22.950000 40.030000 23.270000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950000 40.460000 23.270000 40.780000 ;
      LAYER met4 ;
        RECT 22.950000 40.460000 23.270000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950000 40.890000 23.270000 41.210000 ;
      LAYER met4 ;
        RECT 22.950000 40.890000 23.270000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950000 41.320000 23.270000 41.640000 ;
      LAYER met4 ;
        RECT 22.950000 41.320000 23.270000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950000 41.750000 23.270000 42.070000 ;
      LAYER met4 ;
        RECT 22.950000 41.750000 23.270000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950000 42.180000 23.270000 42.500000 ;
      LAYER met4 ;
        RECT 22.950000 42.180000 23.270000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950000 42.610000 23.270000 42.930000 ;
      LAYER met4 ;
        RECT 22.950000 42.610000 23.270000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950000 43.040000 23.270000 43.360000 ;
      LAYER met4 ;
        RECT 22.950000 43.040000 23.270000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950000 43.470000 23.270000 43.790000 ;
      LAYER met4 ;
        RECT 22.950000 43.470000 23.270000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950000 43.900000 23.270000 44.220000 ;
      LAYER met4 ;
        RECT 22.950000 43.900000 23.270000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.350000 39.600000 23.670000 39.920000 ;
      LAYER met4 ;
        RECT 23.350000 39.600000 23.670000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.350000 40.030000 23.670000 40.350000 ;
      LAYER met4 ;
        RECT 23.350000 40.030000 23.670000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.350000 40.460000 23.670000 40.780000 ;
      LAYER met4 ;
        RECT 23.350000 40.460000 23.670000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.350000 40.890000 23.670000 41.210000 ;
      LAYER met4 ;
        RECT 23.350000 40.890000 23.670000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.350000 41.320000 23.670000 41.640000 ;
      LAYER met4 ;
        RECT 23.350000 41.320000 23.670000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.350000 41.750000 23.670000 42.070000 ;
      LAYER met4 ;
        RECT 23.350000 41.750000 23.670000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.350000 42.180000 23.670000 42.500000 ;
      LAYER met4 ;
        RECT 23.350000 42.180000 23.670000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.350000 42.610000 23.670000 42.930000 ;
      LAYER met4 ;
        RECT 23.350000 42.610000 23.670000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.350000 43.040000 23.670000 43.360000 ;
      LAYER met4 ;
        RECT 23.350000 43.040000 23.670000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.350000 43.470000 23.670000 43.790000 ;
      LAYER met4 ;
        RECT 23.350000 43.470000 23.670000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.350000 43.900000 23.670000 44.220000 ;
      LAYER met4 ;
        RECT 23.350000 43.900000 23.670000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.750000 39.600000 24.070000 39.920000 ;
      LAYER met4 ;
        RECT 23.750000 39.600000 24.070000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.750000 40.030000 24.070000 40.350000 ;
      LAYER met4 ;
        RECT 23.750000 40.030000 24.070000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.750000 40.460000 24.070000 40.780000 ;
      LAYER met4 ;
        RECT 23.750000 40.460000 24.070000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.750000 40.890000 24.070000 41.210000 ;
      LAYER met4 ;
        RECT 23.750000 40.890000 24.070000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.750000 41.320000 24.070000 41.640000 ;
      LAYER met4 ;
        RECT 23.750000 41.320000 24.070000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.750000 41.750000 24.070000 42.070000 ;
      LAYER met4 ;
        RECT 23.750000 41.750000 24.070000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.750000 42.180000 24.070000 42.500000 ;
      LAYER met4 ;
        RECT 23.750000 42.180000 24.070000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.750000 42.610000 24.070000 42.930000 ;
      LAYER met4 ;
        RECT 23.750000 42.610000 24.070000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.750000 43.040000 24.070000 43.360000 ;
      LAYER met4 ;
        RECT 23.750000 43.040000 24.070000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.750000 43.470000 24.070000 43.790000 ;
      LAYER met4 ;
        RECT 23.750000 43.470000 24.070000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.750000 43.900000 24.070000 44.220000 ;
      LAYER met4 ;
        RECT 23.750000 43.900000 24.070000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 39.600000 24.470000 39.920000 ;
      LAYER met4 ;
        RECT 24.150000 39.600000 24.470000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 40.030000 24.470000 40.350000 ;
      LAYER met4 ;
        RECT 24.150000 40.030000 24.470000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 40.460000 24.470000 40.780000 ;
      LAYER met4 ;
        RECT 24.150000 40.460000 24.470000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 40.890000 24.470000 41.210000 ;
      LAYER met4 ;
        RECT 24.150000 40.890000 24.470000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 41.320000 24.470000 41.640000 ;
      LAYER met4 ;
        RECT 24.150000 41.320000 24.470000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 41.750000 24.470000 42.070000 ;
      LAYER met4 ;
        RECT 24.150000 41.750000 24.470000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 42.180000 24.470000 42.500000 ;
      LAYER met4 ;
        RECT 24.150000 42.180000 24.470000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 42.610000 24.470000 42.930000 ;
      LAYER met4 ;
        RECT 24.150000 42.610000 24.470000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 43.040000 24.470000 43.360000 ;
      LAYER met4 ;
        RECT 24.150000 43.040000 24.470000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 43.470000 24.470000 43.790000 ;
      LAYER met4 ;
        RECT 24.150000 43.470000 24.470000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 43.900000 24.470000 44.220000 ;
      LAYER met4 ;
        RECT 24.150000 43.900000 24.470000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.350000 39.600000 3.670000 39.920000 ;
      LAYER met4 ;
        RECT 3.350000 39.600000 3.670000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.350000 40.030000 3.670000 40.350000 ;
      LAYER met4 ;
        RECT 3.350000 40.030000 3.670000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.350000 40.460000 3.670000 40.780000 ;
      LAYER met4 ;
        RECT 3.350000 40.460000 3.670000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.350000 40.890000 3.670000 41.210000 ;
      LAYER met4 ;
        RECT 3.350000 40.890000 3.670000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.350000 41.320000 3.670000 41.640000 ;
      LAYER met4 ;
        RECT 3.350000 41.320000 3.670000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.350000 41.750000 3.670000 42.070000 ;
      LAYER met4 ;
        RECT 3.350000 41.750000 3.670000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.350000 42.180000 3.670000 42.500000 ;
      LAYER met4 ;
        RECT 3.350000 42.180000 3.670000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.350000 42.610000 3.670000 42.930000 ;
      LAYER met4 ;
        RECT 3.350000 42.610000 3.670000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.350000 43.040000 3.670000 43.360000 ;
      LAYER met4 ;
        RECT 3.350000 43.040000 3.670000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.350000 43.470000 3.670000 43.790000 ;
      LAYER met4 ;
        RECT 3.350000 43.470000 3.670000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.350000 43.900000 3.670000 44.220000 ;
      LAYER met4 ;
        RECT 3.350000 43.900000 3.670000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.750000 39.600000 4.070000 39.920000 ;
      LAYER met4 ;
        RECT 3.750000 39.600000 4.070000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.750000 40.030000 4.070000 40.350000 ;
      LAYER met4 ;
        RECT 3.750000 40.030000 4.070000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.750000 40.460000 4.070000 40.780000 ;
      LAYER met4 ;
        RECT 3.750000 40.460000 4.070000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.750000 40.890000 4.070000 41.210000 ;
      LAYER met4 ;
        RECT 3.750000 40.890000 4.070000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.750000 41.320000 4.070000 41.640000 ;
      LAYER met4 ;
        RECT 3.750000 41.320000 4.070000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.750000 41.750000 4.070000 42.070000 ;
      LAYER met4 ;
        RECT 3.750000 41.750000 4.070000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.750000 42.180000 4.070000 42.500000 ;
      LAYER met4 ;
        RECT 3.750000 42.180000 4.070000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.750000 42.610000 4.070000 42.930000 ;
      LAYER met4 ;
        RECT 3.750000 42.610000 4.070000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.750000 43.040000 4.070000 43.360000 ;
      LAYER met4 ;
        RECT 3.750000 43.040000 4.070000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.750000 43.470000 4.070000 43.790000 ;
      LAYER met4 ;
        RECT 3.750000 43.470000 4.070000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.750000 43.900000 4.070000 44.220000 ;
      LAYER met4 ;
        RECT 3.750000 43.900000 4.070000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.150000 39.600000 4.470000 39.920000 ;
      LAYER met4 ;
        RECT 4.150000 39.600000 4.470000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.150000 40.030000 4.470000 40.350000 ;
      LAYER met4 ;
        RECT 4.150000 40.030000 4.470000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.150000 40.460000 4.470000 40.780000 ;
      LAYER met4 ;
        RECT 4.150000 40.460000 4.470000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.150000 40.890000 4.470000 41.210000 ;
      LAYER met4 ;
        RECT 4.150000 40.890000 4.470000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.150000 41.320000 4.470000 41.640000 ;
      LAYER met4 ;
        RECT 4.150000 41.320000 4.470000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.150000 41.750000 4.470000 42.070000 ;
      LAYER met4 ;
        RECT 4.150000 41.750000 4.470000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.150000 42.180000 4.470000 42.500000 ;
      LAYER met4 ;
        RECT 4.150000 42.180000 4.470000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.150000 42.610000 4.470000 42.930000 ;
      LAYER met4 ;
        RECT 4.150000 42.610000 4.470000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.150000 43.040000 4.470000 43.360000 ;
      LAYER met4 ;
        RECT 4.150000 43.040000 4.470000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.150000 43.470000 4.470000 43.790000 ;
      LAYER met4 ;
        RECT 4.150000 43.470000 4.470000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.150000 43.900000 4.470000 44.220000 ;
      LAYER met4 ;
        RECT 4.150000 43.900000 4.470000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550000 39.600000 4.870000 39.920000 ;
      LAYER met4 ;
        RECT 4.550000 39.600000 4.870000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550000 40.030000 4.870000 40.350000 ;
      LAYER met4 ;
        RECT 4.550000 40.030000 4.870000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550000 40.460000 4.870000 40.780000 ;
      LAYER met4 ;
        RECT 4.550000 40.460000 4.870000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550000 40.890000 4.870000 41.210000 ;
      LAYER met4 ;
        RECT 4.550000 40.890000 4.870000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550000 41.320000 4.870000 41.640000 ;
      LAYER met4 ;
        RECT 4.550000 41.320000 4.870000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550000 41.750000 4.870000 42.070000 ;
      LAYER met4 ;
        RECT 4.550000 41.750000 4.870000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550000 42.180000 4.870000 42.500000 ;
      LAYER met4 ;
        RECT 4.550000 42.180000 4.870000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550000 42.610000 4.870000 42.930000 ;
      LAYER met4 ;
        RECT 4.550000 42.610000 4.870000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550000 43.040000 4.870000 43.360000 ;
      LAYER met4 ;
        RECT 4.550000 43.040000 4.870000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550000 43.470000 4.870000 43.790000 ;
      LAYER met4 ;
        RECT 4.550000 43.470000 4.870000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550000 43.900000 4.870000 44.220000 ;
      LAYER met4 ;
        RECT 4.550000 43.900000 4.870000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.950000 39.600000 5.270000 39.920000 ;
      LAYER met4 ;
        RECT 4.950000 39.600000 5.270000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.950000 40.030000 5.270000 40.350000 ;
      LAYER met4 ;
        RECT 4.950000 40.030000 5.270000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.950000 40.460000 5.270000 40.780000 ;
      LAYER met4 ;
        RECT 4.950000 40.460000 5.270000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.950000 40.890000 5.270000 41.210000 ;
      LAYER met4 ;
        RECT 4.950000 40.890000 5.270000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.950000 41.320000 5.270000 41.640000 ;
      LAYER met4 ;
        RECT 4.950000 41.320000 5.270000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.950000 41.750000 5.270000 42.070000 ;
      LAYER met4 ;
        RECT 4.950000 41.750000 5.270000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.950000 42.180000 5.270000 42.500000 ;
      LAYER met4 ;
        RECT 4.950000 42.180000 5.270000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.950000 42.610000 5.270000 42.930000 ;
      LAYER met4 ;
        RECT 4.950000 42.610000 5.270000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.950000 43.040000 5.270000 43.360000 ;
      LAYER met4 ;
        RECT 4.950000 43.040000 5.270000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.950000 43.470000 5.270000 43.790000 ;
      LAYER met4 ;
        RECT 4.950000 43.470000 5.270000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.950000 43.900000 5.270000 44.220000 ;
      LAYER met4 ;
        RECT 4.950000 43.900000 5.270000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.350000 39.600000 5.670000 39.920000 ;
      LAYER met4 ;
        RECT 5.350000 39.600000 5.670000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.350000 40.030000 5.670000 40.350000 ;
      LAYER met4 ;
        RECT 5.350000 40.030000 5.670000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.350000 40.460000 5.670000 40.780000 ;
      LAYER met4 ;
        RECT 5.350000 40.460000 5.670000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.350000 40.890000 5.670000 41.210000 ;
      LAYER met4 ;
        RECT 5.350000 40.890000 5.670000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.350000 41.320000 5.670000 41.640000 ;
      LAYER met4 ;
        RECT 5.350000 41.320000 5.670000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.350000 41.750000 5.670000 42.070000 ;
      LAYER met4 ;
        RECT 5.350000 41.750000 5.670000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.350000 42.180000 5.670000 42.500000 ;
      LAYER met4 ;
        RECT 5.350000 42.180000 5.670000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.350000 42.610000 5.670000 42.930000 ;
      LAYER met4 ;
        RECT 5.350000 42.610000 5.670000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.350000 43.040000 5.670000 43.360000 ;
      LAYER met4 ;
        RECT 5.350000 43.040000 5.670000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.350000 43.470000 5.670000 43.790000 ;
      LAYER met4 ;
        RECT 5.350000 43.470000 5.670000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.350000 43.900000 5.670000 44.220000 ;
      LAYER met4 ;
        RECT 5.350000 43.900000 5.670000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.750000 39.600000 6.070000 39.920000 ;
      LAYER met4 ;
        RECT 5.750000 39.600000 6.070000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.750000 40.030000 6.070000 40.350000 ;
      LAYER met4 ;
        RECT 5.750000 40.030000 6.070000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.750000 40.460000 6.070000 40.780000 ;
      LAYER met4 ;
        RECT 5.750000 40.460000 6.070000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.750000 40.890000 6.070000 41.210000 ;
      LAYER met4 ;
        RECT 5.750000 40.890000 6.070000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.750000 41.320000 6.070000 41.640000 ;
      LAYER met4 ;
        RECT 5.750000 41.320000 6.070000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.750000 41.750000 6.070000 42.070000 ;
      LAYER met4 ;
        RECT 5.750000 41.750000 6.070000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.750000 42.180000 6.070000 42.500000 ;
      LAYER met4 ;
        RECT 5.750000 42.180000 6.070000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.750000 42.610000 6.070000 42.930000 ;
      LAYER met4 ;
        RECT 5.750000 42.610000 6.070000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.750000 43.040000 6.070000 43.360000 ;
      LAYER met4 ;
        RECT 5.750000 43.040000 6.070000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.750000 43.470000 6.070000 43.790000 ;
      LAYER met4 ;
        RECT 5.750000 43.470000 6.070000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.750000 43.900000 6.070000 44.220000 ;
      LAYER met4 ;
        RECT 5.750000 43.900000 6.070000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 39.600000 51.105000 39.920000 ;
      LAYER met4 ;
        RECT 50.785000 39.600000 51.105000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 40.030000 51.105000 40.350000 ;
      LAYER met4 ;
        RECT 50.785000 40.030000 51.105000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 40.460000 51.105000 40.780000 ;
      LAYER met4 ;
        RECT 50.785000 40.460000 51.105000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 40.890000 51.105000 41.210000 ;
      LAYER met4 ;
        RECT 50.785000 40.890000 51.105000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 41.320000 51.105000 41.640000 ;
      LAYER met4 ;
        RECT 50.785000 41.320000 51.105000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 41.750000 51.105000 42.070000 ;
      LAYER met4 ;
        RECT 50.785000 41.750000 51.105000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 42.180000 51.105000 42.500000 ;
      LAYER met4 ;
        RECT 50.785000 42.180000 51.105000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 42.610000 51.105000 42.930000 ;
      LAYER met4 ;
        RECT 50.785000 42.610000 51.105000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 43.040000 51.105000 43.360000 ;
      LAYER met4 ;
        RECT 50.785000 43.040000 51.105000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 43.470000 51.105000 43.790000 ;
      LAYER met4 ;
        RECT 50.785000 43.470000 51.105000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 43.900000 51.105000 44.220000 ;
      LAYER met4 ;
        RECT 50.785000 43.900000 51.105000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 39.600000 51.515000 39.920000 ;
      LAYER met4 ;
        RECT 51.195000 39.600000 51.515000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 40.030000 51.515000 40.350000 ;
      LAYER met4 ;
        RECT 51.195000 40.030000 51.515000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 40.460000 51.515000 40.780000 ;
      LAYER met4 ;
        RECT 51.195000 40.460000 51.515000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 40.890000 51.515000 41.210000 ;
      LAYER met4 ;
        RECT 51.195000 40.890000 51.515000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 41.320000 51.515000 41.640000 ;
      LAYER met4 ;
        RECT 51.195000 41.320000 51.515000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 41.750000 51.515000 42.070000 ;
      LAYER met4 ;
        RECT 51.195000 41.750000 51.515000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 42.180000 51.515000 42.500000 ;
      LAYER met4 ;
        RECT 51.195000 42.180000 51.515000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 42.610000 51.515000 42.930000 ;
      LAYER met4 ;
        RECT 51.195000 42.610000 51.515000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 43.040000 51.515000 43.360000 ;
      LAYER met4 ;
        RECT 51.195000 43.040000 51.515000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 43.470000 51.515000 43.790000 ;
      LAYER met4 ;
        RECT 51.195000 43.470000 51.515000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 43.900000 51.515000 44.220000 ;
      LAYER met4 ;
        RECT 51.195000 43.900000 51.515000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 39.600000 51.925000 39.920000 ;
      LAYER met4 ;
        RECT 51.605000 39.600000 51.925000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 40.030000 51.925000 40.350000 ;
      LAYER met4 ;
        RECT 51.605000 40.030000 51.925000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 40.460000 51.925000 40.780000 ;
      LAYER met4 ;
        RECT 51.605000 40.460000 51.925000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 40.890000 51.925000 41.210000 ;
      LAYER met4 ;
        RECT 51.605000 40.890000 51.925000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 41.320000 51.925000 41.640000 ;
      LAYER met4 ;
        RECT 51.605000 41.320000 51.925000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 41.750000 51.925000 42.070000 ;
      LAYER met4 ;
        RECT 51.605000 41.750000 51.925000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 42.180000 51.925000 42.500000 ;
      LAYER met4 ;
        RECT 51.605000 42.180000 51.925000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 42.610000 51.925000 42.930000 ;
      LAYER met4 ;
        RECT 51.605000 42.610000 51.925000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 43.040000 51.925000 43.360000 ;
      LAYER met4 ;
        RECT 51.605000 43.040000 51.925000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 43.470000 51.925000 43.790000 ;
      LAYER met4 ;
        RECT 51.605000 43.470000 51.925000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 43.900000 51.925000 44.220000 ;
      LAYER met4 ;
        RECT 51.605000 43.900000 51.925000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 39.600000 52.335000 39.920000 ;
      LAYER met4 ;
        RECT 52.015000 39.600000 52.335000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 40.030000 52.335000 40.350000 ;
      LAYER met4 ;
        RECT 52.015000 40.030000 52.335000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 40.460000 52.335000 40.780000 ;
      LAYER met4 ;
        RECT 52.015000 40.460000 52.335000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 40.890000 52.335000 41.210000 ;
      LAYER met4 ;
        RECT 52.015000 40.890000 52.335000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 41.320000 52.335000 41.640000 ;
      LAYER met4 ;
        RECT 52.015000 41.320000 52.335000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 41.750000 52.335000 42.070000 ;
      LAYER met4 ;
        RECT 52.015000 41.750000 52.335000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 42.180000 52.335000 42.500000 ;
      LAYER met4 ;
        RECT 52.015000 42.180000 52.335000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 42.610000 52.335000 42.930000 ;
      LAYER met4 ;
        RECT 52.015000 42.610000 52.335000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 43.040000 52.335000 43.360000 ;
      LAYER met4 ;
        RECT 52.015000 43.040000 52.335000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 43.470000 52.335000 43.790000 ;
      LAYER met4 ;
        RECT 52.015000 43.470000 52.335000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 43.900000 52.335000 44.220000 ;
      LAYER met4 ;
        RECT 52.015000 43.900000 52.335000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 39.600000 52.745000 39.920000 ;
      LAYER met4 ;
        RECT 52.425000 39.600000 52.745000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 40.030000 52.745000 40.350000 ;
      LAYER met4 ;
        RECT 52.425000 40.030000 52.745000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 40.460000 52.745000 40.780000 ;
      LAYER met4 ;
        RECT 52.425000 40.460000 52.745000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 40.890000 52.745000 41.210000 ;
      LAYER met4 ;
        RECT 52.425000 40.890000 52.745000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 41.320000 52.745000 41.640000 ;
      LAYER met4 ;
        RECT 52.425000 41.320000 52.745000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 41.750000 52.745000 42.070000 ;
      LAYER met4 ;
        RECT 52.425000 41.750000 52.745000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 42.180000 52.745000 42.500000 ;
      LAYER met4 ;
        RECT 52.425000 42.180000 52.745000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 42.610000 52.745000 42.930000 ;
      LAYER met4 ;
        RECT 52.425000 42.610000 52.745000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 43.040000 52.745000 43.360000 ;
      LAYER met4 ;
        RECT 52.425000 43.040000 52.745000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 43.470000 52.745000 43.790000 ;
      LAYER met4 ;
        RECT 52.425000 43.470000 52.745000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 43.900000 52.745000 44.220000 ;
      LAYER met4 ;
        RECT 52.425000 43.900000 52.745000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 39.600000 53.155000 39.920000 ;
      LAYER met4 ;
        RECT 52.835000 39.600000 53.155000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 40.030000 53.155000 40.350000 ;
      LAYER met4 ;
        RECT 52.835000 40.030000 53.155000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 40.460000 53.155000 40.780000 ;
      LAYER met4 ;
        RECT 52.835000 40.460000 53.155000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 40.890000 53.155000 41.210000 ;
      LAYER met4 ;
        RECT 52.835000 40.890000 53.155000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 41.320000 53.155000 41.640000 ;
      LAYER met4 ;
        RECT 52.835000 41.320000 53.155000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 41.750000 53.155000 42.070000 ;
      LAYER met4 ;
        RECT 52.835000 41.750000 53.155000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 42.180000 53.155000 42.500000 ;
      LAYER met4 ;
        RECT 52.835000 42.180000 53.155000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 42.610000 53.155000 42.930000 ;
      LAYER met4 ;
        RECT 52.835000 42.610000 53.155000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 43.040000 53.155000 43.360000 ;
      LAYER met4 ;
        RECT 52.835000 43.040000 53.155000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 43.470000 53.155000 43.790000 ;
      LAYER met4 ;
        RECT 52.835000 43.470000 53.155000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 43.900000 53.155000 44.220000 ;
      LAYER met4 ;
        RECT 52.835000 43.900000 53.155000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 39.600000 53.565000 39.920000 ;
      LAYER met4 ;
        RECT 53.245000 39.600000 53.565000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 40.030000 53.565000 40.350000 ;
      LAYER met4 ;
        RECT 53.245000 40.030000 53.565000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 40.460000 53.565000 40.780000 ;
      LAYER met4 ;
        RECT 53.245000 40.460000 53.565000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 40.890000 53.565000 41.210000 ;
      LAYER met4 ;
        RECT 53.245000 40.890000 53.565000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 41.320000 53.565000 41.640000 ;
      LAYER met4 ;
        RECT 53.245000 41.320000 53.565000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 41.750000 53.565000 42.070000 ;
      LAYER met4 ;
        RECT 53.245000 41.750000 53.565000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 42.180000 53.565000 42.500000 ;
      LAYER met4 ;
        RECT 53.245000 42.180000 53.565000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 42.610000 53.565000 42.930000 ;
      LAYER met4 ;
        RECT 53.245000 42.610000 53.565000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 43.040000 53.565000 43.360000 ;
      LAYER met4 ;
        RECT 53.245000 43.040000 53.565000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 43.470000 53.565000 43.790000 ;
      LAYER met4 ;
        RECT 53.245000 43.470000 53.565000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 43.900000 53.565000 44.220000 ;
      LAYER met4 ;
        RECT 53.245000 43.900000 53.565000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 39.600000 53.975000 39.920000 ;
      LAYER met4 ;
        RECT 53.655000 39.600000 53.975000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 40.030000 53.975000 40.350000 ;
      LAYER met4 ;
        RECT 53.655000 40.030000 53.975000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 40.460000 53.975000 40.780000 ;
      LAYER met4 ;
        RECT 53.655000 40.460000 53.975000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 40.890000 53.975000 41.210000 ;
      LAYER met4 ;
        RECT 53.655000 40.890000 53.975000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 41.320000 53.975000 41.640000 ;
      LAYER met4 ;
        RECT 53.655000 41.320000 53.975000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 41.750000 53.975000 42.070000 ;
      LAYER met4 ;
        RECT 53.655000 41.750000 53.975000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 42.180000 53.975000 42.500000 ;
      LAYER met4 ;
        RECT 53.655000 42.180000 53.975000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 42.610000 53.975000 42.930000 ;
      LAYER met4 ;
        RECT 53.655000 42.610000 53.975000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 43.040000 53.975000 43.360000 ;
      LAYER met4 ;
        RECT 53.655000 43.040000 53.975000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 43.470000 53.975000 43.790000 ;
      LAYER met4 ;
        RECT 53.655000 43.470000 53.975000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 43.900000 53.975000 44.220000 ;
      LAYER met4 ;
        RECT 53.655000 43.900000 53.975000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 39.600000 54.385000 39.920000 ;
      LAYER met4 ;
        RECT 54.065000 39.600000 54.385000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 40.030000 54.385000 40.350000 ;
      LAYER met4 ;
        RECT 54.065000 40.030000 54.385000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 40.460000 54.385000 40.780000 ;
      LAYER met4 ;
        RECT 54.065000 40.460000 54.385000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 40.890000 54.385000 41.210000 ;
      LAYER met4 ;
        RECT 54.065000 40.890000 54.385000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 41.320000 54.385000 41.640000 ;
      LAYER met4 ;
        RECT 54.065000 41.320000 54.385000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 41.750000 54.385000 42.070000 ;
      LAYER met4 ;
        RECT 54.065000 41.750000 54.385000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 42.180000 54.385000 42.500000 ;
      LAYER met4 ;
        RECT 54.065000 42.180000 54.385000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 42.610000 54.385000 42.930000 ;
      LAYER met4 ;
        RECT 54.065000 42.610000 54.385000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 43.040000 54.385000 43.360000 ;
      LAYER met4 ;
        RECT 54.065000 43.040000 54.385000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 43.470000 54.385000 43.790000 ;
      LAYER met4 ;
        RECT 54.065000 43.470000 54.385000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 43.900000 54.385000 44.220000 ;
      LAYER met4 ;
        RECT 54.065000 43.900000 54.385000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 39.600000 54.795000 39.920000 ;
      LAYER met4 ;
        RECT 54.475000 39.600000 54.795000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 40.030000 54.795000 40.350000 ;
      LAYER met4 ;
        RECT 54.475000 40.030000 54.795000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 40.460000 54.795000 40.780000 ;
      LAYER met4 ;
        RECT 54.475000 40.460000 54.795000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 40.890000 54.795000 41.210000 ;
      LAYER met4 ;
        RECT 54.475000 40.890000 54.795000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 41.320000 54.795000 41.640000 ;
      LAYER met4 ;
        RECT 54.475000 41.320000 54.795000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 41.750000 54.795000 42.070000 ;
      LAYER met4 ;
        RECT 54.475000 41.750000 54.795000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 42.180000 54.795000 42.500000 ;
      LAYER met4 ;
        RECT 54.475000 42.180000 54.795000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 42.610000 54.795000 42.930000 ;
      LAYER met4 ;
        RECT 54.475000 42.610000 54.795000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 43.040000 54.795000 43.360000 ;
      LAYER met4 ;
        RECT 54.475000 43.040000 54.795000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 43.470000 54.795000 43.790000 ;
      LAYER met4 ;
        RECT 54.475000 43.470000 54.795000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 43.900000 54.795000 44.220000 ;
      LAYER met4 ;
        RECT 54.475000 43.900000 54.795000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 39.600000 55.205000 39.920000 ;
      LAYER met4 ;
        RECT 54.885000 39.600000 55.205000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 40.030000 55.205000 40.350000 ;
      LAYER met4 ;
        RECT 54.885000 40.030000 55.205000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 40.460000 55.205000 40.780000 ;
      LAYER met4 ;
        RECT 54.885000 40.460000 55.205000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 40.890000 55.205000 41.210000 ;
      LAYER met4 ;
        RECT 54.885000 40.890000 55.205000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 41.320000 55.205000 41.640000 ;
      LAYER met4 ;
        RECT 54.885000 41.320000 55.205000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 41.750000 55.205000 42.070000 ;
      LAYER met4 ;
        RECT 54.885000 41.750000 55.205000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 42.180000 55.205000 42.500000 ;
      LAYER met4 ;
        RECT 54.885000 42.180000 55.205000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 42.610000 55.205000 42.930000 ;
      LAYER met4 ;
        RECT 54.885000 42.610000 55.205000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 43.040000 55.205000 43.360000 ;
      LAYER met4 ;
        RECT 54.885000 43.040000 55.205000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 43.470000 55.205000 43.790000 ;
      LAYER met4 ;
        RECT 54.885000 43.470000 55.205000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 43.900000 55.205000 44.220000 ;
      LAYER met4 ;
        RECT 54.885000 43.900000 55.205000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 39.600000 55.615000 39.920000 ;
      LAYER met4 ;
        RECT 55.295000 39.600000 55.615000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 40.030000 55.615000 40.350000 ;
      LAYER met4 ;
        RECT 55.295000 40.030000 55.615000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 40.460000 55.615000 40.780000 ;
      LAYER met4 ;
        RECT 55.295000 40.460000 55.615000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 40.890000 55.615000 41.210000 ;
      LAYER met4 ;
        RECT 55.295000 40.890000 55.615000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 41.320000 55.615000 41.640000 ;
      LAYER met4 ;
        RECT 55.295000 41.320000 55.615000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 41.750000 55.615000 42.070000 ;
      LAYER met4 ;
        RECT 55.295000 41.750000 55.615000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 42.180000 55.615000 42.500000 ;
      LAYER met4 ;
        RECT 55.295000 42.180000 55.615000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 42.610000 55.615000 42.930000 ;
      LAYER met4 ;
        RECT 55.295000 42.610000 55.615000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 43.040000 55.615000 43.360000 ;
      LAYER met4 ;
        RECT 55.295000 43.040000 55.615000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 43.470000 55.615000 43.790000 ;
      LAYER met4 ;
        RECT 55.295000 43.470000 55.615000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 43.900000 55.615000 44.220000 ;
      LAYER met4 ;
        RECT 55.295000 43.900000 55.615000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 39.600000 56.025000 39.920000 ;
      LAYER met4 ;
        RECT 55.705000 39.600000 56.025000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 40.030000 56.025000 40.350000 ;
      LAYER met4 ;
        RECT 55.705000 40.030000 56.025000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 40.460000 56.025000 40.780000 ;
      LAYER met4 ;
        RECT 55.705000 40.460000 56.025000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 40.890000 56.025000 41.210000 ;
      LAYER met4 ;
        RECT 55.705000 40.890000 56.025000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 41.320000 56.025000 41.640000 ;
      LAYER met4 ;
        RECT 55.705000 41.320000 56.025000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 41.750000 56.025000 42.070000 ;
      LAYER met4 ;
        RECT 55.705000 41.750000 56.025000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 42.180000 56.025000 42.500000 ;
      LAYER met4 ;
        RECT 55.705000 42.180000 56.025000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 42.610000 56.025000 42.930000 ;
      LAYER met4 ;
        RECT 55.705000 42.610000 56.025000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 43.040000 56.025000 43.360000 ;
      LAYER met4 ;
        RECT 55.705000 43.040000 56.025000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 43.470000 56.025000 43.790000 ;
      LAYER met4 ;
        RECT 55.705000 43.470000 56.025000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 43.900000 56.025000 44.220000 ;
      LAYER met4 ;
        RECT 55.705000 43.900000 56.025000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 39.600000 56.435000 39.920000 ;
      LAYER met4 ;
        RECT 56.115000 39.600000 56.435000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 40.030000 56.435000 40.350000 ;
      LAYER met4 ;
        RECT 56.115000 40.030000 56.435000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 40.460000 56.435000 40.780000 ;
      LAYER met4 ;
        RECT 56.115000 40.460000 56.435000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 40.890000 56.435000 41.210000 ;
      LAYER met4 ;
        RECT 56.115000 40.890000 56.435000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 41.320000 56.435000 41.640000 ;
      LAYER met4 ;
        RECT 56.115000 41.320000 56.435000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 41.750000 56.435000 42.070000 ;
      LAYER met4 ;
        RECT 56.115000 41.750000 56.435000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 42.180000 56.435000 42.500000 ;
      LAYER met4 ;
        RECT 56.115000 42.180000 56.435000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 42.610000 56.435000 42.930000 ;
      LAYER met4 ;
        RECT 56.115000 42.610000 56.435000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 43.040000 56.435000 43.360000 ;
      LAYER met4 ;
        RECT 56.115000 43.040000 56.435000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 43.470000 56.435000 43.790000 ;
      LAYER met4 ;
        RECT 56.115000 43.470000 56.435000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 43.900000 56.435000 44.220000 ;
      LAYER met4 ;
        RECT 56.115000 43.900000 56.435000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 39.600000 56.845000 39.920000 ;
      LAYER met4 ;
        RECT 56.525000 39.600000 56.845000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 40.030000 56.845000 40.350000 ;
      LAYER met4 ;
        RECT 56.525000 40.030000 56.845000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 40.460000 56.845000 40.780000 ;
      LAYER met4 ;
        RECT 56.525000 40.460000 56.845000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 40.890000 56.845000 41.210000 ;
      LAYER met4 ;
        RECT 56.525000 40.890000 56.845000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 41.320000 56.845000 41.640000 ;
      LAYER met4 ;
        RECT 56.525000 41.320000 56.845000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 41.750000 56.845000 42.070000 ;
      LAYER met4 ;
        RECT 56.525000 41.750000 56.845000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 42.180000 56.845000 42.500000 ;
      LAYER met4 ;
        RECT 56.525000 42.180000 56.845000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 42.610000 56.845000 42.930000 ;
      LAYER met4 ;
        RECT 56.525000 42.610000 56.845000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 43.040000 56.845000 43.360000 ;
      LAYER met4 ;
        RECT 56.525000 43.040000 56.845000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 43.470000 56.845000 43.790000 ;
      LAYER met4 ;
        RECT 56.525000 43.470000 56.845000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 43.900000 56.845000 44.220000 ;
      LAYER met4 ;
        RECT 56.525000 43.900000 56.845000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.935000 39.600000 57.255000 39.920000 ;
      LAYER met4 ;
        RECT 56.935000 39.600000 57.255000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.935000 40.030000 57.255000 40.350000 ;
      LAYER met4 ;
        RECT 56.935000 40.030000 57.255000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.935000 40.460000 57.255000 40.780000 ;
      LAYER met4 ;
        RECT 56.935000 40.460000 57.255000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.935000 40.890000 57.255000 41.210000 ;
      LAYER met4 ;
        RECT 56.935000 40.890000 57.255000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.935000 41.320000 57.255000 41.640000 ;
      LAYER met4 ;
        RECT 56.935000 41.320000 57.255000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.935000 41.750000 57.255000 42.070000 ;
      LAYER met4 ;
        RECT 56.935000 41.750000 57.255000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.935000 42.180000 57.255000 42.500000 ;
      LAYER met4 ;
        RECT 56.935000 42.180000 57.255000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.935000 42.610000 57.255000 42.930000 ;
      LAYER met4 ;
        RECT 56.935000 42.610000 57.255000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.935000 43.040000 57.255000 43.360000 ;
      LAYER met4 ;
        RECT 56.935000 43.040000 57.255000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.935000 43.470000 57.255000 43.790000 ;
      LAYER met4 ;
        RECT 56.935000 43.470000 57.255000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.935000 43.900000 57.255000 44.220000 ;
      LAYER met4 ;
        RECT 56.935000 43.900000 57.255000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.340000 39.600000 57.660000 39.920000 ;
      LAYER met4 ;
        RECT 57.340000 39.600000 57.660000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.340000 40.030000 57.660000 40.350000 ;
      LAYER met4 ;
        RECT 57.340000 40.030000 57.660000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.340000 40.460000 57.660000 40.780000 ;
      LAYER met4 ;
        RECT 57.340000 40.460000 57.660000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.340000 40.890000 57.660000 41.210000 ;
      LAYER met4 ;
        RECT 57.340000 40.890000 57.660000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.340000 41.320000 57.660000 41.640000 ;
      LAYER met4 ;
        RECT 57.340000 41.320000 57.660000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.340000 41.750000 57.660000 42.070000 ;
      LAYER met4 ;
        RECT 57.340000 41.750000 57.660000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.340000 42.180000 57.660000 42.500000 ;
      LAYER met4 ;
        RECT 57.340000 42.180000 57.660000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.340000 42.610000 57.660000 42.930000 ;
      LAYER met4 ;
        RECT 57.340000 42.610000 57.660000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.340000 43.040000 57.660000 43.360000 ;
      LAYER met4 ;
        RECT 57.340000 43.040000 57.660000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.340000 43.470000 57.660000 43.790000 ;
      LAYER met4 ;
        RECT 57.340000 43.470000 57.660000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.340000 43.900000 57.660000 44.220000 ;
      LAYER met4 ;
        RECT 57.340000 43.900000 57.660000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.745000 39.600000 58.065000 39.920000 ;
      LAYER met4 ;
        RECT 57.745000 39.600000 58.065000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.745000 40.030000 58.065000 40.350000 ;
      LAYER met4 ;
        RECT 57.745000 40.030000 58.065000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.745000 40.460000 58.065000 40.780000 ;
      LAYER met4 ;
        RECT 57.745000 40.460000 58.065000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.745000 40.890000 58.065000 41.210000 ;
      LAYER met4 ;
        RECT 57.745000 40.890000 58.065000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.745000 41.320000 58.065000 41.640000 ;
      LAYER met4 ;
        RECT 57.745000 41.320000 58.065000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.745000 41.750000 58.065000 42.070000 ;
      LAYER met4 ;
        RECT 57.745000 41.750000 58.065000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.745000 42.180000 58.065000 42.500000 ;
      LAYER met4 ;
        RECT 57.745000 42.180000 58.065000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.745000 42.610000 58.065000 42.930000 ;
      LAYER met4 ;
        RECT 57.745000 42.610000 58.065000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.745000 43.040000 58.065000 43.360000 ;
      LAYER met4 ;
        RECT 57.745000 43.040000 58.065000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.745000 43.470000 58.065000 43.790000 ;
      LAYER met4 ;
        RECT 57.745000 43.470000 58.065000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.745000 43.900000 58.065000 44.220000 ;
      LAYER met4 ;
        RECT 57.745000 43.900000 58.065000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 39.600000 58.470000 39.920000 ;
      LAYER met4 ;
        RECT 58.150000 39.600000 58.470000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 40.030000 58.470000 40.350000 ;
      LAYER met4 ;
        RECT 58.150000 40.030000 58.470000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 40.460000 58.470000 40.780000 ;
      LAYER met4 ;
        RECT 58.150000 40.460000 58.470000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 40.890000 58.470000 41.210000 ;
      LAYER met4 ;
        RECT 58.150000 40.890000 58.470000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 41.320000 58.470000 41.640000 ;
      LAYER met4 ;
        RECT 58.150000 41.320000 58.470000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 41.750000 58.470000 42.070000 ;
      LAYER met4 ;
        RECT 58.150000 41.750000 58.470000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 42.180000 58.470000 42.500000 ;
      LAYER met4 ;
        RECT 58.150000 42.180000 58.470000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 42.610000 58.470000 42.930000 ;
      LAYER met4 ;
        RECT 58.150000 42.610000 58.470000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 43.040000 58.470000 43.360000 ;
      LAYER met4 ;
        RECT 58.150000 43.040000 58.470000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 43.470000 58.470000 43.790000 ;
      LAYER met4 ;
        RECT 58.150000 43.470000 58.470000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 43.900000 58.470000 44.220000 ;
      LAYER met4 ;
        RECT 58.150000 43.900000 58.470000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.555000 39.600000 58.875000 39.920000 ;
      LAYER met4 ;
        RECT 58.555000 39.600000 58.875000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.555000 40.030000 58.875000 40.350000 ;
      LAYER met4 ;
        RECT 58.555000 40.030000 58.875000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.555000 40.460000 58.875000 40.780000 ;
      LAYER met4 ;
        RECT 58.555000 40.460000 58.875000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.555000 40.890000 58.875000 41.210000 ;
      LAYER met4 ;
        RECT 58.555000 40.890000 58.875000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.555000 41.320000 58.875000 41.640000 ;
      LAYER met4 ;
        RECT 58.555000 41.320000 58.875000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.555000 41.750000 58.875000 42.070000 ;
      LAYER met4 ;
        RECT 58.555000 41.750000 58.875000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.555000 42.180000 58.875000 42.500000 ;
      LAYER met4 ;
        RECT 58.555000 42.180000 58.875000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.555000 42.610000 58.875000 42.930000 ;
      LAYER met4 ;
        RECT 58.555000 42.610000 58.875000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.555000 43.040000 58.875000 43.360000 ;
      LAYER met4 ;
        RECT 58.555000 43.040000 58.875000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.555000 43.470000 58.875000 43.790000 ;
      LAYER met4 ;
        RECT 58.555000 43.470000 58.875000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.555000 43.900000 58.875000 44.220000 ;
      LAYER met4 ;
        RECT 58.555000 43.900000 58.875000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.960000 39.600000 59.280000 39.920000 ;
      LAYER met4 ;
        RECT 58.960000 39.600000 59.280000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.960000 40.030000 59.280000 40.350000 ;
      LAYER met4 ;
        RECT 58.960000 40.030000 59.280000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.960000 40.460000 59.280000 40.780000 ;
      LAYER met4 ;
        RECT 58.960000 40.460000 59.280000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.960000 40.890000 59.280000 41.210000 ;
      LAYER met4 ;
        RECT 58.960000 40.890000 59.280000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.960000 41.320000 59.280000 41.640000 ;
      LAYER met4 ;
        RECT 58.960000 41.320000 59.280000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.960000 41.750000 59.280000 42.070000 ;
      LAYER met4 ;
        RECT 58.960000 41.750000 59.280000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.960000 42.180000 59.280000 42.500000 ;
      LAYER met4 ;
        RECT 58.960000 42.180000 59.280000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.960000 42.610000 59.280000 42.930000 ;
      LAYER met4 ;
        RECT 58.960000 42.610000 59.280000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.960000 43.040000 59.280000 43.360000 ;
      LAYER met4 ;
        RECT 58.960000 43.040000 59.280000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.960000 43.470000 59.280000 43.790000 ;
      LAYER met4 ;
        RECT 58.960000 43.470000 59.280000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.960000 43.900000 59.280000 44.220000 ;
      LAYER met4 ;
        RECT 58.960000 43.900000 59.280000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.365000 39.600000 59.685000 39.920000 ;
      LAYER met4 ;
        RECT 59.365000 39.600000 59.685000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.365000 40.030000 59.685000 40.350000 ;
      LAYER met4 ;
        RECT 59.365000 40.030000 59.685000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.365000 40.460000 59.685000 40.780000 ;
      LAYER met4 ;
        RECT 59.365000 40.460000 59.685000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.365000 40.890000 59.685000 41.210000 ;
      LAYER met4 ;
        RECT 59.365000 40.890000 59.685000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.365000 41.320000 59.685000 41.640000 ;
      LAYER met4 ;
        RECT 59.365000 41.320000 59.685000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.365000 41.750000 59.685000 42.070000 ;
      LAYER met4 ;
        RECT 59.365000 41.750000 59.685000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.365000 42.180000 59.685000 42.500000 ;
      LAYER met4 ;
        RECT 59.365000 42.180000 59.685000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.365000 42.610000 59.685000 42.930000 ;
      LAYER met4 ;
        RECT 59.365000 42.610000 59.685000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.365000 43.040000 59.685000 43.360000 ;
      LAYER met4 ;
        RECT 59.365000 43.040000 59.685000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.365000 43.470000 59.685000 43.790000 ;
      LAYER met4 ;
        RECT 59.365000 43.470000 59.685000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.365000 43.900000 59.685000 44.220000 ;
      LAYER met4 ;
        RECT 59.365000 43.900000 59.685000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.770000 39.600000 60.090000 39.920000 ;
      LAYER met4 ;
        RECT 59.770000 39.600000 60.090000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.770000 40.030000 60.090000 40.350000 ;
      LAYER met4 ;
        RECT 59.770000 40.030000 60.090000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.770000 40.460000 60.090000 40.780000 ;
      LAYER met4 ;
        RECT 59.770000 40.460000 60.090000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.770000 40.890000 60.090000 41.210000 ;
      LAYER met4 ;
        RECT 59.770000 40.890000 60.090000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.770000 41.320000 60.090000 41.640000 ;
      LAYER met4 ;
        RECT 59.770000 41.320000 60.090000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.770000 41.750000 60.090000 42.070000 ;
      LAYER met4 ;
        RECT 59.770000 41.750000 60.090000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.770000 42.180000 60.090000 42.500000 ;
      LAYER met4 ;
        RECT 59.770000 42.180000 60.090000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.770000 42.610000 60.090000 42.930000 ;
      LAYER met4 ;
        RECT 59.770000 42.610000 60.090000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.770000 43.040000 60.090000 43.360000 ;
      LAYER met4 ;
        RECT 59.770000 43.040000 60.090000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.770000 43.470000 60.090000 43.790000 ;
      LAYER met4 ;
        RECT 59.770000 43.470000 60.090000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.770000 43.900000 60.090000 44.220000 ;
      LAYER met4 ;
        RECT 59.770000 43.900000 60.090000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.150000 39.600000 6.470000 39.920000 ;
      LAYER met4 ;
        RECT 6.150000 39.600000 6.470000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.150000 40.030000 6.470000 40.350000 ;
      LAYER met4 ;
        RECT 6.150000 40.030000 6.470000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.150000 40.460000 6.470000 40.780000 ;
      LAYER met4 ;
        RECT 6.150000 40.460000 6.470000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.150000 40.890000 6.470000 41.210000 ;
      LAYER met4 ;
        RECT 6.150000 40.890000 6.470000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.150000 41.320000 6.470000 41.640000 ;
      LAYER met4 ;
        RECT 6.150000 41.320000 6.470000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.150000 41.750000 6.470000 42.070000 ;
      LAYER met4 ;
        RECT 6.150000 41.750000 6.470000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.150000 42.180000 6.470000 42.500000 ;
      LAYER met4 ;
        RECT 6.150000 42.180000 6.470000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.150000 42.610000 6.470000 42.930000 ;
      LAYER met4 ;
        RECT 6.150000 42.610000 6.470000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.150000 43.040000 6.470000 43.360000 ;
      LAYER met4 ;
        RECT 6.150000 43.040000 6.470000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.150000 43.470000 6.470000 43.790000 ;
      LAYER met4 ;
        RECT 6.150000 43.470000 6.470000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.150000 43.900000 6.470000 44.220000 ;
      LAYER met4 ;
        RECT 6.150000 43.900000 6.470000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.550000 39.600000 6.870000 39.920000 ;
      LAYER met4 ;
        RECT 6.550000 39.600000 6.870000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.550000 40.030000 6.870000 40.350000 ;
      LAYER met4 ;
        RECT 6.550000 40.030000 6.870000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.550000 40.460000 6.870000 40.780000 ;
      LAYER met4 ;
        RECT 6.550000 40.460000 6.870000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.550000 40.890000 6.870000 41.210000 ;
      LAYER met4 ;
        RECT 6.550000 40.890000 6.870000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.550000 41.320000 6.870000 41.640000 ;
      LAYER met4 ;
        RECT 6.550000 41.320000 6.870000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.550000 41.750000 6.870000 42.070000 ;
      LAYER met4 ;
        RECT 6.550000 41.750000 6.870000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.550000 42.180000 6.870000 42.500000 ;
      LAYER met4 ;
        RECT 6.550000 42.180000 6.870000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.550000 42.610000 6.870000 42.930000 ;
      LAYER met4 ;
        RECT 6.550000 42.610000 6.870000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.550000 43.040000 6.870000 43.360000 ;
      LAYER met4 ;
        RECT 6.550000 43.040000 6.870000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.550000 43.470000 6.870000 43.790000 ;
      LAYER met4 ;
        RECT 6.550000 43.470000 6.870000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.550000 43.900000 6.870000 44.220000 ;
      LAYER met4 ;
        RECT 6.550000 43.900000 6.870000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.950000 39.600000 7.270000 39.920000 ;
      LAYER met4 ;
        RECT 6.950000 39.600000 7.270000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.950000 40.030000 7.270000 40.350000 ;
      LAYER met4 ;
        RECT 6.950000 40.030000 7.270000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.950000 40.460000 7.270000 40.780000 ;
      LAYER met4 ;
        RECT 6.950000 40.460000 7.270000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.950000 40.890000 7.270000 41.210000 ;
      LAYER met4 ;
        RECT 6.950000 40.890000 7.270000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.950000 41.320000 7.270000 41.640000 ;
      LAYER met4 ;
        RECT 6.950000 41.320000 7.270000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.950000 41.750000 7.270000 42.070000 ;
      LAYER met4 ;
        RECT 6.950000 41.750000 7.270000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.950000 42.180000 7.270000 42.500000 ;
      LAYER met4 ;
        RECT 6.950000 42.180000 7.270000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.950000 42.610000 7.270000 42.930000 ;
      LAYER met4 ;
        RECT 6.950000 42.610000 7.270000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.950000 43.040000 7.270000 43.360000 ;
      LAYER met4 ;
        RECT 6.950000 43.040000 7.270000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.950000 43.470000 7.270000 43.790000 ;
      LAYER met4 ;
        RECT 6.950000 43.470000 7.270000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.950000 43.900000 7.270000 44.220000 ;
      LAYER met4 ;
        RECT 6.950000 43.900000 7.270000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.175000 39.600000 60.495000 39.920000 ;
      LAYER met4 ;
        RECT 60.175000 39.600000 60.495000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.175000 40.030000 60.495000 40.350000 ;
      LAYER met4 ;
        RECT 60.175000 40.030000 60.495000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.175000 40.460000 60.495000 40.780000 ;
      LAYER met4 ;
        RECT 60.175000 40.460000 60.495000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.175000 40.890000 60.495000 41.210000 ;
      LAYER met4 ;
        RECT 60.175000 40.890000 60.495000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.175000 41.320000 60.495000 41.640000 ;
      LAYER met4 ;
        RECT 60.175000 41.320000 60.495000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.175000 41.750000 60.495000 42.070000 ;
      LAYER met4 ;
        RECT 60.175000 41.750000 60.495000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.175000 42.180000 60.495000 42.500000 ;
      LAYER met4 ;
        RECT 60.175000 42.180000 60.495000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.175000 42.610000 60.495000 42.930000 ;
      LAYER met4 ;
        RECT 60.175000 42.610000 60.495000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.175000 43.040000 60.495000 43.360000 ;
      LAYER met4 ;
        RECT 60.175000 43.040000 60.495000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.175000 43.470000 60.495000 43.790000 ;
      LAYER met4 ;
        RECT 60.175000 43.470000 60.495000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.175000 43.900000 60.495000 44.220000 ;
      LAYER met4 ;
        RECT 60.175000 43.900000 60.495000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.580000 39.600000 60.900000 39.920000 ;
      LAYER met4 ;
        RECT 60.580000 39.600000 60.900000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.580000 40.030000 60.900000 40.350000 ;
      LAYER met4 ;
        RECT 60.580000 40.030000 60.900000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.580000 40.460000 60.900000 40.780000 ;
      LAYER met4 ;
        RECT 60.580000 40.460000 60.900000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.580000 40.890000 60.900000 41.210000 ;
      LAYER met4 ;
        RECT 60.580000 40.890000 60.900000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.580000 41.320000 60.900000 41.640000 ;
      LAYER met4 ;
        RECT 60.580000 41.320000 60.900000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.580000 41.750000 60.900000 42.070000 ;
      LAYER met4 ;
        RECT 60.580000 41.750000 60.900000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.580000 42.180000 60.900000 42.500000 ;
      LAYER met4 ;
        RECT 60.580000 42.180000 60.900000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.580000 42.610000 60.900000 42.930000 ;
      LAYER met4 ;
        RECT 60.580000 42.610000 60.900000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.580000 43.040000 60.900000 43.360000 ;
      LAYER met4 ;
        RECT 60.580000 43.040000 60.900000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.580000 43.470000 60.900000 43.790000 ;
      LAYER met4 ;
        RECT 60.580000 43.470000 60.900000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.580000 43.900000 60.900000 44.220000 ;
      LAYER met4 ;
        RECT 60.580000 43.900000 60.900000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.985000 39.600000 61.305000 39.920000 ;
      LAYER met4 ;
        RECT 60.985000 39.600000 61.305000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.985000 40.030000 61.305000 40.350000 ;
      LAYER met4 ;
        RECT 60.985000 40.030000 61.305000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.985000 40.460000 61.305000 40.780000 ;
      LAYER met4 ;
        RECT 60.985000 40.460000 61.305000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.985000 40.890000 61.305000 41.210000 ;
      LAYER met4 ;
        RECT 60.985000 40.890000 61.305000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.985000 41.320000 61.305000 41.640000 ;
      LAYER met4 ;
        RECT 60.985000 41.320000 61.305000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.985000 41.750000 61.305000 42.070000 ;
      LAYER met4 ;
        RECT 60.985000 41.750000 61.305000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.985000 42.180000 61.305000 42.500000 ;
      LAYER met4 ;
        RECT 60.985000 42.180000 61.305000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.985000 42.610000 61.305000 42.930000 ;
      LAYER met4 ;
        RECT 60.985000 42.610000 61.305000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.985000 43.040000 61.305000 43.360000 ;
      LAYER met4 ;
        RECT 60.985000 43.040000 61.305000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.985000 43.470000 61.305000 43.790000 ;
      LAYER met4 ;
        RECT 60.985000 43.470000 61.305000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.985000 43.900000 61.305000 44.220000 ;
      LAYER met4 ;
        RECT 60.985000 43.900000 61.305000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.390000 39.600000 61.710000 39.920000 ;
      LAYER met4 ;
        RECT 61.390000 39.600000 61.710000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.390000 40.030000 61.710000 40.350000 ;
      LAYER met4 ;
        RECT 61.390000 40.030000 61.710000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.390000 40.460000 61.710000 40.780000 ;
      LAYER met4 ;
        RECT 61.390000 40.460000 61.710000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.390000 40.890000 61.710000 41.210000 ;
      LAYER met4 ;
        RECT 61.390000 40.890000 61.710000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.390000 41.320000 61.710000 41.640000 ;
      LAYER met4 ;
        RECT 61.390000 41.320000 61.710000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.390000 41.750000 61.710000 42.070000 ;
      LAYER met4 ;
        RECT 61.390000 41.750000 61.710000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.390000 42.180000 61.710000 42.500000 ;
      LAYER met4 ;
        RECT 61.390000 42.180000 61.710000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.390000 42.610000 61.710000 42.930000 ;
      LAYER met4 ;
        RECT 61.390000 42.610000 61.710000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.390000 43.040000 61.710000 43.360000 ;
      LAYER met4 ;
        RECT 61.390000 43.040000 61.710000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.390000 43.470000 61.710000 43.790000 ;
      LAYER met4 ;
        RECT 61.390000 43.470000 61.710000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.390000 43.900000 61.710000 44.220000 ;
      LAYER met4 ;
        RECT 61.390000 43.900000 61.710000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.795000 39.600000 62.115000 39.920000 ;
      LAYER met4 ;
        RECT 61.795000 39.600000 62.115000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.795000 40.030000 62.115000 40.350000 ;
      LAYER met4 ;
        RECT 61.795000 40.030000 62.115000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.795000 40.460000 62.115000 40.780000 ;
      LAYER met4 ;
        RECT 61.795000 40.460000 62.115000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.795000 40.890000 62.115000 41.210000 ;
      LAYER met4 ;
        RECT 61.795000 40.890000 62.115000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.795000 41.320000 62.115000 41.640000 ;
      LAYER met4 ;
        RECT 61.795000 41.320000 62.115000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.795000 41.750000 62.115000 42.070000 ;
      LAYER met4 ;
        RECT 61.795000 41.750000 62.115000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.795000 42.180000 62.115000 42.500000 ;
      LAYER met4 ;
        RECT 61.795000 42.180000 62.115000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.795000 42.610000 62.115000 42.930000 ;
      LAYER met4 ;
        RECT 61.795000 42.610000 62.115000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.795000 43.040000 62.115000 43.360000 ;
      LAYER met4 ;
        RECT 61.795000 43.040000 62.115000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.795000 43.470000 62.115000 43.790000 ;
      LAYER met4 ;
        RECT 61.795000 43.470000 62.115000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.795000 43.900000 62.115000 44.220000 ;
      LAYER met4 ;
        RECT 61.795000 43.900000 62.115000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.200000 39.600000 62.520000 39.920000 ;
      LAYER met4 ;
        RECT 62.200000 39.600000 62.520000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.200000 40.030000 62.520000 40.350000 ;
      LAYER met4 ;
        RECT 62.200000 40.030000 62.520000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.200000 40.460000 62.520000 40.780000 ;
      LAYER met4 ;
        RECT 62.200000 40.460000 62.520000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.200000 40.890000 62.520000 41.210000 ;
      LAYER met4 ;
        RECT 62.200000 40.890000 62.520000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.200000 41.320000 62.520000 41.640000 ;
      LAYER met4 ;
        RECT 62.200000 41.320000 62.520000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.200000 41.750000 62.520000 42.070000 ;
      LAYER met4 ;
        RECT 62.200000 41.750000 62.520000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.200000 42.180000 62.520000 42.500000 ;
      LAYER met4 ;
        RECT 62.200000 42.180000 62.520000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.200000 42.610000 62.520000 42.930000 ;
      LAYER met4 ;
        RECT 62.200000 42.610000 62.520000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.200000 43.040000 62.520000 43.360000 ;
      LAYER met4 ;
        RECT 62.200000 43.040000 62.520000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.200000 43.470000 62.520000 43.790000 ;
      LAYER met4 ;
        RECT 62.200000 43.470000 62.520000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.200000 43.900000 62.520000 44.220000 ;
      LAYER met4 ;
        RECT 62.200000 43.900000 62.520000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.605000 39.600000 62.925000 39.920000 ;
      LAYER met4 ;
        RECT 62.605000 39.600000 62.925000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.605000 40.030000 62.925000 40.350000 ;
      LAYER met4 ;
        RECT 62.605000 40.030000 62.925000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.605000 40.460000 62.925000 40.780000 ;
      LAYER met4 ;
        RECT 62.605000 40.460000 62.925000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.605000 40.890000 62.925000 41.210000 ;
      LAYER met4 ;
        RECT 62.605000 40.890000 62.925000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.605000 41.320000 62.925000 41.640000 ;
      LAYER met4 ;
        RECT 62.605000 41.320000 62.925000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.605000 41.750000 62.925000 42.070000 ;
      LAYER met4 ;
        RECT 62.605000 41.750000 62.925000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.605000 42.180000 62.925000 42.500000 ;
      LAYER met4 ;
        RECT 62.605000 42.180000 62.925000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.605000 42.610000 62.925000 42.930000 ;
      LAYER met4 ;
        RECT 62.605000 42.610000 62.925000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.605000 43.040000 62.925000 43.360000 ;
      LAYER met4 ;
        RECT 62.605000 43.040000 62.925000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.605000 43.470000 62.925000 43.790000 ;
      LAYER met4 ;
        RECT 62.605000 43.470000 62.925000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.605000 43.900000 62.925000 44.220000 ;
      LAYER met4 ;
        RECT 62.605000 43.900000 62.925000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010000 39.600000 63.330000 39.920000 ;
      LAYER met4 ;
        RECT 63.010000 39.600000 63.330000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010000 40.030000 63.330000 40.350000 ;
      LAYER met4 ;
        RECT 63.010000 40.030000 63.330000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010000 40.460000 63.330000 40.780000 ;
      LAYER met4 ;
        RECT 63.010000 40.460000 63.330000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010000 40.890000 63.330000 41.210000 ;
      LAYER met4 ;
        RECT 63.010000 40.890000 63.330000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010000 41.320000 63.330000 41.640000 ;
      LAYER met4 ;
        RECT 63.010000 41.320000 63.330000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010000 41.750000 63.330000 42.070000 ;
      LAYER met4 ;
        RECT 63.010000 41.750000 63.330000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010000 42.180000 63.330000 42.500000 ;
      LAYER met4 ;
        RECT 63.010000 42.180000 63.330000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010000 42.610000 63.330000 42.930000 ;
      LAYER met4 ;
        RECT 63.010000 42.610000 63.330000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010000 43.040000 63.330000 43.360000 ;
      LAYER met4 ;
        RECT 63.010000 43.040000 63.330000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010000 43.470000 63.330000 43.790000 ;
      LAYER met4 ;
        RECT 63.010000 43.470000 63.330000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010000 43.900000 63.330000 44.220000 ;
      LAYER met4 ;
        RECT 63.010000 43.900000 63.330000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.415000 39.600000 63.735000 39.920000 ;
      LAYER met4 ;
        RECT 63.415000 39.600000 63.735000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.415000 40.030000 63.735000 40.350000 ;
      LAYER met4 ;
        RECT 63.415000 40.030000 63.735000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.415000 40.460000 63.735000 40.780000 ;
      LAYER met4 ;
        RECT 63.415000 40.460000 63.735000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.415000 40.890000 63.735000 41.210000 ;
      LAYER met4 ;
        RECT 63.415000 40.890000 63.735000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.415000 41.320000 63.735000 41.640000 ;
      LAYER met4 ;
        RECT 63.415000 41.320000 63.735000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.415000 41.750000 63.735000 42.070000 ;
      LAYER met4 ;
        RECT 63.415000 41.750000 63.735000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.415000 42.180000 63.735000 42.500000 ;
      LAYER met4 ;
        RECT 63.415000 42.180000 63.735000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.415000 42.610000 63.735000 42.930000 ;
      LAYER met4 ;
        RECT 63.415000 42.610000 63.735000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.415000 43.040000 63.735000 43.360000 ;
      LAYER met4 ;
        RECT 63.415000 43.040000 63.735000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.415000 43.470000 63.735000 43.790000 ;
      LAYER met4 ;
        RECT 63.415000 43.470000 63.735000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.415000 43.900000 63.735000 44.220000 ;
      LAYER met4 ;
        RECT 63.415000 43.900000 63.735000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.820000 39.600000 64.140000 39.920000 ;
      LAYER met4 ;
        RECT 63.820000 39.600000 64.140000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.820000 40.030000 64.140000 40.350000 ;
      LAYER met4 ;
        RECT 63.820000 40.030000 64.140000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.820000 40.460000 64.140000 40.780000 ;
      LAYER met4 ;
        RECT 63.820000 40.460000 64.140000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.820000 40.890000 64.140000 41.210000 ;
      LAYER met4 ;
        RECT 63.820000 40.890000 64.140000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.820000 41.320000 64.140000 41.640000 ;
      LAYER met4 ;
        RECT 63.820000 41.320000 64.140000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.820000 41.750000 64.140000 42.070000 ;
      LAYER met4 ;
        RECT 63.820000 41.750000 64.140000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.820000 42.180000 64.140000 42.500000 ;
      LAYER met4 ;
        RECT 63.820000 42.180000 64.140000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.820000 42.610000 64.140000 42.930000 ;
      LAYER met4 ;
        RECT 63.820000 42.610000 64.140000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.820000 43.040000 64.140000 43.360000 ;
      LAYER met4 ;
        RECT 63.820000 43.040000 64.140000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.820000 43.470000 64.140000 43.790000 ;
      LAYER met4 ;
        RECT 63.820000 43.470000 64.140000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.820000 43.900000 64.140000 44.220000 ;
      LAYER met4 ;
        RECT 63.820000 43.900000 64.140000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.225000 39.600000 64.545000 39.920000 ;
      LAYER met4 ;
        RECT 64.225000 39.600000 64.545000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.225000 40.030000 64.545000 40.350000 ;
      LAYER met4 ;
        RECT 64.225000 40.030000 64.545000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.225000 40.460000 64.545000 40.780000 ;
      LAYER met4 ;
        RECT 64.225000 40.460000 64.545000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.225000 40.890000 64.545000 41.210000 ;
      LAYER met4 ;
        RECT 64.225000 40.890000 64.545000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.225000 41.320000 64.545000 41.640000 ;
      LAYER met4 ;
        RECT 64.225000 41.320000 64.545000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.225000 41.750000 64.545000 42.070000 ;
      LAYER met4 ;
        RECT 64.225000 41.750000 64.545000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.225000 42.180000 64.545000 42.500000 ;
      LAYER met4 ;
        RECT 64.225000 42.180000 64.545000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.225000 42.610000 64.545000 42.930000 ;
      LAYER met4 ;
        RECT 64.225000 42.610000 64.545000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.225000 43.040000 64.545000 43.360000 ;
      LAYER met4 ;
        RECT 64.225000 43.040000 64.545000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.225000 43.470000 64.545000 43.790000 ;
      LAYER met4 ;
        RECT 64.225000 43.470000 64.545000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.225000 43.900000 64.545000 44.220000 ;
      LAYER met4 ;
        RECT 64.225000 43.900000 64.545000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.630000 39.600000 64.950000 39.920000 ;
      LAYER met4 ;
        RECT 64.630000 39.600000 64.950000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.630000 40.030000 64.950000 40.350000 ;
      LAYER met4 ;
        RECT 64.630000 40.030000 64.950000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.630000 40.460000 64.950000 40.780000 ;
      LAYER met4 ;
        RECT 64.630000 40.460000 64.950000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.630000 40.890000 64.950000 41.210000 ;
      LAYER met4 ;
        RECT 64.630000 40.890000 64.950000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.630000 41.320000 64.950000 41.640000 ;
      LAYER met4 ;
        RECT 64.630000 41.320000 64.950000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.630000 41.750000 64.950000 42.070000 ;
      LAYER met4 ;
        RECT 64.630000 41.750000 64.950000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.630000 42.180000 64.950000 42.500000 ;
      LAYER met4 ;
        RECT 64.630000 42.180000 64.950000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.630000 42.610000 64.950000 42.930000 ;
      LAYER met4 ;
        RECT 64.630000 42.610000 64.950000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.630000 43.040000 64.950000 43.360000 ;
      LAYER met4 ;
        RECT 64.630000 43.040000 64.950000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.630000 43.470000 64.950000 43.790000 ;
      LAYER met4 ;
        RECT 64.630000 43.470000 64.950000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.630000 43.900000 64.950000 44.220000 ;
      LAYER met4 ;
        RECT 64.630000 43.900000 64.950000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.035000 39.600000 65.355000 39.920000 ;
      LAYER met4 ;
        RECT 65.035000 39.600000 65.355000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.035000 40.030000 65.355000 40.350000 ;
      LAYER met4 ;
        RECT 65.035000 40.030000 65.355000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.035000 40.460000 65.355000 40.780000 ;
      LAYER met4 ;
        RECT 65.035000 40.460000 65.355000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.035000 40.890000 65.355000 41.210000 ;
      LAYER met4 ;
        RECT 65.035000 40.890000 65.355000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.035000 41.320000 65.355000 41.640000 ;
      LAYER met4 ;
        RECT 65.035000 41.320000 65.355000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.035000 41.750000 65.355000 42.070000 ;
      LAYER met4 ;
        RECT 65.035000 41.750000 65.355000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.035000 42.180000 65.355000 42.500000 ;
      LAYER met4 ;
        RECT 65.035000 42.180000 65.355000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.035000 42.610000 65.355000 42.930000 ;
      LAYER met4 ;
        RECT 65.035000 42.610000 65.355000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.035000 43.040000 65.355000 43.360000 ;
      LAYER met4 ;
        RECT 65.035000 43.040000 65.355000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.035000 43.470000 65.355000 43.790000 ;
      LAYER met4 ;
        RECT 65.035000 43.470000 65.355000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.035000 43.900000 65.355000 44.220000 ;
      LAYER met4 ;
        RECT 65.035000 43.900000 65.355000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.440000 39.600000 65.760000 39.920000 ;
      LAYER met4 ;
        RECT 65.440000 39.600000 65.760000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.440000 40.030000 65.760000 40.350000 ;
      LAYER met4 ;
        RECT 65.440000 40.030000 65.760000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.440000 40.460000 65.760000 40.780000 ;
      LAYER met4 ;
        RECT 65.440000 40.460000 65.760000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.440000 40.890000 65.760000 41.210000 ;
      LAYER met4 ;
        RECT 65.440000 40.890000 65.760000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.440000 41.320000 65.760000 41.640000 ;
      LAYER met4 ;
        RECT 65.440000 41.320000 65.760000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.440000 41.750000 65.760000 42.070000 ;
      LAYER met4 ;
        RECT 65.440000 41.750000 65.760000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.440000 42.180000 65.760000 42.500000 ;
      LAYER met4 ;
        RECT 65.440000 42.180000 65.760000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.440000 42.610000 65.760000 42.930000 ;
      LAYER met4 ;
        RECT 65.440000 42.610000 65.760000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.440000 43.040000 65.760000 43.360000 ;
      LAYER met4 ;
        RECT 65.440000 43.040000 65.760000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.440000 43.470000 65.760000 43.790000 ;
      LAYER met4 ;
        RECT 65.440000 43.470000 65.760000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.440000 43.900000 65.760000 44.220000 ;
      LAYER met4 ;
        RECT 65.440000 43.900000 65.760000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.845000 39.600000 66.165000 39.920000 ;
      LAYER met4 ;
        RECT 65.845000 39.600000 66.165000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.845000 40.030000 66.165000 40.350000 ;
      LAYER met4 ;
        RECT 65.845000 40.030000 66.165000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.845000 40.460000 66.165000 40.780000 ;
      LAYER met4 ;
        RECT 65.845000 40.460000 66.165000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.845000 40.890000 66.165000 41.210000 ;
      LAYER met4 ;
        RECT 65.845000 40.890000 66.165000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.845000 41.320000 66.165000 41.640000 ;
      LAYER met4 ;
        RECT 65.845000 41.320000 66.165000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.845000 41.750000 66.165000 42.070000 ;
      LAYER met4 ;
        RECT 65.845000 41.750000 66.165000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.845000 42.180000 66.165000 42.500000 ;
      LAYER met4 ;
        RECT 65.845000 42.180000 66.165000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.845000 42.610000 66.165000 42.930000 ;
      LAYER met4 ;
        RECT 65.845000 42.610000 66.165000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.845000 43.040000 66.165000 43.360000 ;
      LAYER met4 ;
        RECT 65.845000 43.040000 66.165000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.845000 43.470000 66.165000 43.790000 ;
      LAYER met4 ;
        RECT 65.845000 43.470000 66.165000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.845000 43.900000 66.165000 44.220000 ;
      LAYER met4 ;
        RECT 65.845000 43.900000 66.165000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.250000 39.600000 66.570000 39.920000 ;
      LAYER met4 ;
        RECT 66.250000 39.600000 66.570000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.250000 40.030000 66.570000 40.350000 ;
      LAYER met4 ;
        RECT 66.250000 40.030000 66.570000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.250000 40.460000 66.570000 40.780000 ;
      LAYER met4 ;
        RECT 66.250000 40.460000 66.570000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.250000 40.890000 66.570000 41.210000 ;
      LAYER met4 ;
        RECT 66.250000 40.890000 66.570000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.250000 41.320000 66.570000 41.640000 ;
      LAYER met4 ;
        RECT 66.250000 41.320000 66.570000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.250000 41.750000 66.570000 42.070000 ;
      LAYER met4 ;
        RECT 66.250000 41.750000 66.570000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.250000 42.180000 66.570000 42.500000 ;
      LAYER met4 ;
        RECT 66.250000 42.180000 66.570000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.250000 42.610000 66.570000 42.930000 ;
      LAYER met4 ;
        RECT 66.250000 42.610000 66.570000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.250000 43.040000 66.570000 43.360000 ;
      LAYER met4 ;
        RECT 66.250000 43.040000 66.570000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.250000 43.470000 66.570000 43.790000 ;
      LAYER met4 ;
        RECT 66.250000 43.470000 66.570000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.250000 43.900000 66.570000 44.220000 ;
      LAYER met4 ;
        RECT 66.250000 43.900000 66.570000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.655000 39.600000 66.975000 39.920000 ;
      LAYER met4 ;
        RECT 66.655000 39.600000 66.975000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.655000 40.030000 66.975000 40.350000 ;
      LAYER met4 ;
        RECT 66.655000 40.030000 66.975000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.655000 40.460000 66.975000 40.780000 ;
      LAYER met4 ;
        RECT 66.655000 40.460000 66.975000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.655000 40.890000 66.975000 41.210000 ;
      LAYER met4 ;
        RECT 66.655000 40.890000 66.975000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.655000 41.320000 66.975000 41.640000 ;
      LAYER met4 ;
        RECT 66.655000 41.320000 66.975000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.655000 41.750000 66.975000 42.070000 ;
      LAYER met4 ;
        RECT 66.655000 41.750000 66.975000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.655000 42.180000 66.975000 42.500000 ;
      LAYER met4 ;
        RECT 66.655000 42.180000 66.975000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.655000 42.610000 66.975000 42.930000 ;
      LAYER met4 ;
        RECT 66.655000 42.610000 66.975000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.655000 43.040000 66.975000 43.360000 ;
      LAYER met4 ;
        RECT 66.655000 43.040000 66.975000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.655000 43.470000 66.975000 43.790000 ;
      LAYER met4 ;
        RECT 66.655000 43.470000 66.975000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.655000 43.900000 66.975000 44.220000 ;
      LAYER met4 ;
        RECT 66.655000 43.900000 66.975000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060000 39.600000 67.380000 39.920000 ;
      LAYER met4 ;
        RECT 67.060000 39.600000 67.380000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060000 40.030000 67.380000 40.350000 ;
      LAYER met4 ;
        RECT 67.060000 40.030000 67.380000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060000 40.460000 67.380000 40.780000 ;
      LAYER met4 ;
        RECT 67.060000 40.460000 67.380000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060000 40.890000 67.380000 41.210000 ;
      LAYER met4 ;
        RECT 67.060000 40.890000 67.380000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060000 41.320000 67.380000 41.640000 ;
      LAYER met4 ;
        RECT 67.060000 41.320000 67.380000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060000 41.750000 67.380000 42.070000 ;
      LAYER met4 ;
        RECT 67.060000 41.750000 67.380000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060000 42.180000 67.380000 42.500000 ;
      LAYER met4 ;
        RECT 67.060000 42.180000 67.380000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060000 42.610000 67.380000 42.930000 ;
      LAYER met4 ;
        RECT 67.060000 42.610000 67.380000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060000 43.040000 67.380000 43.360000 ;
      LAYER met4 ;
        RECT 67.060000 43.040000 67.380000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060000 43.470000 67.380000 43.790000 ;
      LAYER met4 ;
        RECT 67.060000 43.470000 67.380000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060000 43.900000 67.380000 44.220000 ;
      LAYER met4 ;
        RECT 67.060000 43.900000 67.380000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.465000 39.600000 67.785000 39.920000 ;
      LAYER met4 ;
        RECT 67.465000 39.600000 67.785000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.465000 40.030000 67.785000 40.350000 ;
      LAYER met4 ;
        RECT 67.465000 40.030000 67.785000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.465000 40.460000 67.785000 40.780000 ;
      LAYER met4 ;
        RECT 67.465000 40.460000 67.785000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.465000 40.890000 67.785000 41.210000 ;
      LAYER met4 ;
        RECT 67.465000 40.890000 67.785000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.465000 41.320000 67.785000 41.640000 ;
      LAYER met4 ;
        RECT 67.465000 41.320000 67.785000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.465000 41.750000 67.785000 42.070000 ;
      LAYER met4 ;
        RECT 67.465000 41.750000 67.785000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.465000 42.180000 67.785000 42.500000 ;
      LAYER met4 ;
        RECT 67.465000 42.180000 67.785000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.465000 42.610000 67.785000 42.930000 ;
      LAYER met4 ;
        RECT 67.465000 42.610000 67.785000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.465000 43.040000 67.785000 43.360000 ;
      LAYER met4 ;
        RECT 67.465000 43.040000 67.785000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.465000 43.470000 67.785000 43.790000 ;
      LAYER met4 ;
        RECT 67.465000 43.470000 67.785000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.465000 43.900000 67.785000 44.220000 ;
      LAYER met4 ;
        RECT 67.465000 43.900000 67.785000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.870000 39.600000 68.190000 39.920000 ;
      LAYER met4 ;
        RECT 67.870000 39.600000 68.190000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.870000 40.030000 68.190000 40.350000 ;
      LAYER met4 ;
        RECT 67.870000 40.030000 68.190000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.870000 40.460000 68.190000 40.780000 ;
      LAYER met4 ;
        RECT 67.870000 40.460000 68.190000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.870000 40.890000 68.190000 41.210000 ;
      LAYER met4 ;
        RECT 67.870000 40.890000 68.190000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.870000 41.320000 68.190000 41.640000 ;
      LAYER met4 ;
        RECT 67.870000 41.320000 68.190000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.870000 41.750000 68.190000 42.070000 ;
      LAYER met4 ;
        RECT 67.870000 41.750000 68.190000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.870000 42.180000 68.190000 42.500000 ;
      LAYER met4 ;
        RECT 67.870000 42.180000 68.190000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.870000 42.610000 68.190000 42.930000 ;
      LAYER met4 ;
        RECT 67.870000 42.610000 68.190000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.870000 43.040000 68.190000 43.360000 ;
      LAYER met4 ;
        RECT 67.870000 43.040000 68.190000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.870000 43.470000 68.190000 43.790000 ;
      LAYER met4 ;
        RECT 67.870000 43.470000 68.190000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.870000 43.900000 68.190000 44.220000 ;
      LAYER met4 ;
        RECT 67.870000 43.900000 68.190000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.275000 39.600000 68.595000 39.920000 ;
      LAYER met4 ;
        RECT 68.275000 39.600000 68.595000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.275000 40.030000 68.595000 40.350000 ;
      LAYER met4 ;
        RECT 68.275000 40.030000 68.595000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.275000 40.460000 68.595000 40.780000 ;
      LAYER met4 ;
        RECT 68.275000 40.460000 68.595000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.275000 40.890000 68.595000 41.210000 ;
      LAYER met4 ;
        RECT 68.275000 40.890000 68.595000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.275000 41.320000 68.595000 41.640000 ;
      LAYER met4 ;
        RECT 68.275000 41.320000 68.595000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.275000 41.750000 68.595000 42.070000 ;
      LAYER met4 ;
        RECT 68.275000 41.750000 68.595000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.275000 42.180000 68.595000 42.500000 ;
      LAYER met4 ;
        RECT 68.275000 42.180000 68.595000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.275000 42.610000 68.595000 42.930000 ;
      LAYER met4 ;
        RECT 68.275000 42.610000 68.595000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.275000 43.040000 68.595000 43.360000 ;
      LAYER met4 ;
        RECT 68.275000 43.040000 68.595000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.275000 43.470000 68.595000 43.790000 ;
      LAYER met4 ;
        RECT 68.275000 43.470000 68.595000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.275000 43.900000 68.595000 44.220000 ;
      LAYER met4 ;
        RECT 68.275000 43.900000 68.595000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.680000 39.600000 69.000000 39.920000 ;
      LAYER met4 ;
        RECT 68.680000 39.600000 69.000000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.680000 40.030000 69.000000 40.350000 ;
      LAYER met4 ;
        RECT 68.680000 40.030000 69.000000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.680000 40.460000 69.000000 40.780000 ;
      LAYER met4 ;
        RECT 68.680000 40.460000 69.000000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.680000 40.890000 69.000000 41.210000 ;
      LAYER met4 ;
        RECT 68.680000 40.890000 69.000000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.680000 41.320000 69.000000 41.640000 ;
      LAYER met4 ;
        RECT 68.680000 41.320000 69.000000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.680000 41.750000 69.000000 42.070000 ;
      LAYER met4 ;
        RECT 68.680000 41.750000 69.000000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.680000 42.180000 69.000000 42.500000 ;
      LAYER met4 ;
        RECT 68.680000 42.180000 69.000000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.680000 42.610000 69.000000 42.930000 ;
      LAYER met4 ;
        RECT 68.680000 42.610000 69.000000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.680000 43.040000 69.000000 43.360000 ;
      LAYER met4 ;
        RECT 68.680000 43.040000 69.000000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.680000 43.470000 69.000000 43.790000 ;
      LAYER met4 ;
        RECT 68.680000 43.470000 69.000000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.680000 43.900000 69.000000 44.220000 ;
      LAYER met4 ;
        RECT 68.680000 43.900000 69.000000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.085000 39.600000 69.405000 39.920000 ;
      LAYER met4 ;
        RECT 69.085000 39.600000 69.405000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.085000 40.030000 69.405000 40.350000 ;
      LAYER met4 ;
        RECT 69.085000 40.030000 69.405000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.085000 40.460000 69.405000 40.780000 ;
      LAYER met4 ;
        RECT 69.085000 40.460000 69.405000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.085000 40.890000 69.405000 41.210000 ;
      LAYER met4 ;
        RECT 69.085000 40.890000 69.405000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.085000 41.320000 69.405000 41.640000 ;
      LAYER met4 ;
        RECT 69.085000 41.320000 69.405000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.085000 41.750000 69.405000 42.070000 ;
      LAYER met4 ;
        RECT 69.085000 41.750000 69.405000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.085000 42.180000 69.405000 42.500000 ;
      LAYER met4 ;
        RECT 69.085000 42.180000 69.405000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.085000 42.610000 69.405000 42.930000 ;
      LAYER met4 ;
        RECT 69.085000 42.610000 69.405000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.085000 43.040000 69.405000 43.360000 ;
      LAYER met4 ;
        RECT 69.085000 43.040000 69.405000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.085000 43.470000 69.405000 43.790000 ;
      LAYER met4 ;
        RECT 69.085000 43.470000 69.405000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.085000 43.900000 69.405000 44.220000 ;
      LAYER met4 ;
        RECT 69.085000 43.900000 69.405000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.490000 39.600000 69.810000 39.920000 ;
      LAYER met4 ;
        RECT 69.490000 39.600000 69.810000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.490000 40.030000 69.810000 40.350000 ;
      LAYER met4 ;
        RECT 69.490000 40.030000 69.810000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.490000 40.460000 69.810000 40.780000 ;
      LAYER met4 ;
        RECT 69.490000 40.460000 69.810000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.490000 40.890000 69.810000 41.210000 ;
      LAYER met4 ;
        RECT 69.490000 40.890000 69.810000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.490000 41.320000 69.810000 41.640000 ;
      LAYER met4 ;
        RECT 69.490000 41.320000 69.810000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.490000 41.750000 69.810000 42.070000 ;
      LAYER met4 ;
        RECT 69.490000 41.750000 69.810000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.490000 42.180000 69.810000 42.500000 ;
      LAYER met4 ;
        RECT 69.490000 42.180000 69.810000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.490000 42.610000 69.810000 42.930000 ;
      LAYER met4 ;
        RECT 69.490000 42.610000 69.810000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.490000 43.040000 69.810000 43.360000 ;
      LAYER met4 ;
        RECT 69.490000 43.040000 69.810000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.490000 43.470000 69.810000 43.790000 ;
      LAYER met4 ;
        RECT 69.490000 43.470000 69.810000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.490000 43.900000 69.810000 44.220000 ;
      LAYER met4 ;
        RECT 69.490000 43.900000 69.810000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.895000 39.600000 70.215000 39.920000 ;
      LAYER met4 ;
        RECT 69.895000 39.600000 70.215000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.895000 40.030000 70.215000 40.350000 ;
      LAYER met4 ;
        RECT 69.895000 40.030000 70.215000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.895000 40.460000 70.215000 40.780000 ;
      LAYER met4 ;
        RECT 69.895000 40.460000 70.215000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.895000 40.890000 70.215000 41.210000 ;
      LAYER met4 ;
        RECT 69.895000 40.890000 70.215000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.895000 41.320000 70.215000 41.640000 ;
      LAYER met4 ;
        RECT 69.895000 41.320000 70.215000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.895000 41.750000 70.215000 42.070000 ;
      LAYER met4 ;
        RECT 69.895000 41.750000 70.215000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.895000 42.180000 70.215000 42.500000 ;
      LAYER met4 ;
        RECT 69.895000 42.180000 70.215000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.895000 42.610000 70.215000 42.930000 ;
      LAYER met4 ;
        RECT 69.895000 42.610000 70.215000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.895000 43.040000 70.215000 43.360000 ;
      LAYER met4 ;
        RECT 69.895000 43.040000 70.215000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.895000 43.470000 70.215000 43.790000 ;
      LAYER met4 ;
        RECT 69.895000 43.470000 70.215000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.895000 43.900000 70.215000 44.220000 ;
      LAYER met4 ;
        RECT 69.895000 43.900000 70.215000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.350000 39.600000 7.670000 39.920000 ;
      LAYER met4 ;
        RECT 7.350000 39.600000 7.670000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.350000 40.030000 7.670000 40.350000 ;
      LAYER met4 ;
        RECT 7.350000 40.030000 7.670000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.350000 40.460000 7.670000 40.780000 ;
      LAYER met4 ;
        RECT 7.350000 40.460000 7.670000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.350000 40.890000 7.670000 41.210000 ;
      LAYER met4 ;
        RECT 7.350000 40.890000 7.670000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.350000 41.320000 7.670000 41.640000 ;
      LAYER met4 ;
        RECT 7.350000 41.320000 7.670000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.350000 41.750000 7.670000 42.070000 ;
      LAYER met4 ;
        RECT 7.350000 41.750000 7.670000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.350000 42.180000 7.670000 42.500000 ;
      LAYER met4 ;
        RECT 7.350000 42.180000 7.670000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.350000 42.610000 7.670000 42.930000 ;
      LAYER met4 ;
        RECT 7.350000 42.610000 7.670000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.350000 43.040000 7.670000 43.360000 ;
      LAYER met4 ;
        RECT 7.350000 43.040000 7.670000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.350000 43.470000 7.670000 43.790000 ;
      LAYER met4 ;
        RECT 7.350000 43.470000 7.670000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.350000 43.900000 7.670000 44.220000 ;
      LAYER met4 ;
        RECT 7.350000 43.900000 7.670000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.750000 39.600000 8.070000 39.920000 ;
      LAYER met4 ;
        RECT 7.750000 39.600000 8.070000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.750000 40.030000 8.070000 40.350000 ;
      LAYER met4 ;
        RECT 7.750000 40.030000 8.070000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.750000 40.460000 8.070000 40.780000 ;
      LAYER met4 ;
        RECT 7.750000 40.460000 8.070000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.750000 40.890000 8.070000 41.210000 ;
      LAYER met4 ;
        RECT 7.750000 40.890000 8.070000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.750000 41.320000 8.070000 41.640000 ;
      LAYER met4 ;
        RECT 7.750000 41.320000 8.070000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.750000 41.750000 8.070000 42.070000 ;
      LAYER met4 ;
        RECT 7.750000 41.750000 8.070000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.750000 42.180000 8.070000 42.500000 ;
      LAYER met4 ;
        RECT 7.750000 42.180000 8.070000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.750000 42.610000 8.070000 42.930000 ;
      LAYER met4 ;
        RECT 7.750000 42.610000 8.070000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.750000 43.040000 8.070000 43.360000 ;
      LAYER met4 ;
        RECT 7.750000 43.040000 8.070000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.750000 43.470000 8.070000 43.790000 ;
      LAYER met4 ;
        RECT 7.750000 43.470000 8.070000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.750000 43.900000 8.070000 44.220000 ;
      LAYER met4 ;
        RECT 7.750000 43.900000 8.070000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.300000 39.600000 70.620000 39.920000 ;
      LAYER met4 ;
        RECT 70.300000 39.600000 70.620000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.300000 40.030000 70.620000 40.350000 ;
      LAYER met4 ;
        RECT 70.300000 40.030000 70.620000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.300000 40.460000 70.620000 40.780000 ;
      LAYER met4 ;
        RECT 70.300000 40.460000 70.620000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.300000 40.890000 70.620000 41.210000 ;
      LAYER met4 ;
        RECT 70.300000 40.890000 70.620000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.300000 41.320000 70.620000 41.640000 ;
      LAYER met4 ;
        RECT 70.300000 41.320000 70.620000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.300000 41.750000 70.620000 42.070000 ;
      LAYER met4 ;
        RECT 70.300000 41.750000 70.620000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.300000 42.180000 70.620000 42.500000 ;
      LAYER met4 ;
        RECT 70.300000 42.180000 70.620000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.300000 42.610000 70.620000 42.930000 ;
      LAYER met4 ;
        RECT 70.300000 42.610000 70.620000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.300000 43.040000 70.620000 43.360000 ;
      LAYER met4 ;
        RECT 70.300000 43.040000 70.620000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.300000 43.470000 70.620000 43.790000 ;
      LAYER met4 ;
        RECT 70.300000 43.470000 70.620000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.300000 43.900000 70.620000 44.220000 ;
      LAYER met4 ;
        RECT 70.300000 43.900000 70.620000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.705000 39.600000 71.025000 39.920000 ;
      LAYER met4 ;
        RECT 70.705000 39.600000 71.025000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.705000 40.030000 71.025000 40.350000 ;
      LAYER met4 ;
        RECT 70.705000 40.030000 71.025000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.705000 40.460000 71.025000 40.780000 ;
      LAYER met4 ;
        RECT 70.705000 40.460000 71.025000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.705000 40.890000 71.025000 41.210000 ;
      LAYER met4 ;
        RECT 70.705000 40.890000 71.025000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.705000 41.320000 71.025000 41.640000 ;
      LAYER met4 ;
        RECT 70.705000 41.320000 71.025000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.705000 41.750000 71.025000 42.070000 ;
      LAYER met4 ;
        RECT 70.705000 41.750000 71.025000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.705000 42.180000 71.025000 42.500000 ;
      LAYER met4 ;
        RECT 70.705000 42.180000 71.025000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.705000 42.610000 71.025000 42.930000 ;
      LAYER met4 ;
        RECT 70.705000 42.610000 71.025000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.705000 43.040000 71.025000 43.360000 ;
      LAYER met4 ;
        RECT 70.705000 43.040000 71.025000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.705000 43.470000 71.025000 43.790000 ;
      LAYER met4 ;
        RECT 70.705000 43.470000 71.025000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.705000 43.900000 71.025000 44.220000 ;
      LAYER met4 ;
        RECT 70.705000 43.900000 71.025000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.110000 39.600000 71.430000 39.920000 ;
      LAYER met4 ;
        RECT 71.110000 39.600000 71.430000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.110000 40.030000 71.430000 40.350000 ;
      LAYER met4 ;
        RECT 71.110000 40.030000 71.430000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.110000 40.460000 71.430000 40.780000 ;
      LAYER met4 ;
        RECT 71.110000 40.460000 71.430000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.110000 40.890000 71.430000 41.210000 ;
      LAYER met4 ;
        RECT 71.110000 40.890000 71.430000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.110000 41.320000 71.430000 41.640000 ;
      LAYER met4 ;
        RECT 71.110000 41.320000 71.430000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.110000 41.750000 71.430000 42.070000 ;
      LAYER met4 ;
        RECT 71.110000 41.750000 71.430000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.110000 42.180000 71.430000 42.500000 ;
      LAYER met4 ;
        RECT 71.110000 42.180000 71.430000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.110000 42.610000 71.430000 42.930000 ;
      LAYER met4 ;
        RECT 71.110000 42.610000 71.430000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.110000 43.040000 71.430000 43.360000 ;
      LAYER met4 ;
        RECT 71.110000 43.040000 71.430000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.110000 43.470000 71.430000 43.790000 ;
      LAYER met4 ;
        RECT 71.110000 43.470000 71.430000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.110000 43.900000 71.430000 44.220000 ;
      LAYER met4 ;
        RECT 71.110000 43.900000 71.430000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.515000 39.600000 71.835000 39.920000 ;
      LAYER met4 ;
        RECT 71.515000 39.600000 71.835000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.515000 40.030000 71.835000 40.350000 ;
      LAYER met4 ;
        RECT 71.515000 40.030000 71.835000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.515000 40.460000 71.835000 40.780000 ;
      LAYER met4 ;
        RECT 71.515000 40.460000 71.835000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.515000 40.890000 71.835000 41.210000 ;
      LAYER met4 ;
        RECT 71.515000 40.890000 71.835000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.515000 41.320000 71.835000 41.640000 ;
      LAYER met4 ;
        RECT 71.515000 41.320000 71.835000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.515000 41.750000 71.835000 42.070000 ;
      LAYER met4 ;
        RECT 71.515000 41.750000 71.835000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.515000 42.180000 71.835000 42.500000 ;
      LAYER met4 ;
        RECT 71.515000 42.180000 71.835000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.515000 42.610000 71.835000 42.930000 ;
      LAYER met4 ;
        RECT 71.515000 42.610000 71.835000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.515000 43.040000 71.835000 43.360000 ;
      LAYER met4 ;
        RECT 71.515000 43.040000 71.835000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.515000 43.470000 71.835000 43.790000 ;
      LAYER met4 ;
        RECT 71.515000 43.470000 71.835000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.515000 43.900000 71.835000 44.220000 ;
      LAYER met4 ;
        RECT 71.515000 43.900000 71.835000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 39.600000 72.240000 39.920000 ;
      LAYER met4 ;
        RECT 71.920000 39.600000 72.240000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 40.030000 72.240000 40.350000 ;
      LAYER met4 ;
        RECT 71.920000 40.030000 72.240000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 40.460000 72.240000 40.780000 ;
      LAYER met4 ;
        RECT 71.920000 40.460000 72.240000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 40.890000 72.240000 41.210000 ;
      LAYER met4 ;
        RECT 71.920000 40.890000 72.240000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 41.320000 72.240000 41.640000 ;
      LAYER met4 ;
        RECT 71.920000 41.320000 72.240000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 41.750000 72.240000 42.070000 ;
      LAYER met4 ;
        RECT 71.920000 41.750000 72.240000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 42.180000 72.240000 42.500000 ;
      LAYER met4 ;
        RECT 71.920000 42.180000 72.240000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 42.610000 72.240000 42.930000 ;
      LAYER met4 ;
        RECT 71.920000 42.610000 72.240000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 43.040000 72.240000 43.360000 ;
      LAYER met4 ;
        RECT 71.920000 43.040000 72.240000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 43.470000 72.240000 43.790000 ;
      LAYER met4 ;
        RECT 71.920000 43.470000 72.240000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 43.900000 72.240000 44.220000 ;
      LAYER met4 ;
        RECT 71.920000 43.900000 72.240000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.325000 39.600000 72.645000 39.920000 ;
      LAYER met4 ;
        RECT 72.325000 39.600000 72.645000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.325000 40.030000 72.645000 40.350000 ;
      LAYER met4 ;
        RECT 72.325000 40.030000 72.645000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.325000 40.460000 72.645000 40.780000 ;
      LAYER met4 ;
        RECT 72.325000 40.460000 72.645000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.325000 40.890000 72.645000 41.210000 ;
      LAYER met4 ;
        RECT 72.325000 40.890000 72.645000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.325000 41.320000 72.645000 41.640000 ;
      LAYER met4 ;
        RECT 72.325000 41.320000 72.645000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.325000 41.750000 72.645000 42.070000 ;
      LAYER met4 ;
        RECT 72.325000 41.750000 72.645000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.325000 42.180000 72.645000 42.500000 ;
      LAYER met4 ;
        RECT 72.325000 42.180000 72.645000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.325000 42.610000 72.645000 42.930000 ;
      LAYER met4 ;
        RECT 72.325000 42.610000 72.645000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.325000 43.040000 72.645000 43.360000 ;
      LAYER met4 ;
        RECT 72.325000 43.040000 72.645000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.325000 43.470000 72.645000 43.790000 ;
      LAYER met4 ;
        RECT 72.325000 43.470000 72.645000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.325000 43.900000 72.645000 44.220000 ;
      LAYER met4 ;
        RECT 72.325000 43.900000 72.645000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 39.600000 73.050000 39.920000 ;
      LAYER met4 ;
        RECT 72.730000 39.600000 73.050000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 40.030000 73.050000 40.350000 ;
      LAYER met4 ;
        RECT 72.730000 40.030000 73.050000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 40.460000 73.050000 40.780000 ;
      LAYER met4 ;
        RECT 72.730000 40.460000 73.050000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 40.890000 73.050000 41.210000 ;
      LAYER met4 ;
        RECT 72.730000 40.890000 73.050000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 41.320000 73.050000 41.640000 ;
      LAYER met4 ;
        RECT 72.730000 41.320000 73.050000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 41.750000 73.050000 42.070000 ;
      LAYER met4 ;
        RECT 72.730000 41.750000 73.050000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 42.180000 73.050000 42.500000 ;
      LAYER met4 ;
        RECT 72.730000 42.180000 73.050000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 42.610000 73.050000 42.930000 ;
      LAYER met4 ;
        RECT 72.730000 42.610000 73.050000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 43.040000 73.050000 43.360000 ;
      LAYER met4 ;
        RECT 72.730000 43.040000 73.050000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 43.470000 73.050000 43.790000 ;
      LAYER met4 ;
        RECT 72.730000 43.470000 73.050000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730000 43.900000 73.050000 44.220000 ;
      LAYER met4 ;
        RECT 72.730000 43.900000 73.050000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135000 39.600000 73.455000 39.920000 ;
      LAYER met4 ;
        RECT 73.135000 39.600000 73.455000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135000 40.030000 73.455000 40.350000 ;
      LAYER met4 ;
        RECT 73.135000 40.030000 73.455000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135000 40.460000 73.455000 40.780000 ;
      LAYER met4 ;
        RECT 73.135000 40.460000 73.455000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135000 40.890000 73.455000 41.210000 ;
      LAYER met4 ;
        RECT 73.135000 40.890000 73.455000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135000 41.320000 73.455000 41.640000 ;
      LAYER met4 ;
        RECT 73.135000 41.320000 73.455000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135000 41.750000 73.455000 42.070000 ;
      LAYER met4 ;
        RECT 73.135000 41.750000 73.455000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135000 42.180000 73.455000 42.500000 ;
      LAYER met4 ;
        RECT 73.135000 42.180000 73.455000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135000 42.610000 73.455000 42.930000 ;
      LAYER met4 ;
        RECT 73.135000 42.610000 73.455000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135000 43.040000 73.455000 43.360000 ;
      LAYER met4 ;
        RECT 73.135000 43.040000 73.455000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135000 43.470000 73.455000 43.790000 ;
      LAYER met4 ;
        RECT 73.135000 43.470000 73.455000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135000 43.900000 73.455000 44.220000 ;
      LAYER met4 ;
        RECT 73.135000 43.900000 73.455000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.540000 39.600000 73.860000 39.920000 ;
      LAYER met4 ;
        RECT 73.540000 39.600000 73.860000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.540000 40.030000 73.860000 40.350000 ;
      LAYER met4 ;
        RECT 73.540000 40.030000 73.860000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.540000 40.460000 73.860000 40.780000 ;
      LAYER met4 ;
        RECT 73.540000 40.460000 73.860000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.540000 40.890000 73.860000 41.210000 ;
      LAYER met4 ;
        RECT 73.540000 40.890000 73.860000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.540000 41.320000 73.860000 41.640000 ;
      LAYER met4 ;
        RECT 73.540000 41.320000 73.860000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.540000 41.750000 73.860000 42.070000 ;
      LAYER met4 ;
        RECT 73.540000 41.750000 73.860000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.540000 42.180000 73.860000 42.500000 ;
      LAYER met4 ;
        RECT 73.540000 42.180000 73.860000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.540000 42.610000 73.860000 42.930000 ;
      LAYER met4 ;
        RECT 73.540000 42.610000 73.860000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.540000 43.040000 73.860000 43.360000 ;
      LAYER met4 ;
        RECT 73.540000 43.040000 73.860000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.540000 43.470000 73.860000 43.790000 ;
      LAYER met4 ;
        RECT 73.540000 43.470000 73.860000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.540000 43.900000 73.860000 44.220000 ;
      LAYER met4 ;
        RECT 73.540000 43.900000 73.860000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.945000 39.600000 74.265000 39.920000 ;
      LAYER met4 ;
        RECT 73.945000 39.600000 74.265000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.945000 40.030000 74.265000 40.350000 ;
      LAYER met4 ;
        RECT 73.945000 40.030000 74.265000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.945000 40.460000 74.265000 40.780000 ;
      LAYER met4 ;
        RECT 73.945000 40.460000 74.265000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.945000 40.890000 74.265000 41.210000 ;
      LAYER met4 ;
        RECT 73.945000 40.890000 74.265000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.945000 41.320000 74.265000 41.640000 ;
      LAYER met4 ;
        RECT 73.945000 41.320000 74.265000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.945000 41.750000 74.265000 42.070000 ;
      LAYER met4 ;
        RECT 73.945000 41.750000 74.265000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.945000 42.180000 74.265000 42.500000 ;
      LAYER met4 ;
        RECT 73.945000 42.180000 74.265000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.945000 42.610000 74.265000 42.930000 ;
      LAYER met4 ;
        RECT 73.945000 42.610000 74.265000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.945000 43.040000 74.265000 43.360000 ;
      LAYER met4 ;
        RECT 73.945000 43.040000 74.265000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.945000 43.470000 74.265000 43.790000 ;
      LAYER met4 ;
        RECT 73.945000 43.470000 74.265000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.945000 43.900000 74.265000 44.220000 ;
      LAYER met4 ;
        RECT 73.945000 43.900000 74.265000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.350000 39.600000 74.670000 39.920000 ;
      LAYER met4 ;
        RECT 74.350000 39.600000 74.670000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.350000 40.030000 74.670000 40.350000 ;
      LAYER met4 ;
        RECT 74.350000 40.030000 74.670000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.350000 40.460000 74.670000 40.780000 ;
      LAYER met4 ;
        RECT 74.350000 40.460000 74.670000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.350000 40.890000 74.670000 41.210000 ;
      LAYER met4 ;
        RECT 74.350000 40.890000 74.670000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.350000 41.320000 74.670000 41.640000 ;
      LAYER met4 ;
        RECT 74.350000 41.320000 74.670000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.350000 41.750000 74.670000 42.070000 ;
      LAYER met4 ;
        RECT 74.350000 41.750000 74.670000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.350000 42.180000 74.670000 42.500000 ;
      LAYER met4 ;
        RECT 74.350000 42.180000 74.670000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.350000 42.610000 74.670000 42.930000 ;
      LAYER met4 ;
        RECT 74.350000 42.610000 74.670000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.350000 43.040000 74.670000 43.360000 ;
      LAYER met4 ;
        RECT 74.350000 43.040000 74.670000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.350000 43.470000 74.670000 43.790000 ;
      LAYER met4 ;
        RECT 74.350000 43.470000 74.670000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.350000 43.900000 74.670000 44.220000 ;
      LAYER met4 ;
        RECT 74.350000 43.900000 74.670000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150000 39.600000 8.470000 39.920000 ;
      LAYER met4 ;
        RECT 8.150000 39.600000 8.470000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150000 40.030000 8.470000 40.350000 ;
      LAYER met4 ;
        RECT 8.150000 40.030000 8.470000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150000 40.460000 8.470000 40.780000 ;
      LAYER met4 ;
        RECT 8.150000 40.460000 8.470000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150000 40.890000 8.470000 41.210000 ;
      LAYER met4 ;
        RECT 8.150000 40.890000 8.470000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150000 41.320000 8.470000 41.640000 ;
      LAYER met4 ;
        RECT 8.150000 41.320000 8.470000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150000 41.750000 8.470000 42.070000 ;
      LAYER met4 ;
        RECT 8.150000 41.750000 8.470000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150000 42.180000 8.470000 42.500000 ;
      LAYER met4 ;
        RECT 8.150000 42.180000 8.470000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150000 42.610000 8.470000 42.930000 ;
      LAYER met4 ;
        RECT 8.150000 42.610000 8.470000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150000 43.040000 8.470000 43.360000 ;
      LAYER met4 ;
        RECT 8.150000 43.040000 8.470000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150000 43.470000 8.470000 43.790000 ;
      LAYER met4 ;
        RECT 8.150000 43.470000 8.470000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150000 43.900000 8.470000 44.220000 ;
      LAYER met4 ;
        RECT 8.150000 43.900000 8.470000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.550000 39.600000 8.870000 39.920000 ;
      LAYER met4 ;
        RECT 8.550000 39.600000 8.870000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.550000 40.030000 8.870000 40.350000 ;
      LAYER met4 ;
        RECT 8.550000 40.030000 8.870000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.550000 40.460000 8.870000 40.780000 ;
      LAYER met4 ;
        RECT 8.550000 40.460000 8.870000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.550000 40.890000 8.870000 41.210000 ;
      LAYER met4 ;
        RECT 8.550000 40.890000 8.870000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.550000 41.320000 8.870000 41.640000 ;
      LAYER met4 ;
        RECT 8.550000 41.320000 8.870000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.550000 41.750000 8.870000 42.070000 ;
      LAYER met4 ;
        RECT 8.550000 41.750000 8.870000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.550000 42.180000 8.870000 42.500000 ;
      LAYER met4 ;
        RECT 8.550000 42.180000 8.870000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.550000 42.610000 8.870000 42.930000 ;
      LAYER met4 ;
        RECT 8.550000 42.610000 8.870000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.550000 43.040000 8.870000 43.360000 ;
      LAYER met4 ;
        RECT 8.550000 43.040000 8.870000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.550000 43.470000 8.870000 43.790000 ;
      LAYER met4 ;
        RECT 8.550000 43.470000 8.870000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.550000 43.900000 8.870000 44.220000 ;
      LAYER met4 ;
        RECT 8.550000 43.900000 8.870000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.950000 39.600000 9.270000 39.920000 ;
      LAYER met4 ;
        RECT 8.950000 39.600000 9.270000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.950000 40.030000 9.270000 40.350000 ;
      LAYER met4 ;
        RECT 8.950000 40.030000 9.270000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.950000 40.460000 9.270000 40.780000 ;
      LAYER met4 ;
        RECT 8.950000 40.460000 9.270000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.950000 40.890000 9.270000 41.210000 ;
      LAYER met4 ;
        RECT 8.950000 40.890000 9.270000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.950000 41.320000 9.270000 41.640000 ;
      LAYER met4 ;
        RECT 8.950000 41.320000 9.270000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.950000 41.750000 9.270000 42.070000 ;
      LAYER met4 ;
        RECT 8.950000 41.750000 9.270000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.950000 42.180000 9.270000 42.500000 ;
      LAYER met4 ;
        RECT 8.950000 42.180000 9.270000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.950000 42.610000 9.270000 42.930000 ;
      LAYER met4 ;
        RECT 8.950000 42.610000 9.270000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.950000 43.040000 9.270000 43.360000 ;
      LAYER met4 ;
        RECT 8.950000 43.040000 9.270000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.950000 43.470000 9.270000 43.790000 ;
      LAYER met4 ;
        RECT 8.950000 43.470000 9.270000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.950000 43.900000 9.270000 44.220000 ;
      LAYER met4 ;
        RECT 8.950000 43.900000 9.270000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.350000 39.600000 9.670000 39.920000 ;
      LAYER met4 ;
        RECT 9.350000 39.600000 9.670000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.350000 40.030000 9.670000 40.350000 ;
      LAYER met4 ;
        RECT 9.350000 40.030000 9.670000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.350000 40.460000 9.670000 40.780000 ;
      LAYER met4 ;
        RECT 9.350000 40.460000 9.670000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.350000 40.890000 9.670000 41.210000 ;
      LAYER met4 ;
        RECT 9.350000 40.890000 9.670000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.350000 41.320000 9.670000 41.640000 ;
      LAYER met4 ;
        RECT 9.350000 41.320000 9.670000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.350000 41.750000 9.670000 42.070000 ;
      LAYER met4 ;
        RECT 9.350000 41.750000 9.670000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.350000 42.180000 9.670000 42.500000 ;
      LAYER met4 ;
        RECT 9.350000 42.180000 9.670000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.350000 42.610000 9.670000 42.930000 ;
      LAYER met4 ;
        RECT 9.350000 42.610000 9.670000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.350000 43.040000 9.670000 43.360000 ;
      LAYER met4 ;
        RECT 9.350000 43.040000 9.670000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.350000 43.470000 9.670000 43.790000 ;
      LAYER met4 ;
        RECT 9.350000 43.470000 9.670000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.350000 43.900000 9.670000 44.220000 ;
      LAYER met4 ;
        RECT 9.350000 43.900000 9.670000 44.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.750000 39.600000 10.070000 39.920000 ;
      LAYER met4 ;
        RECT 9.750000 39.600000 10.070000 39.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.750000 40.030000 10.070000 40.350000 ;
      LAYER met4 ;
        RECT 9.750000 40.030000 10.070000 40.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.750000 40.460000 10.070000 40.780000 ;
      LAYER met4 ;
        RECT 9.750000 40.460000 10.070000 40.780000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.750000 40.890000 10.070000 41.210000 ;
      LAYER met4 ;
        RECT 9.750000 40.890000 10.070000 41.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.750000 41.320000 10.070000 41.640000 ;
      LAYER met4 ;
        RECT 9.750000 41.320000 10.070000 41.640000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.750000 41.750000 10.070000 42.070000 ;
      LAYER met4 ;
        RECT 9.750000 41.750000 10.070000 42.070000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.750000 42.180000 10.070000 42.500000 ;
      LAYER met4 ;
        RECT 9.750000 42.180000 10.070000 42.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.750000 42.610000 10.070000 42.930000 ;
      LAYER met4 ;
        RECT 9.750000 42.610000 10.070000 42.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.750000 43.040000 10.070000 43.360000 ;
      LAYER met4 ;
        RECT 9.750000 43.040000 10.070000 43.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.750000 43.470000 10.070000 43.790000 ;
      LAYER met4 ;
        RECT 9.750000 43.470000 10.070000 43.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.750000 43.900000 10.070000 44.220000 ;
      LAYER met4 ;
        RECT 9.750000 43.900000 10.070000 44.220000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met3 ;
      RECT 0.500000 39.590000 74.700000 44.230000 ;
    LAYER met4 ;
      RECT 0.000000  0.035000 75.000000  45.965000 ;
      RECT 0.000000 49.745000 75.000000  50.725000 ;
      RECT 0.000000 54.505000 75.000000 198.000000 ;
    LAYER met5 ;
      RECT 0.000000  0.135000 72.130000  13.035000 ;
      RECT 0.000000 13.035000 72.435000  17.885000 ;
      RECT 0.000000 17.885000 75.000000  22.335000 ;
      RECT 0.000000 22.335000 72.130000  34.835000 ;
      RECT 0.000000 34.835000 75.000000  44.135000 ;
      RECT 0.000000 44.135000 72.130000  94.585000 ;
      RECT 0.000000 94.585000 75.000000 198.000000 ;
  END
END sky130_fd_io__overlay_vssd_lvc
END LIBRARY
