# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_io__overlay_vccd_lvc
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 198 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 1.270000 54.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 1.270000 49.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.600000 6.890000 24.500000 11.530000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000 6.890000 74.655000 11.530000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 6.885000 24.475000 11.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.780000 6.885000 75.000000 11.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 6.985000 1.270000 11.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.690000  6.960000  0.890000  7.160000 ;
        RECT  0.690000  7.390000  0.890000  7.590000 ;
        RECT  0.690000  7.820000  0.890000  8.020000 ;
        RECT  0.690000  8.250000  0.890000  8.450000 ;
        RECT  0.690000  8.680000  0.890000  8.880000 ;
        RECT  0.690000  9.110000  0.890000  9.310000 ;
        RECT  0.690000  9.540000  0.890000  9.740000 ;
        RECT  0.690000  9.970000  0.890000 10.170000 ;
        RECT  0.690000 10.400000  0.890000 10.600000 ;
        RECT  0.690000 10.830000  0.890000 11.030000 ;
        RECT  0.690000 11.260000  0.890000 11.460000 ;
        RECT  1.100000  6.960000  1.300000  7.160000 ;
        RECT  1.100000  7.390000  1.300000  7.590000 ;
        RECT  1.100000  7.820000  1.300000  8.020000 ;
        RECT  1.100000  8.250000  1.300000  8.450000 ;
        RECT  1.100000  8.680000  1.300000  8.880000 ;
        RECT  1.100000  9.110000  1.300000  9.310000 ;
        RECT  1.100000  9.540000  1.300000  9.740000 ;
        RECT  1.100000  9.970000  1.300000 10.170000 ;
        RECT  1.100000 10.400000  1.300000 10.600000 ;
        RECT  1.100000 10.830000  1.300000 11.030000 ;
        RECT  1.100000 11.260000  1.300000 11.460000 ;
        RECT  1.510000  6.960000  1.710000  7.160000 ;
        RECT  1.510000  7.390000  1.710000  7.590000 ;
        RECT  1.510000  7.820000  1.710000  8.020000 ;
        RECT  1.510000  8.250000  1.710000  8.450000 ;
        RECT  1.510000  8.680000  1.710000  8.880000 ;
        RECT  1.510000  9.110000  1.710000  9.310000 ;
        RECT  1.510000  9.540000  1.710000  9.740000 ;
        RECT  1.510000  9.970000  1.710000 10.170000 ;
        RECT  1.510000 10.400000  1.710000 10.600000 ;
        RECT  1.510000 10.830000  1.710000 11.030000 ;
        RECT  1.510000 11.260000  1.710000 11.460000 ;
        RECT  1.920000  6.960000  2.120000  7.160000 ;
        RECT  1.920000  7.390000  2.120000  7.590000 ;
        RECT  1.920000  7.820000  2.120000  8.020000 ;
        RECT  1.920000  8.250000  2.120000  8.450000 ;
        RECT  1.920000  8.680000  2.120000  8.880000 ;
        RECT  1.920000  9.110000  2.120000  9.310000 ;
        RECT  1.920000  9.540000  2.120000  9.740000 ;
        RECT  1.920000  9.970000  2.120000 10.170000 ;
        RECT  1.920000 10.400000  2.120000 10.600000 ;
        RECT  1.920000 10.830000  2.120000 11.030000 ;
        RECT  1.920000 11.260000  2.120000 11.460000 ;
        RECT  2.330000  6.960000  2.530000  7.160000 ;
        RECT  2.330000  7.390000  2.530000  7.590000 ;
        RECT  2.330000  7.820000  2.530000  8.020000 ;
        RECT  2.330000  8.250000  2.530000  8.450000 ;
        RECT  2.330000  8.680000  2.530000  8.880000 ;
        RECT  2.330000  9.110000  2.530000  9.310000 ;
        RECT  2.330000  9.540000  2.530000  9.740000 ;
        RECT  2.330000  9.970000  2.530000 10.170000 ;
        RECT  2.330000 10.400000  2.530000 10.600000 ;
        RECT  2.330000 10.830000  2.530000 11.030000 ;
        RECT  2.330000 11.260000  2.530000 11.460000 ;
        RECT  2.740000  6.960000  2.940000  7.160000 ;
        RECT  2.740000  7.390000  2.940000  7.590000 ;
        RECT  2.740000  7.820000  2.940000  8.020000 ;
        RECT  2.740000  8.250000  2.940000  8.450000 ;
        RECT  2.740000  8.680000  2.940000  8.880000 ;
        RECT  2.740000  9.110000  2.940000  9.310000 ;
        RECT  2.740000  9.540000  2.940000  9.740000 ;
        RECT  2.740000  9.970000  2.940000 10.170000 ;
        RECT  2.740000 10.400000  2.940000 10.600000 ;
        RECT  2.740000 10.830000  2.940000 11.030000 ;
        RECT  2.740000 11.260000  2.940000 11.460000 ;
        RECT  3.150000  6.960000  3.350000  7.160000 ;
        RECT  3.150000  7.390000  3.350000  7.590000 ;
        RECT  3.150000  7.820000  3.350000  8.020000 ;
        RECT  3.150000  8.250000  3.350000  8.450000 ;
        RECT  3.150000  8.680000  3.350000  8.880000 ;
        RECT  3.150000  9.110000  3.350000  9.310000 ;
        RECT  3.150000  9.540000  3.350000  9.740000 ;
        RECT  3.150000  9.970000  3.350000 10.170000 ;
        RECT  3.150000 10.400000  3.350000 10.600000 ;
        RECT  3.150000 10.830000  3.350000 11.030000 ;
        RECT  3.150000 11.260000  3.350000 11.460000 ;
        RECT  3.555000  6.960000  3.755000  7.160000 ;
        RECT  3.555000  7.390000  3.755000  7.590000 ;
        RECT  3.555000  7.820000  3.755000  8.020000 ;
        RECT  3.555000  8.250000  3.755000  8.450000 ;
        RECT  3.555000  8.680000  3.755000  8.880000 ;
        RECT  3.555000  9.110000  3.755000  9.310000 ;
        RECT  3.555000  9.540000  3.755000  9.740000 ;
        RECT  3.555000  9.970000  3.755000 10.170000 ;
        RECT  3.555000 10.400000  3.755000 10.600000 ;
        RECT  3.555000 10.830000  3.755000 11.030000 ;
        RECT  3.555000 11.260000  3.755000 11.460000 ;
        RECT  3.960000  6.960000  4.160000  7.160000 ;
        RECT  3.960000  7.390000  4.160000  7.590000 ;
        RECT  3.960000  7.820000  4.160000  8.020000 ;
        RECT  3.960000  8.250000  4.160000  8.450000 ;
        RECT  3.960000  8.680000  4.160000  8.880000 ;
        RECT  3.960000  9.110000  4.160000  9.310000 ;
        RECT  3.960000  9.540000  4.160000  9.740000 ;
        RECT  3.960000  9.970000  4.160000 10.170000 ;
        RECT  3.960000 10.400000  4.160000 10.600000 ;
        RECT  3.960000 10.830000  4.160000 11.030000 ;
        RECT  3.960000 11.260000  4.160000 11.460000 ;
        RECT  4.365000  6.960000  4.565000  7.160000 ;
        RECT  4.365000  7.390000  4.565000  7.590000 ;
        RECT  4.365000  7.820000  4.565000  8.020000 ;
        RECT  4.365000  8.250000  4.565000  8.450000 ;
        RECT  4.365000  8.680000  4.565000  8.880000 ;
        RECT  4.365000  9.110000  4.565000  9.310000 ;
        RECT  4.365000  9.540000  4.565000  9.740000 ;
        RECT  4.365000  9.970000  4.565000 10.170000 ;
        RECT  4.365000 10.400000  4.565000 10.600000 ;
        RECT  4.365000 10.830000  4.565000 11.030000 ;
        RECT  4.365000 11.260000  4.565000 11.460000 ;
        RECT  4.770000  6.960000  4.970000  7.160000 ;
        RECT  4.770000  7.390000  4.970000  7.590000 ;
        RECT  4.770000  7.820000  4.970000  8.020000 ;
        RECT  4.770000  8.250000  4.970000  8.450000 ;
        RECT  4.770000  8.680000  4.970000  8.880000 ;
        RECT  4.770000  9.110000  4.970000  9.310000 ;
        RECT  4.770000  9.540000  4.970000  9.740000 ;
        RECT  4.770000  9.970000  4.970000 10.170000 ;
        RECT  4.770000 10.400000  4.970000 10.600000 ;
        RECT  4.770000 10.830000  4.970000 11.030000 ;
        RECT  4.770000 11.260000  4.970000 11.460000 ;
        RECT  5.175000  6.960000  5.375000  7.160000 ;
        RECT  5.175000  7.390000  5.375000  7.590000 ;
        RECT  5.175000  7.820000  5.375000  8.020000 ;
        RECT  5.175000  8.250000  5.375000  8.450000 ;
        RECT  5.175000  8.680000  5.375000  8.880000 ;
        RECT  5.175000  9.110000  5.375000  9.310000 ;
        RECT  5.175000  9.540000  5.375000  9.740000 ;
        RECT  5.175000  9.970000  5.375000 10.170000 ;
        RECT  5.175000 10.400000  5.375000 10.600000 ;
        RECT  5.175000 10.830000  5.375000 11.030000 ;
        RECT  5.175000 11.260000  5.375000 11.460000 ;
        RECT  5.580000  6.960000  5.780000  7.160000 ;
        RECT  5.580000  7.390000  5.780000  7.590000 ;
        RECT  5.580000  7.820000  5.780000  8.020000 ;
        RECT  5.580000  8.250000  5.780000  8.450000 ;
        RECT  5.580000  8.680000  5.780000  8.880000 ;
        RECT  5.580000  9.110000  5.780000  9.310000 ;
        RECT  5.580000  9.540000  5.780000  9.740000 ;
        RECT  5.580000  9.970000  5.780000 10.170000 ;
        RECT  5.580000 10.400000  5.780000 10.600000 ;
        RECT  5.580000 10.830000  5.780000 11.030000 ;
        RECT  5.580000 11.260000  5.780000 11.460000 ;
        RECT  5.985000  6.960000  6.185000  7.160000 ;
        RECT  5.985000  7.390000  6.185000  7.590000 ;
        RECT  5.985000  7.820000  6.185000  8.020000 ;
        RECT  5.985000  8.250000  6.185000  8.450000 ;
        RECT  5.985000  8.680000  6.185000  8.880000 ;
        RECT  5.985000  9.110000  6.185000  9.310000 ;
        RECT  5.985000  9.540000  6.185000  9.740000 ;
        RECT  5.985000  9.970000  6.185000 10.170000 ;
        RECT  5.985000 10.400000  6.185000 10.600000 ;
        RECT  5.985000 10.830000  6.185000 11.030000 ;
        RECT  5.985000 11.260000  6.185000 11.460000 ;
        RECT  6.390000  6.960000  6.590000  7.160000 ;
        RECT  6.390000  7.390000  6.590000  7.590000 ;
        RECT  6.390000  7.820000  6.590000  8.020000 ;
        RECT  6.390000  8.250000  6.590000  8.450000 ;
        RECT  6.390000  8.680000  6.590000  8.880000 ;
        RECT  6.390000  9.110000  6.590000  9.310000 ;
        RECT  6.390000  9.540000  6.590000  9.740000 ;
        RECT  6.390000  9.970000  6.590000 10.170000 ;
        RECT  6.390000 10.400000  6.590000 10.600000 ;
        RECT  6.390000 10.830000  6.590000 11.030000 ;
        RECT  6.390000 11.260000  6.590000 11.460000 ;
        RECT  6.795000  6.960000  6.995000  7.160000 ;
        RECT  6.795000  7.390000  6.995000  7.590000 ;
        RECT  6.795000  7.820000  6.995000  8.020000 ;
        RECT  6.795000  8.250000  6.995000  8.450000 ;
        RECT  6.795000  8.680000  6.995000  8.880000 ;
        RECT  6.795000  9.110000  6.995000  9.310000 ;
        RECT  6.795000  9.540000  6.995000  9.740000 ;
        RECT  6.795000  9.970000  6.995000 10.170000 ;
        RECT  6.795000 10.400000  6.995000 10.600000 ;
        RECT  6.795000 10.830000  6.995000 11.030000 ;
        RECT  6.795000 11.260000  6.995000 11.460000 ;
        RECT  7.200000  6.960000  7.400000  7.160000 ;
        RECT  7.200000  7.390000  7.400000  7.590000 ;
        RECT  7.200000  7.820000  7.400000  8.020000 ;
        RECT  7.200000  8.250000  7.400000  8.450000 ;
        RECT  7.200000  8.680000  7.400000  8.880000 ;
        RECT  7.200000  9.110000  7.400000  9.310000 ;
        RECT  7.200000  9.540000  7.400000  9.740000 ;
        RECT  7.200000  9.970000  7.400000 10.170000 ;
        RECT  7.200000 10.400000  7.400000 10.600000 ;
        RECT  7.200000 10.830000  7.400000 11.030000 ;
        RECT  7.200000 11.260000  7.400000 11.460000 ;
        RECT  7.605000  6.960000  7.805000  7.160000 ;
        RECT  7.605000  7.390000  7.805000  7.590000 ;
        RECT  7.605000  7.820000  7.805000  8.020000 ;
        RECT  7.605000  8.250000  7.805000  8.450000 ;
        RECT  7.605000  8.680000  7.805000  8.880000 ;
        RECT  7.605000  9.110000  7.805000  9.310000 ;
        RECT  7.605000  9.540000  7.805000  9.740000 ;
        RECT  7.605000  9.970000  7.805000 10.170000 ;
        RECT  7.605000 10.400000  7.805000 10.600000 ;
        RECT  7.605000 10.830000  7.805000 11.030000 ;
        RECT  7.605000 11.260000  7.805000 11.460000 ;
        RECT  8.010000  6.960000  8.210000  7.160000 ;
        RECT  8.010000  7.390000  8.210000  7.590000 ;
        RECT  8.010000  7.820000  8.210000  8.020000 ;
        RECT  8.010000  8.250000  8.210000  8.450000 ;
        RECT  8.010000  8.680000  8.210000  8.880000 ;
        RECT  8.010000  9.110000  8.210000  9.310000 ;
        RECT  8.010000  9.540000  8.210000  9.740000 ;
        RECT  8.010000  9.970000  8.210000 10.170000 ;
        RECT  8.010000 10.400000  8.210000 10.600000 ;
        RECT  8.010000 10.830000  8.210000 11.030000 ;
        RECT  8.010000 11.260000  8.210000 11.460000 ;
        RECT  8.415000  6.960000  8.615000  7.160000 ;
        RECT  8.415000  7.390000  8.615000  7.590000 ;
        RECT  8.415000  7.820000  8.615000  8.020000 ;
        RECT  8.415000  8.250000  8.615000  8.450000 ;
        RECT  8.415000  8.680000  8.615000  8.880000 ;
        RECT  8.415000  9.110000  8.615000  9.310000 ;
        RECT  8.415000  9.540000  8.615000  9.740000 ;
        RECT  8.415000  9.970000  8.615000 10.170000 ;
        RECT  8.415000 10.400000  8.615000 10.600000 ;
        RECT  8.415000 10.830000  8.615000 11.030000 ;
        RECT  8.415000 11.260000  8.615000 11.460000 ;
        RECT  8.820000  6.960000  9.020000  7.160000 ;
        RECT  8.820000  7.390000  9.020000  7.590000 ;
        RECT  8.820000  7.820000  9.020000  8.020000 ;
        RECT  8.820000  8.250000  9.020000  8.450000 ;
        RECT  8.820000  8.680000  9.020000  8.880000 ;
        RECT  8.820000  9.110000  9.020000  9.310000 ;
        RECT  8.820000  9.540000  9.020000  9.740000 ;
        RECT  8.820000  9.970000  9.020000 10.170000 ;
        RECT  8.820000 10.400000  9.020000 10.600000 ;
        RECT  8.820000 10.830000  9.020000 11.030000 ;
        RECT  8.820000 11.260000  9.020000 11.460000 ;
        RECT  9.225000  6.960000  9.425000  7.160000 ;
        RECT  9.225000  7.390000  9.425000  7.590000 ;
        RECT  9.225000  7.820000  9.425000  8.020000 ;
        RECT  9.225000  8.250000  9.425000  8.450000 ;
        RECT  9.225000  8.680000  9.425000  8.880000 ;
        RECT  9.225000  9.110000  9.425000  9.310000 ;
        RECT  9.225000  9.540000  9.425000  9.740000 ;
        RECT  9.225000  9.970000  9.425000 10.170000 ;
        RECT  9.225000 10.400000  9.425000 10.600000 ;
        RECT  9.225000 10.830000  9.425000 11.030000 ;
        RECT  9.225000 11.260000  9.425000 11.460000 ;
        RECT  9.630000  6.960000  9.830000  7.160000 ;
        RECT  9.630000  7.390000  9.830000  7.590000 ;
        RECT  9.630000  7.820000  9.830000  8.020000 ;
        RECT  9.630000  8.250000  9.830000  8.450000 ;
        RECT  9.630000  8.680000  9.830000  8.880000 ;
        RECT  9.630000  9.110000  9.830000  9.310000 ;
        RECT  9.630000  9.540000  9.830000  9.740000 ;
        RECT  9.630000  9.970000  9.830000 10.170000 ;
        RECT  9.630000 10.400000  9.830000 10.600000 ;
        RECT  9.630000 10.830000  9.830000 11.030000 ;
        RECT  9.630000 11.260000  9.830000 11.460000 ;
        RECT 10.035000  6.960000 10.235000  7.160000 ;
        RECT 10.035000  7.390000 10.235000  7.590000 ;
        RECT 10.035000  7.820000 10.235000  8.020000 ;
        RECT 10.035000  8.250000 10.235000  8.450000 ;
        RECT 10.035000  8.680000 10.235000  8.880000 ;
        RECT 10.035000  9.110000 10.235000  9.310000 ;
        RECT 10.035000  9.540000 10.235000  9.740000 ;
        RECT 10.035000  9.970000 10.235000 10.170000 ;
        RECT 10.035000 10.400000 10.235000 10.600000 ;
        RECT 10.035000 10.830000 10.235000 11.030000 ;
        RECT 10.035000 11.260000 10.235000 11.460000 ;
        RECT 10.440000  6.960000 10.640000  7.160000 ;
        RECT 10.440000  7.390000 10.640000  7.590000 ;
        RECT 10.440000  7.820000 10.640000  8.020000 ;
        RECT 10.440000  8.250000 10.640000  8.450000 ;
        RECT 10.440000  8.680000 10.640000  8.880000 ;
        RECT 10.440000  9.110000 10.640000  9.310000 ;
        RECT 10.440000  9.540000 10.640000  9.740000 ;
        RECT 10.440000  9.970000 10.640000 10.170000 ;
        RECT 10.440000 10.400000 10.640000 10.600000 ;
        RECT 10.440000 10.830000 10.640000 11.030000 ;
        RECT 10.440000 11.260000 10.640000 11.460000 ;
        RECT 10.845000  6.960000 11.045000  7.160000 ;
        RECT 10.845000  7.390000 11.045000  7.590000 ;
        RECT 10.845000  7.820000 11.045000  8.020000 ;
        RECT 10.845000  8.250000 11.045000  8.450000 ;
        RECT 10.845000  8.680000 11.045000  8.880000 ;
        RECT 10.845000  9.110000 11.045000  9.310000 ;
        RECT 10.845000  9.540000 11.045000  9.740000 ;
        RECT 10.845000  9.970000 11.045000 10.170000 ;
        RECT 10.845000 10.400000 11.045000 10.600000 ;
        RECT 10.845000 10.830000 11.045000 11.030000 ;
        RECT 10.845000 11.260000 11.045000 11.460000 ;
        RECT 11.250000  6.960000 11.450000  7.160000 ;
        RECT 11.250000  7.390000 11.450000  7.590000 ;
        RECT 11.250000  7.820000 11.450000  8.020000 ;
        RECT 11.250000  8.250000 11.450000  8.450000 ;
        RECT 11.250000  8.680000 11.450000  8.880000 ;
        RECT 11.250000  9.110000 11.450000  9.310000 ;
        RECT 11.250000  9.540000 11.450000  9.740000 ;
        RECT 11.250000  9.970000 11.450000 10.170000 ;
        RECT 11.250000 10.400000 11.450000 10.600000 ;
        RECT 11.250000 10.830000 11.450000 11.030000 ;
        RECT 11.250000 11.260000 11.450000 11.460000 ;
        RECT 11.655000  6.960000 11.855000  7.160000 ;
        RECT 11.655000  7.390000 11.855000  7.590000 ;
        RECT 11.655000  7.820000 11.855000  8.020000 ;
        RECT 11.655000  8.250000 11.855000  8.450000 ;
        RECT 11.655000  8.680000 11.855000  8.880000 ;
        RECT 11.655000  9.110000 11.855000  9.310000 ;
        RECT 11.655000  9.540000 11.855000  9.740000 ;
        RECT 11.655000  9.970000 11.855000 10.170000 ;
        RECT 11.655000 10.400000 11.855000 10.600000 ;
        RECT 11.655000 10.830000 11.855000 11.030000 ;
        RECT 11.655000 11.260000 11.855000 11.460000 ;
        RECT 12.060000  6.960000 12.260000  7.160000 ;
        RECT 12.060000  7.390000 12.260000  7.590000 ;
        RECT 12.060000  7.820000 12.260000  8.020000 ;
        RECT 12.060000  8.250000 12.260000  8.450000 ;
        RECT 12.060000  8.680000 12.260000  8.880000 ;
        RECT 12.060000  9.110000 12.260000  9.310000 ;
        RECT 12.060000  9.540000 12.260000  9.740000 ;
        RECT 12.060000  9.970000 12.260000 10.170000 ;
        RECT 12.060000 10.400000 12.260000 10.600000 ;
        RECT 12.060000 10.830000 12.260000 11.030000 ;
        RECT 12.060000 11.260000 12.260000 11.460000 ;
        RECT 12.465000  6.960000 12.665000  7.160000 ;
        RECT 12.465000  7.390000 12.665000  7.590000 ;
        RECT 12.465000  7.820000 12.665000  8.020000 ;
        RECT 12.465000  8.250000 12.665000  8.450000 ;
        RECT 12.465000  8.680000 12.665000  8.880000 ;
        RECT 12.465000  9.110000 12.665000  9.310000 ;
        RECT 12.465000  9.540000 12.665000  9.740000 ;
        RECT 12.465000  9.970000 12.665000 10.170000 ;
        RECT 12.465000 10.400000 12.665000 10.600000 ;
        RECT 12.465000 10.830000 12.665000 11.030000 ;
        RECT 12.465000 11.260000 12.665000 11.460000 ;
        RECT 12.870000  6.960000 13.070000  7.160000 ;
        RECT 12.870000  7.390000 13.070000  7.590000 ;
        RECT 12.870000  7.820000 13.070000  8.020000 ;
        RECT 12.870000  8.250000 13.070000  8.450000 ;
        RECT 12.870000  8.680000 13.070000  8.880000 ;
        RECT 12.870000  9.110000 13.070000  9.310000 ;
        RECT 12.870000  9.540000 13.070000  9.740000 ;
        RECT 12.870000  9.970000 13.070000 10.170000 ;
        RECT 12.870000 10.400000 13.070000 10.600000 ;
        RECT 12.870000 10.830000 13.070000 11.030000 ;
        RECT 12.870000 11.260000 13.070000 11.460000 ;
        RECT 13.275000  6.960000 13.475000  7.160000 ;
        RECT 13.275000  7.390000 13.475000  7.590000 ;
        RECT 13.275000  7.820000 13.475000  8.020000 ;
        RECT 13.275000  8.250000 13.475000  8.450000 ;
        RECT 13.275000  8.680000 13.475000  8.880000 ;
        RECT 13.275000  9.110000 13.475000  9.310000 ;
        RECT 13.275000  9.540000 13.475000  9.740000 ;
        RECT 13.275000  9.970000 13.475000 10.170000 ;
        RECT 13.275000 10.400000 13.475000 10.600000 ;
        RECT 13.275000 10.830000 13.475000 11.030000 ;
        RECT 13.275000 11.260000 13.475000 11.460000 ;
        RECT 13.680000  6.960000 13.880000  7.160000 ;
        RECT 13.680000  7.390000 13.880000  7.590000 ;
        RECT 13.680000  7.820000 13.880000  8.020000 ;
        RECT 13.680000  8.250000 13.880000  8.450000 ;
        RECT 13.680000  8.680000 13.880000  8.880000 ;
        RECT 13.680000  9.110000 13.880000  9.310000 ;
        RECT 13.680000  9.540000 13.880000  9.740000 ;
        RECT 13.680000  9.970000 13.880000 10.170000 ;
        RECT 13.680000 10.400000 13.880000 10.600000 ;
        RECT 13.680000 10.830000 13.880000 11.030000 ;
        RECT 13.680000 11.260000 13.880000 11.460000 ;
        RECT 14.085000  6.960000 14.285000  7.160000 ;
        RECT 14.085000  7.390000 14.285000  7.590000 ;
        RECT 14.085000  7.820000 14.285000  8.020000 ;
        RECT 14.085000  8.250000 14.285000  8.450000 ;
        RECT 14.085000  8.680000 14.285000  8.880000 ;
        RECT 14.085000  9.110000 14.285000  9.310000 ;
        RECT 14.085000  9.540000 14.285000  9.740000 ;
        RECT 14.085000  9.970000 14.285000 10.170000 ;
        RECT 14.085000 10.400000 14.285000 10.600000 ;
        RECT 14.085000 10.830000 14.285000 11.030000 ;
        RECT 14.085000 11.260000 14.285000 11.460000 ;
        RECT 14.490000  6.960000 14.690000  7.160000 ;
        RECT 14.490000  7.390000 14.690000  7.590000 ;
        RECT 14.490000  7.820000 14.690000  8.020000 ;
        RECT 14.490000  8.250000 14.690000  8.450000 ;
        RECT 14.490000  8.680000 14.690000  8.880000 ;
        RECT 14.490000  9.110000 14.690000  9.310000 ;
        RECT 14.490000  9.540000 14.690000  9.740000 ;
        RECT 14.490000  9.970000 14.690000 10.170000 ;
        RECT 14.490000 10.400000 14.690000 10.600000 ;
        RECT 14.490000 10.830000 14.690000 11.030000 ;
        RECT 14.490000 11.260000 14.690000 11.460000 ;
        RECT 14.895000  6.960000 15.095000  7.160000 ;
        RECT 14.895000  7.390000 15.095000  7.590000 ;
        RECT 14.895000  7.820000 15.095000  8.020000 ;
        RECT 14.895000  8.250000 15.095000  8.450000 ;
        RECT 14.895000  8.680000 15.095000  8.880000 ;
        RECT 14.895000  9.110000 15.095000  9.310000 ;
        RECT 14.895000  9.540000 15.095000  9.740000 ;
        RECT 14.895000  9.970000 15.095000 10.170000 ;
        RECT 14.895000 10.400000 15.095000 10.600000 ;
        RECT 14.895000 10.830000 15.095000 11.030000 ;
        RECT 14.895000 11.260000 15.095000 11.460000 ;
        RECT 15.300000  6.960000 15.500000  7.160000 ;
        RECT 15.300000  7.390000 15.500000  7.590000 ;
        RECT 15.300000  7.820000 15.500000  8.020000 ;
        RECT 15.300000  8.250000 15.500000  8.450000 ;
        RECT 15.300000  8.680000 15.500000  8.880000 ;
        RECT 15.300000  9.110000 15.500000  9.310000 ;
        RECT 15.300000  9.540000 15.500000  9.740000 ;
        RECT 15.300000  9.970000 15.500000 10.170000 ;
        RECT 15.300000 10.400000 15.500000 10.600000 ;
        RECT 15.300000 10.830000 15.500000 11.030000 ;
        RECT 15.300000 11.260000 15.500000 11.460000 ;
        RECT 15.705000  6.960000 15.905000  7.160000 ;
        RECT 15.705000  7.390000 15.905000  7.590000 ;
        RECT 15.705000  7.820000 15.905000  8.020000 ;
        RECT 15.705000  8.250000 15.905000  8.450000 ;
        RECT 15.705000  8.680000 15.905000  8.880000 ;
        RECT 15.705000  9.110000 15.905000  9.310000 ;
        RECT 15.705000  9.540000 15.905000  9.740000 ;
        RECT 15.705000  9.970000 15.905000 10.170000 ;
        RECT 15.705000 10.400000 15.905000 10.600000 ;
        RECT 15.705000 10.830000 15.905000 11.030000 ;
        RECT 15.705000 11.260000 15.905000 11.460000 ;
        RECT 16.110000  6.960000 16.310000  7.160000 ;
        RECT 16.110000  7.390000 16.310000  7.590000 ;
        RECT 16.110000  7.820000 16.310000  8.020000 ;
        RECT 16.110000  8.250000 16.310000  8.450000 ;
        RECT 16.110000  8.680000 16.310000  8.880000 ;
        RECT 16.110000  9.110000 16.310000  9.310000 ;
        RECT 16.110000  9.540000 16.310000  9.740000 ;
        RECT 16.110000  9.970000 16.310000 10.170000 ;
        RECT 16.110000 10.400000 16.310000 10.600000 ;
        RECT 16.110000 10.830000 16.310000 11.030000 ;
        RECT 16.110000 11.260000 16.310000 11.460000 ;
        RECT 16.515000  6.960000 16.715000  7.160000 ;
        RECT 16.515000  7.390000 16.715000  7.590000 ;
        RECT 16.515000  7.820000 16.715000  8.020000 ;
        RECT 16.515000  8.250000 16.715000  8.450000 ;
        RECT 16.515000  8.680000 16.715000  8.880000 ;
        RECT 16.515000  9.110000 16.715000  9.310000 ;
        RECT 16.515000  9.540000 16.715000  9.740000 ;
        RECT 16.515000  9.970000 16.715000 10.170000 ;
        RECT 16.515000 10.400000 16.715000 10.600000 ;
        RECT 16.515000 10.830000 16.715000 11.030000 ;
        RECT 16.515000 11.260000 16.715000 11.460000 ;
        RECT 16.920000  6.960000 17.120000  7.160000 ;
        RECT 16.920000  7.390000 17.120000  7.590000 ;
        RECT 16.920000  7.820000 17.120000  8.020000 ;
        RECT 16.920000  8.250000 17.120000  8.450000 ;
        RECT 16.920000  8.680000 17.120000  8.880000 ;
        RECT 16.920000  9.110000 17.120000  9.310000 ;
        RECT 16.920000  9.540000 17.120000  9.740000 ;
        RECT 16.920000  9.970000 17.120000 10.170000 ;
        RECT 16.920000 10.400000 17.120000 10.600000 ;
        RECT 16.920000 10.830000 17.120000 11.030000 ;
        RECT 16.920000 11.260000 17.120000 11.460000 ;
        RECT 17.325000  6.960000 17.525000  7.160000 ;
        RECT 17.325000  7.390000 17.525000  7.590000 ;
        RECT 17.325000  7.820000 17.525000  8.020000 ;
        RECT 17.325000  8.250000 17.525000  8.450000 ;
        RECT 17.325000  8.680000 17.525000  8.880000 ;
        RECT 17.325000  9.110000 17.525000  9.310000 ;
        RECT 17.325000  9.540000 17.525000  9.740000 ;
        RECT 17.325000  9.970000 17.525000 10.170000 ;
        RECT 17.325000 10.400000 17.525000 10.600000 ;
        RECT 17.325000 10.830000 17.525000 11.030000 ;
        RECT 17.325000 11.260000 17.525000 11.460000 ;
        RECT 17.730000  6.960000 17.930000  7.160000 ;
        RECT 17.730000  7.390000 17.930000  7.590000 ;
        RECT 17.730000  7.820000 17.930000  8.020000 ;
        RECT 17.730000  8.250000 17.930000  8.450000 ;
        RECT 17.730000  8.680000 17.930000  8.880000 ;
        RECT 17.730000  9.110000 17.930000  9.310000 ;
        RECT 17.730000  9.540000 17.930000  9.740000 ;
        RECT 17.730000  9.970000 17.930000 10.170000 ;
        RECT 17.730000 10.400000 17.930000 10.600000 ;
        RECT 17.730000 10.830000 17.930000 11.030000 ;
        RECT 17.730000 11.260000 17.930000 11.460000 ;
        RECT 18.135000  6.960000 18.335000  7.160000 ;
        RECT 18.135000  7.390000 18.335000  7.590000 ;
        RECT 18.135000  7.820000 18.335000  8.020000 ;
        RECT 18.135000  8.250000 18.335000  8.450000 ;
        RECT 18.135000  8.680000 18.335000  8.880000 ;
        RECT 18.135000  9.110000 18.335000  9.310000 ;
        RECT 18.135000  9.540000 18.335000  9.740000 ;
        RECT 18.135000  9.970000 18.335000 10.170000 ;
        RECT 18.135000 10.400000 18.335000 10.600000 ;
        RECT 18.135000 10.830000 18.335000 11.030000 ;
        RECT 18.135000 11.260000 18.335000 11.460000 ;
        RECT 18.540000  6.960000 18.740000  7.160000 ;
        RECT 18.540000  7.390000 18.740000  7.590000 ;
        RECT 18.540000  7.820000 18.740000  8.020000 ;
        RECT 18.540000  8.250000 18.740000  8.450000 ;
        RECT 18.540000  8.680000 18.740000  8.880000 ;
        RECT 18.540000  9.110000 18.740000  9.310000 ;
        RECT 18.540000  9.540000 18.740000  9.740000 ;
        RECT 18.540000  9.970000 18.740000 10.170000 ;
        RECT 18.540000 10.400000 18.740000 10.600000 ;
        RECT 18.540000 10.830000 18.740000 11.030000 ;
        RECT 18.540000 11.260000 18.740000 11.460000 ;
        RECT 18.945000  6.960000 19.145000  7.160000 ;
        RECT 18.945000  7.390000 19.145000  7.590000 ;
        RECT 18.945000  7.820000 19.145000  8.020000 ;
        RECT 18.945000  8.250000 19.145000  8.450000 ;
        RECT 18.945000  8.680000 19.145000  8.880000 ;
        RECT 18.945000  9.110000 19.145000  9.310000 ;
        RECT 18.945000  9.540000 19.145000  9.740000 ;
        RECT 18.945000  9.970000 19.145000 10.170000 ;
        RECT 18.945000 10.400000 19.145000 10.600000 ;
        RECT 18.945000 10.830000 19.145000 11.030000 ;
        RECT 18.945000 11.260000 19.145000 11.460000 ;
        RECT 19.350000  6.960000 19.550000  7.160000 ;
        RECT 19.350000  7.390000 19.550000  7.590000 ;
        RECT 19.350000  7.820000 19.550000  8.020000 ;
        RECT 19.350000  8.250000 19.550000  8.450000 ;
        RECT 19.350000  8.680000 19.550000  8.880000 ;
        RECT 19.350000  9.110000 19.550000  9.310000 ;
        RECT 19.350000  9.540000 19.550000  9.740000 ;
        RECT 19.350000  9.970000 19.550000 10.170000 ;
        RECT 19.350000 10.400000 19.550000 10.600000 ;
        RECT 19.350000 10.830000 19.550000 11.030000 ;
        RECT 19.350000 11.260000 19.550000 11.460000 ;
        RECT 19.755000  6.960000 19.955000  7.160000 ;
        RECT 19.755000  7.390000 19.955000  7.590000 ;
        RECT 19.755000  7.820000 19.955000  8.020000 ;
        RECT 19.755000  8.250000 19.955000  8.450000 ;
        RECT 19.755000  8.680000 19.955000  8.880000 ;
        RECT 19.755000  9.110000 19.955000  9.310000 ;
        RECT 19.755000  9.540000 19.955000  9.740000 ;
        RECT 19.755000  9.970000 19.955000 10.170000 ;
        RECT 19.755000 10.400000 19.955000 10.600000 ;
        RECT 19.755000 10.830000 19.955000 11.030000 ;
        RECT 19.755000 11.260000 19.955000 11.460000 ;
        RECT 20.160000  6.960000 20.360000  7.160000 ;
        RECT 20.160000  7.390000 20.360000  7.590000 ;
        RECT 20.160000  7.820000 20.360000  8.020000 ;
        RECT 20.160000  8.250000 20.360000  8.450000 ;
        RECT 20.160000  8.680000 20.360000  8.880000 ;
        RECT 20.160000  9.110000 20.360000  9.310000 ;
        RECT 20.160000  9.540000 20.360000  9.740000 ;
        RECT 20.160000  9.970000 20.360000 10.170000 ;
        RECT 20.160000 10.400000 20.360000 10.600000 ;
        RECT 20.160000 10.830000 20.360000 11.030000 ;
        RECT 20.160000 11.260000 20.360000 11.460000 ;
        RECT 20.565000  6.960000 20.765000  7.160000 ;
        RECT 20.565000  7.390000 20.765000  7.590000 ;
        RECT 20.565000  7.820000 20.765000  8.020000 ;
        RECT 20.565000  8.250000 20.765000  8.450000 ;
        RECT 20.565000  8.680000 20.765000  8.880000 ;
        RECT 20.565000  9.110000 20.765000  9.310000 ;
        RECT 20.565000  9.540000 20.765000  9.740000 ;
        RECT 20.565000  9.970000 20.765000 10.170000 ;
        RECT 20.565000 10.400000 20.765000 10.600000 ;
        RECT 20.565000 10.830000 20.765000 11.030000 ;
        RECT 20.565000 11.260000 20.765000 11.460000 ;
        RECT 20.970000  6.960000 21.170000  7.160000 ;
        RECT 20.970000  7.390000 21.170000  7.590000 ;
        RECT 20.970000  7.820000 21.170000  8.020000 ;
        RECT 20.970000  8.250000 21.170000  8.450000 ;
        RECT 20.970000  8.680000 21.170000  8.880000 ;
        RECT 20.970000  9.110000 21.170000  9.310000 ;
        RECT 20.970000  9.540000 21.170000  9.740000 ;
        RECT 20.970000  9.970000 21.170000 10.170000 ;
        RECT 20.970000 10.400000 21.170000 10.600000 ;
        RECT 20.970000 10.830000 21.170000 11.030000 ;
        RECT 20.970000 11.260000 21.170000 11.460000 ;
        RECT 21.375000  6.960000 21.575000  7.160000 ;
        RECT 21.375000  7.390000 21.575000  7.590000 ;
        RECT 21.375000  7.820000 21.575000  8.020000 ;
        RECT 21.375000  8.250000 21.575000  8.450000 ;
        RECT 21.375000  8.680000 21.575000  8.880000 ;
        RECT 21.375000  9.110000 21.575000  9.310000 ;
        RECT 21.375000  9.540000 21.575000  9.740000 ;
        RECT 21.375000  9.970000 21.575000 10.170000 ;
        RECT 21.375000 10.400000 21.575000 10.600000 ;
        RECT 21.375000 10.830000 21.575000 11.030000 ;
        RECT 21.375000 11.260000 21.575000 11.460000 ;
        RECT 21.780000  6.960000 21.980000  7.160000 ;
        RECT 21.780000  7.390000 21.980000  7.590000 ;
        RECT 21.780000  7.820000 21.980000  8.020000 ;
        RECT 21.780000  8.250000 21.980000  8.450000 ;
        RECT 21.780000  8.680000 21.980000  8.880000 ;
        RECT 21.780000  9.110000 21.980000  9.310000 ;
        RECT 21.780000  9.540000 21.980000  9.740000 ;
        RECT 21.780000  9.970000 21.980000 10.170000 ;
        RECT 21.780000 10.400000 21.980000 10.600000 ;
        RECT 21.780000 10.830000 21.980000 11.030000 ;
        RECT 21.780000 11.260000 21.980000 11.460000 ;
        RECT 22.185000  6.960000 22.385000  7.160000 ;
        RECT 22.185000  7.390000 22.385000  7.590000 ;
        RECT 22.185000  7.820000 22.385000  8.020000 ;
        RECT 22.185000  8.250000 22.385000  8.450000 ;
        RECT 22.185000  8.680000 22.385000  8.880000 ;
        RECT 22.185000  9.110000 22.385000  9.310000 ;
        RECT 22.185000  9.540000 22.385000  9.740000 ;
        RECT 22.185000  9.970000 22.385000 10.170000 ;
        RECT 22.185000 10.400000 22.385000 10.600000 ;
        RECT 22.185000 10.830000 22.385000 11.030000 ;
        RECT 22.185000 11.260000 22.385000 11.460000 ;
        RECT 22.590000  6.960000 22.790000  7.160000 ;
        RECT 22.590000  7.390000 22.790000  7.590000 ;
        RECT 22.590000  7.820000 22.790000  8.020000 ;
        RECT 22.590000  8.250000 22.790000  8.450000 ;
        RECT 22.590000  8.680000 22.790000  8.880000 ;
        RECT 22.590000  9.110000 22.790000  9.310000 ;
        RECT 22.590000  9.540000 22.790000  9.740000 ;
        RECT 22.590000  9.970000 22.790000 10.170000 ;
        RECT 22.590000 10.400000 22.790000 10.600000 ;
        RECT 22.590000 10.830000 22.790000 11.030000 ;
        RECT 22.590000 11.260000 22.790000 11.460000 ;
        RECT 22.995000  6.960000 23.195000  7.160000 ;
        RECT 22.995000  7.390000 23.195000  7.590000 ;
        RECT 22.995000  7.820000 23.195000  8.020000 ;
        RECT 22.995000  8.250000 23.195000  8.450000 ;
        RECT 22.995000  8.680000 23.195000  8.880000 ;
        RECT 22.995000  9.110000 23.195000  9.310000 ;
        RECT 22.995000  9.540000 23.195000  9.740000 ;
        RECT 22.995000  9.970000 23.195000 10.170000 ;
        RECT 22.995000 10.400000 23.195000 10.600000 ;
        RECT 22.995000 10.830000 23.195000 11.030000 ;
        RECT 22.995000 11.260000 23.195000 11.460000 ;
        RECT 23.400000  6.960000 23.600000  7.160000 ;
        RECT 23.400000  7.390000 23.600000  7.590000 ;
        RECT 23.400000  7.820000 23.600000  8.020000 ;
        RECT 23.400000  8.250000 23.600000  8.450000 ;
        RECT 23.400000  8.680000 23.600000  8.880000 ;
        RECT 23.400000  9.110000 23.600000  9.310000 ;
        RECT 23.400000  9.540000 23.600000  9.740000 ;
        RECT 23.400000  9.970000 23.600000 10.170000 ;
        RECT 23.400000 10.400000 23.600000 10.600000 ;
        RECT 23.400000 10.830000 23.600000 11.030000 ;
        RECT 23.400000 11.260000 23.600000 11.460000 ;
        RECT 23.805000  6.960000 24.005000  7.160000 ;
        RECT 23.805000  7.390000 24.005000  7.590000 ;
        RECT 23.805000  7.820000 24.005000  8.020000 ;
        RECT 23.805000  8.250000 24.005000  8.450000 ;
        RECT 23.805000  8.680000 24.005000  8.880000 ;
        RECT 23.805000  9.110000 24.005000  9.310000 ;
        RECT 23.805000  9.540000 24.005000  9.740000 ;
        RECT 23.805000  9.970000 24.005000 10.170000 ;
        RECT 23.805000 10.400000 24.005000 10.600000 ;
        RECT 23.805000 10.830000 24.005000 11.030000 ;
        RECT 23.805000 11.260000 24.005000 11.460000 ;
        RECT 24.210000  6.960000 24.410000  7.160000 ;
        RECT 24.210000  7.390000 24.410000  7.590000 ;
        RECT 24.210000  7.820000 24.410000  8.020000 ;
        RECT 24.210000  8.250000 24.410000  8.450000 ;
        RECT 24.210000  8.680000 24.410000  8.880000 ;
        RECT 24.210000  9.110000 24.410000  9.310000 ;
        RECT 24.210000  9.540000 24.410000  9.740000 ;
        RECT 24.210000  9.970000 24.410000 10.170000 ;
        RECT 24.210000 10.400000 24.410000 10.600000 ;
        RECT 24.210000 10.830000 24.410000 11.030000 ;
        RECT 24.210000 11.260000 24.410000 11.460000 ;
        RECT 50.845000  6.960000 51.045000  7.160000 ;
        RECT 50.845000  7.390000 51.045000  7.590000 ;
        RECT 50.845000  7.820000 51.045000  8.020000 ;
        RECT 50.845000  8.250000 51.045000  8.450000 ;
        RECT 50.845000  8.680000 51.045000  8.880000 ;
        RECT 50.845000  9.110000 51.045000  9.310000 ;
        RECT 50.845000  9.540000 51.045000  9.740000 ;
        RECT 50.845000  9.970000 51.045000 10.170000 ;
        RECT 50.845000 10.400000 51.045000 10.600000 ;
        RECT 50.845000 10.830000 51.045000 11.030000 ;
        RECT 50.845000 11.260000 51.045000 11.460000 ;
        RECT 51.255000  6.960000 51.455000  7.160000 ;
        RECT 51.255000  7.390000 51.455000  7.590000 ;
        RECT 51.255000  7.820000 51.455000  8.020000 ;
        RECT 51.255000  8.250000 51.455000  8.450000 ;
        RECT 51.255000  8.680000 51.455000  8.880000 ;
        RECT 51.255000  9.110000 51.455000  9.310000 ;
        RECT 51.255000  9.540000 51.455000  9.740000 ;
        RECT 51.255000  9.970000 51.455000 10.170000 ;
        RECT 51.255000 10.400000 51.455000 10.600000 ;
        RECT 51.255000 10.830000 51.455000 11.030000 ;
        RECT 51.255000 11.260000 51.455000 11.460000 ;
        RECT 51.665000  6.960000 51.865000  7.160000 ;
        RECT 51.665000  7.390000 51.865000  7.590000 ;
        RECT 51.665000  7.820000 51.865000  8.020000 ;
        RECT 51.665000  8.250000 51.865000  8.450000 ;
        RECT 51.665000  8.680000 51.865000  8.880000 ;
        RECT 51.665000  9.110000 51.865000  9.310000 ;
        RECT 51.665000  9.540000 51.865000  9.740000 ;
        RECT 51.665000  9.970000 51.865000 10.170000 ;
        RECT 51.665000 10.400000 51.865000 10.600000 ;
        RECT 51.665000 10.830000 51.865000 11.030000 ;
        RECT 51.665000 11.260000 51.865000 11.460000 ;
        RECT 52.075000  6.960000 52.275000  7.160000 ;
        RECT 52.075000  7.390000 52.275000  7.590000 ;
        RECT 52.075000  7.820000 52.275000  8.020000 ;
        RECT 52.075000  8.250000 52.275000  8.450000 ;
        RECT 52.075000  8.680000 52.275000  8.880000 ;
        RECT 52.075000  9.110000 52.275000  9.310000 ;
        RECT 52.075000  9.540000 52.275000  9.740000 ;
        RECT 52.075000  9.970000 52.275000 10.170000 ;
        RECT 52.075000 10.400000 52.275000 10.600000 ;
        RECT 52.075000 10.830000 52.275000 11.030000 ;
        RECT 52.075000 11.260000 52.275000 11.460000 ;
        RECT 52.485000  6.960000 52.685000  7.160000 ;
        RECT 52.485000  7.390000 52.685000  7.590000 ;
        RECT 52.485000  7.820000 52.685000  8.020000 ;
        RECT 52.485000  8.250000 52.685000  8.450000 ;
        RECT 52.485000  8.680000 52.685000  8.880000 ;
        RECT 52.485000  9.110000 52.685000  9.310000 ;
        RECT 52.485000  9.540000 52.685000  9.740000 ;
        RECT 52.485000  9.970000 52.685000 10.170000 ;
        RECT 52.485000 10.400000 52.685000 10.600000 ;
        RECT 52.485000 10.830000 52.685000 11.030000 ;
        RECT 52.485000 11.260000 52.685000 11.460000 ;
        RECT 52.895000  6.960000 53.095000  7.160000 ;
        RECT 52.895000  7.390000 53.095000  7.590000 ;
        RECT 52.895000  7.820000 53.095000  8.020000 ;
        RECT 52.895000  8.250000 53.095000  8.450000 ;
        RECT 52.895000  8.680000 53.095000  8.880000 ;
        RECT 52.895000  9.110000 53.095000  9.310000 ;
        RECT 52.895000  9.540000 53.095000  9.740000 ;
        RECT 52.895000  9.970000 53.095000 10.170000 ;
        RECT 52.895000 10.400000 53.095000 10.600000 ;
        RECT 52.895000 10.830000 53.095000 11.030000 ;
        RECT 52.895000 11.260000 53.095000 11.460000 ;
        RECT 53.305000  6.960000 53.505000  7.160000 ;
        RECT 53.305000  7.390000 53.505000  7.590000 ;
        RECT 53.305000  7.820000 53.505000  8.020000 ;
        RECT 53.305000  8.250000 53.505000  8.450000 ;
        RECT 53.305000  8.680000 53.505000  8.880000 ;
        RECT 53.305000  9.110000 53.505000  9.310000 ;
        RECT 53.305000  9.540000 53.505000  9.740000 ;
        RECT 53.305000  9.970000 53.505000 10.170000 ;
        RECT 53.305000 10.400000 53.505000 10.600000 ;
        RECT 53.305000 10.830000 53.505000 11.030000 ;
        RECT 53.305000 11.260000 53.505000 11.460000 ;
        RECT 53.710000  6.960000 53.910000  7.160000 ;
        RECT 53.710000  7.390000 53.910000  7.590000 ;
        RECT 53.710000  7.820000 53.910000  8.020000 ;
        RECT 53.710000  8.250000 53.910000  8.450000 ;
        RECT 53.710000  8.680000 53.910000  8.880000 ;
        RECT 53.710000  9.110000 53.910000  9.310000 ;
        RECT 53.710000  9.540000 53.910000  9.740000 ;
        RECT 53.710000  9.970000 53.910000 10.170000 ;
        RECT 53.710000 10.400000 53.910000 10.600000 ;
        RECT 53.710000 10.830000 53.910000 11.030000 ;
        RECT 53.710000 11.260000 53.910000 11.460000 ;
        RECT 54.115000  6.960000 54.315000  7.160000 ;
        RECT 54.115000  7.390000 54.315000  7.590000 ;
        RECT 54.115000  7.820000 54.315000  8.020000 ;
        RECT 54.115000  8.250000 54.315000  8.450000 ;
        RECT 54.115000  8.680000 54.315000  8.880000 ;
        RECT 54.115000  9.110000 54.315000  9.310000 ;
        RECT 54.115000  9.540000 54.315000  9.740000 ;
        RECT 54.115000  9.970000 54.315000 10.170000 ;
        RECT 54.115000 10.400000 54.315000 10.600000 ;
        RECT 54.115000 10.830000 54.315000 11.030000 ;
        RECT 54.115000 11.260000 54.315000 11.460000 ;
        RECT 54.520000  6.960000 54.720000  7.160000 ;
        RECT 54.520000  7.390000 54.720000  7.590000 ;
        RECT 54.520000  7.820000 54.720000  8.020000 ;
        RECT 54.520000  8.250000 54.720000  8.450000 ;
        RECT 54.520000  8.680000 54.720000  8.880000 ;
        RECT 54.520000  9.110000 54.720000  9.310000 ;
        RECT 54.520000  9.540000 54.720000  9.740000 ;
        RECT 54.520000  9.970000 54.720000 10.170000 ;
        RECT 54.520000 10.400000 54.720000 10.600000 ;
        RECT 54.520000 10.830000 54.720000 11.030000 ;
        RECT 54.520000 11.260000 54.720000 11.460000 ;
        RECT 54.925000  6.960000 55.125000  7.160000 ;
        RECT 54.925000  7.390000 55.125000  7.590000 ;
        RECT 54.925000  7.820000 55.125000  8.020000 ;
        RECT 54.925000  8.250000 55.125000  8.450000 ;
        RECT 54.925000  8.680000 55.125000  8.880000 ;
        RECT 54.925000  9.110000 55.125000  9.310000 ;
        RECT 54.925000  9.540000 55.125000  9.740000 ;
        RECT 54.925000  9.970000 55.125000 10.170000 ;
        RECT 54.925000 10.400000 55.125000 10.600000 ;
        RECT 54.925000 10.830000 55.125000 11.030000 ;
        RECT 54.925000 11.260000 55.125000 11.460000 ;
        RECT 55.330000  6.960000 55.530000  7.160000 ;
        RECT 55.330000  7.390000 55.530000  7.590000 ;
        RECT 55.330000  7.820000 55.530000  8.020000 ;
        RECT 55.330000  8.250000 55.530000  8.450000 ;
        RECT 55.330000  8.680000 55.530000  8.880000 ;
        RECT 55.330000  9.110000 55.530000  9.310000 ;
        RECT 55.330000  9.540000 55.530000  9.740000 ;
        RECT 55.330000  9.970000 55.530000 10.170000 ;
        RECT 55.330000 10.400000 55.530000 10.600000 ;
        RECT 55.330000 10.830000 55.530000 11.030000 ;
        RECT 55.330000 11.260000 55.530000 11.460000 ;
        RECT 55.735000  6.960000 55.935000  7.160000 ;
        RECT 55.735000  7.390000 55.935000  7.590000 ;
        RECT 55.735000  7.820000 55.935000  8.020000 ;
        RECT 55.735000  8.250000 55.935000  8.450000 ;
        RECT 55.735000  8.680000 55.935000  8.880000 ;
        RECT 55.735000  9.110000 55.935000  9.310000 ;
        RECT 55.735000  9.540000 55.935000  9.740000 ;
        RECT 55.735000  9.970000 55.935000 10.170000 ;
        RECT 55.735000 10.400000 55.935000 10.600000 ;
        RECT 55.735000 10.830000 55.935000 11.030000 ;
        RECT 55.735000 11.260000 55.935000 11.460000 ;
        RECT 56.140000  6.960000 56.340000  7.160000 ;
        RECT 56.140000  7.390000 56.340000  7.590000 ;
        RECT 56.140000  7.820000 56.340000  8.020000 ;
        RECT 56.140000  8.250000 56.340000  8.450000 ;
        RECT 56.140000  8.680000 56.340000  8.880000 ;
        RECT 56.140000  9.110000 56.340000  9.310000 ;
        RECT 56.140000  9.540000 56.340000  9.740000 ;
        RECT 56.140000  9.970000 56.340000 10.170000 ;
        RECT 56.140000 10.400000 56.340000 10.600000 ;
        RECT 56.140000 10.830000 56.340000 11.030000 ;
        RECT 56.140000 11.260000 56.340000 11.460000 ;
        RECT 56.545000  6.960000 56.745000  7.160000 ;
        RECT 56.545000  7.390000 56.745000  7.590000 ;
        RECT 56.545000  7.820000 56.745000  8.020000 ;
        RECT 56.545000  8.250000 56.745000  8.450000 ;
        RECT 56.545000  8.680000 56.745000  8.880000 ;
        RECT 56.545000  9.110000 56.745000  9.310000 ;
        RECT 56.545000  9.540000 56.745000  9.740000 ;
        RECT 56.545000  9.970000 56.745000 10.170000 ;
        RECT 56.545000 10.400000 56.745000 10.600000 ;
        RECT 56.545000 10.830000 56.745000 11.030000 ;
        RECT 56.545000 11.260000 56.745000 11.460000 ;
        RECT 56.950000  6.960000 57.150000  7.160000 ;
        RECT 56.950000  7.390000 57.150000  7.590000 ;
        RECT 56.950000  7.820000 57.150000  8.020000 ;
        RECT 56.950000  8.250000 57.150000  8.450000 ;
        RECT 56.950000  8.680000 57.150000  8.880000 ;
        RECT 56.950000  9.110000 57.150000  9.310000 ;
        RECT 56.950000  9.540000 57.150000  9.740000 ;
        RECT 56.950000  9.970000 57.150000 10.170000 ;
        RECT 56.950000 10.400000 57.150000 10.600000 ;
        RECT 56.950000 10.830000 57.150000 11.030000 ;
        RECT 56.950000 11.260000 57.150000 11.460000 ;
        RECT 57.355000  6.960000 57.555000  7.160000 ;
        RECT 57.355000  7.390000 57.555000  7.590000 ;
        RECT 57.355000  7.820000 57.555000  8.020000 ;
        RECT 57.355000  8.250000 57.555000  8.450000 ;
        RECT 57.355000  8.680000 57.555000  8.880000 ;
        RECT 57.355000  9.110000 57.555000  9.310000 ;
        RECT 57.355000  9.540000 57.555000  9.740000 ;
        RECT 57.355000  9.970000 57.555000 10.170000 ;
        RECT 57.355000 10.400000 57.555000 10.600000 ;
        RECT 57.355000 10.830000 57.555000 11.030000 ;
        RECT 57.355000 11.260000 57.555000 11.460000 ;
        RECT 57.760000  6.960000 57.960000  7.160000 ;
        RECT 57.760000  7.390000 57.960000  7.590000 ;
        RECT 57.760000  7.820000 57.960000  8.020000 ;
        RECT 57.760000  8.250000 57.960000  8.450000 ;
        RECT 57.760000  8.680000 57.960000  8.880000 ;
        RECT 57.760000  9.110000 57.960000  9.310000 ;
        RECT 57.760000  9.540000 57.960000  9.740000 ;
        RECT 57.760000  9.970000 57.960000 10.170000 ;
        RECT 57.760000 10.400000 57.960000 10.600000 ;
        RECT 57.760000 10.830000 57.960000 11.030000 ;
        RECT 57.760000 11.260000 57.960000 11.460000 ;
        RECT 58.165000  6.960000 58.365000  7.160000 ;
        RECT 58.165000  7.390000 58.365000  7.590000 ;
        RECT 58.165000  7.820000 58.365000  8.020000 ;
        RECT 58.165000  8.250000 58.365000  8.450000 ;
        RECT 58.165000  8.680000 58.365000  8.880000 ;
        RECT 58.165000  9.110000 58.365000  9.310000 ;
        RECT 58.165000  9.540000 58.365000  9.740000 ;
        RECT 58.165000  9.970000 58.365000 10.170000 ;
        RECT 58.165000 10.400000 58.365000 10.600000 ;
        RECT 58.165000 10.830000 58.365000 11.030000 ;
        RECT 58.165000 11.260000 58.365000 11.460000 ;
        RECT 58.570000  6.960000 58.770000  7.160000 ;
        RECT 58.570000  7.390000 58.770000  7.590000 ;
        RECT 58.570000  7.820000 58.770000  8.020000 ;
        RECT 58.570000  8.250000 58.770000  8.450000 ;
        RECT 58.570000  8.680000 58.770000  8.880000 ;
        RECT 58.570000  9.110000 58.770000  9.310000 ;
        RECT 58.570000  9.540000 58.770000  9.740000 ;
        RECT 58.570000  9.970000 58.770000 10.170000 ;
        RECT 58.570000 10.400000 58.770000 10.600000 ;
        RECT 58.570000 10.830000 58.770000 11.030000 ;
        RECT 58.570000 11.260000 58.770000 11.460000 ;
        RECT 58.975000  6.960000 59.175000  7.160000 ;
        RECT 58.975000  7.390000 59.175000  7.590000 ;
        RECT 58.975000  7.820000 59.175000  8.020000 ;
        RECT 58.975000  8.250000 59.175000  8.450000 ;
        RECT 58.975000  8.680000 59.175000  8.880000 ;
        RECT 58.975000  9.110000 59.175000  9.310000 ;
        RECT 58.975000  9.540000 59.175000  9.740000 ;
        RECT 58.975000  9.970000 59.175000 10.170000 ;
        RECT 58.975000 10.400000 59.175000 10.600000 ;
        RECT 58.975000 10.830000 59.175000 11.030000 ;
        RECT 58.975000 11.260000 59.175000 11.460000 ;
        RECT 59.380000  6.960000 59.580000  7.160000 ;
        RECT 59.380000  7.390000 59.580000  7.590000 ;
        RECT 59.380000  7.820000 59.580000  8.020000 ;
        RECT 59.380000  8.250000 59.580000  8.450000 ;
        RECT 59.380000  8.680000 59.580000  8.880000 ;
        RECT 59.380000  9.110000 59.580000  9.310000 ;
        RECT 59.380000  9.540000 59.580000  9.740000 ;
        RECT 59.380000  9.970000 59.580000 10.170000 ;
        RECT 59.380000 10.400000 59.580000 10.600000 ;
        RECT 59.380000 10.830000 59.580000 11.030000 ;
        RECT 59.380000 11.260000 59.580000 11.460000 ;
        RECT 59.785000  6.960000 59.985000  7.160000 ;
        RECT 59.785000  7.390000 59.985000  7.590000 ;
        RECT 59.785000  7.820000 59.985000  8.020000 ;
        RECT 59.785000  8.250000 59.985000  8.450000 ;
        RECT 59.785000  8.680000 59.985000  8.880000 ;
        RECT 59.785000  9.110000 59.985000  9.310000 ;
        RECT 59.785000  9.540000 59.985000  9.740000 ;
        RECT 59.785000  9.970000 59.985000 10.170000 ;
        RECT 59.785000 10.400000 59.985000 10.600000 ;
        RECT 59.785000 10.830000 59.985000 11.030000 ;
        RECT 59.785000 11.260000 59.985000 11.460000 ;
        RECT 60.190000  6.960000 60.390000  7.160000 ;
        RECT 60.190000  7.390000 60.390000  7.590000 ;
        RECT 60.190000  7.820000 60.390000  8.020000 ;
        RECT 60.190000  8.250000 60.390000  8.450000 ;
        RECT 60.190000  8.680000 60.390000  8.880000 ;
        RECT 60.190000  9.110000 60.390000  9.310000 ;
        RECT 60.190000  9.540000 60.390000  9.740000 ;
        RECT 60.190000  9.970000 60.390000 10.170000 ;
        RECT 60.190000 10.400000 60.390000 10.600000 ;
        RECT 60.190000 10.830000 60.390000 11.030000 ;
        RECT 60.190000 11.260000 60.390000 11.460000 ;
        RECT 60.595000  6.960000 60.795000  7.160000 ;
        RECT 60.595000  7.390000 60.795000  7.590000 ;
        RECT 60.595000  7.820000 60.795000  8.020000 ;
        RECT 60.595000  8.250000 60.795000  8.450000 ;
        RECT 60.595000  8.680000 60.795000  8.880000 ;
        RECT 60.595000  9.110000 60.795000  9.310000 ;
        RECT 60.595000  9.540000 60.795000  9.740000 ;
        RECT 60.595000  9.970000 60.795000 10.170000 ;
        RECT 60.595000 10.400000 60.795000 10.600000 ;
        RECT 60.595000 10.830000 60.795000 11.030000 ;
        RECT 60.595000 11.260000 60.795000 11.460000 ;
        RECT 61.000000  6.960000 61.200000  7.160000 ;
        RECT 61.000000  7.390000 61.200000  7.590000 ;
        RECT 61.000000  7.820000 61.200000  8.020000 ;
        RECT 61.000000  8.250000 61.200000  8.450000 ;
        RECT 61.000000  8.680000 61.200000  8.880000 ;
        RECT 61.000000  9.110000 61.200000  9.310000 ;
        RECT 61.000000  9.540000 61.200000  9.740000 ;
        RECT 61.000000  9.970000 61.200000 10.170000 ;
        RECT 61.000000 10.400000 61.200000 10.600000 ;
        RECT 61.000000 10.830000 61.200000 11.030000 ;
        RECT 61.000000 11.260000 61.200000 11.460000 ;
        RECT 61.405000  6.960000 61.605000  7.160000 ;
        RECT 61.405000  7.390000 61.605000  7.590000 ;
        RECT 61.405000  7.820000 61.605000  8.020000 ;
        RECT 61.405000  8.250000 61.605000  8.450000 ;
        RECT 61.405000  8.680000 61.605000  8.880000 ;
        RECT 61.405000  9.110000 61.605000  9.310000 ;
        RECT 61.405000  9.540000 61.605000  9.740000 ;
        RECT 61.405000  9.970000 61.605000 10.170000 ;
        RECT 61.405000 10.400000 61.605000 10.600000 ;
        RECT 61.405000 10.830000 61.605000 11.030000 ;
        RECT 61.405000 11.260000 61.605000 11.460000 ;
        RECT 61.810000  6.960000 62.010000  7.160000 ;
        RECT 61.810000  7.390000 62.010000  7.590000 ;
        RECT 61.810000  7.820000 62.010000  8.020000 ;
        RECT 61.810000  8.250000 62.010000  8.450000 ;
        RECT 61.810000  8.680000 62.010000  8.880000 ;
        RECT 61.810000  9.110000 62.010000  9.310000 ;
        RECT 61.810000  9.540000 62.010000  9.740000 ;
        RECT 61.810000  9.970000 62.010000 10.170000 ;
        RECT 61.810000 10.400000 62.010000 10.600000 ;
        RECT 61.810000 10.830000 62.010000 11.030000 ;
        RECT 61.810000 11.260000 62.010000 11.460000 ;
        RECT 62.215000  6.960000 62.415000  7.160000 ;
        RECT 62.215000  7.390000 62.415000  7.590000 ;
        RECT 62.215000  7.820000 62.415000  8.020000 ;
        RECT 62.215000  8.250000 62.415000  8.450000 ;
        RECT 62.215000  8.680000 62.415000  8.880000 ;
        RECT 62.215000  9.110000 62.415000  9.310000 ;
        RECT 62.215000  9.540000 62.415000  9.740000 ;
        RECT 62.215000  9.970000 62.415000 10.170000 ;
        RECT 62.215000 10.400000 62.415000 10.600000 ;
        RECT 62.215000 10.830000 62.415000 11.030000 ;
        RECT 62.215000 11.260000 62.415000 11.460000 ;
        RECT 62.620000  6.960000 62.820000  7.160000 ;
        RECT 62.620000  7.390000 62.820000  7.590000 ;
        RECT 62.620000  7.820000 62.820000  8.020000 ;
        RECT 62.620000  8.250000 62.820000  8.450000 ;
        RECT 62.620000  8.680000 62.820000  8.880000 ;
        RECT 62.620000  9.110000 62.820000  9.310000 ;
        RECT 62.620000  9.540000 62.820000  9.740000 ;
        RECT 62.620000  9.970000 62.820000 10.170000 ;
        RECT 62.620000 10.400000 62.820000 10.600000 ;
        RECT 62.620000 10.830000 62.820000 11.030000 ;
        RECT 62.620000 11.260000 62.820000 11.460000 ;
        RECT 63.025000  6.960000 63.225000  7.160000 ;
        RECT 63.025000  7.390000 63.225000  7.590000 ;
        RECT 63.025000  7.820000 63.225000  8.020000 ;
        RECT 63.025000  8.250000 63.225000  8.450000 ;
        RECT 63.025000  8.680000 63.225000  8.880000 ;
        RECT 63.025000  9.110000 63.225000  9.310000 ;
        RECT 63.025000  9.540000 63.225000  9.740000 ;
        RECT 63.025000  9.970000 63.225000 10.170000 ;
        RECT 63.025000 10.400000 63.225000 10.600000 ;
        RECT 63.025000 10.830000 63.225000 11.030000 ;
        RECT 63.025000 11.260000 63.225000 11.460000 ;
        RECT 63.430000  6.960000 63.630000  7.160000 ;
        RECT 63.430000  7.390000 63.630000  7.590000 ;
        RECT 63.430000  7.820000 63.630000  8.020000 ;
        RECT 63.430000  8.250000 63.630000  8.450000 ;
        RECT 63.430000  8.680000 63.630000  8.880000 ;
        RECT 63.430000  9.110000 63.630000  9.310000 ;
        RECT 63.430000  9.540000 63.630000  9.740000 ;
        RECT 63.430000  9.970000 63.630000 10.170000 ;
        RECT 63.430000 10.400000 63.630000 10.600000 ;
        RECT 63.430000 10.830000 63.630000 11.030000 ;
        RECT 63.430000 11.260000 63.630000 11.460000 ;
        RECT 63.835000  6.960000 64.035000  7.160000 ;
        RECT 63.835000  7.390000 64.035000  7.590000 ;
        RECT 63.835000  7.820000 64.035000  8.020000 ;
        RECT 63.835000  8.250000 64.035000  8.450000 ;
        RECT 63.835000  8.680000 64.035000  8.880000 ;
        RECT 63.835000  9.110000 64.035000  9.310000 ;
        RECT 63.835000  9.540000 64.035000  9.740000 ;
        RECT 63.835000  9.970000 64.035000 10.170000 ;
        RECT 63.835000 10.400000 64.035000 10.600000 ;
        RECT 63.835000 10.830000 64.035000 11.030000 ;
        RECT 63.835000 11.260000 64.035000 11.460000 ;
        RECT 64.240000  6.960000 64.440000  7.160000 ;
        RECT 64.240000  7.390000 64.440000  7.590000 ;
        RECT 64.240000  7.820000 64.440000  8.020000 ;
        RECT 64.240000  8.250000 64.440000  8.450000 ;
        RECT 64.240000  8.680000 64.440000  8.880000 ;
        RECT 64.240000  9.110000 64.440000  9.310000 ;
        RECT 64.240000  9.540000 64.440000  9.740000 ;
        RECT 64.240000  9.970000 64.440000 10.170000 ;
        RECT 64.240000 10.400000 64.440000 10.600000 ;
        RECT 64.240000 10.830000 64.440000 11.030000 ;
        RECT 64.240000 11.260000 64.440000 11.460000 ;
        RECT 64.645000  6.960000 64.845000  7.160000 ;
        RECT 64.645000  7.390000 64.845000  7.590000 ;
        RECT 64.645000  7.820000 64.845000  8.020000 ;
        RECT 64.645000  8.250000 64.845000  8.450000 ;
        RECT 64.645000  8.680000 64.845000  8.880000 ;
        RECT 64.645000  9.110000 64.845000  9.310000 ;
        RECT 64.645000  9.540000 64.845000  9.740000 ;
        RECT 64.645000  9.970000 64.845000 10.170000 ;
        RECT 64.645000 10.400000 64.845000 10.600000 ;
        RECT 64.645000 10.830000 64.845000 11.030000 ;
        RECT 64.645000 11.260000 64.845000 11.460000 ;
        RECT 65.050000  6.960000 65.250000  7.160000 ;
        RECT 65.050000  7.390000 65.250000  7.590000 ;
        RECT 65.050000  7.820000 65.250000  8.020000 ;
        RECT 65.050000  8.250000 65.250000  8.450000 ;
        RECT 65.050000  8.680000 65.250000  8.880000 ;
        RECT 65.050000  9.110000 65.250000  9.310000 ;
        RECT 65.050000  9.540000 65.250000  9.740000 ;
        RECT 65.050000  9.970000 65.250000 10.170000 ;
        RECT 65.050000 10.400000 65.250000 10.600000 ;
        RECT 65.050000 10.830000 65.250000 11.030000 ;
        RECT 65.050000 11.260000 65.250000 11.460000 ;
        RECT 65.455000  6.960000 65.655000  7.160000 ;
        RECT 65.455000  7.390000 65.655000  7.590000 ;
        RECT 65.455000  7.820000 65.655000  8.020000 ;
        RECT 65.455000  8.250000 65.655000  8.450000 ;
        RECT 65.455000  8.680000 65.655000  8.880000 ;
        RECT 65.455000  9.110000 65.655000  9.310000 ;
        RECT 65.455000  9.540000 65.655000  9.740000 ;
        RECT 65.455000  9.970000 65.655000 10.170000 ;
        RECT 65.455000 10.400000 65.655000 10.600000 ;
        RECT 65.455000 10.830000 65.655000 11.030000 ;
        RECT 65.455000 11.260000 65.655000 11.460000 ;
        RECT 65.860000  6.960000 66.060000  7.160000 ;
        RECT 65.860000  7.390000 66.060000  7.590000 ;
        RECT 65.860000  7.820000 66.060000  8.020000 ;
        RECT 65.860000  8.250000 66.060000  8.450000 ;
        RECT 65.860000  8.680000 66.060000  8.880000 ;
        RECT 65.860000  9.110000 66.060000  9.310000 ;
        RECT 65.860000  9.540000 66.060000  9.740000 ;
        RECT 65.860000  9.970000 66.060000 10.170000 ;
        RECT 65.860000 10.400000 66.060000 10.600000 ;
        RECT 65.860000 10.830000 66.060000 11.030000 ;
        RECT 65.860000 11.260000 66.060000 11.460000 ;
        RECT 66.265000  6.960000 66.465000  7.160000 ;
        RECT 66.265000  7.390000 66.465000  7.590000 ;
        RECT 66.265000  7.820000 66.465000  8.020000 ;
        RECT 66.265000  8.250000 66.465000  8.450000 ;
        RECT 66.265000  8.680000 66.465000  8.880000 ;
        RECT 66.265000  9.110000 66.465000  9.310000 ;
        RECT 66.265000  9.540000 66.465000  9.740000 ;
        RECT 66.265000  9.970000 66.465000 10.170000 ;
        RECT 66.265000 10.400000 66.465000 10.600000 ;
        RECT 66.265000 10.830000 66.465000 11.030000 ;
        RECT 66.265000 11.260000 66.465000 11.460000 ;
        RECT 66.670000  6.960000 66.870000  7.160000 ;
        RECT 66.670000  7.390000 66.870000  7.590000 ;
        RECT 66.670000  7.820000 66.870000  8.020000 ;
        RECT 66.670000  8.250000 66.870000  8.450000 ;
        RECT 66.670000  8.680000 66.870000  8.880000 ;
        RECT 66.670000  9.110000 66.870000  9.310000 ;
        RECT 66.670000  9.540000 66.870000  9.740000 ;
        RECT 66.670000  9.970000 66.870000 10.170000 ;
        RECT 66.670000 10.400000 66.870000 10.600000 ;
        RECT 66.670000 10.830000 66.870000 11.030000 ;
        RECT 66.670000 11.260000 66.870000 11.460000 ;
        RECT 67.075000  6.960000 67.275000  7.160000 ;
        RECT 67.075000  7.390000 67.275000  7.590000 ;
        RECT 67.075000  7.820000 67.275000  8.020000 ;
        RECT 67.075000  8.250000 67.275000  8.450000 ;
        RECT 67.075000  8.680000 67.275000  8.880000 ;
        RECT 67.075000  9.110000 67.275000  9.310000 ;
        RECT 67.075000  9.540000 67.275000  9.740000 ;
        RECT 67.075000  9.970000 67.275000 10.170000 ;
        RECT 67.075000 10.400000 67.275000 10.600000 ;
        RECT 67.075000 10.830000 67.275000 11.030000 ;
        RECT 67.075000 11.260000 67.275000 11.460000 ;
        RECT 67.480000  6.960000 67.680000  7.160000 ;
        RECT 67.480000  7.390000 67.680000  7.590000 ;
        RECT 67.480000  7.820000 67.680000  8.020000 ;
        RECT 67.480000  8.250000 67.680000  8.450000 ;
        RECT 67.480000  8.680000 67.680000  8.880000 ;
        RECT 67.480000  9.110000 67.680000  9.310000 ;
        RECT 67.480000  9.540000 67.680000  9.740000 ;
        RECT 67.480000  9.970000 67.680000 10.170000 ;
        RECT 67.480000 10.400000 67.680000 10.600000 ;
        RECT 67.480000 10.830000 67.680000 11.030000 ;
        RECT 67.480000 11.260000 67.680000 11.460000 ;
        RECT 67.885000  6.960000 68.085000  7.160000 ;
        RECT 67.885000  7.390000 68.085000  7.590000 ;
        RECT 67.885000  7.820000 68.085000  8.020000 ;
        RECT 67.885000  8.250000 68.085000  8.450000 ;
        RECT 67.885000  8.680000 68.085000  8.880000 ;
        RECT 67.885000  9.110000 68.085000  9.310000 ;
        RECT 67.885000  9.540000 68.085000  9.740000 ;
        RECT 67.885000  9.970000 68.085000 10.170000 ;
        RECT 67.885000 10.400000 68.085000 10.600000 ;
        RECT 67.885000 10.830000 68.085000 11.030000 ;
        RECT 67.885000 11.260000 68.085000 11.460000 ;
        RECT 68.290000  6.960000 68.490000  7.160000 ;
        RECT 68.290000  7.390000 68.490000  7.590000 ;
        RECT 68.290000  7.820000 68.490000  8.020000 ;
        RECT 68.290000  8.250000 68.490000  8.450000 ;
        RECT 68.290000  8.680000 68.490000  8.880000 ;
        RECT 68.290000  9.110000 68.490000  9.310000 ;
        RECT 68.290000  9.540000 68.490000  9.740000 ;
        RECT 68.290000  9.970000 68.490000 10.170000 ;
        RECT 68.290000 10.400000 68.490000 10.600000 ;
        RECT 68.290000 10.830000 68.490000 11.030000 ;
        RECT 68.290000 11.260000 68.490000 11.460000 ;
        RECT 68.695000  6.960000 68.895000  7.160000 ;
        RECT 68.695000  7.390000 68.895000  7.590000 ;
        RECT 68.695000  7.820000 68.895000  8.020000 ;
        RECT 68.695000  8.250000 68.895000  8.450000 ;
        RECT 68.695000  8.680000 68.895000  8.880000 ;
        RECT 68.695000  9.110000 68.895000  9.310000 ;
        RECT 68.695000  9.540000 68.895000  9.740000 ;
        RECT 68.695000  9.970000 68.895000 10.170000 ;
        RECT 68.695000 10.400000 68.895000 10.600000 ;
        RECT 68.695000 10.830000 68.895000 11.030000 ;
        RECT 68.695000 11.260000 68.895000 11.460000 ;
        RECT 69.100000  6.960000 69.300000  7.160000 ;
        RECT 69.100000  7.390000 69.300000  7.590000 ;
        RECT 69.100000  7.820000 69.300000  8.020000 ;
        RECT 69.100000  8.250000 69.300000  8.450000 ;
        RECT 69.100000  8.680000 69.300000  8.880000 ;
        RECT 69.100000  9.110000 69.300000  9.310000 ;
        RECT 69.100000  9.540000 69.300000  9.740000 ;
        RECT 69.100000  9.970000 69.300000 10.170000 ;
        RECT 69.100000 10.400000 69.300000 10.600000 ;
        RECT 69.100000 10.830000 69.300000 11.030000 ;
        RECT 69.100000 11.260000 69.300000 11.460000 ;
        RECT 69.505000  6.960000 69.705000  7.160000 ;
        RECT 69.505000  7.390000 69.705000  7.590000 ;
        RECT 69.505000  7.820000 69.705000  8.020000 ;
        RECT 69.505000  8.250000 69.705000  8.450000 ;
        RECT 69.505000  8.680000 69.705000  8.880000 ;
        RECT 69.505000  9.110000 69.705000  9.310000 ;
        RECT 69.505000  9.540000 69.705000  9.740000 ;
        RECT 69.505000  9.970000 69.705000 10.170000 ;
        RECT 69.505000 10.400000 69.705000 10.600000 ;
        RECT 69.505000 10.830000 69.705000 11.030000 ;
        RECT 69.505000 11.260000 69.705000 11.460000 ;
        RECT 69.910000  6.960000 70.110000  7.160000 ;
        RECT 69.910000  7.390000 70.110000  7.590000 ;
        RECT 69.910000  7.820000 70.110000  8.020000 ;
        RECT 69.910000  8.250000 70.110000  8.450000 ;
        RECT 69.910000  8.680000 70.110000  8.880000 ;
        RECT 69.910000  9.110000 70.110000  9.310000 ;
        RECT 69.910000  9.540000 70.110000  9.740000 ;
        RECT 69.910000  9.970000 70.110000 10.170000 ;
        RECT 69.910000 10.400000 70.110000 10.600000 ;
        RECT 69.910000 10.830000 70.110000 11.030000 ;
        RECT 69.910000 11.260000 70.110000 11.460000 ;
        RECT 70.315000  6.960000 70.515000  7.160000 ;
        RECT 70.315000  7.390000 70.515000  7.590000 ;
        RECT 70.315000  7.820000 70.515000  8.020000 ;
        RECT 70.315000  8.250000 70.515000  8.450000 ;
        RECT 70.315000  8.680000 70.515000  8.880000 ;
        RECT 70.315000  9.110000 70.515000  9.310000 ;
        RECT 70.315000  9.540000 70.515000  9.740000 ;
        RECT 70.315000  9.970000 70.515000 10.170000 ;
        RECT 70.315000 10.400000 70.515000 10.600000 ;
        RECT 70.315000 10.830000 70.515000 11.030000 ;
        RECT 70.315000 11.260000 70.515000 11.460000 ;
        RECT 70.720000  6.960000 70.920000  7.160000 ;
        RECT 70.720000  7.390000 70.920000  7.590000 ;
        RECT 70.720000  7.820000 70.920000  8.020000 ;
        RECT 70.720000  8.250000 70.920000  8.450000 ;
        RECT 70.720000  8.680000 70.920000  8.880000 ;
        RECT 70.720000  9.110000 70.920000  9.310000 ;
        RECT 70.720000  9.540000 70.920000  9.740000 ;
        RECT 70.720000  9.970000 70.920000 10.170000 ;
        RECT 70.720000 10.400000 70.920000 10.600000 ;
        RECT 70.720000 10.830000 70.920000 11.030000 ;
        RECT 70.720000 11.260000 70.920000 11.460000 ;
        RECT 71.125000  6.960000 71.325000  7.160000 ;
        RECT 71.125000  7.390000 71.325000  7.590000 ;
        RECT 71.125000  7.820000 71.325000  8.020000 ;
        RECT 71.125000  8.250000 71.325000  8.450000 ;
        RECT 71.125000  8.680000 71.325000  8.880000 ;
        RECT 71.125000  9.110000 71.325000  9.310000 ;
        RECT 71.125000  9.540000 71.325000  9.740000 ;
        RECT 71.125000  9.970000 71.325000 10.170000 ;
        RECT 71.125000 10.400000 71.325000 10.600000 ;
        RECT 71.125000 10.830000 71.325000 11.030000 ;
        RECT 71.125000 11.260000 71.325000 11.460000 ;
        RECT 71.530000  6.960000 71.730000  7.160000 ;
        RECT 71.530000  7.390000 71.730000  7.590000 ;
        RECT 71.530000  7.820000 71.730000  8.020000 ;
        RECT 71.530000  8.250000 71.730000  8.450000 ;
        RECT 71.530000  8.680000 71.730000  8.880000 ;
        RECT 71.530000  9.110000 71.730000  9.310000 ;
        RECT 71.530000  9.540000 71.730000  9.740000 ;
        RECT 71.530000  9.970000 71.730000 10.170000 ;
        RECT 71.530000 10.400000 71.730000 10.600000 ;
        RECT 71.530000 10.830000 71.730000 11.030000 ;
        RECT 71.530000 11.260000 71.730000 11.460000 ;
        RECT 71.935000  6.960000 72.135000  7.160000 ;
        RECT 71.935000  7.390000 72.135000  7.590000 ;
        RECT 71.935000  7.820000 72.135000  8.020000 ;
        RECT 71.935000  8.250000 72.135000  8.450000 ;
        RECT 71.935000  8.680000 72.135000  8.880000 ;
        RECT 71.935000  9.110000 72.135000  9.310000 ;
        RECT 71.935000  9.540000 72.135000  9.740000 ;
        RECT 71.935000  9.970000 72.135000 10.170000 ;
        RECT 71.935000 10.400000 72.135000 10.600000 ;
        RECT 71.935000 10.830000 72.135000 11.030000 ;
        RECT 71.935000 11.260000 72.135000 11.460000 ;
        RECT 72.340000  6.960000 72.540000  7.160000 ;
        RECT 72.340000  7.390000 72.540000  7.590000 ;
        RECT 72.340000  7.820000 72.540000  8.020000 ;
        RECT 72.340000  8.250000 72.540000  8.450000 ;
        RECT 72.340000  8.680000 72.540000  8.880000 ;
        RECT 72.340000  9.110000 72.540000  9.310000 ;
        RECT 72.340000  9.540000 72.540000  9.740000 ;
        RECT 72.340000  9.970000 72.540000 10.170000 ;
        RECT 72.340000 10.400000 72.540000 10.600000 ;
        RECT 72.340000 10.830000 72.540000 11.030000 ;
        RECT 72.340000 11.260000 72.540000 11.460000 ;
        RECT 72.745000  6.960000 72.945000  7.160000 ;
        RECT 72.745000  7.390000 72.945000  7.590000 ;
        RECT 72.745000  7.820000 72.945000  8.020000 ;
        RECT 72.745000  8.250000 72.945000  8.450000 ;
        RECT 72.745000  8.680000 72.945000  8.880000 ;
        RECT 72.745000  9.110000 72.945000  9.310000 ;
        RECT 72.745000  9.540000 72.945000  9.740000 ;
        RECT 72.745000  9.970000 72.945000 10.170000 ;
        RECT 72.745000 10.400000 72.945000 10.600000 ;
        RECT 72.745000 10.830000 72.945000 11.030000 ;
        RECT 72.745000 11.260000 72.945000 11.460000 ;
        RECT 73.150000  6.960000 73.350000  7.160000 ;
        RECT 73.150000  7.390000 73.350000  7.590000 ;
        RECT 73.150000  7.820000 73.350000  8.020000 ;
        RECT 73.150000  8.250000 73.350000  8.450000 ;
        RECT 73.150000  8.680000 73.350000  8.880000 ;
        RECT 73.150000  9.110000 73.350000  9.310000 ;
        RECT 73.150000  9.540000 73.350000  9.740000 ;
        RECT 73.150000  9.970000 73.350000 10.170000 ;
        RECT 73.150000 10.400000 73.350000 10.600000 ;
        RECT 73.150000 10.830000 73.350000 11.030000 ;
        RECT 73.150000 11.260000 73.350000 11.460000 ;
        RECT 73.555000  6.960000 73.755000  7.160000 ;
        RECT 73.555000  7.390000 73.755000  7.590000 ;
        RECT 73.555000  7.820000 73.755000  8.020000 ;
        RECT 73.555000  8.250000 73.755000  8.450000 ;
        RECT 73.555000  8.680000 73.755000  8.880000 ;
        RECT 73.555000  9.110000 73.755000  9.310000 ;
        RECT 73.555000  9.540000 73.755000  9.740000 ;
        RECT 73.555000  9.970000 73.755000 10.170000 ;
        RECT 73.555000 10.400000 73.755000 10.600000 ;
        RECT 73.555000 10.830000 73.755000 11.030000 ;
        RECT 73.555000 11.260000 73.755000 11.460000 ;
        RECT 73.960000  6.960000 74.160000  7.160000 ;
        RECT 73.960000  7.390000 74.160000  7.590000 ;
        RECT 73.960000  7.820000 74.160000  8.020000 ;
        RECT 73.960000  8.250000 74.160000  8.450000 ;
        RECT 73.960000  8.680000 74.160000  8.880000 ;
        RECT 73.960000  9.110000 74.160000  9.310000 ;
        RECT 73.960000  9.540000 74.160000  9.740000 ;
        RECT 73.960000  9.970000 74.160000 10.170000 ;
        RECT 73.960000 10.400000 74.160000 10.600000 ;
        RECT 73.960000 10.830000 74.160000 11.030000 ;
        RECT 73.960000 11.260000 74.160000 11.460000 ;
        RECT 74.365000  6.960000 74.565000  7.160000 ;
        RECT 74.365000  7.390000 74.565000  7.590000 ;
        RECT 74.365000  7.820000 74.565000  8.020000 ;
        RECT 74.365000  8.250000 74.565000  8.450000 ;
        RECT 74.365000  8.680000 74.565000  8.880000 ;
        RECT 74.365000  9.110000 74.565000  9.310000 ;
        RECT 74.365000  9.540000 74.565000  9.740000 ;
        RECT 74.365000  9.970000 74.565000 10.170000 ;
        RECT 74.365000 10.400000 74.565000 10.600000 ;
        RECT 74.365000 10.830000 74.565000 11.030000 ;
        RECT 74.365000 11.260000 74.565000 11.460000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 0.035000 1.270000 5.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 0.035000 75.000000 5.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 0.135000 1.270000 5.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 12.935000 0.965000 16.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 12.935000 75.000000 16.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 13.035000 0.965000 16.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 17.785000 1.270000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 68.035000 1.270000 93.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 17.785000 75.000000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 68.035000 75.000000 93.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 17.885000 1.270000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 68.035000 1.270000 92.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 17.885000 75.000000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 62.085000 1.270000 66.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 62.085000 75.000000 66.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 62.185000 1.270000 66.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 34.735000 1.270000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 45.735000 1.270000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 49.645000 1.270000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 54.405000 1.270000 54.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 34.735000 75.000000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 45.735000 75.000000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 49.645000 75.000000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 54.405000 75.000000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 34.840000 1.270000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 45.735000 1.270000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 34.840000 75.000000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 39.585000 1.270000 44.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 39.585000 75.000000 44.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 39.685000 1.270000 44.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 23.835000 1.270000 28.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 23.835000 75.000000 28.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 23.935000 1.270000 28.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 56.235000 1.270000 60.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.235000 75.000000 60.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 56.335000 1.270000 60.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 29.885000 1.270000 33.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 29.885000 75.000000 33.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 29.985000 1.270000 33.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 198.000000 ;
  END
END sky130_fd_io__overlay_vccd_lvc
END LIBRARY
