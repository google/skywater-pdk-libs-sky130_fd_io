# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__top_sio_macro
  CLASS BLOCK ;
  FOREIGN sky130_fd_io__top_sio_macro ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  480.0000 BY  253.7150 ;
  SYMMETRY R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 106.840000 480.000000 109.820000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 102.080000 480.000000 105.060000 ;
    END
  END AMUXBUS_B
  PIN DFT_REFGEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.655000 0.000000 451.915000 236.650000 ;
    END
  END DFT_REFGEN
  PIN DM0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.380000 0.000000 156.640000 28.955000 ;
    END
  END DM0[0]
  PIN DM0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.980000 0.000000 156.240000 33.225000 ;
    END
  END DM0[1]
  PIN DM0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.810000 0.000000 154.070000 42.095000 ;
    END
  END DM0[2]
  PIN DM1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.365000 0.000000 233.625000 28.955000 ;
    END
  END DM1[0]
  PIN DM1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.765000 0.000000 234.025000 33.225000 ;
    END
  END DM1[1]
  PIN DM1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.935000 0.000000 236.195000 42.095000 ;
    END
  END DM1[2]
  PIN ENABLE_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.335000 0.000000 236.595000 2.190000 ;
    END
    PORT
      LAYER met2 ;
        RECT 236.335000 0.000000 236.595000 2.210000 ;
    END
    PORT
      LAYER met2 ;
        RECT 236.335000 2.210000 236.615000 2.230000 ;
    END
    PORT
      LAYER met2 ;
        RECT 236.335000 2.235000 236.640000 3.005000 ;
    END
    PORT
      LAYER met2 ;
        RECT 236.335000 2.960000 236.595000 3.050000 ;
    END
    PORT
      LAYER met2 ;
        RECT 236.335000 3.005000 236.620000 3.025000 ;
    END
    PORT
      LAYER met2 ;
        RECT 236.335000 3.050000 236.595000 34.945000 ;
    END
    PORT
      LAYER met2 ;
        RECT 236.595000 2.190000 236.640000 2.235000 ;
    END
    PORT
      LAYER met2 ;
        RECT 236.595000 3.005000 236.640000 3.050000 ;
    END
  END ENABLE_H
  PIN ENABLE_VDDA_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.405000 0.000000 452.665000 234.180000 ;
    END
  END ENABLE_VDDA_H
  PIN HLD_H_N[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.575000 0.000000 135.835000 36.690000 ;
    END
  END HLD_H_N[0]
  PIN HLD_H_N[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.170000 0.000000 254.430000 36.690000 ;
    END
  END HLD_H_N[1]
  PIN HLD_H_N_REFGEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.995000 0.000000 405.255000 14.810000 ;
    END
  END HLD_H_N_REFGEN
  PIN HLD_OVR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.200000 0.000000 141.545000 2.085000 ;
    END
  END HLD_OVR[0]
  PIN HLD_OVR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.460000 0.000000 248.805000 2.085000 ;
    END
  END HLD_OVR[1]
  PIN IBUF_SEL[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.175000 0.000000 135.435000 28.950000 ;
    END
  END IBUF_SEL[0]
  PIN IBUF_SEL[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.570000 0.000000 254.830000 28.950000 ;
    END
  END IBUF_SEL[1]
  PIN IBUF_SEL_REFGEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.690000 0.000000 422.950000 22.530000 ;
    END
  END IBUF_SEL_REFGEN
  PIN IN[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.005000 0.000000 142.265000 6.970000 ;
    END
  END IN[0]
  PIN IN[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.740000 0.000000 248.000000 6.970000 ;
    END
  END IN[1]
  PIN INP_DIS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.710000 0.000000 106.970000 1.350000 ;
    END
  END INP_DIS[0]
  PIN INP_DIS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.035000 0.000000 283.295000 1.350000 ;
    END
  END INP_DIS[1]
  PIN IN_H[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.405000 0.000000 142.665000 9.980000 ;
    END
  END IN_H[0]
  PIN IN_H[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.340000 0.000000 247.600000 9.980000 ;
    END
  END IN_H[1]
  PIN OE_N[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.215000 0.000000 147.475000 26.920000 ;
    END
  END OE_N[0]
  PIN OE_N[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.530000 0.000000 242.790000 26.920000 ;
    END
  END OE_N[1]
  PIN OUT[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.455000 0.000000 121.715000 46.020000 ;
    END
  END OUT[0]
  PIN OUT[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.290000 0.000000 268.550000 46.020000 ;
    END
  END OUT[1]
  PIN PAD[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 107.190000 131.985000 169.890000 194.600000 ;
    END
  END PAD[0]
  PIN PAD[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 220.115000 131.985000 282.815000 194.600000 ;
    END
  END PAD[1]
  PIN PAD_A_ESD_0_H[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.260000 0.000000 86.105000 29.615000 ;
    END
  END PAD_A_ESD_0_H[0]
  PIN PAD_A_ESD_0_H[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.900000 0.000000 304.745000 29.615000 ;
    END
  END PAD_A_ESD_0_H[1]
  PIN PAD_A_ESD_1_H[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.990000 0.000000 178.990000 23.820000 ;
    END
  END PAD_A_ESD_1_H[0]
  PIN PAD_A_ESD_1_H[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.015000 0.000000 213.015000 23.820000 ;
    END
  END PAD_A_ESD_1_H[1]
  PIN PAD_A_NOESD_H[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.245000 0.000000 87.095000 24.475000 ;
    END
  END PAD_A_NOESD_H[0]
  PIN PAD_A_NOESD_H[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.910000 0.000000 303.760000 24.475000 ;
    END
  END PAD_A_NOESD_H[1]
  PIN SLOW[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.615000 0.000000 147.875000 45.525000 ;
    END
  END SLOW[0]
  PIN SLOW[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.130000 0.000000 242.390000 45.525000 ;
    END
  END SLOW[1]
  PIN TIE_LO_ESD[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.090000 0.000000 110.350000 17.465000 ;
    END
  END TIE_LO_ESD[0]
  PIN TIE_LO_ESD[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.655000 0.000000 279.915000 17.465000 ;
    END
  END TIE_LO_ESD[1]
  PIN VINREF_DFT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.030000 0.000000 466.670000 49.025000 ;
    END
  END VINREF_DFT
  PIN VOHREF
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.445000 0.000000 419.705000 4.425000 ;
    END
  END VOHREF
  PIN VOH_SEL[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.405000 0.000000 449.665000 83.625000 ;
    END
  END VOH_SEL[0]
  PIN VOH_SEL[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.155000 0.000000 450.415000 236.010000 ;
    END
  END VOH_SEL[1]
  PIN VOH_SEL[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.905000 0.000000 451.165000 236.330000 ;
    END
  END VOH_SEL[2]
  PIN VOUTREF_DFT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.530000 0.000000 465.170000 45.435000 ;
    END
  END VOUTREF_DFT
  PIN VREF_SEL[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.155000 0.000000 453.415000 15.430000 ;
    END
  END VREF_SEL[0]
  PIN VREF_SEL[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.905000 0.000000 454.165000 16.050000 ;
    END
  END VREF_SEL[1]
  PIN VREG_EN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.805000 0.000000 150.065000 28.250000 ;
    END
  END VREG_EN[0]
  PIN VREG_EN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.940000 0.000000 240.200000 28.250000 ;
    END
  END VREG_EN[1]
  PIN VREG_EN_REFGEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.840000 0.000000 445.100000 16.795000 ;
    END
  END VREG_EN_REFGEN
  PIN VTRIP_SEL[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.125000 0.000000 128.385000 10.175000 ;
    END
  END VTRIP_SEL[0]
  PIN VTRIP_SEL[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.620000 0.000000 261.880000 10.175000 ;
    END
  END VTRIP_SEL[1]
  PIN VTRIP_SEL_REFGEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.840000 0.000000 403.100000 22.530000 ;
    END
  END VTRIP_SEL_REFGEN
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000000 62.700000 480.000000 67.150000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000000 55.850000 480.000000 61.100000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000000 68.750000 480.000000 72.000000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000000 73.600000 480.000000 78.050000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000000 117.900000 480.000000 122.150000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000000 90.550000 480.000000 93.800000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000000 95.400000 480.000000 99.850000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000000 79.650000 480.000000 84.100000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000000 112.050000 480.000000 116.300000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000000 85.700000 480.000000 88.950000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT 1.120000 0.130000 477.515000 253.585000 ;
    LAYER met1 ;
      RECT 1.460000 0.070000 477.545000 253.645000 ;
    LAYER met2 ;
      RECT   1.505000   0.000000  84.980000  29.895000 ;
      RECT   1.505000  29.895000 121.175000  46.300000 ;
      RECT   1.505000  46.300000 449.125000  83.905000 ;
      RECT   1.505000  83.905000 449.875000 236.290000 ;
      RECT   1.505000 236.290000 450.625000 236.610000 ;
      RECT   1.505000 236.610000 451.375000 236.930000 ;
      RECT   1.505000 236.930000 478.500000 253.400000 ;
      RECT  86.385000  24.755000 121.175000  29.895000 ;
      RECT  87.375000   0.000000 106.430000   1.630000 ;
      RECT  87.375000   1.630000 109.810000  17.745000 ;
      RECT  87.375000  17.745000 121.175000  24.755000 ;
      RECT 107.250000   0.000000 109.810000   1.630000 ;
      RECT 110.630000   0.000000 121.175000  17.745000 ;
      RECT 121.995000   0.000000 127.845000  10.455000 ;
      RECT 121.995000  10.455000 134.895000  29.230000 ;
      RECT 121.995000  29.230000 135.295000  36.970000 ;
      RECT 121.995000  36.970000 147.335000  45.805000 ;
      RECT 121.995000  45.805000 268.010000  46.300000 ;
      RECT 128.665000   0.000000 134.895000  10.455000 ;
      RECT 136.115000   0.000000 140.920000   2.365000 ;
      RECT 136.115000   2.365000 141.725000   7.250000 ;
      RECT 136.115000   7.250000 142.125000  10.260000 ;
      RECT 136.115000  10.260000 146.935000  27.200000 ;
      RECT 136.115000  27.200000 147.335000  36.970000 ;
      RECT 142.945000   0.000000 146.935000  10.260000 ;
      RECT 148.155000   0.000000 149.525000  28.530000 ;
      RECT 148.155000  28.530000 153.530000  42.375000 ;
      RECT 148.155000  42.375000 241.850000  45.805000 ;
      RECT 150.345000   0.000000 153.530000  28.530000 ;
      RECT 154.350000   0.000000 155.700000  33.505000 ;
      RECT 154.350000  33.505000 235.655000  42.375000 ;
      RECT 156.520000  29.235000 233.485000  33.505000 ;
      RECT 156.920000   0.000000 176.710000  24.100000 ;
      RECT 156.920000  24.100000 233.085000  29.235000 ;
      RECT 179.270000   0.000000 210.735000  24.100000 ;
      RECT 213.295000   0.000000 233.085000  24.100000 ;
      RECT 234.305000   0.000000 235.655000  33.505000 ;
      RECT 236.475000  35.225000 241.850000  42.375000 ;
      RECT 236.875000   0.000000 239.660000   1.910000 ;
      RECT 236.875000   3.330000 239.660000  28.530000 ;
      RECT 236.875000  28.530000 241.850000  35.225000 ;
      RECT 236.920000   1.910000 239.660000   3.330000 ;
      RECT 240.480000   0.000000 241.850000  28.530000 ;
      RECT 242.670000  27.200000 253.890000  36.970000 ;
      RECT 242.670000  36.970000 268.010000  45.805000 ;
      RECT 243.070000   0.000000 247.060000  10.260000 ;
      RECT 243.070000  10.260000 253.890000  27.200000 ;
      RECT 247.880000   7.250000 253.890000  10.260000 ;
      RECT 248.280000   2.365000 253.890000   7.250000 ;
      RECT 249.085000   0.000000 253.890000   2.365000 ;
      RECT 254.710000  29.230000 268.010000  36.970000 ;
      RECT 255.110000   0.000000 261.340000  10.455000 ;
      RECT 255.110000  10.455000 268.010000  29.230000 ;
      RECT 262.160000   0.000000 268.010000  10.455000 ;
      RECT 268.830000   0.000000 279.375000  17.745000 ;
      RECT 268.830000  17.745000 302.630000  24.755000 ;
      RECT 268.830000  24.755000 303.620000  29.895000 ;
      RECT 268.830000  29.895000 449.125000  46.300000 ;
      RECT 280.195000   0.000000 282.755000   1.630000 ;
      RECT 280.195000   1.630000 302.630000  17.745000 ;
      RECT 283.575000   0.000000 302.630000   1.630000 ;
      RECT 305.025000   0.000000 402.560000  22.810000 ;
      RECT 305.025000  22.810000 449.125000  29.895000 ;
      RECT 403.380000   0.000000 404.715000  15.090000 ;
      RECT 403.380000  15.090000 422.410000  22.810000 ;
      RECT 405.535000   0.000000 419.165000   4.705000 ;
      RECT 405.535000   4.705000 422.410000  15.090000 ;
      RECT 419.985000   0.000000 422.410000   4.705000 ;
      RECT 423.230000   0.000000 444.560000  17.075000 ;
      RECT 423.230000  17.075000 449.125000  22.810000 ;
      RECT 445.380000   0.000000 449.125000  17.075000 ;
      RECT 452.195000 234.460000 478.500000 236.930000 ;
      RECT 452.945000  15.710000 453.625000  16.330000 ;
      RECT 452.945000  16.330000 464.250000  45.715000 ;
      RECT 452.945000  45.715000 465.750000  49.305000 ;
      RECT 452.945000  49.305000 478.500000 234.460000 ;
      RECT 454.445000   0.000000 464.250000  16.330000 ;
      RECT 465.450000   0.000000 465.750000  45.715000 ;
      RECT 466.950000   0.000000 478.500000  49.305000 ;
    LAYER met3 ;
      RECT 0.300000 2.255000 479.700000 253.715000 ;
    LAYER met4 ;
      RECT 0.000000  55.750000 480.000000 101.680000 ;
      RECT 0.000000 105.460000 480.000000 106.440000 ;
      RECT 0.000000 110.220000 480.000000 253.715000 ;
    LAYER met5 ;
      RECT   0.000000 101.450000 480.000000 110.450000 ;
      RECT   0.000000 123.750000 480.000000 130.385000 ;
      RECT   0.000000 130.385000 105.590000 196.200000 ;
      RECT   0.000000 196.200000 480.000000 253.715000 ;
      RECT 171.490000 130.385000 218.515000 196.200000 ;
      RECT 284.415000 130.385000 480.000000 196.200000 ;
  END
END sky130_fd_io__top_sio_macro
END LIBRARY
