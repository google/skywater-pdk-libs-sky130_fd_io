/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_IO__TOP_POWER_LVC_WPAD_PP_SYMBOL_V
`define SKY130_FD_IO__TOP_POWER_LVC_WPAD_PP_SYMBOL_V

/**
 * top_power_lvc_wpad: A power pad with an ESD low-voltage clamp.
 *
 * Verilog stub (with power pins) for graphical symbol definition
 * generation.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_io__top_power_lvc_wpad (
           //# {{data|Data Signals}}
           inout P_PAD       ,

           //# {{control|Control Signals}}
           inout AMUXBUS_A   ,
           inout AMUXBUS_B   ,

           //# {{power|Power}}
           inout BDY2_B2B    ,
           inout VSWITCH     ,
           inout P_CORE      ,
           inout VCCD        ,
           inout VCCHIB      ,
           inout VDDA        ,
           inout VDDIO       ,
           inout VDDIO_Q     ,
           inout DRN_LVC1    ,
           inout DRN_LVC2    ,
           inout OGC_LVC     ,
           inout SRC_BDY_LVC1,
           inout SRC_BDY_LVC2,
           inout VSSA        ,
           inout VSSD        ,
           inout VSSIO       ,
           inout VSSIO_Q
       );
endmodule

`default_nettype wire
`endif  // SKY130_FD_IO__TOP_POWER_LVC_WPAD_PP_SYMBOL_V
