# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__overlay_vssio_lvc
  CLASS BLOCK ;
  FOREIGN sky130_fd_io__overlay_vssio_lvc ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  75.00000 BY  198.0000 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.530000 23.850000 0.850000 24.170000 ;
      LAYER met4 ;
        RECT 0.530000 23.850000 0.850000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 24.280000 0.850000 24.600000 ;
      LAYER met4 ;
        RECT 0.530000 24.280000 0.850000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 24.710000 0.850000 25.030000 ;
      LAYER met4 ;
        RECT 0.530000 24.710000 0.850000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 25.140000 0.850000 25.460000 ;
      LAYER met4 ;
        RECT 0.530000 25.140000 0.850000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 25.570000 0.850000 25.890000 ;
      LAYER met4 ;
        RECT 0.530000 25.570000 0.850000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 26.000000 0.850000 26.320000 ;
      LAYER met4 ;
        RECT 0.530000 26.000000 0.850000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 26.430000 0.850000 26.750000 ;
      LAYER met4 ;
        RECT 0.530000 26.430000 0.850000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 26.860000 0.850000 27.180000 ;
      LAYER met4 ;
        RECT 0.530000 26.860000 0.850000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 27.290000 0.850000 27.610000 ;
      LAYER met4 ;
        RECT 0.530000 27.290000 0.850000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 27.720000 0.850000 28.040000 ;
      LAYER met4 ;
        RECT 0.530000 27.720000 0.850000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 28.150000 0.850000 28.470000 ;
      LAYER met4 ;
        RECT 0.530000 28.150000 0.850000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 173.840000 12.875000 181.360000 ;
      LAYER met4 ;
        RECT 0.555000 173.840000 12.875000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 181.445000 0.875000 181.765000 ;
      LAYER met4 ;
        RECT 0.555000 181.445000 0.875000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 181.850000 0.875000 182.170000 ;
      LAYER met4 ;
        RECT 0.555000 181.850000 0.875000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 182.255000 0.875000 182.575000 ;
      LAYER met4 ;
        RECT 0.555000 182.255000 0.875000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 182.660000 0.875000 182.980000 ;
      LAYER met4 ;
        RECT 0.555000 182.660000 0.875000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 183.065000 0.875000 183.385000 ;
      LAYER met4 ;
        RECT 0.555000 183.065000 0.875000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 183.470000 0.875000 183.790000 ;
      LAYER met4 ;
        RECT 0.555000 183.470000 0.875000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 183.875000 0.875000 184.195000 ;
      LAYER met4 ;
        RECT 0.555000 183.875000 0.875000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 184.280000 0.875000 184.600000 ;
      LAYER met4 ;
        RECT 0.555000 184.280000 0.875000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 184.685000 0.875000 185.005000 ;
      LAYER met4 ;
        RECT 0.555000 184.685000 0.875000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 185.090000 0.875000 185.410000 ;
      LAYER met4 ;
        RECT 0.555000 185.090000 0.875000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 185.495000 0.875000 185.815000 ;
      LAYER met4 ;
        RECT 0.555000 185.495000 0.875000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 185.900000 0.875000 186.220000 ;
      LAYER met4 ;
        RECT 0.555000 185.900000 0.875000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 186.305000 0.875000 186.625000 ;
      LAYER met4 ;
        RECT 0.555000 186.305000 0.875000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 186.710000 0.875000 187.030000 ;
      LAYER met4 ;
        RECT 0.555000 186.710000 0.875000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 187.115000 0.875000 187.435000 ;
      LAYER met4 ;
        RECT 0.555000 187.115000 0.875000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 187.520000 0.875000 187.840000 ;
      LAYER met4 ;
        RECT 0.555000 187.520000 0.875000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 187.925000 0.875000 188.245000 ;
      LAYER met4 ;
        RECT 0.555000 187.925000 0.875000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 188.330000 0.875000 188.650000 ;
      LAYER met4 ;
        RECT 0.555000 188.330000 0.875000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 188.735000 0.875000 189.055000 ;
      LAYER met4 ;
        RECT 0.555000 188.735000 0.875000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 189.140000 0.875000 189.460000 ;
      LAYER met4 ;
        RECT 0.555000 189.140000 0.875000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 189.545000 0.875000 189.865000 ;
      LAYER met4 ;
        RECT 0.555000 189.545000 0.875000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 189.950000 0.875000 190.270000 ;
      LAYER met4 ;
        RECT 0.555000 189.950000 0.875000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 190.355000 0.875000 190.675000 ;
      LAYER met4 ;
        RECT 0.555000 190.355000 0.875000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 190.760000 0.875000 191.080000 ;
      LAYER met4 ;
        RECT 0.555000 190.760000 0.875000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 191.165000 0.875000 191.485000 ;
      LAYER met4 ;
        RECT 0.555000 191.165000 0.875000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 191.570000 0.875000 191.890000 ;
      LAYER met4 ;
        RECT 0.555000 191.570000 0.875000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 191.975000 0.875000 192.295000 ;
      LAYER met4 ;
        RECT 0.555000 191.975000 0.875000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 192.380000 0.875000 192.700000 ;
      LAYER met4 ;
        RECT 0.555000 192.380000 0.875000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 192.785000 0.875000 193.105000 ;
      LAYER met4 ;
        RECT 0.555000 192.785000 0.875000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 193.190000 0.875000 193.510000 ;
      LAYER met4 ;
        RECT 0.555000 193.190000 0.875000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 193.595000 0.875000 193.915000 ;
      LAYER met4 ;
        RECT 0.555000 193.595000 0.875000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 194.000000 0.875000 194.320000 ;
      LAYER met4 ;
        RECT 0.555000 194.000000 0.875000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 194.405000 0.875000 194.725000 ;
      LAYER met4 ;
        RECT 0.555000 194.405000 0.875000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 194.810000 0.875000 195.130000 ;
      LAYER met4 ;
        RECT 0.555000 194.810000 0.875000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 195.215000 0.875000 195.535000 ;
      LAYER met4 ;
        RECT 0.555000 195.215000 0.875000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 195.620000 0.875000 195.940000 ;
      LAYER met4 ;
        RECT 0.555000 195.620000 0.875000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 196.025000 0.875000 196.345000 ;
      LAYER met4 ;
        RECT 0.555000 196.025000 0.875000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 196.430000 0.875000 196.750000 ;
      LAYER met4 ;
        RECT 0.555000 196.430000 0.875000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 196.835000 0.875000 197.155000 ;
      LAYER met4 ;
        RECT 0.555000 196.835000 0.875000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 197.240000 0.875000 197.560000 ;
      LAYER met4 ;
        RECT 0.555000 197.240000 0.875000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555000 197.645000 0.875000 197.965000 ;
      LAYER met4 ;
        RECT 0.555000 197.645000 0.875000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.615000 173.900000 0.815000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.615000 174.300000 0.815000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.615000 174.700000 0.815000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.615000 175.100000 0.815000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.615000 175.500000 0.815000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.615000 175.900000 0.815000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.615000 176.300000 0.815000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.615000 176.700000 0.815000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.615000 177.100000 0.815000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.615000 177.500000 0.815000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.615000 177.900000 0.815000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.615000 178.300000 0.815000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.615000 178.700000 0.815000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.615000 179.100000 0.815000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.615000 179.500000 0.815000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.615000 179.900000 0.815000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.615000 180.300000 0.815000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.615000 180.700000 0.815000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.615000 181.100000 0.815000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 23.850000 1.260000 24.170000 ;
      LAYER met4 ;
        RECT 0.940000 23.850000 1.260000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 24.280000 1.260000 24.600000 ;
      LAYER met4 ;
        RECT 0.940000 24.280000 1.260000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 24.710000 1.260000 25.030000 ;
      LAYER met4 ;
        RECT 0.940000 24.710000 1.260000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 25.140000 1.260000 25.460000 ;
      LAYER met4 ;
        RECT 0.940000 25.140000 1.260000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 25.570000 1.260000 25.890000 ;
      LAYER met4 ;
        RECT 0.940000 25.570000 1.260000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 26.000000 1.260000 26.320000 ;
      LAYER met4 ;
        RECT 0.940000 26.000000 1.260000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 26.430000 1.260000 26.750000 ;
      LAYER met4 ;
        RECT 0.940000 26.430000 1.260000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 26.860000 1.260000 27.180000 ;
      LAYER met4 ;
        RECT 0.940000 26.860000 1.260000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 27.290000 1.260000 27.610000 ;
      LAYER met4 ;
        RECT 0.940000 27.290000 1.260000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 27.720000 1.260000 28.040000 ;
      LAYER met4 ;
        RECT 0.940000 27.720000 1.260000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 28.150000 1.260000 28.470000 ;
      LAYER met4 ;
        RECT 0.940000 28.150000 1.260000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 181.445000 1.275000 181.765000 ;
      LAYER met4 ;
        RECT 0.955000 181.445000 1.275000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 181.850000 1.275000 182.170000 ;
      LAYER met4 ;
        RECT 0.955000 181.850000 1.275000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 182.255000 1.275000 182.575000 ;
      LAYER met4 ;
        RECT 0.955000 182.255000 1.275000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 182.660000 1.275000 182.980000 ;
      LAYER met4 ;
        RECT 0.955000 182.660000 1.275000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 183.065000 1.275000 183.385000 ;
      LAYER met4 ;
        RECT 0.955000 183.065000 1.275000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 183.470000 1.275000 183.790000 ;
      LAYER met4 ;
        RECT 0.955000 183.470000 1.275000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 183.875000 1.275000 184.195000 ;
      LAYER met4 ;
        RECT 0.955000 183.875000 1.275000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 184.280000 1.275000 184.600000 ;
      LAYER met4 ;
        RECT 0.955000 184.280000 1.275000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 184.685000 1.275000 185.005000 ;
      LAYER met4 ;
        RECT 0.955000 184.685000 1.275000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 185.090000 1.275000 185.410000 ;
      LAYER met4 ;
        RECT 0.955000 185.090000 1.275000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 185.495000 1.275000 185.815000 ;
      LAYER met4 ;
        RECT 0.955000 185.495000 1.275000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 185.900000 1.275000 186.220000 ;
      LAYER met4 ;
        RECT 0.955000 185.900000 1.275000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 186.305000 1.275000 186.625000 ;
      LAYER met4 ;
        RECT 0.955000 186.305000 1.275000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 186.710000 1.275000 187.030000 ;
      LAYER met4 ;
        RECT 0.955000 186.710000 1.275000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 187.115000 1.275000 187.435000 ;
      LAYER met4 ;
        RECT 0.955000 187.115000 1.275000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 187.520000 1.275000 187.840000 ;
      LAYER met4 ;
        RECT 0.955000 187.520000 1.275000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 187.925000 1.275000 188.245000 ;
      LAYER met4 ;
        RECT 0.955000 187.925000 1.275000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 188.330000 1.275000 188.650000 ;
      LAYER met4 ;
        RECT 0.955000 188.330000 1.275000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 188.735000 1.275000 189.055000 ;
      LAYER met4 ;
        RECT 0.955000 188.735000 1.275000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 189.140000 1.275000 189.460000 ;
      LAYER met4 ;
        RECT 0.955000 189.140000 1.275000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 189.545000 1.275000 189.865000 ;
      LAYER met4 ;
        RECT 0.955000 189.545000 1.275000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 189.950000 1.275000 190.270000 ;
      LAYER met4 ;
        RECT 0.955000 189.950000 1.275000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 190.355000 1.275000 190.675000 ;
      LAYER met4 ;
        RECT 0.955000 190.355000 1.275000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 190.760000 1.275000 191.080000 ;
      LAYER met4 ;
        RECT 0.955000 190.760000 1.275000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 191.165000 1.275000 191.485000 ;
      LAYER met4 ;
        RECT 0.955000 191.165000 1.275000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 191.570000 1.275000 191.890000 ;
      LAYER met4 ;
        RECT 0.955000 191.570000 1.275000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 191.975000 1.275000 192.295000 ;
      LAYER met4 ;
        RECT 0.955000 191.975000 1.275000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 192.380000 1.275000 192.700000 ;
      LAYER met4 ;
        RECT 0.955000 192.380000 1.275000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 192.785000 1.275000 193.105000 ;
      LAYER met4 ;
        RECT 0.955000 192.785000 1.275000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 193.190000 1.275000 193.510000 ;
      LAYER met4 ;
        RECT 0.955000 193.190000 1.275000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 193.595000 1.275000 193.915000 ;
      LAYER met4 ;
        RECT 0.955000 193.595000 1.275000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 194.000000 1.275000 194.320000 ;
      LAYER met4 ;
        RECT 0.955000 194.000000 1.275000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 194.405000 1.275000 194.725000 ;
      LAYER met4 ;
        RECT 0.955000 194.405000 1.275000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 194.810000 1.275000 195.130000 ;
      LAYER met4 ;
        RECT 0.955000 194.810000 1.275000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 195.215000 1.275000 195.535000 ;
      LAYER met4 ;
        RECT 0.955000 195.215000 1.275000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 195.620000 1.275000 195.940000 ;
      LAYER met4 ;
        RECT 0.955000 195.620000 1.275000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 196.025000 1.275000 196.345000 ;
      LAYER met4 ;
        RECT 0.955000 196.025000 1.275000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 196.430000 1.275000 196.750000 ;
      LAYER met4 ;
        RECT 0.955000 196.430000 1.275000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 196.835000 1.275000 197.155000 ;
      LAYER met4 ;
        RECT 0.955000 196.835000 1.275000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 197.240000 1.275000 197.560000 ;
      LAYER met4 ;
        RECT 0.955000 197.240000 1.275000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955000 197.645000 1.275000 197.965000 ;
      LAYER met4 ;
        RECT 0.955000 197.645000 1.275000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.015000 173.900000 1.215000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.015000 174.300000 1.215000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.015000 174.700000 1.215000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.015000 175.100000 1.215000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.015000 175.500000 1.215000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.015000 175.900000 1.215000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.015000 176.300000 1.215000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.015000 176.700000 1.215000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.015000 177.100000 1.215000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.015000 177.500000 1.215000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.015000 177.900000 1.215000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.015000 178.300000 1.215000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.015000 178.700000 1.215000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.015000 179.100000 1.215000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.015000 179.500000 1.215000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.015000 179.900000 1.215000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.015000 180.300000 1.215000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.015000 180.700000 1.215000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.015000 181.100000 1.215000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 23.850000 1.670000 24.170000 ;
      LAYER met4 ;
        RECT 1.350000 23.850000 1.670000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 24.280000 1.670000 24.600000 ;
      LAYER met4 ;
        RECT 1.350000 24.280000 1.670000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 24.710000 1.670000 25.030000 ;
      LAYER met4 ;
        RECT 1.350000 24.710000 1.670000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 25.140000 1.670000 25.460000 ;
      LAYER met4 ;
        RECT 1.350000 25.140000 1.670000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 25.570000 1.670000 25.890000 ;
      LAYER met4 ;
        RECT 1.350000 25.570000 1.670000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 26.000000 1.670000 26.320000 ;
      LAYER met4 ;
        RECT 1.350000 26.000000 1.670000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 26.430000 1.670000 26.750000 ;
      LAYER met4 ;
        RECT 1.350000 26.430000 1.670000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 26.860000 1.670000 27.180000 ;
      LAYER met4 ;
        RECT 1.350000 26.860000 1.670000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 27.290000 1.670000 27.610000 ;
      LAYER met4 ;
        RECT 1.350000 27.290000 1.670000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 27.720000 1.670000 28.040000 ;
      LAYER met4 ;
        RECT 1.350000 27.720000 1.670000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 28.150000 1.670000 28.470000 ;
      LAYER met4 ;
        RECT 1.350000 28.150000 1.670000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 181.445000 1.675000 181.765000 ;
      LAYER met4 ;
        RECT 1.355000 181.445000 1.675000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 181.850000 1.675000 182.170000 ;
      LAYER met4 ;
        RECT 1.355000 181.850000 1.675000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 182.255000 1.675000 182.575000 ;
      LAYER met4 ;
        RECT 1.355000 182.255000 1.675000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 182.660000 1.675000 182.980000 ;
      LAYER met4 ;
        RECT 1.355000 182.660000 1.675000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 183.065000 1.675000 183.385000 ;
      LAYER met4 ;
        RECT 1.355000 183.065000 1.675000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 183.470000 1.675000 183.790000 ;
      LAYER met4 ;
        RECT 1.355000 183.470000 1.675000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 183.875000 1.675000 184.195000 ;
      LAYER met4 ;
        RECT 1.355000 183.875000 1.675000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 184.280000 1.675000 184.600000 ;
      LAYER met4 ;
        RECT 1.355000 184.280000 1.675000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 184.685000 1.675000 185.005000 ;
      LAYER met4 ;
        RECT 1.355000 184.685000 1.675000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 185.090000 1.675000 185.410000 ;
      LAYER met4 ;
        RECT 1.355000 185.090000 1.675000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 185.495000 1.675000 185.815000 ;
      LAYER met4 ;
        RECT 1.355000 185.495000 1.675000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 185.900000 1.675000 186.220000 ;
      LAYER met4 ;
        RECT 1.355000 185.900000 1.675000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 186.305000 1.675000 186.625000 ;
      LAYER met4 ;
        RECT 1.355000 186.305000 1.675000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 186.710000 1.675000 187.030000 ;
      LAYER met4 ;
        RECT 1.355000 186.710000 1.675000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 187.115000 1.675000 187.435000 ;
      LAYER met4 ;
        RECT 1.355000 187.115000 1.675000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 187.520000 1.675000 187.840000 ;
      LAYER met4 ;
        RECT 1.355000 187.520000 1.675000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 187.925000 1.675000 188.245000 ;
      LAYER met4 ;
        RECT 1.355000 187.925000 1.675000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 188.330000 1.675000 188.650000 ;
      LAYER met4 ;
        RECT 1.355000 188.330000 1.675000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 188.735000 1.675000 189.055000 ;
      LAYER met4 ;
        RECT 1.355000 188.735000 1.675000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 189.140000 1.675000 189.460000 ;
      LAYER met4 ;
        RECT 1.355000 189.140000 1.675000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 189.545000 1.675000 189.865000 ;
      LAYER met4 ;
        RECT 1.355000 189.545000 1.675000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 189.950000 1.675000 190.270000 ;
      LAYER met4 ;
        RECT 1.355000 189.950000 1.675000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 190.355000 1.675000 190.675000 ;
      LAYER met4 ;
        RECT 1.355000 190.355000 1.675000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 190.760000 1.675000 191.080000 ;
      LAYER met4 ;
        RECT 1.355000 190.760000 1.675000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 191.165000 1.675000 191.485000 ;
      LAYER met4 ;
        RECT 1.355000 191.165000 1.675000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 191.570000 1.675000 191.890000 ;
      LAYER met4 ;
        RECT 1.355000 191.570000 1.675000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 191.975000 1.675000 192.295000 ;
      LAYER met4 ;
        RECT 1.355000 191.975000 1.675000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 192.380000 1.675000 192.700000 ;
      LAYER met4 ;
        RECT 1.355000 192.380000 1.675000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 192.785000 1.675000 193.105000 ;
      LAYER met4 ;
        RECT 1.355000 192.785000 1.675000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 193.190000 1.675000 193.510000 ;
      LAYER met4 ;
        RECT 1.355000 193.190000 1.675000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 193.595000 1.675000 193.915000 ;
      LAYER met4 ;
        RECT 1.355000 193.595000 1.675000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 194.000000 1.675000 194.320000 ;
      LAYER met4 ;
        RECT 1.355000 194.000000 1.675000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 194.405000 1.675000 194.725000 ;
      LAYER met4 ;
        RECT 1.355000 194.405000 1.675000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 194.810000 1.675000 195.130000 ;
      LAYER met4 ;
        RECT 1.355000 194.810000 1.675000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 195.215000 1.675000 195.535000 ;
      LAYER met4 ;
        RECT 1.355000 195.215000 1.675000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 195.620000 1.675000 195.940000 ;
      LAYER met4 ;
        RECT 1.355000 195.620000 1.675000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 196.025000 1.675000 196.345000 ;
      LAYER met4 ;
        RECT 1.355000 196.025000 1.675000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 196.430000 1.675000 196.750000 ;
      LAYER met4 ;
        RECT 1.355000 196.430000 1.675000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 196.835000 1.675000 197.155000 ;
      LAYER met4 ;
        RECT 1.355000 196.835000 1.675000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 197.240000 1.675000 197.560000 ;
      LAYER met4 ;
        RECT 1.355000 197.240000 1.675000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355000 197.645000 1.675000 197.965000 ;
      LAYER met4 ;
        RECT 1.355000 197.645000 1.675000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.415000 173.900000 1.615000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.415000 174.300000 1.615000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.415000 174.700000 1.615000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.415000 175.100000 1.615000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.415000 175.500000 1.615000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.415000 175.900000 1.615000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.415000 176.300000 1.615000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.415000 176.700000 1.615000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.415000 177.100000 1.615000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.415000 177.500000 1.615000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.415000 177.900000 1.615000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.415000 178.300000 1.615000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.415000 178.700000 1.615000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.415000 179.100000 1.615000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.415000 179.500000 1.615000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.415000 179.900000 1.615000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.415000 180.300000 1.615000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.415000 180.700000 1.615000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.415000 181.100000 1.615000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 181.445000 2.075000 181.765000 ;
      LAYER met4 ;
        RECT 1.755000 181.445000 2.075000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 181.850000 2.075000 182.170000 ;
      LAYER met4 ;
        RECT 1.755000 181.850000 2.075000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 182.255000 2.075000 182.575000 ;
      LAYER met4 ;
        RECT 1.755000 182.255000 2.075000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 182.660000 2.075000 182.980000 ;
      LAYER met4 ;
        RECT 1.755000 182.660000 2.075000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 183.065000 2.075000 183.385000 ;
      LAYER met4 ;
        RECT 1.755000 183.065000 2.075000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 183.470000 2.075000 183.790000 ;
      LAYER met4 ;
        RECT 1.755000 183.470000 2.075000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 183.875000 2.075000 184.195000 ;
      LAYER met4 ;
        RECT 1.755000 183.875000 2.075000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 184.280000 2.075000 184.600000 ;
      LAYER met4 ;
        RECT 1.755000 184.280000 2.075000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 184.685000 2.075000 185.005000 ;
      LAYER met4 ;
        RECT 1.755000 184.685000 2.075000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 185.090000 2.075000 185.410000 ;
      LAYER met4 ;
        RECT 1.755000 185.090000 2.075000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 185.495000 2.075000 185.815000 ;
      LAYER met4 ;
        RECT 1.755000 185.495000 2.075000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 185.900000 2.075000 186.220000 ;
      LAYER met4 ;
        RECT 1.755000 185.900000 2.075000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 186.305000 2.075000 186.625000 ;
      LAYER met4 ;
        RECT 1.755000 186.305000 2.075000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 186.710000 2.075000 187.030000 ;
      LAYER met4 ;
        RECT 1.755000 186.710000 2.075000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 187.115000 2.075000 187.435000 ;
      LAYER met4 ;
        RECT 1.755000 187.115000 2.075000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 187.520000 2.075000 187.840000 ;
      LAYER met4 ;
        RECT 1.755000 187.520000 2.075000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 187.925000 2.075000 188.245000 ;
      LAYER met4 ;
        RECT 1.755000 187.925000 2.075000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 188.330000 2.075000 188.650000 ;
      LAYER met4 ;
        RECT 1.755000 188.330000 2.075000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 188.735000 2.075000 189.055000 ;
      LAYER met4 ;
        RECT 1.755000 188.735000 2.075000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 189.140000 2.075000 189.460000 ;
      LAYER met4 ;
        RECT 1.755000 189.140000 2.075000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 189.545000 2.075000 189.865000 ;
      LAYER met4 ;
        RECT 1.755000 189.545000 2.075000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 189.950000 2.075000 190.270000 ;
      LAYER met4 ;
        RECT 1.755000 189.950000 2.075000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 190.355000 2.075000 190.675000 ;
      LAYER met4 ;
        RECT 1.755000 190.355000 2.075000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 190.760000 2.075000 191.080000 ;
      LAYER met4 ;
        RECT 1.755000 190.760000 2.075000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 191.165000 2.075000 191.485000 ;
      LAYER met4 ;
        RECT 1.755000 191.165000 2.075000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 191.570000 2.075000 191.890000 ;
      LAYER met4 ;
        RECT 1.755000 191.570000 2.075000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 191.975000 2.075000 192.295000 ;
      LAYER met4 ;
        RECT 1.755000 191.975000 2.075000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 192.380000 2.075000 192.700000 ;
      LAYER met4 ;
        RECT 1.755000 192.380000 2.075000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 192.785000 2.075000 193.105000 ;
      LAYER met4 ;
        RECT 1.755000 192.785000 2.075000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 193.190000 2.075000 193.510000 ;
      LAYER met4 ;
        RECT 1.755000 193.190000 2.075000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 193.595000 2.075000 193.915000 ;
      LAYER met4 ;
        RECT 1.755000 193.595000 2.075000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 194.000000 2.075000 194.320000 ;
      LAYER met4 ;
        RECT 1.755000 194.000000 2.075000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 194.405000 2.075000 194.725000 ;
      LAYER met4 ;
        RECT 1.755000 194.405000 2.075000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 194.810000 2.075000 195.130000 ;
      LAYER met4 ;
        RECT 1.755000 194.810000 2.075000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 195.215000 2.075000 195.535000 ;
      LAYER met4 ;
        RECT 1.755000 195.215000 2.075000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 195.620000 2.075000 195.940000 ;
      LAYER met4 ;
        RECT 1.755000 195.620000 2.075000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 196.025000 2.075000 196.345000 ;
      LAYER met4 ;
        RECT 1.755000 196.025000 2.075000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 196.430000 2.075000 196.750000 ;
      LAYER met4 ;
        RECT 1.755000 196.430000 2.075000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 196.835000 2.075000 197.155000 ;
      LAYER met4 ;
        RECT 1.755000 196.835000 2.075000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 197.240000 2.075000 197.560000 ;
      LAYER met4 ;
        RECT 1.755000 197.240000 2.075000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 197.645000 2.075000 197.965000 ;
      LAYER met4 ;
        RECT 1.755000 197.645000 2.075000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 23.850000 2.080000 24.170000 ;
      LAYER met4 ;
        RECT 1.760000 23.850000 2.080000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 24.280000 2.080000 24.600000 ;
      LAYER met4 ;
        RECT 1.760000 24.280000 2.080000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 24.710000 2.080000 25.030000 ;
      LAYER met4 ;
        RECT 1.760000 24.710000 2.080000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 25.140000 2.080000 25.460000 ;
      LAYER met4 ;
        RECT 1.760000 25.140000 2.080000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 25.570000 2.080000 25.890000 ;
      LAYER met4 ;
        RECT 1.760000 25.570000 2.080000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 26.000000 2.080000 26.320000 ;
      LAYER met4 ;
        RECT 1.760000 26.000000 2.080000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 26.430000 2.080000 26.750000 ;
      LAYER met4 ;
        RECT 1.760000 26.430000 2.080000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 26.860000 2.080000 27.180000 ;
      LAYER met4 ;
        RECT 1.760000 26.860000 2.080000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 27.290000 2.080000 27.610000 ;
      LAYER met4 ;
        RECT 1.760000 27.290000 2.080000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 27.720000 2.080000 28.040000 ;
      LAYER met4 ;
        RECT 1.760000 27.720000 2.080000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 28.150000 2.080000 28.470000 ;
      LAYER met4 ;
        RECT 1.760000 28.150000 2.080000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815000 173.900000 2.015000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815000 174.300000 2.015000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815000 174.700000 2.015000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815000 175.100000 2.015000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815000 175.500000 2.015000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815000 175.900000 2.015000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815000 176.300000 2.015000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815000 176.700000 2.015000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815000 177.100000 2.015000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815000 177.500000 2.015000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815000 177.900000 2.015000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815000 178.300000 2.015000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815000 178.700000 2.015000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815000 179.100000 2.015000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815000 179.500000 2.015000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815000 179.900000 2.015000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815000 180.300000 2.015000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815000 180.700000 2.015000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815000 181.100000 2.015000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 181.445000 10.475000 181.765000 ;
      LAYER met4 ;
        RECT 10.155000 181.445000 10.475000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 181.850000 10.475000 182.170000 ;
      LAYER met4 ;
        RECT 10.155000 181.850000 10.475000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 182.255000 10.475000 182.575000 ;
      LAYER met4 ;
        RECT 10.155000 182.255000 10.475000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 182.660000 10.475000 182.980000 ;
      LAYER met4 ;
        RECT 10.155000 182.660000 10.475000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 183.065000 10.475000 183.385000 ;
      LAYER met4 ;
        RECT 10.155000 183.065000 10.475000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 183.470000 10.475000 183.790000 ;
      LAYER met4 ;
        RECT 10.155000 183.470000 10.475000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 183.875000 10.475000 184.195000 ;
      LAYER met4 ;
        RECT 10.155000 183.875000 10.475000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 184.280000 10.475000 184.600000 ;
      LAYER met4 ;
        RECT 10.155000 184.280000 10.475000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 184.685000 10.475000 185.005000 ;
      LAYER met4 ;
        RECT 10.155000 184.685000 10.475000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 185.090000 10.475000 185.410000 ;
      LAYER met4 ;
        RECT 10.155000 185.090000 10.475000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 185.495000 10.475000 185.815000 ;
      LAYER met4 ;
        RECT 10.155000 185.495000 10.475000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 185.900000 10.475000 186.220000 ;
      LAYER met4 ;
        RECT 10.155000 185.900000 10.475000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 186.305000 10.475000 186.625000 ;
      LAYER met4 ;
        RECT 10.155000 186.305000 10.475000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 186.710000 10.475000 187.030000 ;
      LAYER met4 ;
        RECT 10.155000 186.710000 10.475000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 187.115000 10.475000 187.435000 ;
      LAYER met4 ;
        RECT 10.155000 187.115000 10.475000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 187.520000 10.475000 187.840000 ;
      LAYER met4 ;
        RECT 10.155000 187.520000 10.475000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 187.925000 10.475000 188.245000 ;
      LAYER met4 ;
        RECT 10.155000 187.925000 10.475000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 188.330000 10.475000 188.650000 ;
      LAYER met4 ;
        RECT 10.155000 188.330000 10.475000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 188.735000 10.475000 189.055000 ;
      LAYER met4 ;
        RECT 10.155000 188.735000 10.475000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 189.140000 10.475000 189.460000 ;
      LAYER met4 ;
        RECT 10.155000 189.140000 10.475000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 189.545000 10.475000 189.865000 ;
      LAYER met4 ;
        RECT 10.155000 189.545000 10.475000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 189.950000 10.475000 190.270000 ;
      LAYER met4 ;
        RECT 10.155000 189.950000 10.475000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 190.355000 10.475000 190.675000 ;
      LAYER met4 ;
        RECT 10.155000 190.355000 10.475000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 190.760000 10.475000 191.080000 ;
      LAYER met4 ;
        RECT 10.155000 190.760000 10.475000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 191.165000 10.475000 191.485000 ;
      LAYER met4 ;
        RECT 10.155000 191.165000 10.475000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 191.570000 10.475000 191.890000 ;
      LAYER met4 ;
        RECT 10.155000 191.570000 10.475000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 191.975000 10.475000 192.295000 ;
      LAYER met4 ;
        RECT 10.155000 191.975000 10.475000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 192.380000 10.475000 192.700000 ;
      LAYER met4 ;
        RECT 10.155000 192.380000 10.475000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 192.785000 10.475000 193.105000 ;
      LAYER met4 ;
        RECT 10.155000 192.785000 10.475000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 193.190000 10.475000 193.510000 ;
      LAYER met4 ;
        RECT 10.155000 193.190000 10.475000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 193.595000 10.475000 193.915000 ;
      LAYER met4 ;
        RECT 10.155000 193.595000 10.475000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 194.000000 10.475000 194.320000 ;
      LAYER met4 ;
        RECT 10.155000 194.000000 10.475000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 194.405000 10.475000 194.725000 ;
      LAYER met4 ;
        RECT 10.155000 194.405000 10.475000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 194.810000 10.475000 195.130000 ;
      LAYER met4 ;
        RECT 10.155000 194.810000 10.475000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 195.215000 10.475000 195.535000 ;
      LAYER met4 ;
        RECT 10.155000 195.215000 10.475000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 195.620000 10.475000 195.940000 ;
      LAYER met4 ;
        RECT 10.155000 195.620000 10.475000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 196.025000 10.475000 196.345000 ;
      LAYER met4 ;
        RECT 10.155000 196.025000 10.475000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 196.430000 10.475000 196.750000 ;
      LAYER met4 ;
        RECT 10.155000 196.430000 10.475000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 196.835000 10.475000 197.155000 ;
      LAYER met4 ;
        RECT 10.155000 196.835000 10.475000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 197.240000 10.475000 197.560000 ;
      LAYER met4 ;
        RECT 10.155000 197.240000 10.475000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155000 197.645000 10.475000 197.965000 ;
      LAYER met4 ;
        RECT 10.155000 197.645000 10.475000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.215000 173.900000 10.415000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.215000 174.300000 10.415000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.215000 174.700000 10.415000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.215000 175.100000 10.415000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.215000 175.500000 10.415000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.215000 175.900000 10.415000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.215000 176.300000 10.415000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.215000 176.700000 10.415000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.215000 177.100000 10.415000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.215000 177.500000 10.415000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.215000 177.900000 10.415000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.215000 178.300000 10.415000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.215000 178.700000 10.415000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.215000 179.100000 10.415000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.215000 179.500000 10.415000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.215000 179.900000 10.415000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.215000 180.300000 10.415000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.215000 180.700000 10.415000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.215000 181.100000 10.415000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 23.850000 10.600000 24.170000 ;
      LAYER met4 ;
        RECT 10.280000 23.850000 10.600000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 24.280000 10.600000 24.600000 ;
      LAYER met4 ;
        RECT 10.280000 24.280000 10.600000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 24.710000 10.600000 25.030000 ;
      LAYER met4 ;
        RECT 10.280000 24.710000 10.600000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 25.140000 10.600000 25.460000 ;
      LAYER met4 ;
        RECT 10.280000 25.140000 10.600000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 25.570000 10.600000 25.890000 ;
      LAYER met4 ;
        RECT 10.280000 25.570000 10.600000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 26.000000 10.600000 26.320000 ;
      LAYER met4 ;
        RECT 10.280000 26.000000 10.600000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 26.430000 10.600000 26.750000 ;
      LAYER met4 ;
        RECT 10.280000 26.430000 10.600000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 26.860000 10.600000 27.180000 ;
      LAYER met4 ;
        RECT 10.280000 26.860000 10.600000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 27.290000 10.600000 27.610000 ;
      LAYER met4 ;
        RECT 10.280000 27.290000 10.600000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 27.720000 10.600000 28.040000 ;
      LAYER met4 ;
        RECT 10.280000 27.720000 10.600000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 28.150000 10.600000 28.470000 ;
      LAYER met4 ;
        RECT 10.280000 28.150000 10.600000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 181.445000 10.875000 181.765000 ;
      LAYER met4 ;
        RECT 10.555000 181.445000 10.875000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 181.850000 10.875000 182.170000 ;
      LAYER met4 ;
        RECT 10.555000 181.850000 10.875000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 182.255000 10.875000 182.575000 ;
      LAYER met4 ;
        RECT 10.555000 182.255000 10.875000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 182.660000 10.875000 182.980000 ;
      LAYER met4 ;
        RECT 10.555000 182.660000 10.875000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 183.065000 10.875000 183.385000 ;
      LAYER met4 ;
        RECT 10.555000 183.065000 10.875000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 183.470000 10.875000 183.790000 ;
      LAYER met4 ;
        RECT 10.555000 183.470000 10.875000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 183.875000 10.875000 184.195000 ;
      LAYER met4 ;
        RECT 10.555000 183.875000 10.875000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 184.280000 10.875000 184.600000 ;
      LAYER met4 ;
        RECT 10.555000 184.280000 10.875000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 184.685000 10.875000 185.005000 ;
      LAYER met4 ;
        RECT 10.555000 184.685000 10.875000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 185.090000 10.875000 185.410000 ;
      LAYER met4 ;
        RECT 10.555000 185.090000 10.875000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 185.495000 10.875000 185.815000 ;
      LAYER met4 ;
        RECT 10.555000 185.495000 10.875000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 185.900000 10.875000 186.220000 ;
      LAYER met4 ;
        RECT 10.555000 185.900000 10.875000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 186.305000 10.875000 186.625000 ;
      LAYER met4 ;
        RECT 10.555000 186.305000 10.875000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 186.710000 10.875000 187.030000 ;
      LAYER met4 ;
        RECT 10.555000 186.710000 10.875000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 187.115000 10.875000 187.435000 ;
      LAYER met4 ;
        RECT 10.555000 187.115000 10.875000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 187.520000 10.875000 187.840000 ;
      LAYER met4 ;
        RECT 10.555000 187.520000 10.875000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 187.925000 10.875000 188.245000 ;
      LAYER met4 ;
        RECT 10.555000 187.925000 10.875000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 188.330000 10.875000 188.650000 ;
      LAYER met4 ;
        RECT 10.555000 188.330000 10.875000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 188.735000 10.875000 189.055000 ;
      LAYER met4 ;
        RECT 10.555000 188.735000 10.875000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 189.140000 10.875000 189.460000 ;
      LAYER met4 ;
        RECT 10.555000 189.140000 10.875000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 189.545000 10.875000 189.865000 ;
      LAYER met4 ;
        RECT 10.555000 189.545000 10.875000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 189.950000 10.875000 190.270000 ;
      LAYER met4 ;
        RECT 10.555000 189.950000 10.875000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 190.355000 10.875000 190.675000 ;
      LAYER met4 ;
        RECT 10.555000 190.355000 10.875000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 190.760000 10.875000 191.080000 ;
      LAYER met4 ;
        RECT 10.555000 190.760000 10.875000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 191.165000 10.875000 191.485000 ;
      LAYER met4 ;
        RECT 10.555000 191.165000 10.875000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 191.570000 10.875000 191.890000 ;
      LAYER met4 ;
        RECT 10.555000 191.570000 10.875000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 191.975000 10.875000 192.295000 ;
      LAYER met4 ;
        RECT 10.555000 191.975000 10.875000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 192.380000 10.875000 192.700000 ;
      LAYER met4 ;
        RECT 10.555000 192.380000 10.875000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 192.785000 10.875000 193.105000 ;
      LAYER met4 ;
        RECT 10.555000 192.785000 10.875000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 193.190000 10.875000 193.510000 ;
      LAYER met4 ;
        RECT 10.555000 193.190000 10.875000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 193.595000 10.875000 193.915000 ;
      LAYER met4 ;
        RECT 10.555000 193.595000 10.875000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 194.000000 10.875000 194.320000 ;
      LAYER met4 ;
        RECT 10.555000 194.000000 10.875000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 194.405000 10.875000 194.725000 ;
      LAYER met4 ;
        RECT 10.555000 194.405000 10.875000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 194.810000 10.875000 195.130000 ;
      LAYER met4 ;
        RECT 10.555000 194.810000 10.875000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 195.215000 10.875000 195.535000 ;
      LAYER met4 ;
        RECT 10.555000 195.215000 10.875000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 195.620000 10.875000 195.940000 ;
      LAYER met4 ;
        RECT 10.555000 195.620000 10.875000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 196.025000 10.875000 196.345000 ;
      LAYER met4 ;
        RECT 10.555000 196.025000 10.875000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 196.430000 10.875000 196.750000 ;
      LAYER met4 ;
        RECT 10.555000 196.430000 10.875000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 196.835000 10.875000 197.155000 ;
      LAYER met4 ;
        RECT 10.555000 196.835000 10.875000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 197.240000 10.875000 197.560000 ;
      LAYER met4 ;
        RECT 10.555000 197.240000 10.875000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555000 197.645000 10.875000 197.965000 ;
      LAYER met4 ;
        RECT 10.555000 197.645000 10.875000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.615000 173.900000 10.815000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.615000 174.300000 10.815000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.615000 174.700000 10.815000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.615000 175.100000 10.815000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.615000 175.500000 10.815000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.615000 175.900000 10.815000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.615000 176.300000 10.815000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.615000 176.700000 10.815000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.615000 177.100000 10.815000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.615000 177.500000 10.815000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.615000 177.900000 10.815000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.615000 178.300000 10.815000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.615000 178.700000 10.815000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.615000 179.100000 10.815000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.615000 179.500000 10.815000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.615000 179.900000 10.815000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.615000 180.300000 10.815000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.615000 180.700000 10.815000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.615000 181.100000 10.815000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 23.850000 11.005000 24.170000 ;
      LAYER met4 ;
        RECT 10.685000 23.850000 11.005000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 24.280000 11.005000 24.600000 ;
      LAYER met4 ;
        RECT 10.685000 24.280000 11.005000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 24.710000 11.005000 25.030000 ;
      LAYER met4 ;
        RECT 10.685000 24.710000 11.005000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 25.140000 11.005000 25.460000 ;
      LAYER met4 ;
        RECT 10.685000 25.140000 11.005000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 25.570000 11.005000 25.890000 ;
      LAYER met4 ;
        RECT 10.685000 25.570000 11.005000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 26.000000 11.005000 26.320000 ;
      LAYER met4 ;
        RECT 10.685000 26.000000 11.005000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 26.430000 11.005000 26.750000 ;
      LAYER met4 ;
        RECT 10.685000 26.430000 11.005000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 26.860000 11.005000 27.180000 ;
      LAYER met4 ;
        RECT 10.685000 26.860000 11.005000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 27.290000 11.005000 27.610000 ;
      LAYER met4 ;
        RECT 10.685000 27.290000 11.005000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 27.720000 11.005000 28.040000 ;
      LAYER met4 ;
        RECT 10.685000 27.720000 11.005000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 28.150000 11.005000 28.470000 ;
      LAYER met4 ;
        RECT 10.685000 28.150000 11.005000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 181.445000 11.275000 181.765000 ;
      LAYER met4 ;
        RECT 10.955000 181.445000 11.275000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 181.850000 11.275000 182.170000 ;
      LAYER met4 ;
        RECT 10.955000 181.850000 11.275000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 182.255000 11.275000 182.575000 ;
      LAYER met4 ;
        RECT 10.955000 182.255000 11.275000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 182.660000 11.275000 182.980000 ;
      LAYER met4 ;
        RECT 10.955000 182.660000 11.275000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 183.065000 11.275000 183.385000 ;
      LAYER met4 ;
        RECT 10.955000 183.065000 11.275000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 183.470000 11.275000 183.790000 ;
      LAYER met4 ;
        RECT 10.955000 183.470000 11.275000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 183.875000 11.275000 184.195000 ;
      LAYER met4 ;
        RECT 10.955000 183.875000 11.275000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 184.280000 11.275000 184.600000 ;
      LAYER met4 ;
        RECT 10.955000 184.280000 11.275000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 184.685000 11.275000 185.005000 ;
      LAYER met4 ;
        RECT 10.955000 184.685000 11.275000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 185.090000 11.275000 185.410000 ;
      LAYER met4 ;
        RECT 10.955000 185.090000 11.275000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 185.495000 11.275000 185.815000 ;
      LAYER met4 ;
        RECT 10.955000 185.495000 11.275000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 185.900000 11.275000 186.220000 ;
      LAYER met4 ;
        RECT 10.955000 185.900000 11.275000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 186.305000 11.275000 186.625000 ;
      LAYER met4 ;
        RECT 10.955000 186.305000 11.275000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 186.710000 11.275000 187.030000 ;
      LAYER met4 ;
        RECT 10.955000 186.710000 11.275000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 187.115000 11.275000 187.435000 ;
      LAYER met4 ;
        RECT 10.955000 187.115000 11.275000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 187.520000 11.275000 187.840000 ;
      LAYER met4 ;
        RECT 10.955000 187.520000 11.275000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 187.925000 11.275000 188.245000 ;
      LAYER met4 ;
        RECT 10.955000 187.925000 11.275000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 188.330000 11.275000 188.650000 ;
      LAYER met4 ;
        RECT 10.955000 188.330000 11.275000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 188.735000 11.275000 189.055000 ;
      LAYER met4 ;
        RECT 10.955000 188.735000 11.275000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 189.140000 11.275000 189.460000 ;
      LAYER met4 ;
        RECT 10.955000 189.140000 11.275000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 189.545000 11.275000 189.865000 ;
      LAYER met4 ;
        RECT 10.955000 189.545000 11.275000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 189.950000 11.275000 190.270000 ;
      LAYER met4 ;
        RECT 10.955000 189.950000 11.275000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 190.355000 11.275000 190.675000 ;
      LAYER met4 ;
        RECT 10.955000 190.355000 11.275000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 190.760000 11.275000 191.080000 ;
      LAYER met4 ;
        RECT 10.955000 190.760000 11.275000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 191.165000 11.275000 191.485000 ;
      LAYER met4 ;
        RECT 10.955000 191.165000 11.275000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 191.570000 11.275000 191.890000 ;
      LAYER met4 ;
        RECT 10.955000 191.570000 11.275000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 191.975000 11.275000 192.295000 ;
      LAYER met4 ;
        RECT 10.955000 191.975000 11.275000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 192.380000 11.275000 192.700000 ;
      LAYER met4 ;
        RECT 10.955000 192.380000 11.275000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 192.785000 11.275000 193.105000 ;
      LAYER met4 ;
        RECT 10.955000 192.785000 11.275000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 193.190000 11.275000 193.510000 ;
      LAYER met4 ;
        RECT 10.955000 193.190000 11.275000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 193.595000 11.275000 193.915000 ;
      LAYER met4 ;
        RECT 10.955000 193.595000 11.275000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 194.000000 11.275000 194.320000 ;
      LAYER met4 ;
        RECT 10.955000 194.000000 11.275000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 194.405000 11.275000 194.725000 ;
      LAYER met4 ;
        RECT 10.955000 194.405000 11.275000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 194.810000 11.275000 195.130000 ;
      LAYER met4 ;
        RECT 10.955000 194.810000 11.275000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 195.215000 11.275000 195.535000 ;
      LAYER met4 ;
        RECT 10.955000 195.215000 11.275000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 195.620000 11.275000 195.940000 ;
      LAYER met4 ;
        RECT 10.955000 195.620000 11.275000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 196.025000 11.275000 196.345000 ;
      LAYER met4 ;
        RECT 10.955000 196.025000 11.275000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 196.430000 11.275000 196.750000 ;
      LAYER met4 ;
        RECT 10.955000 196.430000 11.275000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 196.835000 11.275000 197.155000 ;
      LAYER met4 ;
        RECT 10.955000 196.835000 11.275000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 197.240000 11.275000 197.560000 ;
      LAYER met4 ;
        RECT 10.955000 197.240000 11.275000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955000 197.645000 11.275000 197.965000 ;
      LAYER met4 ;
        RECT 10.955000 197.645000 11.275000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.015000 173.900000 11.215000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.015000 174.300000 11.215000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.015000 174.700000 11.215000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.015000 175.100000 11.215000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.015000 175.500000 11.215000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.015000 175.900000 11.215000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.015000 176.300000 11.215000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.015000 176.700000 11.215000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.015000 177.100000 11.215000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.015000 177.500000 11.215000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.015000 177.900000 11.215000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.015000 178.300000 11.215000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.015000 178.700000 11.215000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.015000 179.100000 11.215000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.015000 179.500000 11.215000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.015000 179.900000 11.215000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.015000 180.300000 11.215000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.015000 180.700000 11.215000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.015000 181.100000 11.215000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 23.850000 11.410000 24.170000 ;
      LAYER met4 ;
        RECT 11.090000 23.850000 11.410000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 24.280000 11.410000 24.600000 ;
      LAYER met4 ;
        RECT 11.090000 24.280000 11.410000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 24.710000 11.410000 25.030000 ;
      LAYER met4 ;
        RECT 11.090000 24.710000 11.410000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 25.140000 11.410000 25.460000 ;
      LAYER met4 ;
        RECT 11.090000 25.140000 11.410000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 25.570000 11.410000 25.890000 ;
      LAYER met4 ;
        RECT 11.090000 25.570000 11.410000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 26.000000 11.410000 26.320000 ;
      LAYER met4 ;
        RECT 11.090000 26.000000 11.410000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 26.430000 11.410000 26.750000 ;
      LAYER met4 ;
        RECT 11.090000 26.430000 11.410000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 26.860000 11.410000 27.180000 ;
      LAYER met4 ;
        RECT 11.090000 26.860000 11.410000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 27.290000 11.410000 27.610000 ;
      LAYER met4 ;
        RECT 11.090000 27.290000 11.410000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 27.720000 11.410000 28.040000 ;
      LAYER met4 ;
        RECT 11.090000 27.720000 11.410000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 28.150000 11.410000 28.470000 ;
      LAYER met4 ;
        RECT 11.090000 28.150000 11.410000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 181.445000 11.675000 181.765000 ;
      LAYER met4 ;
        RECT 11.355000 181.445000 11.675000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 181.850000 11.675000 182.170000 ;
      LAYER met4 ;
        RECT 11.355000 181.850000 11.675000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 182.255000 11.675000 182.575000 ;
      LAYER met4 ;
        RECT 11.355000 182.255000 11.675000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 182.660000 11.675000 182.980000 ;
      LAYER met4 ;
        RECT 11.355000 182.660000 11.675000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 183.065000 11.675000 183.385000 ;
      LAYER met4 ;
        RECT 11.355000 183.065000 11.675000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 183.470000 11.675000 183.790000 ;
      LAYER met4 ;
        RECT 11.355000 183.470000 11.675000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 183.875000 11.675000 184.195000 ;
      LAYER met4 ;
        RECT 11.355000 183.875000 11.675000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 184.280000 11.675000 184.600000 ;
      LAYER met4 ;
        RECT 11.355000 184.280000 11.675000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 184.685000 11.675000 185.005000 ;
      LAYER met4 ;
        RECT 11.355000 184.685000 11.675000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 185.090000 11.675000 185.410000 ;
      LAYER met4 ;
        RECT 11.355000 185.090000 11.675000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 185.495000 11.675000 185.815000 ;
      LAYER met4 ;
        RECT 11.355000 185.495000 11.675000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 185.900000 11.675000 186.220000 ;
      LAYER met4 ;
        RECT 11.355000 185.900000 11.675000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 186.305000 11.675000 186.625000 ;
      LAYER met4 ;
        RECT 11.355000 186.305000 11.675000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 186.710000 11.675000 187.030000 ;
      LAYER met4 ;
        RECT 11.355000 186.710000 11.675000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 187.115000 11.675000 187.435000 ;
      LAYER met4 ;
        RECT 11.355000 187.115000 11.675000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 187.520000 11.675000 187.840000 ;
      LAYER met4 ;
        RECT 11.355000 187.520000 11.675000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 187.925000 11.675000 188.245000 ;
      LAYER met4 ;
        RECT 11.355000 187.925000 11.675000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 188.330000 11.675000 188.650000 ;
      LAYER met4 ;
        RECT 11.355000 188.330000 11.675000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 188.735000 11.675000 189.055000 ;
      LAYER met4 ;
        RECT 11.355000 188.735000 11.675000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 189.140000 11.675000 189.460000 ;
      LAYER met4 ;
        RECT 11.355000 189.140000 11.675000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 189.545000 11.675000 189.865000 ;
      LAYER met4 ;
        RECT 11.355000 189.545000 11.675000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 189.950000 11.675000 190.270000 ;
      LAYER met4 ;
        RECT 11.355000 189.950000 11.675000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 190.355000 11.675000 190.675000 ;
      LAYER met4 ;
        RECT 11.355000 190.355000 11.675000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 190.760000 11.675000 191.080000 ;
      LAYER met4 ;
        RECT 11.355000 190.760000 11.675000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 191.165000 11.675000 191.485000 ;
      LAYER met4 ;
        RECT 11.355000 191.165000 11.675000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 191.570000 11.675000 191.890000 ;
      LAYER met4 ;
        RECT 11.355000 191.570000 11.675000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 191.975000 11.675000 192.295000 ;
      LAYER met4 ;
        RECT 11.355000 191.975000 11.675000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 192.380000 11.675000 192.700000 ;
      LAYER met4 ;
        RECT 11.355000 192.380000 11.675000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 192.785000 11.675000 193.105000 ;
      LAYER met4 ;
        RECT 11.355000 192.785000 11.675000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 193.190000 11.675000 193.510000 ;
      LAYER met4 ;
        RECT 11.355000 193.190000 11.675000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 193.595000 11.675000 193.915000 ;
      LAYER met4 ;
        RECT 11.355000 193.595000 11.675000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 194.000000 11.675000 194.320000 ;
      LAYER met4 ;
        RECT 11.355000 194.000000 11.675000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 194.405000 11.675000 194.725000 ;
      LAYER met4 ;
        RECT 11.355000 194.405000 11.675000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 194.810000 11.675000 195.130000 ;
      LAYER met4 ;
        RECT 11.355000 194.810000 11.675000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 195.215000 11.675000 195.535000 ;
      LAYER met4 ;
        RECT 11.355000 195.215000 11.675000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 195.620000 11.675000 195.940000 ;
      LAYER met4 ;
        RECT 11.355000 195.620000 11.675000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 196.025000 11.675000 196.345000 ;
      LAYER met4 ;
        RECT 11.355000 196.025000 11.675000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 196.430000 11.675000 196.750000 ;
      LAYER met4 ;
        RECT 11.355000 196.430000 11.675000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 196.835000 11.675000 197.155000 ;
      LAYER met4 ;
        RECT 11.355000 196.835000 11.675000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 197.240000 11.675000 197.560000 ;
      LAYER met4 ;
        RECT 11.355000 197.240000 11.675000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355000 197.645000 11.675000 197.965000 ;
      LAYER met4 ;
        RECT 11.355000 197.645000 11.675000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.415000 173.900000 11.615000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.415000 174.300000 11.615000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.415000 174.700000 11.615000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.415000 175.100000 11.615000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.415000 175.500000 11.615000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.415000 175.900000 11.615000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.415000 176.300000 11.615000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.415000 176.700000 11.615000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.415000 177.100000 11.615000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.415000 177.500000 11.615000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.415000 177.900000 11.615000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.415000 178.300000 11.615000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.415000 178.700000 11.615000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.415000 179.100000 11.615000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.415000 179.500000 11.615000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.415000 179.900000 11.615000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.415000 180.300000 11.615000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.415000 180.700000 11.615000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.415000 181.100000 11.615000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 23.850000 11.815000 24.170000 ;
      LAYER met4 ;
        RECT 11.495000 23.850000 11.815000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 24.280000 11.815000 24.600000 ;
      LAYER met4 ;
        RECT 11.495000 24.280000 11.815000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 24.710000 11.815000 25.030000 ;
      LAYER met4 ;
        RECT 11.495000 24.710000 11.815000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 25.140000 11.815000 25.460000 ;
      LAYER met4 ;
        RECT 11.495000 25.140000 11.815000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 25.570000 11.815000 25.890000 ;
      LAYER met4 ;
        RECT 11.495000 25.570000 11.815000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 26.000000 11.815000 26.320000 ;
      LAYER met4 ;
        RECT 11.495000 26.000000 11.815000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 26.430000 11.815000 26.750000 ;
      LAYER met4 ;
        RECT 11.495000 26.430000 11.815000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 26.860000 11.815000 27.180000 ;
      LAYER met4 ;
        RECT 11.495000 26.860000 11.815000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 27.290000 11.815000 27.610000 ;
      LAYER met4 ;
        RECT 11.495000 27.290000 11.815000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 27.720000 11.815000 28.040000 ;
      LAYER met4 ;
        RECT 11.495000 27.720000 11.815000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 28.150000 11.815000 28.470000 ;
      LAYER met4 ;
        RECT 11.495000 28.150000 11.815000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 181.445000 12.075000 181.765000 ;
      LAYER met4 ;
        RECT 11.755000 181.445000 12.075000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 181.850000 12.075000 182.170000 ;
      LAYER met4 ;
        RECT 11.755000 181.850000 12.075000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 182.255000 12.075000 182.575000 ;
      LAYER met4 ;
        RECT 11.755000 182.255000 12.075000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 182.660000 12.075000 182.980000 ;
      LAYER met4 ;
        RECT 11.755000 182.660000 12.075000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 183.065000 12.075000 183.385000 ;
      LAYER met4 ;
        RECT 11.755000 183.065000 12.075000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 183.470000 12.075000 183.790000 ;
      LAYER met4 ;
        RECT 11.755000 183.470000 12.075000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 183.875000 12.075000 184.195000 ;
      LAYER met4 ;
        RECT 11.755000 183.875000 12.075000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 184.280000 12.075000 184.600000 ;
      LAYER met4 ;
        RECT 11.755000 184.280000 12.075000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 184.685000 12.075000 185.005000 ;
      LAYER met4 ;
        RECT 11.755000 184.685000 12.075000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 185.090000 12.075000 185.410000 ;
      LAYER met4 ;
        RECT 11.755000 185.090000 12.075000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 185.495000 12.075000 185.815000 ;
      LAYER met4 ;
        RECT 11.755000 185.495000 12.075000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 185.900000 12.075000 186.220000 ;
      LAYER met4 ;
        RECT 11.755000 185.900000 12.075000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 186.305000 12.075000 186.625000 ;
      LAYER met4 ;
        RECT 11.755000 186.305000 12.075000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 186.710000 12.075000 187.030000 ;
      LAYER met4 ;
        RECT 11.755000 186.710000 12.075000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 187.115000 12.075000 187.435000 ;
      LAYER met4 ;
        RECT 11.755000 187.115000 12.075000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 187.520000 12.075000 187.840000 ;
      LAYER met4 ;
        RECT 11.755000 187.520000 12.075000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 187.925000 12.075000 188.245000 ;
      LAYER met4 ;
        RECT 11.755000 187.925000 12.075000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 188.330000 12.075000 188.650000 ;
      LAYER met4 ;
        RECT 11.755000 188.330000 12.075000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 188.735000 12.075000 189.055000 ;
      LAYER met4 ;
        RECT 11.755000 188.735000 12.075000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 189.140000 12.075000 189.460000 ;
      LAYER met4 ;
        RECT 11.755000 189.140000 12.075000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 189.545000 12.075000 189.865000 ;
      LAYER met4 ;
        RECT 11.755000 189.545000 12.075000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 189.950000 12.075000 190.270000 ;
      LAYER met4 ;
        RECT 11.755000 189.950000 12.075000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 190.355000 12.075000 190.675000 ;
      LAYER met4 ;
        RECT 11.755000 190.355000 12.075000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 190.760000 12.075000 191.080000 ;
      LAYER met4 ;
        RECT 11.755000 190.760000 12.075000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 191.165000 12.075000 191.485000 ;
      LAYER met4 ;
        RECT 11.755000 191.165000 12.075000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 191.570000 12.075000 191.890000 ;
      LAYER met4 ;
        RECT 11.755000 191.570000 12.075000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 191.975000 12.075000 192.295000 ;
      LAYER met4 ;
        RECT 11.755000 191.975000 12.075000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 192.380000 12.075000 192.700000 ;
      LAYER met4 ;
        RECT 11.755000 192.380000 12.075000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 192.785000 12.075000 193.105000 ;
      LAYER met4 ;
        RECT 11.755000 192.785000 12.075000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 193.190000 12.075000 193.510000 ;
      LAYER met4 ;
        RECT 11.755000 193.190000 12.075000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 193.595000 12.075000 193.915000 ;
      LAYER met4 ;
        RECT 11.755000 193.595000 12.075000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 194.000000 12.075000 194.320000 ;
      LAYER met4 ;
        RECT 11.755000 194.000000 12.075000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 194.405000 12.075000 194.725000 ;
      LAYER met4 ;
        RECT 11.755000 194.405000 12.075000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 194.810000 12.075000 195.130000 ;
      LAYER met4 ;
        RECT 11.755000 194.810000 12.075000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 195.215000 12.075000 195.535000 ;
      LAYER met4 ;
        RECT 11.755000 195.215000 12.075000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 195.620000 12.075000 195.940000 ;
      LAYER met4 ;
        RECT 11.755000 195.620000 12.075000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 196.025000 12.075000 196.345000 ;
      LAYER met4 ;
        RECT 11.755000 196.025000 12.075000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 196.430000 12.075000 196.750000 ;
      LAYER met4 ;
        RECT 11.755000 196.430000 12.075000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 196.835000 12.075000 197.155000 ;
      LAYER met4 ;
        RECT 11.755000 196.835000 12.075000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 197.240000 12.075000 197.560000 ;
      LAYER met4 ;
        RECT 11.755000 197.240000 12.075000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755000 197.645000 12.075000 197.965000 ;
      LAYER met4 ;
        RECT 11.755000 197.645000 12.075000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.815000 173.900000 12.015000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.815000 174.300000 12.015000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.815000 174.700000 12.015000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.815000 175.100000 12.015000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.815000 175.500000 12.015000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.815000 175.900000 12.015000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.815000 176.300000 12.015000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.815000 176.700000 12.015000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.815000 177.100000 12.015000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.815000 177.500000 12.015000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.815000 177.900000 12.015000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.815000 178.300000 12.015000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.815000 178.700000 12.015000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.815000 179.100000 12.015000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.815000 179.500000 12.015000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.815000 179.900000 12.015000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.815000 180.300000 12.015000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.815000 180.700000 12.015000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.815000 181.100000 12.015000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 23.850000 12.220000 24.170000 ;
      LAYER met4 ;
        RECT 11.900000 23.850000 12.220000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 24.280000 12.220000 24.600000 ;
      LAYER met4 ;
        RECT 11.900000 24.280000 12.220000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 24.710000 12.220000 25.030000 ;
      LAYER met4 ;
        RECT 11.900000 24.710000 12.220000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 25.140000 12.220000 25.460000 ;
      LAYER met4 ;
        RECT 11.900000 25.140000 12.220000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 25.570000 12.220000 25.890000 ;
      LAYER met4 ;
        RECT 11.900000 25.570000 12.220000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 26.000000 12.220000 26.320000 ;
      LAYER met4 ;
        RECT 11.900000 26.000000 12.220000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 26.430000 12.220000 26.750000 ;
      LAYER met4 ;
        RECT 11.900000 26.430000 12.220000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 26.860000 12.220000 27.180000 ;
      LAYER met4 ;
        RECT 11.900000 26.860000 12.220000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 27.290000 12.220000 27.610000 ;
      LAYER met4 ;
        RECT 11.900000 27.290000 12.220000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 27.720000 12.220000 28.040000 ;
      LAYER met4 ;
        RECT 11.900000 27.720000 12.220000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 28.150000 12.220000 28.470000 ;
      LAYER met4 ;
        RECT 11.900000 28.150000 12.220000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 181.445000 12.475000 181.765000 ;
      LAYER met4 ;
        RECT 12.155000 181.445000 12.475000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 181.850000 12.475000 182.170000 ;
      LAYER met4 ;
        RECT 12.155000 181.850000 12.475000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 182.255000 12.475000 182.575000 ;
      LAYER met4 ;
        RECT 12.155000 182.255000 12.475000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 182.660000 12.475000 182.980000 ;
      LAYER met4 ;
        RECT 12.155000 182.660000 12.475000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 183.065000 12.475000 183.385000 ;
      LAYER met4 ;
        RECT 12.155000 183.065000 12.475000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 183.470000 12.475000 183.790000 ;
      LAYER met4 ;
        RECT 12.155000 183.470000 12.475000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 183.875000 12.475000 184.195000 ;
      LAYER met4 ;
        RECT 12.155000 183.875000 12.475000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 184.280000 12.475000 184.600000 ;
      LAYER met4 ;
        RECT 12.155000 184.280000 12.475000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 184.685000 12.475000 185.005000 ;
      LAYER met4 ;
        RECT 12.155000 184.685000 12.475000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 185.090000 12.475000 185.410000 ;
      LAYER met4 ;
        RECT 12.155000 185.090000 12.475000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 185.495000 12.475000 185.815000 ;
      LAYER met4 ;
        RECT 12.155000 185.495000 12.475000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 185.900000 12.475000 186.220000 ;
      LAYER met4 ;
        RECT 12.155000 185.900000 12.475000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 186.305000 12.475000 186.625000 ;
      LAYER met4 ;
        RECT 12.155000 186.305000 12.475000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 186.710000 12.475000 187.030000 ;
      LAYER met4 ;
        RECT 12.155000 186.710000 12.475000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 187.115000 12.475000 187.435000 ;
      LAYER met4 ;
        RECT 12.155000 187.115000 12.475000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 187.520000 12.475000 187.840000 ;
      LAYER met4 ;
        RECT 12.155000 187.520000 12.475000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 187.925000 12.475000 188.245000 ;
      LAYER met4 ;
        RECT 12.155000 187.925000 12.475000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 188.330000 12.475000 188.650000 ;
      LAYER met4 ;
        RECT 12.155000 188.330000 12.475000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 188.735000 12.475000 189.055000 ;
      LAYER met4 ;
        RECT 12.155000 188.735000 12.475000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 189.140000 12.475000 189.460000 ;
      LAYER met4 ;
        RECT 12.155000 189.140000 12.475000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 189.545000 12.475000 189.865000 ;
      LAYER met4 ;
        RECT 12.155000 189.545000 12.475000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 189.950000 12.475000 190.270000 ;
      LAYER met4 ;
        RECT 12.155000 189.950000 12.475000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 190.355000 12.475000 190.675000 ;
      LAYER met4 ;
        RECT 12.155000 190.355000 12.475000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 190.760000 12.475000 191.080000 ;
      LAYER met4 ;
        RECT 12.155000 190.760000 12.475000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 191.165000 12.475000 191.485000 ;
      LAYER met4 ;
        RECT 12.155000 191.165000 12.475000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 191.570000 12.475000 191.890000 ;
      LAYER met4 ;
        RECT 12.155000 191.570000 12.475000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 191.975000 12.475000 192.295000 ;
      LAYER met4 ;
        RECT 12.155000 191.975000 12.475000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 192.380000 12.475000 192.700000 ;
      LAYER met4 ;
        RECT 12.155000 192.380000 12.475000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 192.785000 12.475000 193.105000 ;
      LAYER met4 ;
        RECT 12.155000 192.785000 12.475000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 193.190000 12.475000 193.510000 ;
      LAYER met4 ;
        RECT 12.155000 193.190000 12.475000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 193.595000 12.475000 193.915000 ;
      LAYER met4 ;
        RECT 12.155000 193.595000 12.475000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 194.000000 12.475000 194.320000 ;
      LAYER met4 ;
        RECT 12.155000 194.000000 12.475000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 194.405000 12.475000 194.725000 ;
      LAYER met4 ;
        RECT 12.155000 194.405000 12.475000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 194.810000 12.475000 195.130000 ;
      LAYER met4 ;
        RECT 12.155000 194.810000 12.475000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 195.215000 12.475000 195.535000 ;
      LAYER met4 ;
        RECT 12.155000 195.215000 12.475000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 195.620000 12.475000 195.940000 ;
      LAYER met4 ;
        RECT 12.155000 195.620000 12.475000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 196.025000 12.475000 196.345000 ;
      LAYER met4 ;
        RECT 12.155000 196.025000 12.475000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 196.430000 12.475000 196.750000 ;
      LAYER met4 ;
        RECT 12.155000 196.430000 12.475000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 196.835000 12.475000 197.155000 ;
      LAYER met4 ;
        RECT 12.155000 196.835000 12.475000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 197.240000 12.475000 197.560000 ;
      LAYER met4 ;
        RECT 12.155000 197.240000 12.475000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 197.645000 12.475000 197.965000 ;
      LAYER met4 ;
        RECT 12.155000 197.645000 12.475000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.215000 173.900000 12.415000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.215000 174.300000 12.415000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.215000 174.700000 12.415000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.215000 175.100000 12.415000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.215000 175.500000 12.415000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.215000 175.900000 12.415000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.215000 176.300000 12.415000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.215000 176.700000 12.415000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.215000 177.100000 12.415000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.215000 177.500000 12.415000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.215000 177.900000 12.415000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.215000 178.300000 12.415000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.215000 178.700000 12.415000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.215000 179.100000 12.415000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.215000 179.500000 12.415000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.215000 179.900000 12.415000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.215000 180.300000 12.415000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.215000 180.700000 12.415000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.215000 181.100000 12.415000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 23.850000 12.625000 24.170000 ;
      LAYER met4 ;
        RECT 12.305000 23.850000 12.625000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 24.280000 12.625000 24.600000 ;
      LAYER met4 ;
        RECT 12.305000 24.280000 12.625000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 24.710000 12.625000 25.030000 ;
      LAYER met4 ;
        RECT 12.305000 24.710000 12.625000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 25.140000 12.625000 25.460000 ;
      LAYER met4 ;
        RECT 12.305000 25.140000 12.625000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 25.570000 12.625000 25.890000 ;
      LAYER met4 ;
        RECT 12.305000 25.570000 12.625000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 26.000000 12.625000 26.320000 ;
      LAYER met4 ;
        RECT 12.305000 26.000000 12.625000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 26.430000 12.625000 26.750000 ;
      LAYER met4 ;
        RECT 12.305000 26.430000 12.625000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 26.860000 12.625000 27.180000 ;
      LAYER met4 ;
        RECT 12.305000 26.860000 12.625000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 27.290000 12.625000 27.610000 ;
      LAYER met4 ;
        RECT 12.305000 27.290000 12.625000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 27.720000 12.625000 28.040000 ;
      LAYER met4 ;
        RECT 12.305000 27.720000 12.625000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 28.150000 12.625000 28.470000 ;
      LAYER met4 ;
        RECT 12.305000 28.150000 12.625000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 181.445000 12.875000 181.765000 ;
      LAYER met4 ;
        RECT 12.555000 181.445000 12.875000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 181.850000 12.875000 182.170000 ;
      LAYER met4 ;
        RECT 12.555000 181.850000 12.875000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 182.255000 12.875000 182.575000 ;
      LAYER met4 ;
        RECT 12.555000 182.255000 12.875000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 182.660000 12.875000 182.980000 ;
      LAYER met4 ;
        RECT 12.555000 182.660000 12.875000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 183.065000 12.875000 183.385000 ;
      LAYER met4 ;
        RECT 12.555000 183.065000 12.875000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 183.470000 12.875000 183.790000 ;
      LAYER met4 ;
        RECT 12.555000 183.470000 12.875000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 183.875000 12.875000 184.195000 ;
      LAYER met4 ;
        RECT 12.555000 183.875000 12.875000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 184.280000 12.875000 184.600000 ;
      LAYER met4 ;
        RECT 12.555000 184.280000 12.875000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 184.685000 12.875000 185.005000 ;
      LAYER met4 ;
        RECT 12.555000 184.685000 12.875000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 185.090000 12.875000 185.410000 ;
      LAYER met4 ;
        RECT 12.555000 185.090000 12.875000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 185.495000 12.875000 185.815000 ;
      LAYER met4 ;
        RECT 12.555000 185.495000 12.875000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 185.900000 12.875000 186.220000 ;
      LAYER met4 ;
        RECT 12.555000 185.900000 12.875000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 186.305000 12.875000 186.625000 ;
      LAYER met4 ;
        RECT 12.555000 186.305000 12.875000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 186.710000 12.875000 187.030000 ;
      LAYER met4 ;
        RECT 12.555000 186.710000 12.875000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 187.115000 12.875000 187.435000 ;
      LAYER met4 ;
        RECT 12.555000 187.115000 12.875000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 187.520000 12.875000 187.840000 ;
      LAYER met4 ;
        RECT 12.555000 187.520000 12.875000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 187.925000 12.875000 188.245000 ;
      LAYER met4 ;
        RECT 12.555000 187.925000 12.875000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 188.330000 12.875000 188.650000 ;
      LAYER met4 ;
        RECT 12.555000 188.330000 12.875000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 188.735000 12.875000 189.055000 ;
      LAYER met4 ;
        RECT 12.555000 188.735000 12.875000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 189.140000 12.875000 189.460000 ;
      LAYER met4 ;
        RECT 12.555000 189.140000 12.875000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 189.545000 12.875000 189.865000 ;
      LAYER met4 ;
        RECT 12.555000 189.545000 12.875000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 189.950000 12.875000 190.270000 ;
      LAYER met4 ;
        RECT 12.555000 189.950000 12.875000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 190.355000 12.875000 190.675000 ;
      LAYER met4 ;
        RECT 12.555000 190.355000 12.875000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 190.760000 12.875000 191.080000 ;
      LAYER met4 ;
        RECT 12.555000 190.760000 12.875000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 191.165000 12.875000 191.485000 ;
      LAYER met4 ;
        RECT 12.555000 191.165000 12.875000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 191.570000 12.875000 191.890000 ;
      LAYER met4 ;
        RECT 12.555000 191.570000 12.875000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 191.975000 12.875000 192.295000 ;
      LAYER met4 ;
        RECT 12.555000 191.975000 12.875000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 192.380000 12.875000 192.700000 ;
      LAYER met4 ;
        RECT 12.555000 192.380000 12.875000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 192.785000 12.875000 193.105000 ;
      LAYER met4 ;
        RECT 12.555000 192.785000 12.875000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 193.190000 12.875000 193.510000 ;
      LAYER met4 ;
        RECT 12.555000 193.190000 12.875000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 193.595000 12.875000 193.915000 ;
      LAYER met4 ;
        RECT 12.555000 193.595000 12.875000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 194.000000 12.875000 194.320000 ;
      LAYER met4 ;
        RECT 12.555000 194.000000 12.875000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 194.405000 12.875000 194.725000 ;
      LAYER met4 ;
        RECT 12.555000 194.405000 12.875000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 194.810000 12.875000 195.130000 ;
      LAYER met4 ;
        RECT 12.555000 194.810000 12.875000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 195.215000 12.875000 195.535000 ;
      LAYER met4 ;
        RECT 12.555000 195.215000 12.875000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 195.620000 12.875000 195.940000 ;
      LAYER met4 ;
        RECT 12.555000 195.620000 12.875000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 196.025000 12.875000 196.345000 ;
      LAYER met4 ;
        RECT 12.555000 196.025000 12.875000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 196.430000 12.875000 196.750000 ;
      LAYER met4 ;
        RECT 12.555000 196.430000 12.875000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 196.835000 12.875000 197.155000 ;
      LAYER met4 ;
        RECT 12.555000 196.835000 12.875000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 197.240000 12.875000 197.560000 ;
      LAYER met4 ;
        RECT 12.555000 197.240000 12.875000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555000 197.645000 12.875000 197.965000 ;
      LAYER met4 ;
        RECT 12.555000 197.645000 12.875000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.615000 173.900000 12.815000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.615000 174.300000 12.815000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.615000 174.700000 12.815000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.615000 175.100000 12.815000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.615000 175.500000 12.815000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.615000 175.900000 12.815000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.615000 176.300000 12.815000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.615000 176.700000 12.815000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.615000 177.100000 12.815000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.615000 177.500000 12.815000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.615000 177.900000 12.815000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.615000 178.300000 12.815000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.615000 178.700000 12.815000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.615000 179.100000 12.815000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.615000 179.500000 12.815000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.615000 179.900000 12.815000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.615000 180.300000 12.815000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.615000 180.700000 12.815000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 23.850000 13.030000 24.170000 ;
      LAYER met4 ;
        RECT 12.710000 23.850000 13.030000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 24.280000 13.030000 24.600000 ;
      LAYER met4 ;
        RECT 12.710000 24.280000 13.030000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 24.710000 13.030000 25.030000 ;
      LAYER met4 ;
        RECT 12.710000 24.710000 13.030000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 25.140000 13.030000 25.460000 ;
      LAYER met4 ;
        RECT 12.710000 25.140000 13.030000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 25.570000 13.030000 25.890000 ;
      LAYER met4 ;
        RECT 12.710000 25.570000 13.030000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 26.000000 13.030000 26.320000 ;
      LAYER met4 ;
        RECT 12.710000 26.000000 13.030000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 26.430000 13.030000 26.750000 ;
      LAYER met4 ;
        RECT 12.710000 26.430000 13.030000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 26.860000 13.030000 27.180000 ;
      LAYER met4 ;
        RECT 12.710000 26.860000 13.030000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 27.290000 13.030000 27.610000 ;
      LAYER met4 ;
        RECT 12.710000 27.290000 13.030000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 27.720000 13.030000 28.040000 ;
      LAYER met4 ;
        RECT 12.710000 27.720000 13.030000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 28.150000 13.030000 28.470000 ;
      LAYER met4 ;
        RECT 12.710000 28.150000 13.030000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 23.850000 13.435000 24.170000 ;
      LAYER met4 ;
        RECT 13.115000 23.850000 13.435000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 24.280000 13.435000 24.600000 ;
      LAYER met4 ;
        RECT 13.115000 24.280000 13.435000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 24.710000 13.435000 25.030000 ;
      LAYER met4 ;
        RECT 13.115000 24.710000 13.435000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 25.140000 13.435000 25.460000 ;
      LAYER met4 ;
        RECT 13.115000 25.140000 13.435000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 25.570000 13.435000 25.890000 ;
      LAYER met4 ;
        RECT 13.115000 25.570000 13.435000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 26.000000 13.435000 26.320000 ;
      LAYER met4 ;
        RECT 13.115000 26.000000 13.435000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 26.430000 13.435000 26.750000 ;
      LAYER met4 ;
        RECT 13.115000 26.430000 13.435000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 26.860000 13.435000 27.180000 ;
      LAYER met4 ;
        RECT 13.115000 26.860000 13.435000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 27.290000 13.435000 27.610000 ;
      LAYER met4 ;
        RECT 13.115000 27.290000 13.435000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 27.720000 13.435000 28.040000 ;
      LAYER met4 ;
        RECT 13.115000 27.720000 13.435000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 28.150000 13.435000 28.470000 ;
      LAYER met4 ;
        RECT 13.115000 28.150000 13.435000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 23.850000 13.840000 24.170000 ;
      LAYER met4 ;
        RECT 13.520000 23.850000 13.840000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 24.280000 13.840000 24.600000 ;
      LAYER met4 ;
        RECT 13.520000 24.280000 13.840000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 24.710000 13.840000 25.030000 ;
      LAYER met4 ;
        RECT 13.520000 24.710000 13.840000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 25.140000 13.840000 25.460000 ;
      LAYER met4 ;
        RECT 13.520000 25.140000 13.840000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 25.570000 13.840000 25.890000 ;
      LAYER met4 ;
        RECT 13.520000 25.570000 13.840000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 26.000000 13.840000 26.320000 ;
      LAYER met4 ;
        RECT 13.520000 26.000000 13.840000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 26.430000 13.840000 26.750000 ;
      LAYER met4 ;
        RECT 13.520000 26.430000 13.840000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 26.860000 13.840000 27.180000 ;
      LAYER met4 ;
        RECT 13.520000 26.860000 13.840000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 27.290000 13.840000 27.610000 ;
      LAYER met4 ;
        RECT 13.520000 27.290000 13.840000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 27.720000 13.840000 28.040000 ;
      LAYER met4 ;
        RECT 13.520000 27.720000 13.840000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 28.150000 13.840000 28.470000 ;
      LAYER met4 ;
        RECT 13.520000 28.150000 13.840000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 23.850000 14.245000 24.170000 ;
      LAYER met4 ;
        RECT 13.925000 23.850000 14.245000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 24.280000 14.245000 24.600000 ;
      LAYER met4 ;
        RECT 13.925000 24.280000 14.245000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 24.710000 14.245000 25.030000 ;
      LAYER met4 ;
        RECT 13.925000 24.710000 14.245000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 25.140000 14.245000 25.460000 ;
      LAYER met4 ;
        RECT 13.925000 25.140000 14.245000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 25.570000 14.245000 25.890000 ;
      LAYER met4 ;
        RECT 13.925000 25.570000 14.245000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 26.000000 14.245000 26.320000 ;
      LAYER met4 ;
        RECT 13.925000 26.000000 14.245000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 26.430000 14.245000 26.750000 ;
      LAYER met4 ;
        RECT 13.925000 26.430000 14.245000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 26.860000 14.245000 27.180000 ;
      LAYER met4 ;
        RECT 13.925000 26.860000 14.245000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 27.290000 14.245000 27.610000 ;
      LAYER met4 ;
        RECT 13.925000 27.290000 14.245000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 27.720000 14.245000 28.040000 ;
      LAYER met4 ;
        RECT 13.925000 27.720000 14.245000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 28.150000 14.245000 28.470000 ;
      LAYER met4 ;
        RECT 13.925000 28.150000 14.245000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 23.850000 14.650000 24.170000 ;
      LAYER met4 ;
        RECT 14.330000 23.850000 14.650000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 24.280000 14.650000 24.600000 ;
      LAYER met4 ;
        RECT 14.330000 24.280000 14.650000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 24.710000 14.650000 25.030000 ;
      LAYER met4 ;
        RECT 14.330000 24.710000 14.650000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 25.140000 14.650000 25.460000 ;
      LAYER met4 ;
        RECT 14.330000 25.140000 14.650000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 25.570000 14.650000 25.890000 ;
      LAYER met4 ;
        RECT 14.330000 25.570000 14.650000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 26.000000 14.650000 26.320000 ;
      LAYER met4 ;
        RECT 14.330000 26.000000 14.650000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 26.430000 14.650000 26.750000 ;
      LAYER met4 ;
        RECT 14.330000 26.430000 14.650000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 26.860000 14.650000 27.180000 ;
      LAYER met4 ;
        RECT 14.330000 26.860000 14.650000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 27.290000 14.650000 27.610000 ;
      LAYER met4 ;
        RECT 14.330000 27.290000 14.650000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 27.720000 14.650000 28.040000 ;
      LAYER met4 ;
        RECT 14.330000 27.720000 14.650000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 28.150000 14.650000 28.470000 ;
      LAYER met4 ;
        RECT 14.330000 28.150000 14.650000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 23.850000 15.055000 24.170000 ;
      LAYER met4 ;
        RECT 14.735000 23.850000 15.055000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 24.280000 15.055000 24.600000 ;
      LAYER met4 ;
        RECT 14.735000 24.280000 15.055000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 24.710000 15.055000 25.030000 ;
      LAYER met4 ;
        RECT 14.735000 24.710000 15.055000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 25.140000 15.055000 25.460000 ;
      LAYER met4 ;
        RECT 14.735000 25.140000 15.055000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 25.570000 15.055000 25.890000 ;
      LAYER met4 ;
        RECT 14.735000 25.570000 15.055000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 26.000000 15.055000 26.320000 ;
      LAYER met4 ;
        RECT 14.735000 26.000000 15.055000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 26.430000 15.055000 26.750000 ;
      LAYER met4 ;
        RECT 14.735000 26.430000 15.055000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 26.860000 15.055000 27.180000 ;
      LAYER met4 ;
        RECT 14.735000 26.860000 15.055000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 27.290000 15.055000 27.610000 ;
      LAYER met4 ;
        RECT 14.735000 27.290000 15.055000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 27.720000 15.055000 28.040000 ;
      LAYER met4 ;
        RECT 14.735000 27.720000 15.055000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 28.150000 15.055000 28.470000 ;
      LAYER met4 ;
        RECT 14.735000 28.150000 15.055000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 23.850000 15.460000 24.170000 ;
      LAYER met4 ;
        RECT 15.140000 23.850000 15.460000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 24.280000 15.460000 24.600000 ;
      LAYER met4 ;
        RECT 15.140000 24.280000 15.460000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 24.710000 15.460000 25.030000 ;
      LAYER met4 ;
        RECT 15.140000 24.710000 15.460000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 25.140000 15.460000 25.460000 ;
      LAYER met4 ;
        RECT 15.140000 25.140000 15.460000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 25.570000 15.460000 25.890000 ;
      LAYER met4 ;
        RECT 15.140000 25.570000 15.460000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 26.000000 15.460000 26.320000 ;
      LAYER met4 ;
        RECT 15.140000 26.000000 15.460000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 26.430000 15.460000 26.750000 ;
      LAYER met4 ;
        RECT 15.140000 26.430000 15.460000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 26.860000 15.460000 27.180000 ;
      LAYER met4 ;
        RECT 15.140000 26.860000 15.460000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 27.290000 15.460000 27.610000 ;
      LAYER met4 ;
        RECT 15.140000 27.290000 15.460000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 27.720000 15.460000 28.040000 ;
      LAYER met4 ;
        RECT 15.140000 27.720000 15.460000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 28.150000 15.460000 28.470000 ;
      LAYER met4 ;
        RECT 15.140000 28.150000 15.460000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 23.850000 15.865000 24.170000 ;
      LAYER met4 ;
        RECT 15.545000 23.850000 15.865000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 24.280000 15.865000 24.600000 ;
      LAYER met4 ;
        RECT 15.545000 24.280000 15.865000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 24.710000 15.865000 25.030000 ;
      LAYER met4 ;
        RECT 15.545000 24.710000 15.865000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 25.140000 15.865000 25.460000 ;
      LAYER met4 ;
        RECT 15.545000 25.140000 15.865000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 25.570000 15.865000 25.890000 ;
      LAYER met4 ;
        RECT 15.545000 25.570000 15.865000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 26.000000 15.865000 26.320000 ;
      LAYER met4 ;
        RECT 15.545000 26.000000 15.865000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 26.430000 15.865000 26.750000 ;
      LAYER met4 ;
        RECT 15.545000 26.430000 15.865000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 26.860000 15.865000 27.180000 ;
      LAYER met4 ;
        RECT 15.545000 26.860000 15.865000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 27.290000 15.865000 27.610000 ;
      LAYER met4 ;
        RECT 15.545000 27.290000 15.865000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 27.720000 15.865000 28.040000 ;
      LAYER met4 ;
        RECT 15.545000 27.720000 15.865000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 28.150000 15.865000 28.470000 ;
      LAYER met4 ;
        RECT 15.545000 28.150000 15.865000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 23.850000 16.270000 24.170000 ;
      LAYER met4 ;
        RECT 15.950000 23.850000 16.270000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 24.280000 16.270000 24.600000 ;
      LAYER met4 ;
        RECT 15.950000 24.280000 16.270000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 24.710000 16.270000 25.030000 ;
      LAYER met4 ;
        RECT 15.950000 24.710000 16.270000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 25.140000 16.270000 25.460000 ;
      LAYER met4 ;
        RECT 15.950000 25.140000 16.270000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 25.570000 16.270000 25.890000 ;
      LAYER met4 ;
        RECT 15.950000 25.570000 16.270000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 26.000000 16.270000 26.320000 ;
      LAYER met4 ;
        RECT 15.950000 26.000000 16.270000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 26.430000 16.270000 26.750000 ;
      LAYER met4 ;
        RECT 15.950000 26.430000 16.270000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 26.860000 16.270000 27.180000 ;
      LAYER met4 ;
        RECT 15.950000 26.860000 16.270000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 27.290000 16.270000 27.610000 ;
      LAYER met4 ;
        RECT 15.950000 27.290000 16.270000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 27.720000 16.270000 28.040000 ;
      LAYER met4 ;
        RECT 15.950000 27.720000 16.270000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 28.150000 16.270000 28.470000 ;
      LAYER met4 ;
        RECT 15.950000 28.150000 16.270000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 23.850000 16.675000 24.170000 ;
      LAYER met4 ;
        RECT 16.355000 23.850000 16.675000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 24.280000 16.675000 24.600000 ;
      LAYER met4 ;
        RECT 16.355000 24.280000 16.675000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 24.710000 16.675000 25.030000 ;
      LAYER met4 ;
        RECT 16.355000 24.710000 16.675000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 25.140000 16.675000 25.460000 ;
      LAYER met4 ;
        RECT 16.355000 25.140000 16.675000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 25.570000 16.675000 25.890000 ;
      LAYER met4 ;
        RECT 16.355000 25.570000 16.675000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 26.000000 16.675000 26.320000 ;
      LAYER met4 ;
        RECT 16.355000 26.000000 16.675000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 26.430000 16.675000 26.750000 ;
      LAYER met4 ;
        RECT 16.355000 26.430000 16.675000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 26.860000 16.675000 27.180000 ;
      LAYER met4 ;
        RECT 16.355000 26.860000 16.675000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 27.290000 16.675000 27.610000 ;
      LAYER met4 ;
        RECT 16.355000 27.290000 16.675000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 27.720000 16.675000 28.040000 ;
      LAYER met4 ;
        RECT 16.355000 27.720000 16.675000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 28.150000 16.675000 28.470000 ;
      LAYER met4 ;
        RECT 16.355000 28.150000 16.675000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 23.850000 17.080000 24.170000 ;
      LAYER met4 ;
        RECT 16.760000 23.850000 17.080000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 24.280000 17.080000 24.600000 ;
      LAYER met4 ;
        RECT 16.760000 24.280000 17.080000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 24.710000 17.080000 25.030000 ;
      LAYER met4 ;
        RECT 16.760000 24.710000 17.080000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 25.140000 17.080000 25.460000 ;
      LAYER met4 ;
        RECT 16.760000 25.140000 17.080000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 25.570000 17.080000 25.890000 ;
      LAYER met4 ;
        RECT 16.760000 25.570000 17.080000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 26.000000 17.080000 26.320000 ;
      LAYER met4 ;
        RECT 16.760000 26.000000 17.080000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 26.430000 17.080000 26.750000 ;
      LAYER met4 ;
        RECT 16.760000 26.430000 17.080000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 26.860000 17.080000 27.180000 ;
      LAYER met4 ;
        RECT 16.760000 26.860000 17.080000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 27.290000 17.080000 27.610000 ;
      LAYER met4 ;
        RECT 16.760000 27.290000 17.080000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 27.720000 17.080000 28.040000 ;
      LAYER met4 ;
        RECT 16.760000 27.720000 17.080000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 28.150000 17.080000 28.470000 ;
      LAYER met4 ;
        RECT 16.760000 28.150000 17.080000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 23.850000 17.485000 24.170000 ;
      LAYER met4 ;
        RECT 17.165000 23.850000 17.485000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 24.280000 17.485000 24.600000 ;
      LAYER met4 ;
        RECT 17.165000 24.280000 17.485000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 24.710000 17.485000 25.030000 ;
      LAYER met4 ;
        RECT 17.165000 24.710000 17.485000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 25.140000 17.485000 25.460000 ;
      LAYER met4 ;
        RECT 17.165000 25.140000 17.485000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 25.570000 17.485000 25.890000 ;
      LAYER met4 ;
        RECT 17.165000 25.570000 17.485000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 26.000000 17.485000 26.320000 ;
      LAYER met4 ;
        RECT 17.165000 26.000000 17.485000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 26.430000 17.485000 26.750000 ;
      LAYER met4 ;
        RECT 17.165000 26.430000 17.485000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 26.860000 17.485000 27.180000 ;
      LAYER met4 ;
        RECT 17.165000 26.860000 17.485000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 27.290000 17.485000 27.610000 ;
      LAYER met4 ;
        RECT 17.165000 27.290000 17.485000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 27.720000 17.485000 28.040000 ;
      LAYER met4 ;
        RECT 17.165000 27.720000 17.485000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 28.150000 17.485000 28.470000 ;
      LAYER met4 ;
        RECT 17.165000 28.150000 17.485000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 23.850000 17.890000 24.170000 ;
      LAYER met4 ;
        RECT 17.570000 23.850000 17.890000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 24.280000 17.890000 24.600000 ;
      LAYER met4 ;
        RECT 17.570000 24.280000 17.890000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 24.710000 17.890000 25.030000 ;
      LAYER met4 ;
        RECT 17.570000 24.710000 17.890000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 25.140000 17.890000 25.460000 ;
      LAYER met4 ;
        RECT 17.570000 25.140000 17.890000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 25.570000 17.890000 25.890000 ;
      LAYER met4 ;
        RECT 17.570000 25.570000 17.890000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 26.000000 17.890000 26.320000 ;
      LAYER met4 ;
        RECT 17.570000 26.000000 17.890000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 26.430000 17.890000 26.750000 ;
      LAYER met4 ;
        RECT 17.570000 26.430000 17.890000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 26.860000 17.890000 27.180000 ;
      LAYER met4 ;
        RECT 17.570000 26.860000 17.890000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 27.290000 17.890000 27.610000 ;
      LAYER met4 ;
        RECT 17.570000 27.290000 17.890000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 27.720000 17.890000 28.040000 ;
      LAYER met4 ;
        RECT 17.570000 27.720000 17.890000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 28.150000 17.890000 28.470000 ;
      LAYER met4 ;
        RECT 17.570000 28.150000 17.890000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 23.850000 18.295000 24.170000 ;
      LAYER met4 ;
        RECT 17.975000 23.850000 18.295000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 24.280000 18.295000 24.600000 ;
      LAYER met4 ;
        RECT 17.975000 24.280000 18.295000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 24.710000 18.295000 25.030000 ;
      LAYER met4 ;
        RECT 17.975000 24.710000 18.295000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 25.140000 18.295000 25.460000 ;
      LAYER met4 ;
        RECT 17.975000 25.140000 18.295000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 25.570000 18.295000 25.890000 ;
      LAYER met4 ;
        RECT 17.975000 25.570000 18.295000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 26.000000 18.295000 26.320000 ;
      LAYER met4 ;
        RECT 17.975000 26.000000 18.295000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 26.430000 18.295000 26.750000 ;
      LAYER met4 ;
        RECT 17.975000 26.430000 18.295000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 26.860000 18.295000 27.180000 ;
      LAYER met4 ;
        RECT 17.975000 26.860000 18.295000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 27.290000 18.295000 27.610000 ;
      LAYER met4 ;
        RECT 17.975000 27.290000 18.295000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 27.720000 18.295000 28.040000 ;
      LAYER met4 ;
        RECT 17.975000 27.720000 18.295000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 28.150000 18.295000 28.470000 ;
      LAYER met4 ;
        RECT 17.975000 28.150000 18.295000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 23.850000 18.700000 24.170000 ;
      LAYER met4 ;
        RECT 18.380000 23.850000 18.700000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 24.280000 18.700000 24.600000 ;
      LAYER met4 ;
        RECT 18.380000 24.280000 18.700000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 24.710000 18.700000 25.030000 ;
      LAYER met4 ;
        RECT 18.380000 24.710000 18.700000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 25.140000 18.700000 25.460000 ;
      LAYER met4 ;
        RECT 18.380000 25.140000 18.700000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 25.570000 18.700000 25.890000 ;
      LAYER met4 ;
        RECT 18.380000 25.570000 18.700000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 26.000000 18.700000 26.320000 ;
      LAYER met4 ;
        RECT 18.380000 26.000000 18.700000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 26.430000 18.700000 26.750000 ;
      LAYER met4 ;
        RECT 18.380000 26.430000 18.700000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 26.860000 18.700000 27.180000 ;
      LAYER met4 ;
        RECT 18.380000 26.860000 18.700000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 27.290000 18.700000 27.610000 ;
      LAYER met4 ;
        RECT 18.380000 27.290000 18.700000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 27.720000 18.700000 28.040000 ;
      LAYER met4 ;
        RECT 18.380000 27.720000 18.700000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 28.150000 18.700000 28.470000 ;
      LAYER met4 ;
        RECT 18.380000 28.150000 18.700000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 23.850000 19.105000 24.170000 ;
      LAYER met4 ;
        RECT 18.785000 23.850000 19.105000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 24.280000 19.105000 24.600000 ;
      LAYER met4 ;
        RECT 18.785000 24.280000 19.105000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 24.710000 19.105000 25.030000 ;
      LAYER met4 ;
        RECT 18.785000 24.710000 19.105000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 25.140000 19.105000 25.460000 ;
      LAYER met4 ;
        RECT 18.785000 25.140000 19.105000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 25.570000 19.105000 25.890000 ;
      LAYER met4 ;
        RECT 18.785000 25.570000 19.105000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 26.000000 19.105000 26.320000 ;
      LAYER met4 ;
        RECT 18.785000 26.000000 19.105000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 26.430000 19.105000 26.750000 ;
      LAYER met4 ;
        RECT 18.785000 26.430000 19.105000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 26.860000 19.105000 27.180000 ;
      LAYER met4 ;
        RECT 18.785000 26.860000 19.105000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 27.290000 19.105000 27.610000 ;
      LAYER met4 ;
        RECT 18.785000 27.290000 19.105000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 27.720000 19.105000 28.040000 ;
      LAYER met4 ;
        RECT 18.785000 27.720000 19.105000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 28.150000 19.105000 28.470000 ;
      LAYER met4 ;
        RECT 18.785000 28.150000 19.105000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 23.850000 19.510000 24.170000 ;
      LAYER met4 ;
        RECT 19.190000 23.850000 19.510000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 24.280000 19.510000 24.600000 ;
      LAYER met4 ;
        RECT 19.190000 24.280000 19.510000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 24.710000 19.510000 25.030000 ;
      LAYER met4 ;
        RECT 19.190000 24.710000 19.510000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 25.140000 19.510000 25.460000 ;
      LAYER met4 ;
        RECT 19.190000 25.140000 19.510000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 25.570000 19.510000 25.890000 ;
      LAYER met4 ;
        RECT 19.190000 25.570000 19.510000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 26.000000 19.510000 26.320000 ;
      LAYER met4 ;
        RECT 19.190000 26.000000 19.510000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 26.430000 19.510000 26.750000 ;
      LAYER met4 ;
        RECT 19.190000 26.430000 19.510000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 26.860000 19.510000 27.180000 ;
      LAYER met4 ;
        RECT 19.190000 26.860000 19.510000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 27.290000 19.510000 27.610000 ;
      LAYER met4 ;
        RECT 19.190000 27.290000 19.510000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 27.720000 19.510000 28.040000 ;
      LAYER met4 ;
        RECT 19.190000 27.720000 19.510000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 28.150000 19.510000 28.470000 ;
      LAYER met4 ;
        RECT 19.190000 28.150000 19.510000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 23.850000 19.915000 24.170000 ;
      LAYER met4 ;
        RECT 19.595000 23.850000 19.915000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 24.280000 19.915000 24.600000 ;
      LAYER met4 ;
        RECT 19.595000 24.280000 19.915000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 24.710000 19.915000 25.030000 ;
      LAYER met4 ;
        RECT 19.595000 24.710000 19.915000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 25.140000 19.915000 25.460000 ;
      LAYER met4 ;
        RECT 19.595000 25.140000 19.915000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 25.570000 19.915000 25.890000 ;
      LAYER met4 ;
        RECT 19.595000 25.570000 19.915000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 26.000000 19.915000 26.320000 ;
      LAYER met4 ;
        RECT 19.595000 26.000000 19.915000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 26.430000 19.915000 26.750000 ;
      LAYER met4 ;
        RECT 19.595000 26.430000 19.915000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 26.860000 19.915000 27.180000 ;
      LAYER met4 ;
        RECT 19.595000 26.860000 19.915000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 27.290000 19.915000 27.610000 ;
      LAYER met4 ;
        RECT 19.595000 27.290000 19.915000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 27.720000 19.915000 28.040000 ;
      LAYER met4 ;
        RECT 19.595000 27.720000 19.915000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 28.150000 19.915000 28.470000 ;
      LAYER met4 ;
        RECT 19.595000 28.150000 19.915000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 181.445000 2.475000 181.765000 ;
      LAYER met4 ;
        RECT 2.155000 181.445000 2.475000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 181.850000 2.475000 182.170000 ;
      LAYER met4 ;
        RECT 2.155000 181.850000 2.475000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 182.255000 2.475000 182.575000 ;
      LAYER met4 ;
        RECT 2.155000 182.255000 2.475000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 182.660000 2.475000 182.980000 ;
      LAYER met4 ;
        RECT 2.155000 182.660000 2.475000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 183.065000 2.475000 183.385000 ;
      LAYER met4 ;
        RECT 2.155000 183.065000 2.475000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 183.470000 2.475000 183.790000 ;
      LAYER met4 ;
        RECT 2.155000 183.470000 2.475000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 183.875000 2.475000 184.195000 ;
      LAYER met4 ;
        RECT 2.155000 183.875000 2.475000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 184.280000 2.475000 184.600000 ;
      LAYER met4 ;
        RECT 2.155000 184.280000 2.475000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 184.685000 2.475000 185.005000 ;
      LAYER met4 ;
        RECT 2.155000 184.685000 2.475000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 185.090000 2.475000 185.410000 ;
      LAYER met4 ;
        RECT 2.155000 185.090000 2.475000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 185.495000 2.475000 185.815000 ;
      LAYER met4 ;
        RECT 2.155000 185.495000 2.475000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 185.900000 2.475000 186.220000 ;
      LAYER met4 ;
        RECT 2.155000 185.900000 2.475000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 186.305000 2.475000 186.625000 ;
      LAYER met4 ;
        RECT 2.155000 186.305000 2.475000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 186.710000 2.475000 187.030000 ;
      LAYER met4 ;
        RECT 2.155000 186.710000 2.475000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 187.115000 2.475000 187.435000 ;
      LAYER met4 ;
        RECT 2.155000 187.115000 2.475000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 187.520000 2.475000 187.840000 ;
      LAYER met4 ;
        RECT 2.155000 187.520000 2.475000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 187.925000 2.475000 188.245000 ;
      LAYER met4 ;
        RECT 2.155000 187.925000 2.475000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 188.330000 2.475000 188.650000 ;
      LAYER met4 ;
        RECT 2.155000 188.330000 2.475000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 188.735000 2.475000 189.055000 ;
      LAYER met4 ;
        RECT 2.155000 188.735000 2.475000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 189.140000 2.475000 189.460000 ;
      LAYER met4 ;
        RECT 2.155000 189.140000 2.475000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 189.545000 2.475000 189.865000 ;
      LAYER met4 ;
        RECT 2.155000 189.545000 2.475000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 189.950000 2.475000 190.270000 ;
      LAYER met4 ;
        RECT 2.155000 189.950000 2.475000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 190.355000 2.475000 190.675000 ;
      LAYER met4 ;
        RECT 2.155000 190.355000 2.475000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 190.760000 2.475000 191.080000 ;
      LAYER met4 ;
        RECT 2.155000 190.760000 2.475000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 191.165000 2.475000 191.485000 ;
      LAYER met4 ;
        RECT 2.155000 191.165000 2.475000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 191.570000 2.475000 191.890000 ;
      LAYER met4 ;
        RECT 2.155000 191.570000 2.475000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 191.975000 2.475000 192.295000 ;
      LAYER met4 ;
        RECT 2.155000 191.975000 2.475000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 192.380000 2.475000 192.700000 ;
      LAYER met4 ;
        RECT 2.155000 192.380000 2.475000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 192.785000 2.475000 193.105000 ;
      LAYER met4 ;
        RECT 2.155000 192.785000 2.475000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 193.190000 2.475000 193.510000 ;
      LAYER met4 ;
        RECT 2.155000 193.190000 2.475000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 193.595000 2.475000 193.915000 ;
      LAYER met4 ;
        RECT 2.155000 193.595000 2.475000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 194.000000 2.475000 194.320000 ;
      LAYER met4 ;
        RECT 2.155000 194.000000 2.475000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 194.405000 2.475000 194.725000 ;
      LAYER met4 ;
        RECT 2.155000 194.405000 2.475000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 194.810000 2.475000 195.130000 ;
      LAYER met4 ;
        RECT 2.155000 194.810000 2.475000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 195.215000 2.475000 195.535000 ;
      LAYER met4 ;
        RECT 2.155000 195.215000 2.475000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 195.620000 2.475000 195.940000 ;
      LAYER met4 ;
        RECT 2.155000 195.620000 2.475000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 196.025000 2.475000 196.345000 ;
      LAYER met4 ;
        RECT 2.155000 196.025000 2.475000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 196.430000 2.475000 196.750000 ;
      LAYER met4 ;
        RECT 2.155000 196.430000 2.475000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 196.835000 2.475000 197.155000 ;
      LAYER met4 ;
        RECT 2.155000 196.835000 2.475000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 197.240000 2.475000 197.560000 ;
      LAYER met4 ;
        RECT 2.155000 197.240000 2.475000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155000 197.645000 2.475000 197.965000 ;
      LAYER met4 ;
        RECT 2.155000 197.645000 2.475000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 23.850000 2.490000 24.170000 ;
      LAYER met4 ;
        RECT 2.170000 23.850000 2.490000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 24.280000 2.490000 24.600000 ;
      LAYER met4 ;
        RECT 2.170000 24.280000 2.490000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 24.710000 2.490000 25.030000 ;
      LAYER met4 ;
        RECT 2.170000 24.710000 2.490000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 25.140000 2.490000 25.460000 ;
      LAYER met4 ;
        RECT 2.170000 25.140000 2.490000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 25.570000 2.490000 25.890000 ;
      LAYER met4 ;
        RECT 2.170000 25.570000 2.490000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 26.000000 2.490000 26.320000 ;
      LAYER met4 ;
        RECT 2.170000 26.000000 2.490000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 26.430000 2.490000 26.750000 ;
      LAYER met4 ;
        RECT 2.170000 26.430000 2.490000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 26.860000 2.490000 27.180000 ;
      LAYER met4 ;
        RECT 2.170000 26.860000 2.490000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 27.290000 2.490000 27.610000 ;
      LAYER met4 ;
        RECT 2.170000 27.290000 2.490000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 27.720000 2.490000 28.040000 ;
      LAYER met4 ;
        RECT 2.170000 27.720000 2.490000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 28.150000 2.490000 28.470000 ;
      LAYER met4 ;
        RECT 2.170000 28.150000 2.490000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 173.900000 2.415000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 174.300000 2.415000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 174.700000 2.415000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 175.100000 2.415000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 175.500000 2.415000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 175.900000 2.415000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 176.300000 2.415000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 176.700000 2.415000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 177.100000 2.415000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 177.500000 2.415000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 177.900000 2.415000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 178.300000 2.415000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 178.700000 2.415000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 179.100000 2.415000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 179.500000 2.415000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 179.900000 2.415000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 180.300000 2.415000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 180.700000 2.415000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 181.100000 2.415000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 181.445000 2.875000 181.765000 ;
      LAYER met4 ;
        RECT 2.555000 181.445000 2.875000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 181.850000 2.875000 182.170000 ;
      LAYER met4 ;
        RECT 2.555000 181.850000 2.875000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 182.255000 2.875000 182.575000 ;
      LAYER met4 ;
        RECT 2.555000 182.255000 2.875000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 182.660000 2.875000 182.980000 ;
      LAYER met4 ;
        RECT 2.555000 182.660000 2.875000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 183.065000 2.875000 183.385000 ;
      LAYER met4 ;
        RECT 2.555000 183.065000 2.875000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 183.470000 2.875000 183.790000 ;
      LAYER met4 ;
        RECT 2.555000 183.470000 2.875000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 183.875000 2.875000 184.195000 ;
      LAYER met4 ;
        RECT 2.555000 183.875000 2.875000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 184.280000 2.875000 184.600000 ;
      LAYER met4 ;
        RECT 2.555000 184.280000 2.875000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 184.685000 2.875000 185.005000 ;
      LAYER met4 ;
        RECT 2.555000 184.685000 2.875000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 185.090000 2.875000 185.410000 ;
      LAYER met4 ;
        RECT 2.555000 185.090000 2.875000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 185.495000 2.875000 185.815000 ;
      LAYER met4 ;
        RECT 2.555000 185.495000 2.875000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 185.900000 2.875000 186.220000 ;
      LAYER met4 ;
        RECT 2.555000 185.900000 2.875000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 186.305000 2.875000 186.625000 ;
      LAYER met4 ;
        RECT 2.555000 186.305000 2.875000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 186.710000 2.875000 187.030000 ;
      LAYER met4 ;
        RECT 2.555000 186.710000 2.875000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 187.115000 2.875000 187.435000 ;
      LAYER met4 ;
        RECT 2.555000 187.115000 2.875000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 187.520000 2.875000 187.840000 ;
      LAYER met4 ;
        RECT 2.555000 187.520000 2.875000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 187.925000 2.875000 188.245000 ;
      LAYER met4 ;
        RECT 2.555000 187.925000 2.875000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 188.330000 2.875000 188.650000 ;
      LAYER met4 ;
        RECT 2.555000 188.330000 2.875000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 188.735000 2.875000 189.055000 ;
      LAYER met4 ;
        RECT 2.555000 188.735000 2.875000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 189.140000 2.875000 189.460000 ;
      LAYER met4 ;
        RECT 2.555000 189.140000 2.875000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 189.545000 2.875000 189.865000 ;
      LAYER met4 ;
        RECT 2.555000 189.545000 2.875000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 189.950000 2.875000 190.270000 ;
      LAYER met4 ;
        RECT 2.555000 189.950000 2.875000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 190.355000 2.875000 190.675000 ;
      LAYER met4 ;
        RECT 2.555000 190.355000 2.875000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 190.760000 2.875000 191.080000 ;
      LAYER met4 ;
        RECT 2.555000 190.760000 2.875000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 191.165000 2.875000 191.485000 ;
      LAYER met4 ;
        RECT 2.555000 191.165000 2.875000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 191.570000 2.875000 191.890000 ;
      LAYER met4 ;
        RECT 2.555000 191.570000 2.875000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 191.975000 2.875000 192.295000 ;
      LAYER met4 ;
        RECT 2.555000 191.975000 2.875000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 192.380000 2.875000 192.700000 ;
      LAYER met4 ;
        RECT 2.555000 192.380000 2.875000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 192.785000 2.875000 193.105000 ;
      LAYER met4 ;
        RECT 2.555000 192.785000 2.875000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 193.190000 2.875000 193.510000 ;
      LAYER met4 ;
        RECT 2.555000 193.190000 2.875000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 193.595000 2.875000 193.915000 ;
      LAYER met4 ;
        RECT 2.555000 193.595000 2.875000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 194.000000 2.875000 194.320000 ;
      LAYER met4 ;
        RECT 2.555000 194.000000 2.875000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 194.405000 2.875000 194.725000 ;
      LAYER met4 ;
        RECT 2.555000 194.405000 2.875000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 194.810000 2.875000 195.130000 ;
      LAYER met4 ;
        RECT 2.555000 194.810000 2.875000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 195.215000 2.875000 195.535000 ;
      LAYER met4 ;
        RECT 2.555000 195.215000 2.875000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 195.620000 2.875000 195.940000 ;
      LAYER met4 ;
        RECT 2.555000 195.620000 2.875000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 196.025000 2.875000 196.345000 ;
      LAYER met4 ;
        RECT 2.555000 196.025000 2.875000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 196.430000 2.875000 196.750000 ;
      LAYER met4 ;
        RECT 2.555000 196.430000 2.875000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 196.835000 2.875000 197.155000 ;
      LAYER met4 ;
        RECT 2.555000 196.835000 2.875000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 197.240000 2.875000 197.560000 ;
      LAYER met4 ;
        RECT 2.555000 197.240000 2.875000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555000 197.645000 2.875000 197.965000 ;
      LAYER met4 ;
        RECT 2.555000 197.645000 2.875000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 23.850000 2.900000 24.170000 ;
      LAYER met4 ;
        RECT 2.580000 23.850000 2.900000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 24.280000 2.900000 24.600000 ;
      LAYER met4 ;
        RECT 2.580000 24.280000 2.900000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 24.710000 2.900000 25.030000 ;
      LAYER met4 ;
        RECT 2.580000 24.710000 2.900000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 25.140000 2.900000 25.460000 ;
      LAYER met4 ;
        RECT 2.580000 25.140000 2.900000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 25.570000 2.900000 25.890000 ;
      LAYER met4 ;
        RECT 2.580000 25.570000 2.900000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 26.000000 2.900000 26.320000 ;
      LAYER met4 ;
        RECT 2.580000 26.000000 2.900000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 26.430000 2.900000 26.750000 ;
      LAYER met4 ;
        RECT 2.580000 26.430000 2.900000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 26.860000 2.900000 27.180000 ;
      LAYER met4 ;
        RECT 2.580000 26.860000 2.900000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 27.290000 2.900000 27.610000 ;
      LAYER met4 ;
        RECT 2.580000 27.290000 2.900000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 27.720000 2.900000 28.040000 ;
      LAYER met4 ;
        RECT 2.580000 27.720000 2.900000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 28.150000 2.900000 28.470000 ;
      LAYER met4 ;
        RECT 2.580000 28.150000 2.900000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.615000 173.900000 2.815000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.615000 174.300000 2.815000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.615000 174.700000 2.815000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.615000 175.100000 2.815000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.615000 175.500000 2.815000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.615000 175.900000 2.815000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.615000 176.300000 2.815000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.615000 176.700000 2.815000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.615000 177.100000 2.815000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.615000 177.500000 2.815000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.615000 177.900000 2.815000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.615000 178.300000 2.815000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.615000 178.700000 2.815000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.615000 179.100000 2.815000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.615000 179.500000 2.815000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.615000 179.900000 2.815000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.615000 180.300000 2.815000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.615000 180.700000 2.815000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.615000 181.100000 2.815000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 181.445000 3.275000 181.765000 ;
      LAYER met4 ;
        RECT 2.955000 181.445000 3.275000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 181.850000 3.275000 182.170000 ;
      LAYER met4 ;
        RECT 2.955000 181.850000 3.275000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 182.255000 3.275000 182.575000 ;
      LAYER met4 ;
        RECT 2.955000 182.255000 3.275000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 182.660000 3.275000 182.980000 ;
      LAYER met4 ;
        RECT 2.955000 182.660000 3.275000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 183.065000 3.275000 183.385000 ;
      LAYER met4 ;
        RECT 2.955000 183.065000 3.275000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 183.470000 3.275000 183.790000 ;
      LAYER met4 ;
        RECT 2.955000 183.470000 3.275000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 183.875000 3.275000 184.195000 ;
      LAYER met4 ;
        RECT 2.955000 183.875000 3.275000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 184.280000 3.275000 184.600000 ;
      LAYER met4 ;
        RECT 2.955000 184.280000 3.275000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 184.685000 3.275000 185.005000 ;
      LAYER met4 ;
        RECT 2.955000 184.685000 3.275000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 185.090000 3.275000 185.410000 ;
      LAYER met4 ;
        RECT 2.955000 185.090000 3.275000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 185.495000 3.275000 185.815000 ;
      LAYER met4 ;
        RECT 2.955000 185.495000 3.275000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 185.900000 3.275000 186.220000 ;
      LAYER met4 ;
        RECT 2.955000 185.900000 3.275000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 186.305000 3.275000 186.625000 ;
      LAYER met4 ;
        RECT 2.955000 186.305000 3.275000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 186.710000 3.275000 187.030000 ;
      LAYER met4 ;
        RECT 2.955000 186.710000 3.275000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 187.115000 3.275000 187.435000 ;
      LAYER met4 ;
        RECT 2.955000 187.115000 3.275000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 187.520000 3.275000 187.840000 ;
      LAYER met4 ;
        RECT 2.955000 187.520000 3.275000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 187.925000 3.275000 188.245000 ;
      LAYER met4 ;
        RECT 2.955000 187.925000 3.275000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 188.330000 3.275000 188.650000 ;
      LAYER met4 ;
        RECT 2.955000 188.330000 3.275000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 188.735000 3.275000 189.055000 ;
      LAYER met4 ;
        RECT 2.955000 188.735000 3.275000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 189.140000 3.275000 189.460000 ;
      LAYER met4 ;
        RECT 2.955000 189.140000 3.275000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 189.545000 3.275000 189.865000 ;
      LAYER met4 ;
        RECT 2.955000 189.545000 3.275000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 189.950000 3.275000 190.270000 ;
      LAYER met4 ;
        RECT 2.955000 189.950000 3.275000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 190.355000 3.275000 190.675000 ;
      LAYER met4 ;
        RECT 2.955000 190.355000 3.275000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 190.760000 3.275000 191.080000 ;
      LAYER met4 ;
        RECT 2.955000 190.760000 3.275000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 191.165000 3.275000 191.485000 ;
      LAYER met4 ;
        RECT 2.955000 191.165000 3.275000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 191.570000 3.275000 191.890000 ;
      LAYER met4 ;
        RECT 2.955000 191.570000 3.275000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 191.975000 3.275000 192.295000 ;
      LAYER met4 ;
        RECT 2.955000 191.975000 3.275000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 192.380000 3.275000 192.700000 ;
      LAYER met4 ;
        RECT 2.955000 192.380000 3.275000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 192.785000 3.275000 193.105000 ;
      LAYER met4 ;
        RECT 2.955000 192.785000 3.275000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 193.190000 3.275000 193.510000 ;
      LAYER met4 ;
        RECT 2.955000 193.190000 3.275000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 193.595000 3.275000 193.915000 ;
      LAYER met4 ;
        RECT 2.955000 193.595000 3.275000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 194.000000 3.275000 194.320000 ;
      LAYER met4 ;
        RECT 2.955000 194.000000 3.275000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 194.405000 3.275000 194.725000 ;
      LAYER met4 ;
        RECT 2.955000 194.405000 3.275000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 194.810000 3.275000 195.130000 ;
      LAYER met4 ;
        RECT 2.955000 194.810000 3.275000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 195.215000 3.275000 195.535000 ;
      LAYER met4 ;
        RECT 2.955000 195.215000 3.275000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 195.620000 3.275000 195.940000 ;
      LAYER met4 ;
        RECT 2.955000 195.620000 3.275000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 196.025000 3.275000 196.345000 ;
      LAYER met4 ;
        RECT 2.955000 196.025000 3.275000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 196.430000 3.275000 196.750000 ;
      LAYER met4 ;
        RECT 2.955000 196.430000 3.275000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 196.835000 3.275000 197.155000 ;
      LAYER met4 ;
        RECT 2.955000 196.835000 3.275000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 197.240000 3.275000 197.560000 ;
      LAYER met4 ;
        RECT 2.955000 197.240000 3.275000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955000 197.645000 3.275000 197.965000 ;
      LAYER met4 ;
        RECT 2.955000 197.645000 3.275000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 23.850000 3.310000 24.170000 ;
      LAYER met4 ;
        RECT 2.990000 23.850000 3.310000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 24.280000 3.310000 24.600000 ;
      LAYER met4 ;
        RECT 2.990000 24.280000 3.310000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 24.710000 3.310000 25.030000 ;
      LAYER met4 ;
        RECT 2.990000 24.710000 3.310000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 25.140000 3.310000 25.460000 ;
      LAYER met4 ;
        RECT 2.990000 25.140000 3.310000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 25.570000 3.310000 25.890000 ;
      LAYER met4 ;
        RECT 2.990000 25.570000 3.310000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 26.000000 3.310000 26.320000 ;
      LAYER met4 ;
        RECT 2.990000 26.000000 3.310000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 26.430000 3.310000 26.750000 ;
      LAYER met4 ;
        RECT 2.990000 26.430000 3.310000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 26.860000 3.310000 27.180000 ;
      LAYER met4 ;
        RECT 2.990000 26.860000 3.310000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 27.290000 3.310000 27.610000 ;
      LAYER met4 ;
        RECT 2.990000 27.290000 3.310000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 27.720000 3.310000 28.040000 ;
      LAYER met4 ;
        RECT 2.990000 27.720000 3.310000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 28.150000 3.310000 28.470000 ;
      LAYER met4 ;
        RECT 2.990000 28.150000 3.310000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 23.850000 20.320000 24.170000 ;
      LAYER met4 ;
        RECT 20.000000 23.850000 20.320000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 24.280000 20.320000 24.600000 ;
      LAYER met4 ;
        RECT 20.000000 24.280000 20.320000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 24.710000 20.320000 25.030000 ;
      LAYER met4 ;
        RECT 20.000000 24.710000 20.320000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 25.140000 20.320000 25.460000 ;
      LAYER met4 ;
        RECT 20.000000 25.140000 20.320000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 25.570000 20.320000 25.890000 ;
      LAYER met4 ;
        RECT 20.000000 25.570000 20.320000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 26.000000 20.320000 26.320000 ;
      LAYER met4 ;
        RECT 20.000000 26.000000 20.320000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 26.430000 20.320000 26.750000 ;
      LAYER met4 ;
        RECT 20.000000 26.430000 20.320000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 26.860000 20.320000 27.180000 ;
      LAYER met4 ;
        RECT 20.000000 26.860000 20.320000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 27.290000 20.320000 27.610000 ;
      LAYER met4 ;
        RECT 20.000000 27.290000 20.320000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 27.720000 20.320000 28.040000 ;
      LAYER met4 ;
        RECT 20.000000 27.720000 20.320000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 28.150000 20.320000 28.470000 ;
      LAYER met4 ;
        RECT 20.000000 28.150000 20.320000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 23.850000 20.725000 24.170000 ;
      LAYER met4 ;
        RECT 20.405000 23.850000 20.725000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 24.280000 20.725000 24.600000 ;
      LAYER met4 ;
        RECT 20.405000 24.280000 20.725000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 24.710000 20.725000 25.030000 ;
      LAYER met4 ;
        RECT 20.405000 24.710000 20.725000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 25.140000 20.725000 25.460000 ;
      LAYER met4 ;
        RECT 20.405000 25.140000 20.725000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 25.570000 20.725000 25.890000 ;
      LAYER met4 ;
        RECT 20.405000 25.570000 20.725000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 26.000000 20.725000 26.320000 ;
      LAYER met4 ;
        RECT 20.405000 26.000000 20.725000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 26.430000 20.725000 26.750000 ;
      LAYER met4 ;
        RECT 20.405000 26.430000 20.725000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 26.860000 20.725000 27.180000 ;
      LAYER met4 ;
        RECT 20.405000 26.860000 20.725000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 27.290000 20.725000 27.610000 ;
      LAYER met4 ;
        RECT 20.405000 27.290000 20.725000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 27.720000 20.725000 28.040000 ;
      LAYER met4 ;
        RECT 20.405000 27.720000 20.725000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 28.150000 20.725000 28.470000 ;
      LAYER met4 ;
        RECT 20.405000 28.150000 20.725000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 23.850000 21.130000 24.170000 ;
      LAYER met4 ;
        RECT 20.810000 23.850000 21.130000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 24.280000 21.130000 24.600000 ;
      LAYER met4 ;
        RECT 20.810000 24.280000 21.130000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 24.710000 21.130000 25.030000 ;
      LAYER met4 ;
        RECT 20.810000 24.710000 21.130000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 25.140000 21.130000 25.460000 ;
      LAYER met4 ;
        RECT 20.810000 25.140000 21.130000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 25.570000 21.130000 25.890000 ;
      LAYER met4 ;
        RECT 20.810000 25.570000 21.130000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 26.000000 21.130000 26.320000 ;
      LAYER met4 ;
        RECT 20.810000 26.000000 21.130000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 26.430000 21.130000 26.750000 ;
      LAYER met4 ;
        RECT 20.810000 26.430000 21.130000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 26.860000 21.130000 27.180000 ;
      LAYER met4 ;
        RECT 20.810000 26.860000 21.130000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 27.290000 21.130000 27.610000 ;
      LAYER met4 ;
        RECT 20.810000 27.290000 21.130000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 27.720000 21.130000 28.040000 ;
      LAYER met4 ;
        RECT 20.810000 27.720000 21.130000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 28.150000 21.130000 28.470000 ;
      LAYER met4 ;
        RECT 20.810000 28.150000 21.130000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 23.850000 21.535000 24.170000 ;
      LAYER met4 ;
        RECT 21.215000 23.850000 21.535000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 24.280000 21.535000 24.600000 ;
      LAYER met4 ;
        RECT 21.215000 24.280000 21.535000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 24.710000 21.535000 25.030000 ;
      LAYER met4 ;
        RECT 21.215000 24.710000 21.535000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 25.140000 21.535000 25.460000 ;
      LAYER met4 ;
        RECT 21.215000 25.140000 21.535000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 25.570000 21.535000 25.890000 ;
      LAYER met4 ;
        RECT 21.215000 25.570000 21.535000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 26.000000 21.535000 26.320000 ;
      LAYER met4 ;
        RECT 21.215000 26.000000 21.535000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 26.430000 21.535000 26.750000 ;
      LAYER met4 ;
        RECT 21.215000 26.430000 21.535000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 26.860000 21.535000 27.180000 ;
      LAYER met4 ;
        RECT 21.215000 26.860000 21.535000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 27.290000 21.535000 27.610000 ;
      LAYER met4 ;
        RECT 21.215000 27.290000 21.535000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 27.720000 21.535000 28.040000 ;
      LAYER met4 ;
        RECT 21.215000 27.720000 21.535000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 28.150000 21.535000 28.470000 ;
      LAYER met4 ;
        RECT 21.215000 28.150000 21.535000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 23.850000 21.940000 24.170000 ;
      LAYER met4 ;
        RECT 21.620000 23.850000 21.940000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 24.280000 21.940000 24.600000 ;
      LAYER met4 ;
        RECT 21.620000 24.280000 21.940000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 24.710000 21.940000 25.030000 ;
      LAYER met4 ;
        RECT 21.620000 24.710000 21.940000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 25.140000 21.940000 25.460000 ;
      LAYER met4 ;
        RECT 21.620000 25.140000 21.940000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 25.570000 21.940000 25.890000 ;
      LAYER met4 ;
        RECT 21.620000 25.570000 21.940000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 26.000000 21.940000 26.320000 ;
      LAYER met4 ;
        RECT 21.620000 26.000000 21.940000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 26.430000 21.940000 26.750000 ;
      LAYER met4 ;
        RECT 21.620000 26.430000 21.940000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 26.860000 21.940000 27.180000 ;
      LAYER met4 ;
        RECT 21.620000 26.860000 21.940000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 27.290000 21.940000 27.610000 ;
      LAYER met4 ;
        RECT 21.620000 27.290000 21.940000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 27.720000 21.940000 28.040000 ;
      LAYER met4 ;
        RECT 21.620000 27.720000 21.940000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 28.150000 21.940000 28.470000 ;
      LAYER met4 ;
        RECT 21.620000 28.150000 21.940000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 23.850000 22.345000 24.170000 ;
      LAYER met4 ;
        RECT 22.025000 23.850000 22.345000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 24.280000 22.345000 24.600000 ;
      LAYER met4 ;
        RECT 22.025000 24.280000 22.345000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 24.710000 22.345000 25.030000 ;
      LAYER met4 ;
        RECT 22.025000 24.710000 22.345000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 25.140000 22.345000 25.460000 ;
      LAYER met4 ;
        RECT 22.025000 25.140000 22.345000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 25.570000 22.345000 25.890000 ;
      LAYER met4 ;
        RECT 22.025000 25.570000 22.345000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 26.000000 22.345000 26.320000 ;
      LAYER met4 ;
        RECT 22.025000 26.000000 22.345000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 26.430000 22.345000 26.750000 ;
      LAYER met4 ;
        RECT 22.025000 26.430000 22.345000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 26.860000 22.345000 27.180000 ;
      LAYER met4 ;
        RECT 22.025000 26.860000 22.345000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 27.290000 22.345000 27.610000 ;
      LAYER met4 ;
        RECT 22.025000 27.290000 22.345000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 27.720000 22.345000 28.040000 ;
      LAYER met4 ;
        RECT 22.025000 27.720000 22.345000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 28.150000 22.345000 28.470000 ;
      LAYER met4 ;
        RECT 22.025000 28.150000 22.345000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 23.850000 22.750000 24.170000 ;
      LAYER met4 ;
        RECT 22.430000 23.850000 22.750000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 24.280000 22.750000 24.600000 ;
      LAYER met4 ;
        RECT 22.430000 24.280000 22.750000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 24.710000 22.750000 25.030000 ;
      LAYER met4 ;
        RECT 22.430000 24.710000 22.750000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 25.140000 22.750000 25.460000 ;
      LAYER met4 ;
        RECT 22.430000 25.140000 22.750000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 25.570000 22.750000 25.890000 ;
      LAYER met4 ;
        RECT 22.430000 25.570000 22.750000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 26.000000 22.750000 26.320000 ;
      LAYER met4 ;
        RECT 22.430000 26.000000 22.750000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 26.430000 22.750000 26.750000 ;
      LAYER met4 ;
        RECT 22.430000 26.430000 22.750000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 26.860000 22.750000 27.180000 ;
      LAYER met4 ;
        RECT 22.430000 26.860000 22.750000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 27.290000 22.750000 27.610000 ;
      LAYER met4 ;
        RECT 22.430000 27.290000 22.750000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 27.720000 22.750000 28.040000 ;
      LAYER met4 ;
        RECT 22.430000 27.720000 22.750000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 28.150000 22.750000 28.470000 ;
      LAYER met4 ;
        RECT 22.430000 28.150000 22.750000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 23.850000 23.155000 24.170000 ;
      LAYER met4 ;
        RECT 22.835000 23.850000 23.155000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 24.280000 23.155000 24.600000 ;
      LAYER met4 ;
        RECT 22.835000 24.280000 23.155000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 24.710000 23.155000 25.030000 ;
      LAYER met4 ;
        RECT 22.835000 24.710000 23.155000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 25.140000 23.155000 25.460000 ;
      LAYER met4 ;
        RECT 22.835000 25.140000 23.155000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 25.570000 23.155000 25.890000 ;
      LAYER met4 ;
        RECT 22.835000 25.570000 23.155000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 26.000000 23.155000 26.320000 ;
      LAYER met4 ;
        RECT 22.835000 26.000000 23.155000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 26.430000 23.155000 26.750000 ;
      LAYER met4 ;
        RECT 22.835000 26.430000 23.155000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 26.860000 23.155000 27.180000 ;
      LAYER met4 ;
        RECT 22.835000 26.860000 23.155000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 27.290000 23.155000 27.610000 ;
      LAYER met4 ;
        RECT 22.835000 27.290000 23.155000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 27.720000 23.155000 28.040000 ;
      LAYER met4 ;
        RECT 22.835000 27.720000 23.155000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 28.150000 23.155000 28.470000 ;
      LAYER met4 ;
        RECT 22.835000 28.150000 23.155000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 23.850000 23.560000 24.170000 ;
      LAYER met4 ;
        RECT 23.240000 23.850000 23.560000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 24.280000 23.560000 24.600000 ;
      LAYER met4 ;
        RECT 23.240000 24.280000 23.560000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 24.710000 23.560000 25.030000 ;
      LAYER met4 ;
        RECT 23.240000 24.710000 23.560000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 25.140000 23.560000 25.460000 ;
      LAYER met4 ;
        RECT 23.240000 25.140000 23.560000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 25.570000 23.560000 25.890000 ;
      LAYER met4 ;
        RECT 23.240000 25.570000 23.560000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 26.000000 23.560000 26.320000 ;
      LAYER met4 ;
        RECT 23.240000 26.000000 23.560000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 26.430000 23.560000 26.750000 ;
      LAYER met4 ;
        RECT 23.240000 26.430000 23.560000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 26.860000 23.560000 27.180000 ;
      LAYER met4 ;
        RECT 23.240000 26.860000 23.560000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 27.290000 23.560000 27.610000 ;
      LAYER met4 ;
        RECT 23.240000 27.290000 23.560000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 27.720000 23.560000 28.040000 ;
      LAYER met4 ;
        RECT 23.240000 27.720000 23.560000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 28.150000 23.560000 28.470000 ;
      LAYER met4 ;
        RECT 23.240000 28.150000 23.560000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 23.850000 23.965000 24.170000 ;
      LAYER met4 ;
        RECT 23.645000 23.850000 23.965000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 24.280000 23.965000 24.600000 ;
      LAYER met4 ;
        RECT 23.645000 24.280000 23.965000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 24.710000 23.965000 25.030000 ;
      LAYER met4 ;
        RECT 23.645000 24.710000 23.965000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 25.140000 23.965000 25.460000 ;
      LAYER met4 ;
        RECT 23.645000 25.140000 23.965000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 25.570000 23.965000 25.890000 ;
      LAYER met4 ;
        RECT 23.645000 25.570000 23.965000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 26.000000 23.965000 26.320000 ;
      LAYER met4 ;
        RECT 23.645000 26.000000 23.965000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 26.430000 23.965000 26.750000 ;
      LAYER met4 ;
        RECT 23.645000 26.430000 23.965000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 26.860000 23.965000 27.180000 ;
      LAYER met4 ;
        RECT 23.645000 26.860000 23.965000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 27.290000 23.965000 27.610000 ;
      LAYER met4 ;
        RECT 23.645000 27.290000 23.965000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 27.720000 23.965000 28.040000 ;
      LAYER met4 ;
        RECT 23.645000 27.720000 23.965000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 28.150000 23.965000 28.470000 ;
      LAYER met4 ;
        RECT 23.645000 28.150000 23.965000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 23.850000 24.370000 24.170000 ;
      LAYER met4 ;
        RECT 24.050000 23.850000 24.370000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 24.280000 24.370000 24.600000 ;
      LAYER met4 ;
        RECT 24.050000 24.280000 24.370000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 24.710000 24.370000 25.030000 ;
      LAYER met4 ;
        RECT 24.050000 24.710000 24.370000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 25.140000 24.370000 25.460000 ;
      LAYER met4 ;
        RECT 24.050000 25.140000 24.370000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 25.570000 24.370000 25.890000 ;
      LAYER met4 ;
        RECT 24.050000 25.570000 24.370000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 26.000000 24.370000 26.320000 ;
      LAYER met4 ;
        RECT 24.050000 26.000000 24.370000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 26.430000 24.370000 26.750000 ;
      LAYER met4 ;
        RECT 24.050000 26.430000 24.370000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 26.860000 24.370000 27.180000 ;
      LAYER met4 ;
        RECT 24.050000 26.860000 24.370000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 27.290000 24.370000 27.610000 ;
      LAYER met4 ;
        RECT 24.050000 27.290000 24.370000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 27.720000 24.370000 28.040000 ;
      LAYER met4 ;
        RECT 24.050000 27.720000 24.370000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 28.150000 24.370000 28.470000 ;
      LAYER met4 ;
        RECT 24.050000 28.150000 24.370000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.015000 173.900000 3.215000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.015000 174.300000 3.215000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.015000 174.700000 3.215000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.015000 175.100000 3.215000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.015000 175.500000 3.215000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.015000 175.900000 3.215000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.015000 176.300000 3.215000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.015000 176.700000 3.215000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.015000 177.100000 3.215000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.015000 177.500000 3.215000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.015000 177.900000 3.215000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.015000 178.300000 3.215000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.015000 178.700000 3.215000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.015000 179.100000 3.215000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.015000 179.500000 3.215000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.015000 179.900000 3.215000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.015000 180.300000 3.215000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.015000 180.700000 3.215000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.015000 181.100000 3.215000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 181.445000 3.675000 181.765000 ;
      LAYER met4 ;
        RECT 3.355000 181.445000 3.675000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 181.850000 3.675000 182.170000 ;
      LAYER met4 ;
        RECT 3.355000 181.850000 3.675000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 182.255000 3.675000 182.575000 ;
      LAYER met4 ;
        RECT 3.355000 182.255000 3.675000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 182.660000 3.675000 182.980000 ;
      LAYER met4 ;
        RECT 3.355000 182.660000 3.675000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 183.065000 3.675000 183.385000 ;
      LAYER met4 ;
        RECT 3.355000 183.065000 3.675000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 183.470000 3.675000 183.790000 ;
      LAYER met4 ;
        RECT 3.355000 183.470000 3.675000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 183.875000 3.675000 184.195000 ;
      LAYER met4 ;
        RECT 3.355000 183.875000 3.675000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 184.280000 3.675000 184.600000 ;
      LAYER met4 ;
        RECT 3.355000 184.280000 3.675000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 184.685000 3.675000 185.005000 ;
      LAYER met4 ;
        RECT 3.355000 184.685000 3.675000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 185.090000 3.675000 185.410000 ;
      LAYER met4 ;
        RECT 3.355000 185.090000 3.675000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 185.495000 3.675000 185.815000 ;
      LAYER met4 ;
        RECT 3.355000 185.495000 3.675000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 185.900000 3.675000 186.220000 ;
      LAYER met4 ;
        RECT 3.355000 185.900000 3.675000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 186.305000 3.675000 186.625000 ;
      LAYER met4 ;
        RECT 3.355000 186.305000 3.675000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 186.710000 3.675000 187.030000 ;
      LAYER met4 ;
        RECT 3.355000 186.710000 3.675000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 187.115000 3.675000 187.435000 ;
      LAYER met4 ;
        RECT 3.355000 187.115000 3.675000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 187.520000 3.675000 187.840000 ;
      LAYER met4 ;
        RECT 3.355000 187.520000 3.675000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 187.925000 3.675000 188.245000 ;
      LAYER met4 ;
        RECT 3.355000 187.925000 3.675000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 188.330000 3.675000 188.650000 ;
      LAYER met4 ;
        RECT 3.355000 188.330000 3.675000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 188.735000 3.675000 189.055000 ;
      LAYER met4 ;
        RECT 3.355000 188.735000 3.675000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 189.140000 3.675000 189.460000 ;
      LAYER met4 ;
        RECT 3.355000 189.140000 3.675000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 189.545000 3.675000 189.865000 ;
      LAYER met4 ;
        RECT 3.355000 189.545000 3.675000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 189.950000 3.675000 190.270000 ;
      LAYER met4 ;
        RECT 3.355000 189.950000 3.675000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 190.355000 3.675000 190.675000 ;
      LAYER met4 ;
        RECT 3.355000 190.355000 3.675000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 190.760000 3.675000 191.080000 ;
      LAYER met4 ;
        RECT 3.355000 190.760000 3.675000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 191.165000 3.675000 191.485000 ;
      LAYER met4 ;
        RECT 3.355000 191.165000 3.675000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 191.570000 3.675000 191.890000 ;
      LAYER met4 ;
        RECT 3.355000 191.570000 3.675000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 191.975000 3.675000 192.295000 ;
      LAYER met4 ;
        RECT 3.355000 191.975000 3.675000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 192.380000 3.675000 192.700000 ;
      LAYER met4 ;
        RECT 3.355000 192.380000 3.675000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 192.785000 3.675000 193.105000 ;
      LAYER met4 ;
        RECT 3.355000 192.785000 3.675000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 193.190000 3.675000 193.510000 ;
      LAYER met4 ;
        RECT 3.355000 193.190000 3.675000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 193.595000 3.675000 193.915000 ;
      LAYER met4 ;
        RECT 3.355000 193.595000 3.675000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 194.000000 3.675000 194.320000 ;
      LAYER met4 ;
        RECT 3.355000 194.000000 3.675000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 194.405000 3.675000 194.725000 ;
      LAYER met4 ;
        RECT 3.355000 194.405000 3.675000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 194.810000 3.675000 195.130000 ;
      LAYER met4 ;
        RECT 3.355000 194.810000 3.675000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 195.215000 3.675000 195.535000 ;
      LAYER met4 ;
        RECT 3.355000 195.215000 3.675000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 195.620000 3.675000 195.940000 ;
      LAYER met4 ;
        RECT 3.355000 195.620000 3.675000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 196.025000 3.675000 196.345000 ;
      LAYER met4 ;
        RECT 3.355000 196.025000 3.675000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 196.430000 3.675000 196.750000 ;
      LAYER met4 ;
        RECT 3.355000 196.430000 3.675000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 196.835000 3.675000 197.155000 ;
      LAYER met4 ;
        RECT 3.355000 196.835000 3.675000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 197.240000 3.675000 197.560000 ;
      LAYER met4 ;
        RECT 3.355000 197.240000 3.675000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355000 197.645000 3.675000 197.965000 ;
      LAYER met4 ;
        RECT 3.355000 197.645000 3.675000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 23.850000 3.715000 24.170000 ;
      LAYER met4 ;
        RECT 3.395000 23.850000 3.715000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 24.280000 3.715000 24.600000 ;
      LAYER met4 ;
        RECT 3.395000 24.280000 3.715000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 24.710000 3.715000 25.030000 ;
      LAYER met4 ;
        RECT 3.395000 24.710000 3.715000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 25.140000 3.715000 25.460000 ;
      LAYER met4 ;
        RECT 3.395000 25.140000 3.715000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 25.570000 3.715000 25.890000 ;
      LAYER met4 ;
        RECT 3.395000 25.570000 3.715000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 26.000000 3.715000 26.320000 ;
      LAYER met4 ;
        RECT 3.395000 26.000000 3.715000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 26.430000 3.715000 26.750000 ;
      LAYER met4 ;
        RECT 3.395000 26.430000 3.715000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 26.860000 3.715000 27.180000 ;
      LAYER met4 ;
        RECT 3.395000 26.860000 3.715000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 27.290000 3.715000 27.610000 ;
      LAYER met4 ;
        RECT 3.395000 27.290000 3.715000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 27.720000 3.715000 28.040000 ;
      LAYER met4 ;
        RECT 3.395000 27.720000 3.715000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 28.150000 3.715000 28.470000 ;
      LAYER met4 ;
        RECT 3.395000 28.150000 3.715000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.415000 173.900000 3.615000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.415000 174.300000 3.615000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.415000 174.700000 3.615000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.415000 175.100000 3.615000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.415000 175.500000 3.615000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.415000 175.900000 3.615000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.415000 176.300000 3.615000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.415000 176.700000 3.615000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.415000 177.100000 3.615000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.415000 177.500000 3.615000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.415000 177.900000 3.615000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.415000 178.300000 3.615000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.415000 178.700000 3.615000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.415000 179.100000 3.615000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.415000 179.500000 3.615000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.415000 179.900000 3.615000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.415000 180.300000 3.615000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.415000 180.700000 3.615000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.415000 181.100000 3.615000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 181.445000 4.075000 181.765000 ;
      LAYER met4 ;
        RECT 3.755000 181.445000 4.075000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 181.850000 4.075000 182.170000 ;
      LAYER met4 ;
        RECT 3.755000 181.850000 4.075000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 182.255000 4.075000 182.575000 ;
      LAYER met4 ;
        RECT 3.755000 182.255000 4.075000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 182.660000 4.075000 182.980000 ;
      LAYER met4 ;
        RECT 3.755000 182.660000 4.075000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 183.065000 4.075000 183.385000 ;
      LAYER met4 ;
        RECT 3.755000 183.065000 4.075000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 183.470000 4.075000 183.790000 ;
      LAYER met4 ;
        RECT 3.755000 183.470000 4.075000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 183.875000 4.075000 184.195000 ;
      LAYER met4 ;
        RECT 3.755000 183.875000 4.075000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 184.280000 4.075000 184.600000 ;
      LAYER met4 ;
        RECT 3.755000 184.280000 4.075000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 184.685000 4.075000 185.005000 ;
      LAYER met4 ;
        RECT 3.755000 184.685000 4.075000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 185.090000 4.075000 185.410000 ;
      LAYER met4 ;
        RECT 3.755000 185.090000 4.075000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 185.495000 4.075000 185.815000 ;
      LAYER met4 ;
        RECT 3.755000 185.495000 4.075000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 185.900000 4.075000 186.220000 ;
      LAYER met4 ;
        RECT 3.755000 185.900000 4.075000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 186.305000 4.075000 186.625000 ;
      LAYER met4 ;
        RECT 3.755000 186.305000 4.075000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 186.710000 4.075000 187.030000 ;
      LAYER met4 ;
        RECT 3.755000 186.710000 4.075000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 187.115000 4.075000 187.435000 ;
      LAYER met4 ;
        RECT 3.755000 187.115000 4.075000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 187.520000 4.075000 187.840000 ;
      LAYER met4 ;
        RECT 3.755000 187.520000 4.075000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 187.925000 4.075000 188.245000 ;
      LAYER met4 ;
        RECT 3.755000 187.925000 4.075000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 188.330000 4.075000 188.650000 ;
      LAYER met4 ;
        RECT 3.755000 188.330000 4.075000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 188.735000 4.075000 189.055000 ;
      LAYER met4 ;
        RECT 3.755000 188.735000 4.075000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 189.140000 4.075000 189.460000 ;
      LAYER met4 ;
        RECT 3.755000 189.140000 4.075000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 189.545000 4.075000 189.865000 ;
      LAYER met4 ;
        RECT 3.755000 189.545000 4.075000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 189.950000 4.075000 190.270000 ;
      LAYER met4 ;
        RECT 3.755000 189.950000 4.075000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 190.355000 4.075000 190.675000 ;
      LAYER met4 ;
        RECT 3.755000 190.355000 4.075000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 190.760000 4.075000 191.080000 ;
      LAYER met4 ;
        RECT 3.755000 190.760000 4.075000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 191.165000 4.075000 191.485000 ;
      LAYER met4 ;
        RECT 3.755000 191.165000 4.075000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 191.570000 4.075000 191.890000 ;
      LAYER met4 ;
        RECT 3.755000 191.570000 4.075000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 191.975000 4.075000 192.295000 ;
      LAYER met4 ;
        RECT 3.755000 191.975000 4.075000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 192.380000 4.075000 192.700000 ;
      LAYER met4 ;
        RECT 3.755000 192.380000 4.075000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 192.785000 4.075000 193.105000 ;
      LAYER met4 ;
        RECT 3.755000 192.785000 4.075000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 193.190000 4.075000 193.510000 ;
      LAYER met4 ;
        RECT 3.755000 193.190000 4.075000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 193.595000 4.075000 193.915000 ;
      LAYER met4 ;
        RECT 3.755000 193.595000 4.075000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 194.000000 4.075000 194.320000 ;
      LAYER met4 ;
        RECT 3.755000 194.000000 4.075000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 194.405000 4.075000 194.725000 ;
      LAYER met4 ;
        RECT 3.755000 194.405000 4.075000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 194.810000 4.075000 195.130000 ;
      LAYER met4 ;
        RECT 3.755000 194.810000 4.075000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 195.215000 4.075000 195.535000 ;
      LAYER met4 ;
        RECT 3.755000 195.215000 4.075000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 195.620000 4.075000 195.940000 ;
      LAYER met4 ;
        RECT 3.755000 195.620000 4.075000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 196.025000 4.075000 196.345000 ;
      LAYER met4 ;
        RECT 3.755000 196.025000 4.075000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 196.430000 4.075000 196.750000 ;
      LAYER met4 ;
        RECT 3.755000 196.430000 4.075000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 196.835000 4.075000 197.155000 ;
      LAYER met4 ;
        RECT 3.755000 196.835000 4.075000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 197.240000 4.075000 197.560000 ;
      LAYER met4 ;
        RECT 3.755000 197.240000 4.075000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755000 197.645000 4.075000 197.965000 ;
      LAYER met4 ;
        RECT 3.755000 197.645000 4.075000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 23.850000 4.120000 24.170000 ;
      LAYER met4 ;
        RECT 3.800000 23.850000 4.120000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 24.280000 4.120000 24.600000 ;
      LAYER met4 ;
        RECT 3.800000 24.280000 4.120000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 24.710000 4.120000 25.030000 ;
      LAYER met4 ;
        RECT 3.800000 24.710000 4.120000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 25.140000 4.120000 25.460000 ;
      LAYER met4 ;
        RECT 3.800000 25.140000 4.120000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 25.570000 4.120000 25.890000 ;
      LAYER met4 ;
        RECT 3.800000 25.570000 4.120000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 26.000000 4.120000 26.320000 ;
      LAYER met4 ;
        RECT 3.800000 26.000000 4.120000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 26.430000 4.120000 26.750000 ;
      LAYER met4 ;
        RECT 3.800000 26.430000 4.120000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 26.860000 4.120000 27.180000 ;
      LAYER met4 ;
        RECT 3.800000 26.860000 4.120000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 27.290000 4.120000 27.610000 ;
      LAYER met4 ;
        RECT 3.800000 27.290000 4.120000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 27.720000 4.120000 28.040000 ;
      LAYER met4 ;
        RECT 3.800000 27.720000 4.120000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 28.150000 4.120000 28.470000 ;
      LAYER met4 ;
        RECT 3.800000 28.150000 4.120000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.815000 173.900000 4.015000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.815000 174.300000 4.015000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.815000 174.700000 4.015000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.815000 175.100000 4.015000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.815000 175.500000 4.015000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.815000 175.900000 4.015000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.815000 176.300000 4.015000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.815000 176.700000 4.015000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.815000 177.100000 4.015000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.815000 177.500000 4.015000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.815000 177.900000 4.015000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.815000 178.300000 4.015000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.815000 178.700000 4.015000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.815000 179.100000 4.015000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.815000 179.500000 4.015000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.815000 179.900000 4.015000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.815000 180.300000 4.015000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.815000 180.700000 4.015000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.815000 181.100000 4.015000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 181.445000 4.475000 181.765000 ;
      LAYER met4 ;
        RECT 4.155000 181.445000 4.475000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 181.850000 4.475000 182.170000 ;
      LAYER met4 ;
        RECT 4.155000 181.850000 4.475000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 182.255000 4.475000 182.575000 ;
      LAYER met4 ;
        RECT 4.155000 182.255000 4.475000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 182.660000 4.475000 182.980000 ;
      LAYER met4 ;
        RECT 4.155000 182.660000 4.475000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 183.065000 4.475000 183.385000 ;
      LAYER met4 ;
        RECT 4.155000 183.065000 4.475000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 183.470000 4.475000 183.790000 ;
      LAYER met4 ;
        RECT 4.155000 183.470000 4.475000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 183.875000 4.475000 184.195000 ;
      LAYER met4 ;
        RECT 4.155000 183.875000 4.475000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 184.280000 4.475000 184.600000 ;
      LAYER met4 ;
        RECT 4.155000 184.280000 4.475000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 184.685000 4.475000 185.005000 ;
      LAYER met4 ;
        RECT 4.155000 184.685000 4.475000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 185.090000 4.475000 185.410000 ;
      LAYER met4 ;
        RECT 4.155000 185.090000 4.475000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 185.495000 4.475000 185.815000 ;
      LAYER met4 ;
        RECT 4.155000 185.495000 4.475000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 185.900000 4.475000 186.220000 ;
      LAYER met4 ;
        RECT 4.155000 185.900000 4.475000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 186.305000 4.475000 186.625000 ;
      LAYER met4 ;
        RECT 4.155000 186.305000 4.475000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 186.710000 4.475000 187.030000 ;
      LAYER met4 ;
        RECT 4.155000 186.710000 4.475000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 187.115000 4.475000 187.435000 ;
      LAYER met4 ;
        RECT 4.155000 187.115000 4.475000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 187.520000 4.475000 187.840000 ;
      LAYER met4 ;
        RECT 4.155000 187.520000 4.475000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 187.925000 4.475000 188.245000 ;
      LAYER met4 ;
        RECT 4.155000 187.925000 4.475000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 188.330000 4.475000 188.650000 ;
      LAYER met4 ;
        RECT 4.155000 188.330000 4.475000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 188.735000 4.475000 189.055000 ;
      LAYER met4 ;
        RECT 4.155000 188.735000 4.475000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 189.140000 4.475000 189.460000 ;
      LAYER met4 ;
        RECT 4.155000 189.140000 4.475000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 189.545000 4.475000 189.865000 ;
      LAYER met4 ;
        RECT 4.155000 189.545000 4.475000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 189.950000 4.475000 190.270000 ;
      LAYER met4 ;
        RECT 4.155000 189.950000 4.475000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 190.355000 4.475000 190.675000 ;
      LAYER met4 ;
        RECT 4.155000 190.355000 4.475000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 190.760000 4.475000 191.080000 ;
      LAYER met4 ;
        RECT 4.155000 190.760000 4.475000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 191.165000 4.475000 191.485000 ;
      LAYER met4 ;
        RECT 4.155000 191.165000 4.475000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 191.570000 4.475000 191.890000 ;
      LAYER met4 ;
        RECT 4.155000 191.570000 4.475000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 191.975000 4.475000 192.295000 ;
      LAYER met4 ;
        RECT 4.155000 191.975000 4.475000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 192.380000 4.475000 192.700000 ;
      LAYER met4 ;
        RECT 4.155000 192.380000 4.475000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 192.785000 4.475000 193.105000 ;
      LAYER met4 ;
        RECT 4.155000 192.785000 4.475000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 193.190000 4.475000 193.510000 ;
      LAYER met4 ;
        RECT 4.155000 193.190000 4.475000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 193.595000 4.475000 193.915000 ;
      LAYER met4 ;
        RECT 4.155000 193.595000 4.475000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 194.000000 4.475000 194.320000 ;
      LAYER met4 ;
        RECT 4.155000 194.000000 4.475000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 194.405000 4.475000 194.725000 ;
      LAYER met4 ;
        RECT 4.155000 194.405000 4.475000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 194.810000 4.475000 195.130000 ;
      LAYER met4 ;
        RECT 4.155000 194.810000 4.475000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 195.215000 4.475000 195.535000 ;
      LAYER met4 ;
        RECT 4.155000 195.215000 4.475000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 195.620000 4.475000 195.940000 ;
      LAYER met4 ;
        RECT 4.155000 195.620000 4.475000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 196.025000 4.475000 196.345000 ;
      LAYER met4 ;
        RECT 4.155000 196.025000 4.475000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 196.430000 4.475000 196.750000 ;
      LAYER met4 ;
        RECT 4.155000 196.430000 4.475000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 196.835000 4.475000 197.155000 ;
      LAYER met4 ;
        RECT 4.155000 196.835000 4.475000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 197.240000 4.475000 197.560000 ;
      LAYER met4 ;
        RECT 4.155000 197.240000 4.475000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155000 197.645000 4.475000 197.965000 ;
      LAYER met4 ;
        RECT 4.155000 197.645000 4.475000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 23.850000 4.525000 24.170000 ;
      LAYER met4 ;
        RECT 4.205000 23.850000 4.525000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 24.280000 4.525000 24.600000 ;
      LAYER met4 ;
        RECT 4.205000 24.280000 4.525000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 24.710000 4.525000 25.030000 ;
      LAYER met4 ;
        RECT 4.205000 24.710000 4.525000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 25.140000 4.525000 25.460000 ;
      LAYER met4 ;
        RECT 4.205000 25.140000 4.525000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 25.570000 4.525000 25.890000 ;
      LAYER met4 ;
        RECT 4.205000 25.570000 4.525000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 26.000000 4.525000 26.320000 ;
      LAYER met4 ;
        RECT 4.205000 26.000000 4.525000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 26.430000 4.525000 26.750000 ;
      LAYER met4 ;
        RECT 4.205000 26.430000 4.525000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 26.860000 4.525000 27.180000 ;
      LAYER met4 ;
        RECT 4.205000 26.860000 4.525000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 27.290000 4.525000 27.610000 ;
      LAYER met4 ;
        RECT 4.205000 27.290000 4.525000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 27.720000 4.525000 28.040000 ;
      LAYER met4 ;
        RECT 4.205000 27.720000 4.525000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 28.150000 4.525000 28.470000 ;
      LAYER met4 ;
        RECT 4.205000 28.150000 4.525000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.215000 173.900000 4.415000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.215000 174.300000 4.415000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.215000 174.700000 4.415000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.215000 175.100000 4.415000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.215000 175.500000 4.415000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.215000 175.900000 4.415000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.215000 176.300000 4.415000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.215000 176.700000 4.415000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.215000 177.100000 4.415000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.215000 177.500000 4.415000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.215000 177.900000 4.415000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.215000 178.300000 4.415000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.215000 178.700000 4.415000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.215000 179.100000 4.415000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.215000 179.500000 4.415000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.215000 179.900000 4.415000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.215000 180.300000 4.415000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.215000 180.700000 4.415000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.215000 181.100000 4.415000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 181.445000 4.875000 181.765000 ;
      LAYER met4 ;
        RECT 4.555000 181.445000 4.875000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 181.850000 4.875000 182.170000 ;
      LAYER met4 ;
        RECT 4.555000 181.850000 4.875000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 182.255000 4.875000 182.575000 ;
      LAYER met4 ;
        RECT 4.555000 182.255000 4.875000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 182.660000 4.875000 182.980000 ;
      LAYER met4 ;
        RECT 4.555000 182.660000 4.875000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 183.065000 4.875000 183.385000 ;
      LAYER met4 ;
        RECT 4.555000 183.065000 4.875000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 183.470000 4.875000 183.790000 ;
      LAYER met4 ;
        RECT 4.555000 183.470000 4.875000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 183.875000 4.875000 184.195000 ;
      LAYER met4 ;
        RECT 4.555000 183.875000 4.875000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 184.280000 4.875000 184.600000 ;
      LAYER met4 ;
        RECT 4.555000 184.280000 4.875000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 184.685000 4.875000 185.005000 ;
      LAYER met4 ;
        RECT 4.555000 184.685000 4.875000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 185.090000 4.875000 185.410000 ;
      LAYER met4 ;
        RECT 4.555000 185.090000 4.875000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 185.495000 4.875000 185.815000 ;
      LAYER met4 ;
        RECT 4.555000 185.495000 4.875000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 185.900000 4.875000 186.220000 ;
      LAYER met4 ;
        RECT 4.555000 185.900000 4.875000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 186.305000 4.875000 186.625000 ;
      LAYER met4 ;
        RECT 4.555000 186.305000 4.875000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 186.710000 4.875000 187.030000 ;
      LAYER met4 ;
        RECT 4.555000 186.710000 4.875000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 187.115000 4.875000 187.435000 ;
      LAYER met4 ;
        RECT 4.555000 187.115000 4.875000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 187.520000 4.875000 187.840000 ;
      LAYER met4 ;
        RECT 4.555000 187.520000 4.875000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 187.925000 4.875000 188.245000 ;
      LAYER met4 ;
        RECT 4.555000 187.925000 4.875000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 188.330000 4.875000 188.650000 ;
      LAYER met4 ;
        RECT 4.555000 188.330000 4.875000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 188.735000 4.875000 189.055000 ;
      LAYER met4 ;
        RECT 4.555000 188.735000 4.875000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 189.140000 4.875000 189.460000 ;
      LAYER met4 ;
        RECT 4.555000 189.140000 4.875000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 189.545000 4.875000 189.865000 ;
      LAYER met4 ;
        RECT 4.555000 189.545000 4.875000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 189.950000 4.875000 190.270000 ;
      LAYER met4 ;
        RECT 4.555000 189.950000 4.875000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 190.355000 4.875000 190.675000 ;
      LAYER met4 ;
        RECT 4.555000 190.355000 4.875000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 190.760000 4.875000 191.080000 ;
      LAYER met4 ;
        RECT 4.555000 190.760000 4.875000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 191.165000 4.875000 191.485000 ;
      LAYER met4 ;
        RECT 4.555000 191.165000 4.875000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 191.570000 4.875000 191.890000 ;
      LAYER met4 ;
        RECT 4.555000 191.570000 4.875000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 191.975000 4.875000 192.295000 ;
      LAYER met4 ;
        RECT 4.555000 191.975000 4.875000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 192.380000 4.875000 192.700000 ;
      LAYER met4 ;
        RECT 4.555000 192.380000 4.875000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 192.785000 4.875000 193.105000 ;
      LAYER met4 ;
        RECT 4.555000 192.785000 4.875000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 193.190000 4.875000 193.510000 ;
      LAYER met4 ;
        RECT 4.555000 193.190000 4.875000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 193.595000 4.875000 193.915000 ;
      LAYER met4 ;
        RECT 4.555000 193.595000 4.875000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 194.000000 4.875000 194.320000 ;
      LAYER met4 ;
        RECT 4.555000 194.000000 4.875000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 194.405000 4.875000 194.725000 ;
      LAYER met4 ;
        RECT 4.555000 194.405000 4.875000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 194.810000 4.875000 195.130000 ;
      LAYER met4 ;
        RECT 4.555000 194.810000 4.875000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 195.215000 4.875000 195.535000 ;
      LAYER met4 ;
        RECT 4.555000 195.215000 4.875000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 195.620000 4.875000 195.940000 ;
      LAYER met4 ;
        RECT 4.555000 195.620000 4.875000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 196.025000 4.875000 196.345000 ;
      LAYER met4 ;
        RECT 4.555000 196.025000 4.875000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 196.430000 4.875000 196.750000 ;
      LAYER met4 ;
        RECT 4.555000 196.430000 4.875000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 196.835000 4.875000 197.155000 ;
      LAYER met4 ;
        RECT 4.555000 196.835000 4.875000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 197.240000 4.875000 197.560000 ;
      LAYER met4 ;
        RECT 4.555000 197.240000 4.875000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555000 197.645000 4.875000 197.965000 ;
      LAYER met4 ;
        RECT 4.555000 197.645000 4.875000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 23.850000 4.930000 24.170000 ;
      LAYER met4 ;
        RECT 4.610000 23.850000 4.930000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 24.280000 4.930000 24.600000 ;
      LAYER met4 ;
        RECT 4.610000 24.280000 4.930000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 24.710000 4.930000 25.030000 ;
      LAYER met4 ;
        RECT 4.610000 24.710000 4.930000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 25.140000 4.930000 25.460000 ;
      LAYER met4 ;
        RECT 4.610000 25.140000 4.930000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 25.570000 4.930000 25.890000 ;
      LAYER met4 ;
        RECT 4.610000 25.570000 4.930000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 26.000000 4.930000 26.320000 ;
      LAYER met4 ;
        RECT 4.610000 26.000000 4.930000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 26.430000 4.930000 26.750000 ;
      LAYER met4 ;
        RECT 4.610000 26.430000 4.930000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 26.860000 4.930000 27.180000 ;
      LAYER met4 ;
        RECT 4.610000 26.860000 4.930000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 27.290000 4.930000 27.610000 ;
      LAYER met4 ;
        RECT 4.610000 27.290000 4.930000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 27.720000 4.930000 28.040000 ;
      LAYER met4 ;
        RECT 4.610000 27.720000 4.930000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 28.150000 4.930000 28.470000 ;
      LAYER met4 ;
        RECT 4.610000 28.150000 4.930000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.615000 173.900000 4.815000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.615000 174.300000 4.815000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.615000 174.700000 4.815000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.615000 175.100000 4.815000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.615000 175.500000 4.815000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.615000 175.900000 4.815000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.615000 176.300000 4.815000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.615000 176.700000 4.815000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.615000 177.100000 4.815000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.615000 177.500000 4.815000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.615000 177.900000 4.815000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.615000 178.300000 4.815000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.615000 178.700000 4.815000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.615000 179.100000 4.815000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.615000 179.500000 4.815000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.615000 179.900000 4.815000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.615000 180.300000 4.815000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.615000 180.700000 4.815000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.615000 181.100000 4.815000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 181.445000 5.275000 181.765000 ;
      LAYER met4 ;
        RECT 4.955000 181.445000 5.275000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 181.850000 5.275000 182.170000 ;
      LAYER met4 ;
        RECT 4.955000 181.850000 5.275000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 182.255000 5.275000 182.575000 ;
      LAYER met4 ;
        RECT 4.955000 182.255000 5.275000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 182.660000 5.275000 182.980000 ;
      LAYER met4 ;
        RECT 4.955000 182.660000 5.275000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 183.065000 5.275000 183.385000 ;
      LAYER met4 ;
        RECT 4.955000 183.065000 5.275000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 183.470000 5.275000 183.790000 ;
      LAYER met4 ;
        RECT 4.955000 183.470000 5.275000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 183.875000 5.275000 184.195000 ;
      LAYER met4 ;
        RECT 4.955000 183.875000 5.275000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 184.280000 5.275000 184.600000 ;
      LAYER met4 ;
        RECT 4.955000 184.280000 5.275000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 184.685000 5.275000 185.005000 ;
      LAYER met4 ;
        RECT 4.955000 184.685000 5.275000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 185.090000 5.275000 185.410000 ;
      LAYER met4 ;
        RECT 4.955000 185.090000 5.275000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 185.495000 5.275000 185.815000 ;
      LAYER met4 ;
        RECT 4.955000 185.495000 5.275000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 185.900000 5.275000 186.220000 ;
      LAYER met4 ;
        RECT 4.955000 185.900000 5.275000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 186.305000 5.275000 186.625000 ;
      LAYER met4 ;
        RECT 4.955000 186.305000 5.275000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 186.710000 5.275000 187.030000 ;
      LAYER met4 ;
        RECT 4.955000 186.710000 5.275000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 187.115000 5.275000 187.435000 ;
      LAYER met4 ;
        RECT 4.955000 187.115000 5.275000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 187.520000 5.275000 187.840000 ;
      LAYER met4 ;
        RECT 4.955000 187.520000 5.275000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 187.925000 5.275000 188.245000 ;
      LAYER met4 ;
        RECT 4.955000 187.925000 5.275000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 188.330000 5.275000 188.650000 ;
      LAYER met4 ;
        RECT 4.955000 188.330000 5.275000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 188.735000 5.275000 189.055000 ;
      LAYER met4 ;
        RECT 4.955000 188.735000 5.275000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 189.140000 5.275000 189.460000 ;
      LAYER met4 ;
        RECT 4.955000 189.140000 5.275000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 189.545000 5.275000 189.865000 ;
      LAYER met4 ;
        RECT 4.955000 189.545000 5.275000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 189.950000 5.275000 190.270000 ;
      LAYER met4 ;
        RECT 4.955000 189.950000 5.275000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 190.355000 5.275000 190.675000 ;
      LAYER met4 ;
        RECT 4.955000 190.355000 5.275000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 190.760000 5.275000 191.080000 ;
      LAYER met4 ;
        RECT 4.955000 190.760000 5.275000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 191.165000 5.275000 191.485000 ;
      LAYER met4 ;
        RECT 4.955000 191.165000 5.275000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 191.570000 5.275000 191.890000 ;
      LAYER met4 ;
        RECT 4.955000 191.570000 5.275000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 191.975000 5.275000 192.295000 ;
      LAYER met4 ;
        RECT 4.955000 191.975000 5.275000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 192.380000 5.275000 192.700000 ;
      LAYER met4 ;
        RECT 4.955000 192.380000 5.275000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 192.785000 5.275000 193.105000 ;
      LAYER met4 ;
        RECT 4.955000 192.785000 5.275000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 193.190000 5.275000 193.510000 ;
      LAYER met4 ;
        RECT 4.955000 193.190000 5.275000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 193.595000 5.275000 193.915000 ;
      LAYER met4 ;
        RECT 4.955000 193.595000 5.275000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 194.000000 5.275000 194.320000 ;
      LAYER met4 ;
        RECT 4.955000 194.000000 5.275000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 194.405000 5.275000 194.725000 ;
      LAYER met4 ;
        RECT 4.955000 194.405000 5.275000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 194.810000 5.275000 195.130000 ;
      LAYER met4 ;
        RECT 4.955000 194.810000 5.275000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 195.215000 5.275000 195.535000 ;
      LAYER met4 ;
        RECT 4.955000 195.215000 5.275000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 195.620000 5.275000 195.940000 ;
      LAYER met4 ;
        RECT 4.955000 195.620000 5.275000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 196.025000 5.275000 196.345000 ;
      LAYER met4 ;
        RECT 4.955000 196.025000 5.275000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 196.430000 5.275000 196.750000 ;
      LAYER met4 ;
        RECT 4.955000 196.430000 5.275000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 196.835000 5.275000 197.155000 ;
      LAYER met4 ;
        RECT 4.955000 196.835000 5.275000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 197.240000 5.275000 197.560000 ;
      LAYER met4 ;
        RECT 4.955000 197.240000 5.275000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955000 197.645000 5.275000 197.965000 ;
      LAYER met4 ;
        RECT 4.955000 197.645000 5.275000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 173.900000 5.215000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 174.300000 5.215000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 174.700000 5.215000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 175.100000 5.215000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 175.500000 5.215000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 175.900000 5.215000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 176.300000 5.215000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 176.700000 5.215000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 177.100000 5.215000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 177.500000 5.215000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 177.900000 5.215000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 178.300000 5.215000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 178.700000 5.215000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 179.100000 5.215000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 179.500000 5.215000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 179.900000 5.215000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 180.300000 5.215000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 180.700000 5.215000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 181.100000 5.215000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 23.850000 5.335000 24.170000 ;
      LAYER met4 ;
        RECT 5.015000 23.850000 5.335000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 24.280000 5.335000 24.600000 ;
      LAYER met4 ;
        RECT 5.015000 24.280000 5.335000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 24.710000 5.335000 25.030000 ;
      LAYER met4 ;
        RECT 5.015000 24.710000 5.335000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 25.140000 5.335000 25.460000 ;
      LAYER met4 ;
        RECT 5.015000 25.140000 5.335000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 25.570000 5.335000 25.890000 ;
      LAYER met4 ;
        RECT 5.015000 25.570000 5.335000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 26.000000 5.335000 26.320000 ;
      LAYER met4 ;
        RECT 5.015000 26.000000 5.335000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 26.430000 5.335000 26.750000 ;
      LAYER met4 ;
        RECT 5.015000 26.430000 5.335000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 26.860000 5.335000 27.180000 ;
      LAYER met4 ;
        RECT 5.015000 26.860000 5.335000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 27.290000 5.335000 27.610000 ;
      LAYER met4 ;
        RECT 5.015000 27.290000 5.335000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 27.720000 5.335000 28.040000 ;
      LAYER met4 ;
        RECT 5.015000 27.720000 5.335000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 28.150000 5.335000 28.470000 ;
      LAYER met4 ;
        RECT 5.015000 28.150000 5.335000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 181.445000 5.675000 181.765000 ;
      LAYER met4 ;
        RECT 5.355000 181.445000 5.675000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 181.850000 5.675000 182.170000 ;
      LAYER met4 ;
        RECT 5.355000 181.850000 5.675000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 182.255000 5.675000 182.575000 ;
      LAYER met4 ;
        RECT 5.355000 182.255000 5.675000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 182.660000 5.675000 182.980000 ;
      LAYER met4 ;
        RECT 5.355000 182.660000 5.675000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 183.065000 5.675000 183.385000 ;
      LAYER met4 ;
        RECT 5.355000 183.065000 5.675000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 183.470000 5.675000 183.790000 ;
      LAYER met4 ;
        RECT 5.355000 183.470000 5.675000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 183.875000 5.675000 184.195000 ;
      LAYER met4 ;
        RECT 5.355000 183.875000 5.675000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 184.280000 5.675000 184.600000 ;
      LAYER met4 ;
        RECT 5.355000 184.280000 5.675000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 184.685000 5.675000 185.005000 ;
      LAYER met4 ;
        RECT 5.355000 184.685000 5.675000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 185.090000 5.675000 185.410000 ;
      LAYER met4 ;
        RECT 5.355000 185.090000 5.675000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 185.495000 5.675000 185.815000 ;
      LAYER met4 ;
        RECT 5.355000 185.495000 5.675000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 185.900000 5.675000 186.220000 ;
      LAYER met4 ;
        RECT 5.355000 185.900000 5.675000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 186.305000 5.675000 186.625000 ;
      LAYER met4 ;
        RECT 5.355000 186.305000 5.675000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 186.710000 5.675000 187.030000 ;
      LAYER met4 ;
        RECT 5.355000 186.710000 5.675000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 187.115000 5.675000 187.435000 ;
      LAYER met4 ;
        RECT 5.355000 187.115000 5.675000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 187.520000 5.675000 187.840000 ;
      LAYER met4 ;
        RECT 5.355000 187.520000 5.675000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 187.925000 5.675000 188.245000 ;
      LAYER met4 ;
        RECT 5.355000 187.925000 5.675000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 188.330000 5.675000 188.650000 ;
      LAYER met4 ;
        RECT 5.355000 188.330000 5.675000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 188.735000 5.675000 189.055000 ;
      LAYER met4 ;
        RECT 5.355000 188.735000 5.675000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 189.140000 5.675000 189.460000 ;
      LAYER met4 ;
        RECT 5.355000 189.140000 5.675000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 189.545000 5.675000 189.865000 ;
      LAYER met4 ;
        RECT 5.355000 189.545000 5.675000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 189.950000 5.675000 190.270000 ;
      LAYER met4 ;
        RECT 5.355000 189.950000 5.675000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 190.355000 5.675000 190.675000 ;
      LAYER met4 ;
        RECT 5.355000 190.355000 5.675000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 190.760000 5.675000 191.080000 ;
      LAYER met4 ;
        RECT 5.355000 190.760000 5.675000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 191.165000 5.675000 191.485000 ;
      LAYER met4 ;
        RECT 5.355000 191.165000 5.675000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 191.570000 5.675000 191.890000 ;
      LAYER met4 ;
        RECT 5.355000 191.570000 5.675000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 191.975000 5.675000 192.295000 ;
      LAYER met4 ;
        RECT 5.355000 191.975000 5.675000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 192.380000 5.675000 192.700000 ;
      LAYER met4 ;
        RECT 5.355000 192.380000 5.675000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 192.785000 5.675000 193.105000 ;
      LAYER met4 ;
        RECT 5.355000 192.785000 5.675000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 193.190000 5.675000 193.510000 ;
      LAYER met4 ;
        RECT 5.355000 193.190000 5.675000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 193.595000 5.675000 193.915000 ;
      LAYER met4 ;
        RECT 5.355000 193.595000 5.675000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 194.000000 5.675000 194.320000 ;
      LAYER met4 ;
        RECT 5.355000 194.000000 5.675000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 194.405000 5.675000 194.725000 ;
      LAYER met4 ;
        RECT 5.355000 194.405000 5.675000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 194.810000 5.675000 195.130000 ;
      LAYER met4 ;
        RECT 5.355000 194.810000 5.675000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 195.215000 5.675000 195.535000 ;
      LAYER met4 ;
        RECT 5.355000 195.215000 5.675000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 195.620000 5.675000 195.940000 ;
      LAYER met4 ;
        RECT 5.355000 195.620000 5.675000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 196.025000 5.675000 196.345000 ;
      LAYER met4 ;
        RECT 5.355000 196.025000 5.675000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 196.430000 5.675000 196.750000 ;
      LAYER met4 ;
        RECT 5.355000 196.430000 5.675000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 196.835000 5.675000 197.155000 ;
      LAYER met4 ;
        RECT 5.355000 196.835000 5.675000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 197.240000 5.675000 197.560000 ;
      LAYER met4 ;
        RECT 5.355000 197.240000 5.675000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355000 197.645000 5.675000 197.965000 ;
      LAYER met4 ;
        RECT 5.355000 197.645000 5.675000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 173.900000 5.615000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 174.300000 5.615000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 174.700000 5.615000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 175.100000 5.615000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 175.500000 5.615000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 175.900000 5.615000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 176.300000 5.615000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 176.700000 5.615000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 177.100000 5.615000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 177.500000 5.615000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 177.900000 5.615000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 178.300000 5.615000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 178.700000 5.615000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 179.100000 5.615000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 179.500000 5.615000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 179.900000 5.615000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 180.300000 5.615000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 180.700000 5.615000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 181.100000 5.615000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 23.850000 5.740000 24.170000 ;
      LAYER met4 ;
        RECT 5.420000 23.850000 5.740000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 24.280000 5.740000 24.600000 ;
      LAYER met4 ;
        RECT 5.420000 24.280000 5.740000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 24.710000 5.740000 25.030000 ;
      LAYER met4 ;
        RECT 5.420000 24.710000 5.740000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 25.140000 5.740000 25.460000 ;
      LAYER met4 ;
        RECT 5.420000 25.140000 5.740000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 25.570000 5.740000 25.890000 ;
      LAYER met4 ;
        RECT 5.420000 25.570000 5.740000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 26.000000 5.740000 26.320000 ;
      LAYER met4 ;
        RECT 5.420000 26.000000 5.740000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 26.430000 5.740000 26.750000 ;
      LAYER met4 ;
        RECT 5.420000 26.430000 5.740000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 26.860000 5.740000 27.180000 ;
      LAYER met4 ;
        RECT 5.420000 26.860000 5.740000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 27.290000 5.740000 27.610000 ;
      LAYER met4 ;
        RECT 5.420000 27.290000 5.740000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 27.720000 5.740000 28.040000 ;
      LAYER met4 ;
        RECT 5.420000 27.720000 5.740000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 28.150000 5.740000 28.470000 ;
      LAYER met4 ;
        RECT 5.420000 28.150000 5.740000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 181.445000 6.075000 181.765000 ;
      LAYER met4 ;
        RECT 5.755000 181.445000 6.075000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 181.850000 6.075000 182.170000 ;
      LAYER met4 ;
        RECT 5.755000 181.850000 6.075000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 182.255000 6.075000 182.575000 ;
      LAYER met4 ;
        RECT 5.755000 182.255000 6.075000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 182.660000 6.075000 182.980000 ;
      LAYER met4 ;
        RECT 5.755000 182.660000 6.075000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 183.065000 6.075000 183.385000 ;
      LAYER met4 ;
        RECT 5.755000 183.065000 6.075000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 183.470000 6.075000 183.790000 ;
      LAYER met4 ;
        RECT 5.755000 183.470000 6.075000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 183.875000 6.075000 184.195000 ;
      LAYER met4 ;
        RECT 5.755000 183.875000 6.075000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 184.280000 6.075000 184.600000 ;
      LAYER met4 ;
        RECT 5.755000 184.280000 6.075000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 184.685000 6.075000 185.005000 ;
      LAYER met4 ;
        RECT 5.755000 184.685000 6.075000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 185.090000 6.075000 185.410000 ;
      LAYER met4 ;
        RECT 5.755000 185.090000 6.075000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 185.495000 6.075000 185.815000 ;
      LAYER met4 ;
        RECT 5.755000 185.495000 6.075000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 185.900000 6.075000 186.220000 ;
      LAYER met4 ;
        RECT 5.755000 185.900000 6.075000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 186.305000 6.075000 186.625000 ;
      LAYER met4 ;
        RECT 5.755000 186.305000 6.075000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 186.710000 6.075000 187.030000 ;
      LAYER met4 ;
        RECT 5.755000 186.710000 6.075000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 187.115000 6.075000 187.435000 ;
      LAYER met4 ;
        RECT 5.755000 187.115000 6.075000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 187.520000 6.075000 187.840000 ;
      LAYER met4 ;
        RECT 5.755000 187.520000 6.075000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 187.925000 6.075000 188.245000 ;
      LAYER met4 ;
        RECT 5.755000 187.925000 6.075000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 188.330000 6.075000 188.650000 ;
      LAYER met4 ;
        RECT 5.755000 188.330000 6.075000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 188.735000 6.075000 189.055000 ;
      LAYER met4 ;
        RECT 5.755000 188.735000 6.075000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 189.140000 6.075000 189.460000 ;
      LAYER met4 ;
        RECT 5.755000 189.140000 6.075000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 189.545000 6.075000 189.865000 ;
      LAYER met4 ;
        RECT 5.755000 189.545000 6.075000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 189.950000 6.075000 190.270000 ;
      LAYER met4 ;
        RECT 5.755000 189.950000 6.075000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 190.355000 6.075000 190.675000 ;
      LAYER met4 ;
        RECT 5.755000 190.355000 6.075000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 190.760000 6.075000 191.080000 ;
      LAYER met4 ;
        RECT 5.755000 190.760000 6.075000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 191.165000 6.075000 191.485000 ;
      LAYER met4 ;
        RECT 5.755000 191.165000 6.075000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 191.570000 6.075000 191.890000 ;
      LAYER met4 ;
        RECT 5.755000 191.570000 6.075000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 191.975000 6.075000 192.295000 ;
      LAYER met4 ;
        RECT 5.755000 191.975000 6.075000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 192.380000 6.075000 192.700000 ;
      LAYER met4 ;
        RECT 5.755000 192.380000 6.075000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 192.785000 6.075000 193.105000 ;
      LAYER met4 ;
        RECT 5.755000 192.785000 6.075000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 193.190000 6.075000 193.510000 ;
      LAYER met4 ;
        RECT 5.755000 193.190000 6.075000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 193.595000 6.075000 193.915000 ;
      LAYER met4 ;
        RECT 5.755000 193.595000 6.075000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 194.000000 6.075000 194.320000 ;
      LAYER met4 ;
        RECT 5.755000 194.000000 6.075000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 194.405000 6.075000 194.725000 ;
      LAYER met4 ;
        RECT 5.755000 194.405000 6.075000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 194.810000 6.075000 195.130000 ;
      LAYER met4 ;
        RECT 5.755000 194.810000 6.075000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 195.215000 6.075000 195.535000 ;
      LAYER met4 ;
        RECT 5.755000 195.215000 6.075000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 195.620000 6.075000 195.940000 ;
      LAYER met4 ;
        RECT 5.755000 195.620000 6.075000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 196.025000 6.075000 196.345000 ;
      LAYER met4 ;
        RECT 5.755000 196.025000 6.075000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 196.430000 6.075000 196.750000 ;
      LAYER met4 ;
        RECT 5.755000 196.430000 6.075000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 196.835000 6.075000 197.155000 ;
      LAYER met4 ;
        RECT 5.755000 196.835000 6.075000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 197.240000 6.075000 197.560000 ;
      LAYER met4 ;
        RECT 5.755000 197.240000 6.075000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755000 197.645000 6.075000 197.965000 ;
      LAYER met4 ;
        RECT 5.755000 197.645000 6.075000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.815000 173.900000 6.015000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.815000 174.300000 6.015000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.815000 174.700000 6.015000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.815000 175.100000 6.015000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.815000 175.500000 6.015000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.815000 175.900000 6.015000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.815000 176.300000 6.015000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.815000 176.700000 6.015000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.815000 177.100000 6.015000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.815000 177.500000 6.015000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.815000 177.900000 6.015000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.815000 178.300000 6.015000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.815000 178.700000 6.015000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.815000 179.100000 6.015000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.815000 179.500000 6.015000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.815000 179.900000 6.015000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.815000 180.300000 6.015000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.815000 180.700000 6.015000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.815000 181.100000 6.015000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 23.850000 6.145000 24.170000 ;
      LAYER met4 ;
        RECT 5.825000 23.850000 6.145000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 24.280000 6.145000 24.600000 ;
      LAYER met4 ;
        RECT 5.825000 24.280000 6.145000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 24.710000 6.145000 25.030000 ;
      LAYER met4 ;
        RECT 5.825000 24.710000 6.145000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 25.140000 6.145000 25.460000 ;
      LAYER met4 ;
        RECT 5.825000 25.140000 6.145000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 25.570000 6.145000 25.890000 ;
      LAYER met4 ;
        RECT 5.825000 25.570000 6.145000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 26.000000 6.145000 26.320000 ;
      LAYER met4 ;
        RECT 5.825000 26.000000 6.145000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 26.430000 6.145000 26.750000 ;
      LAYER met4 ;
        RECT 5.825000 26.430000 6.145000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 26.860000 6.145000 27.180000 ;
      LAYER met4 ;
        RECT 5.825000 26.860000 6.145000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 27.290000 6.145000 27.610000 ;
      LAYER met4 ;
        RECT 5.825000 27.290000 6.145000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 27.720000 6.145000 28.040000 ;
      LAYER met4 ;
        RECT 5.825000 27.720000 6.145000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 28.150000 6.145000 28.470000 ;
      LAYER met4 ;
        RECT 5.825000 28.150000 6.145000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 23.850000 51.105000 24.170000 ;
      LAYER met4 ;
        RECT 50.785000 23.850000 51.105000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 24.280000 51.105000 24.600000 ;
      LAYER met4 ;
        RECT 50.785000 24.280000 51.105000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 24.710000 51.105000 25.030000 ;
      LAYER met4 ;
        RECT 50.785000 24.710000 51.105000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 25.140000 51.105000 25.460000 ;
      LAYER met4 ;
        RECT 50.785000 25.140000 51.105000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 25.570000 51.105000 25.890000 ;
      LAYER met4 ;
        RECT 50.785000 25.570000 51.105000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 26.000000 51.105000 26.320000 ;
      LAYER met4 ;
        RECT 50.785000 26.000000 51.105000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 26.430000 51.105000 26.750000 ;
      LAYER met4 ;
        RECT 50.785000 26.430000 51.105000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 26.860000 51.105000 27.180000 ;
      LAYER met4 ;
        RECT 50.785000 26.860000 51.105000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 27.290000 51.105000 27.610000 ;
      LAYER met4 ;
        RECT 50.785000 27.290000 51.105000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 27.720000 51.105000 28.040000 ;
      LAYER met4 ;
        RECT 50.785000 27.720000 51.105000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 28.150000 51.105000 28.470000 ;
      LAYER met4 ;
        RECT 50.785000 28.150000 51.105000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 23.850000 51.515000 24.170000 ;
      LAYER met4 ;
        RECT 51.195000 23.850000 51.515000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 24.280000 51.515000 24.600000 ;
      LAYER met4 ;
        RECT 51.195000 24.280000 51.515000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 24.710000 51.515000 25.030000 ;
      LAYER met4 ;
        RECT 51.195000 24.710000 51.515000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 25.140000 51.515000 25.460000 ;
      LAYER met4 ;
        RECT 51.195000 25.140000 51.515000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 25.570000 51.515000 25.890000 ;
      LAYER met4 ;
        RECT 51.195000 25.570000 51.515000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 26.000000 51.515000 26.320000 ;
      LAYER met4 ;
        RECT 51.195000 26.000000 51.515000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 26.430000 51.515000 26.750000 ;
      LAYER met4 ;
        RECT 51.195000 26.430000 51.515000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 26.860000 51.515000 27.180000 ;
      LAYER met4 ;
        RECT 51.195000 26.860000 51.515000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 27.290000 51.515000 27.610000 ;
      LAYER met4 ;
        RECT 51.195000 27.290000 51.515000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 27.720000 51.515000 28.040000 ;
      LAYER met4 ;
        RECT 51.195000 27.720000 51.515000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 28.150000 51.515000 28.470000 ;
      LAYER met4 ;
        RECT 51.195000 28.150000 51.515000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 23.850000 51.925000 24.170000 ;
      LAYER met4 ;
        RECT 51.605000 23.850000 51.925000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 24.280000 51.925000 24.600000 ;
      LAYER met4 ;
        RECT 51.605000 24.280000 51.925000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 24.710000 51.925000 25.030000 ;
      LAYER met4 ;
        RECT 51.605000 24.710000 51.925000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 25.140000 51.925000 25.460000 ;
      LAYER met4 ;
        RECT 51.605000 25.140000 51.925000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 25.570000 51.925000 25.890000 ;
      LAYER met4 ;
        RECT 51.605000 25.570000 51.925000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 26.000000 51.925000 26.320000 ;
      LAYER met4 ;
        RECT 51.605000 26.000000 51.925000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 26.430000 51.925000 26.750000 ;
      LAYER met4 ;
        RECT 51.605000 26.430000 51.925000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 26.860000 51.925000 27.180000 ;
      LAYER met4 ;
        RECT 51.605000 26.860000 51.925000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 27.290000 51.925000 27.610000 ;
      LAYER met4 ;
        RECT 51.605000 27.290000 51.925000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 27.720000 51.925000 28.040000 ;
      LAYER met4 ;
        RECT 51.605000 27.720000 51.925000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 28.150000 51.925000 28.470000 ;
      LAYER met4 ;
        RECT 51.605000 28.150000 51.925000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 23.850000 52.335000 24.170000 ;
      LAYER met4 ;
        RECT 52.015000 23.850000 52.335000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 24.280000 52.335000 24.600000 ;
      LAYER met4 ;
        RECT 52.015000 24.280000 52.335000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 24.710000 52.335000 25.030000 ;
      LAYER met4 ;
        RECT 52.015000 24.710000 52.335000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 25.140000 52.335000 25.460000 ;
      LAYER met4 ;
        RECT 52.015000 25.140000 52.335000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 25.570000 52.335000 25.890000 ;
      LAYER met4 ;
        RECT 52.015000 25.570000 52.335000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 26.000000 52.335000 26.320000 ;
      LAYER met4 ;
        RECT 52.015000 26.000000 52.335000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 26.430000 52.335000 26.750000 ;
      LAYER met4 ;
        RECT 52.015000 26.430000 52.335000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 26.860000 52.335000 27.180000 ;
      LAYER met4 ;
        RECT 52.015000 26.860000 52.335000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 27.290000 52.335000 27.610000 ;
      LAYER met4 ;
        RECT 52.015000 27.290000 52.335000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 27.720000 52.335000 28.040000 ;
      LAYER met4 ;
        RECT 52.015000 27.720000 52.335000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 28.150000 52.335000 28.470000 ;
      LAYER met4 ;
        RECT 52.015000 28.150000 52.335000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 23.850000 52.745000 24.170000 ;
      LAYER met4 ;
        RECT 52.425000 23.850000 52.745000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 24.280000 52.745000 24.600000 ;
      LAYER met4 ;
        RECT 52.425000 24.280000 52.745000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 24.710000 52.745000 25.030000 ;
      LAYER met4 ;
        RECT 52.425000 24.710000 52.745000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 25.140000 52.745000 25.460000 ;
      LAYER met4 ;
        RECT 52.425000 25.140000 52.745000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 25.570000 52.745000 25.890000 ;
      LAYER met4 ;
        RECT 52.425000 25.570000 52.745000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 26.000000 52.745000 26.320000 ;
      LAYER met4 ;
        RECT 52.425000 26.000000 52.745000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 26.430000 52.745000 26.750000 ;
      LAYER met4 ;
        RECT 52.425000 26.430000 52.745000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 26.860000 52.745000 27.180000 ;
      LAYER met4 ;
        RECT 52.425000 26.860000 52.745000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 27.290000 52.745000 27.610000 ;
      LAYER met4 ;
        RECT 52.425000 27.290000 52.745000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 27.720000 52.745000 28.040000 ;
      LAYER met4 ;
        RECT 52.425000 27.720000 52.745000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 28.150000 52.745000 28.470000 ;
      LAYER met4 ;
        RECT 52.425000 28.150000 52.745000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 23.850000 53.155000 24.170000 ;
      LAYER met4 ;
        RECT 52.835000 23.850000 53.155000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 24.280000 53.155000 24.600000 ;
      LAYER met4 ;
        RECT 52.835000 24.280000 53.155000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 24.710000 53.155000 25.030000 ;
      LAYER met4 ;
        RECT 52.835000 24.710000 53.155000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 25.140000 53.155000 25.460000 ;
      LAYER met4 ;
        RECT 52.835000 25.140000 53.155000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 25.570000 53.155000 25.890000 ;
      LAYER met4 ;
        RECT 52.835000 25.570000 53.155000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 26.000000 53.155000 26.320000 ;
      LAYER met4 ;
        RECT 52.835000 26.000000 53.155000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 26.430000 53.155000 26.750000 ;
      LAYER met4 ;
        RECT 52.835000 26.430000 53.155000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 26.860000 53.155000 27.180000 ;
      LAYER met4 ;
        RECT 52.835000 26.860000 53.155000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 27.290000 53.155000 27.610000 ;
      LAYER met4 ;
        RECT 52.835000 27.290000 53.155000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 27.720000 53.155000 28.040000 ;
      LAYER met4 ;
        RECT 52.835000 27.720000 53.155000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 28.150000 53.155000 28.470000 ;
      LAYER met4 ;
        RECT 52.835000 28.150000 53.155000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 23.850000 53.565000 24.170000 ;
      LAYER met4 ;
        RECT 53.245000 23.850000 53.565000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 24.280000 53.565000 24.600000 ;
      LAYER met4 ;
        RECT 53.245000 24.280000 53.565000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 24.710000 53.565000 25.030000 ;
      LAYER met4 ;
        RECT 53.245000 24.710000 53.565000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 25.140000 53.565000 25.460000 ;
      LAYER met4 ;
        RECT 53.245000 25.140000 53.565000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 25.570000 53.565000 25.890000 ;
      LAYER met4 ;
        RECT 53.245000 25.570000 53.565000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 26.000000 53.565000 26.320000 ;
      LAYER met4 ;
        RECT 53.245000 26.000000 53.565000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 26.430000 53.565000 26.750000 ;
      LAYER met4 ;
        RECT 53.245000 26.430000 53.565000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 26.860000 53.565000 27.180000 ;
      LAYER met4 ;
        RECT 53.245000 26.860000 53.565000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 27.290000 53.565000 27.610000 ;
      LAYER met4 ;
        RECT 53.245000 27.290000 53.565000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 27.720000 53.565000 28.040000 ;
      LAYER met4 ;
        RECT 53.245000 27.720000 53.565000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 28.150000 53.565000 28.470000 ;
      LAYER met4 ;
        RECT 53.245000 28.150000 53.565000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 23.850000 53.975000 24.170000 ;
      LAYER met4 ;
        RECT 53.655000 23.850000 53.975000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 24.280000 53.975000 24.600000 ;
      LAYER met4 ;
        RECT 53.655000 24.280000 53.975000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 24.710000 53.975000 25.030000 ;
      LAYER met4 ;
        RECT 53.655000 24.710000 53.975000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 25.140000 53.975000 25.460000 ;
      LAYER met4 ;
        RECT 53.655000 25.140000 53.975000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 25.570000 53.975000 25.890000 ;
      LAYER met4 ;
        RECT 53.655000 25.570000 53.975000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 26.000000 53.975000 26.320000 ;
      LAYER met4 ;
        RECT 53.655000 26.000000 53.975000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 26.430000 53.975000 26.750000 ;
      LAYER met4 ;
        RECT 53.655000 26.430000 53.975000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 26.860000 53.975000 27.180000 ;
      LAYER met4 ;
        RECT 53.655000 26.860000 53.975000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 27.290000 53.975000 27.610000 ;
      LAYER met4 ;
        RECT 53.655000 27.290000 53.975000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 27.720000 53.975000 28.040000 ;
      LAYER met4 ;
        RECT 53.655000 27.720000 53.975000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 28.150000 53.975000 28.470000 ;
      LAYER met4 ;
        RECT 53.655000 28.150000 53.975000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 23.850000 54.385000 24.170000 ;
      LAYER met4 ;
        RECT 54.065000 23.850000 54.385000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 24.280000 54.385000 24.600000 ;
      LAYER met4 ;
        RECT 54.065000 24.280000 54.385000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 24.710000 54.385000 25.030000 ;
      LAYER met4 ;
        RECT 54.065000 24.710000 54.385000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 25.140000 54.385000 25.460000 ;
      LAYER met4 ;
        RECT 54.065000 25.140000 54.385000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 25.570000 54.385000 25.890000 ;
      LAYER met4 ;
        RECT 54.065000 25.570000 54.385000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 26.000000 54.385000 26.320000 ;
      LAYER met4 ;
        RECT 54.065000 26.000000 54.385000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 26.430000 54.385000 26.750000 ;
      LAYER met4 ;
        RECT 54.065000 26.430000 54.385000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 26.860000 54.385000 27.180000 ;
      LAYER met4 ;
        RECT 54.065000 26.860000 54.385000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 27.290000 54.385000 27.610000 ;
      LAYER met4 ;
        RECT 54.065000 27.290000 54.385000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 27.720000 54.385000 28.040000 ;
      LAYER met4 ;
        RECT 54.065000 27.720000 54.385000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 28.150000 54.385000 28.470000 ;
      LAYER met4 ;
        RECT 54.065000 28.150000 54.385000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 23.850000 54.795000 24.170000 ;
      LAYER met4 ;
        RECT 54.475000 23.850000 54.795000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 24.280000 54.795000 24.600000 ;
      LAYER met4 ;
        RECT 54.475000 24.280000 54.795000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 24.710000 54.795000 25.030000 ;
      LAYER met4 ;
        RECT 54.475000 24.710000 54.795000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 25.140000 54.795000 25.460000 ;
      LAYER met4 ;
        RECT 54.475000 25.140000 54.795000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 25.570000 54.795000 25.890000 ;
      LAYER met4 ;
        RECT 54.475000 25.570000 54.795000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 26.000000 54.795000 26.320000 ;
      LAYER met4 ;
        RECT 54.475000 26.000000 54.795000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 26.430000 54.795000 26.750000 ;
      LAYER met4 ;
        RECT 54.475000 26.430000 54.795000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 26.860000 54.795000 27.180000 ;
      LAYER met4 ;
        RECT 54.475000 26.860000 54.795000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 27.290000 54.795000 27.610000 ;
      LAYER met4 ;
        RECT 54.475000 27.290000 54.795000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 27.720000 54.795000 28.040000 ;
      LAYER met4 ;
        RECT 54.475000 27.720000 54.795000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 28.150000 54.795000 28.470000 ;
      LAYER met4 ;
        RECT 54.475000 28.150000 54.795000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 23.850000 55.205000 24.170000 ;
      LAYER met4 ;
        RECT 54.885000 23.850000 55.205000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 24.280000 55.205000 24.600000 ;
      LAYER met4 ;
        RECT 54.885000 24.280000 55.205000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 24.710000 55.205000 25.030000 ;
      LAYER met4 ;
        RECT 54.885000 24.710000 55.205000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 25.140000 55.205000 25.460000 ;
      LAYER met4 ;
        RECT 54.885000 25.140000 55.205000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 25.570000 55.205000 25.890000 ;
      LAYER met4 ;
        RECT 54.885000 25.570000 55.205000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 26.000000 55.205000 26.320000 ;
      LAYER met4 ;
        RECT 54.885000 26.000000 55.205000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 26.430000 55.205000 26.750000 ;
      LAYER met4 ;
        RECT 54.885000 26.430000 55.205000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 26.860000 55.205000 27.180000 ;
      LAYER met4 ;
        RECT 54.885000 26.860000 55.205000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 27.290000 55.205000 27.610000 ;
      LAYER met4 ;
        RECT 54.885000 27.290000 55.205000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 27.720000 55.205000 28.040000 ;
      LAYER met4 ;
        RECT 54.885000 27.720000 55.205000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 28.150000 55.205000 28.470000 ;
      LAYER met4 ;
        RECT 54.885000 28.150000 55.205000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 23.850000 55.615000 24.170000 ;
      LAYER met4 ;
        RECT 55.295000 23.850000 55.615000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 24.280000 55.615000 24.600000 ;
      LAYER met4 ;
        RECT 55.295000 24.280000 55.615000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 24.710000 55.615000 25.030000 ;
      LAYER met4 ;
        RECT 55.295000 24.710000 55.615000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 25.140000 55.615000 25.460000 ;
      LAYER met4 ;
        RECT 55.295000 25.140000 55.615000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 25.570000 55.615000 25.890000 ;
      LAYER met4 ;
        RECT 55.295000 25.570000 55.615000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 26.000000 55.615000 26.320000 ;
      LAYER met4 ;
        RECT 55.295000 26.000000 55.615000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 26.430000 55.615000 26.750000 ;
      LAYER met4 ;
        RECT 55.295000 26.430000 55.615000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 26.860000 55.615000 27.180000 ;
      LAYER met4 ;
        RECT 55.295000 26.860000 55.615000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 27.290000 55.615000 27.610000 ;
      LAYER met4 ;
        RECT 55.295000 27.290000 55.615000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 27.720000 55.615000 28.040000 ;
      LAYER met4 ;
        RECT 55.295000 27.720000 55.615000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 28.150000 55.615000 28.470000 ;
      LAYER met4 ;
        RECT 55.295000 28.150000 55.615000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 23.850000 56.025000 24.170000 ;
      LAYER met4 ;
        RECT 55.705000 23.850000 56.025000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 24.280000 56.025000 24.600000 ;
      LAYER met4 ;
        RECT 55.705000 24.280000 56.025000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 24.710000 56.025000 25.030000 ;
      LAYER met4 ;
        RECT 55.705000 24.710000 56.025000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 25.140000 56.025000 25.460000 ;
      LAYER met4 ;
        RECT 55.705000 25.140000 56.025000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 25.570000 56.025000 25.890000 ;
      LAYER met4 ;
        RECT 55.705000 25.570000 56.025000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 26.000000 56.025000 26.320000 ;
      LAYER met4 ;
        RECT 55.705000 26.000000 56.025000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 26.430000 56.025000 26.750000 ;
      LAYER met4 ;
        RECT 55.705000 26.430000 56.025000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 26.860000 56.025000 27.180000 ;
      LAYER met4 ;
        RECT 55.705000 26.860000 56.025000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 27.290000 56.025000 27.610000 ;
      LAYER met4 ;
        RECT 55.705000 27.290000 56.025000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 27.720000 56.025000 28.040000 ;
      LAYER met4 ;
        RECT 55.705000 27.720000 56.025000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 28.150000 56.025000 28.470000 ;
      LAYER met4 ;
        RECT 55.705000 28.150000 56.025000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 23.850000 56.435000 24.170000 ;
      LAYER met4 ;
        RECT 56.115000 23.850000 56.435000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 24.280000 56.435000 24.600000 ;
      LAYER met4 ;
        RECT 56.115000 24.280000 56.435000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 24.710000 56.435000 25.030000 ;
      LAYER met4 ;
        RECT 56.115000 24.710000 56.435000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 25.140000 56.435000 25.460000 ;
      LAYER met4 ;
        RECT 56.115000 25.140000 56.435000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 25.570000 56.435000 25.890000 ;
      LAYER met4 ;
        RECT 56.115000 25.570000 56.435000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 26.000000 56.435000 26.320000 ;
      LAYER met4 ;
        RECT 56.115000 26.000000 56.435000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 26.430000 56.435000 26.750000 ;
      LAYER met4 ;
        RECT 56.115000 26.430000 56.435000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 26.860000 56.435000 27.180000 ;
      LAYER met4 ;
        RECT 56.115000 26.860000 56.435000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 27.290000 56.435000 27.610000 ;
      LAYER met4 ;
        RECT 56.115000 27.290000 56.435000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 27.720000 56.435000 28.040000 ;
      LAYER met4 ;
        RECT 56.115000 27.720000 56.435000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 28.150000 56.435000 28.470000 ;
      LAYER met4 ;
        RECT 56.115000 28.150000 56.435000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 23.850000 56.845000 24.170000 ;
      LAYER met4 ;
        RECT 56.525000 23.850000 56.845000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 24.280000 56.845000 24.600000 ;
      LAYER met4 ;
        RECT 56.525000 24.280000 56.845000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 24.710000 56.845000 25.030000 ;
      LAYER met4 ;
        RECT 56.525000 24.710000 56.845000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 25.140000 56.845000 25.460000 ;
      LAYER met4 ;
        RECT 56.525000 25.140000 56.845000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 25.570000 56.845000 25.890000 ;
      LAYER met4 ;
        RECT 56.525000 25.570000 56.845000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 26.000000 56.845000 26.320000 ;
      LAYER met4 ;
        RECT 56.525000 26.000000 56.845000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 26.430000 56.845000 26.750000 ;
      LAYER met4 ;
        RECT 56.525000 26.430000 56.845000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 26.860000 56.845000 27.180000 ;
      LAYER met4 ;
        RECT 56.525000 26.860000 56.845000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 27.290000 56.845000 27.610000 ;
      LAYER met4 ;
        RECT 56.525000 27.290000 56.845000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 27.720000 56.845000 28.040000 ;
      LAYER met4 ;
        RECT 56.525000 27.720000 56.845000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 28.150000 56.845000 28.470000 ;
      LAYER met4 ;
        RECT 56.525000 28.150000 56.845000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 23.850000 57.250000 24.170000 ;
      LAYER met4 ;
        RECT 56.930000 23.850000 57.250000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 24.280000 57.250000 24.600000 ;
      LAYER met4 ;
        RECT 56.930000 24.280000 57.250000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 24.710000 57.250000 25.030000 ;
      LAYER met4 ;
        RECT 56.930000 24.710000 57.250000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 25.140000 57.250000 25.460000 ;
      LAYER met4 ;
        RECT 56.930000 25.140000 57.250000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 25.570000 57.250000 25.890000 ;
      LAYER met4 ;
        RECT 56.930000 25.570000 57.250000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 26.000000 57.250000 26.320000 ;
      LAYER met4 ;
        RECT 56.930000 26.000000 57.250000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 26.430000 57.250000 26.750000 ;
      LAYER met4 ;
        RECT 56.930000 26.430000 57.250000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 26.860000 57.250000 27.180000 ;
      LAYER met4 ;
        RECT 56.930000 26.860000 57.250000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 27.290000 57.250000 27.610000 ;
      LAYER met4 ;
        RECT 56.930000 27.290000 57.250000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 27.720000 57.250000 28.040000 ;
      LAYER met4 ;
        RECT 56.930000 27.720000 57.250000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 28.150000 57.250000 28.470000 ;
      LAYER met4 ;
        RECT 56.930000 28.150000 57.250000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 23.850000 57.655000 24.170000 ;
      LAYER met4 ;
        RECT 57.335000 23.850000 57.655000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 24.280000 57.655000 24.600000 ;
      LAYER met4 ;
        RECT 57.335000 24.280000 57.655000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 24.710000 57.655000 25.030000 ;
      LAYER met4 ;
        RECT 57.335000 24.710000 57.655000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 25.140000 57.655000 25.460000 ;
      LAYER met4 ;
        RECT 57.335000 25.140000 57.655000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 25.570000 57.655000 25.890000 ;
      LAYER met4 ;
        RECT 57.335000 25.570000 57.655000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 26.000000 57.655000 26.320000 ;
      LAYER met4 ;
        RECT 57.335000 26.000000 57.655000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 26.430000 57.655000 26.750000 ;
      LAYER met4 ;
        RECT 57.335000 26.430000 57.655000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 26.860000 57.655000 27.180000 ;
      LAYER met4 ;
        RECT 57.335000 26.860000 57.655000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 27.290000 57.655000 27.610000 ;
      LAYER met4 ;
        RECT 57.335000 27.290000 57.655000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 27.720000 57.655000 28.040000 ;
      LAYER met4 ;
        RECT 57.335000 27.720000 57.655000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 28.150000 57.655000 28.470000 ;
      LAYER met4 ;
        RECT 57.335000 28.150000 57.655000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 23.850000 58.060000 24.170000 ;
      LAYER met4 ;
        RECT 57.740000 23.850000 58.060000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 24.280000 58.060000 24.600000 ;
      LAYER met4 ;
        RECT 57.740000 24.280000 58.060000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 24.710000 58.060000 25.030000 ;
      LAYER met4 ;
        RECT 57.740000 24.710000 58.060000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 25.140000 58.060000 25.460000 ;
      LAYER met4 ;
        RECT 57.740000 25.140000 58.060000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 25.570000 58.060000 25.890000 ;
      LAYER met4 ;
        RECT 57.740000 25.570000 58.060000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 26.000000 58.060000 26.320000 ;
      LAYER met4 ;
        RECT 57.740000 26.000000 58.060000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 26.430000 58.060000 26.750000 ;
      LAYER met4 ;
        RECT 57.740000 26.430000 58.060000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 26.860000 58.060000 27.180000 ;
      LAYER met4 ;
        RECT 57.740000 26.860000 58.060000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 27.290000 58.060000 27.610000 ;
      LAYER met4 ;
        RECT 57.740000 27.290000 58.060000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 27.720000 58.060000 28.040000 ;
      LAYER met4 ;
        RECT 57.740000 27.720000 58.060000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 28.150000 58.060000 28.470000 ;
      LAYER met4 ;
        RECT 57.740000 28.150000 58.060000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 23.850000 58.465000 24.170000 ;
      LAYER met4 ;
        RECT 58.145000 23.850000 58.465000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 24.280000 58.465000 24.600000 ;
      LAYER met4 ;
        RECT 58.145000 24.280000 58.465000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 24.710000 58.465000 25.030000 ;
      LAYER met4 ;
        RECT 58.145000 24.710000 58.465000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 25.140000 58.465000 25.460000 ;
      LAYER met4 ;
        RECT 58.145000 25.140000 58.465000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 25.570000 58.465000 25.890000 ;
      LAYER met4 ;
        RECT 58.145000 25.570000 58.465000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 26.000000 58.465000 26.320000 ;
      LAYER met4 ;
        RECT 58.145000 26.000000 58.465000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 26.430000 58.465000 26.750000 ;
      LAYER met4 ;
        RECT 58.145000 26.430000 58.465000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 26.860000 58.465000 27.180000 ;
      LAYER met4 ;
        RECT 58.145000 26.860000 58.465000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 27.290000 58.465000 27.610000 ;
      LAYER met4 ;
        RECT 58.145000 27.290000 58.465000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 27.720000 58.465000 28.040000 ;
      LAYER met4 ;
        RECT 58.145000 27.720000 58.465000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 28.150000 58.465000 28.470000 ;
      LAYER met4 ;
        RECT 58.145000 28.150000 58.465000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 23.850000 58.870000 24.170000 ;
      LAYER met4 ;
        RECT 58.550000 23.850000 58.870000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 24.280000 58.870000 24.600000 ;
      LAYER met4 ;
        RECT 58.550000 24.280000 58.870000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 24.710000 58.870000 25.030000 ;
      LAYER met4 ;
        RECT 58.550000 24.710000 58.870000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 25.140000 58.870000 25.460000 ;
      LAYER met4 ;
        RECT 58.550000 25.140000 58.870000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 25.570000 58.870000 25.890000 ;
      LAYER met4 ;
        RECT 58.550000 25.570000 58.870000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 26.000000 58.870000 26.320000 ;
      LAYER met4 ;
        RECT 58.550000 26.000000 58.870000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 26.430000 58.870000 26.750000 ;
      LAYER met4 ;
        RECT 58.550000 26.430000 58.870000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 26.860000 58.870000 27.180000 ;
      LAYER met4 ;
        RECT 58.550000 26.860000 58.870000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 27.290000 58.870000 27.610000 ;
      LAYER met4 ;
        RECT 58.550000 27.290000 58.870000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 27.720000 58.870000 28.040000 ;
      LAYER met4 ;
        RECT 58.550000 27.720000 58.870000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 28.150000 58.870000 28.470000 ;
      LAYER met4 ;
        RECT 58.550000 28.150000 58.870000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 23.850000 59.275000 24.170000 ;
      LAYER met4 ;
        RECT 58.955000 23.850000 59.275000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 24.280000 59.275000 24.600000 ;
      LAYER met4 ;
        RECT 58.955000 24.280000 59.275000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 24.710000 59.275000 25.030000 ;
      LAYER met4 ;
        RECT 58.955000 24.710000 59.275000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 25.140000 59.275000 25.460000 ;
      LAYER met4 ;
        RECT 58.955000 25.140000 59.275000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 25.570000 59.275000 25.890000 ;
      LAYER met4 ;
        RECT 58.955000 25.570000 59.275000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 26.000000 59.275000 26.320000 ;
      LAYER met4 ;
        RECT 58.955000 26.000000 59.275000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 26.430000 59.275000 26.750000 ;
      LAYER met4 ;
        RECT 58.955000 26.430000 59.275000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 26.860000 59.275000 27.180000 ;
      LAYER met4 ;
        RECT 58.955000 26.860000 59.275000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 27.290000 59.275000 27.610000 ;
      LAYER met4 ;
        RECT 58.955000 27.290000 59.275000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 27.720000 59.275000 28.040000 ;
      LAYER met4 ;
        RECT 58.955000 27.720000 59.275000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 28.150000 59.275000 28.470000 ;
      LAYER met4 ;
        RECT 58.955000 28.150000 59.275000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 23.850000 59.680000 24.170000 ;
      LAYER met4 ;
        RECT 59.360000 23.850000 59.680000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 24.280000 59.680000 24.600000 ;
      LAYER met4 ;
        RECT 59.360000 24.280000 59.680000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 24.710000 59.680000 25.030000 ;
      LAYER met4 ;
        RECT 59.360000 24.710000 59.680000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 25.140000 59.680000 25.460000 ;
      LAYER met4 ;
        RECT 59.360000 25.140000 59.680000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 25.570000 59.680000 25.890000 ;
      LAYER met4 ;
        RECT 59.360000 25.570000 59.680000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 26.000000 59.680000 26.320000 ;
      LAYER met4 ;
        RECT 59.360000 26.000000 59.680000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 26.430000 59.680000 26.750000 ;
      LAYER met4 ;
        RECT 59.360000 26.430000 59.680000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 26.860000 59.680000 27.180000 ;
      LAYER met4 ;
        RECT 59.360000 26.860000 59.680000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 27.290000 59.680000 27.610000 ;
      LAYER met4 ;
        RECT 59.360000 27.290000 59.680000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 27.720000 59.680000 28.040000 ;
      LAYER met4 ;
        RECT 59.360000 27.720000 59.680000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 28.150000 59.680000 28.470000 ;
      LAYER met4 ;
        RECT 59.360000 28.150000 59.680000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 23.850000 60.085000 24.170000 ;
      LAYER met4 ;
        RECT 59.765000 23.850000 60.085000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 24.280000 60.085000 24.600000 ;
      LAYER met4 ;
        RECT 59.765000 24.280000 60.085000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 24.710000 60.085000 25.030000 ;
      LAYER met4 ;
        RECT 59.765000 24.710000 60.085000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 25.140000 60.085000 25.460000 ;
      LAYER met4 ;
        RECT 59.765000 25.140000 60.085000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 25.570000 60.085000 25.890000 ;
      LAYER met4 ;
        RECT 59.765000 25.570000 60.085000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 26.000000 60.085000 26.320000 ;
      LAYER met4 ;
        RECT 59.765000 26.000000 60.085000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 26.430000 60.085000 26.750000 ;
      LAYER met4 ;
        RECT 59.765000 26.430000 60.085000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 26.860000 60.085000 27.180000 ;
      LAYER met4 ;
        RECT 59.765000 26.860000 60.085000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 27.290000 60.085000 27.610000 ;
      LAYER met4 ;
        RECT 59.765000 27.290000 60.085000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 27.720000 60.085000 28.040000 ;
      LAYER met4 ;
        RECT 59.765000 27.720000 60.085000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 28.150000 60.085000 28.470000 ;
      LAYER met4 ;
        RECT 59.765000 28.150000 60.085000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 181.445000 6.475000 181.765000 ;
      LAYER met4 ;
        RECT 6.155000 181.445000 6.475000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 181.850000 6.475000 182.170000 ;
      LAYER met4 ;
        RECT 6.155000 181.850000 6.475000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 182.255000 6.475000 182.575000 ;
      LAYER met4 ;
        RECT 6.155000 182.255000 6.475000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 182.660000 6.475000 182.980000 ;
      LAYER met4 ;
        RECT 6.155000 182.660000 6.475000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 183.065000 6.475000 183.385000 ;
      LAYER met4 ;
        RECT 6.155000 183.065000 6.475000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 183.470000 6.475000 183.790000 ;
      LAYER met4 ;
        RECT 6.155000 183.470000 6.475000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 183.875000 6.475000 184.195000 ;
      LAYER met4 ;
        RECT 6.155000 183.875000 6.475000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 184.280000 6.475000 184.600000 ;
      LAYER met4 ;
        RECT 6.155000 184.280000 6.475000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 184.685000 6.475000 185.005000 ;
      LAYER met4 ;
        RECT 6.155000 184.685000 6.475000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 185.090000 6.475000 185.410000 ;
      LAYER met4 ;
        RECT 6.155000 185.090000 6.475000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 185.495000 6.475000 185.815000 ;
      LAYER met4 ;
        RECT 6.155000 185.495000 6.475000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 185.900000 6.475000 186.220000 ;
      LAYER met4 ;
        RECT 6.155000 185.900000 6.475000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 186.305000 6.475000 186.625000 ;
      LAYER met4 ;
        RECT 6.155000 186.305000 6.475000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 186.710000 6.475000 187.030000 ;
      LAYER met4 ;
        RECT 6.155000 186.710000 6.475000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 187.115000 6.475000 187.435000 ;
      LAYER met4 ;
        RECT 6.155000 187.115000 6.475000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 187.520000 6.475000 187.840000 ;
      LAYER met4 ;
        RECT 6.155000 187.520000 6.475000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 187.925000 6.475000 188.245000 ;
      LAYER met4 ;
        RECT 6.155000 187.925000 6.475000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 188.330000 6.475000 188.650000 ;
      LAYER met4 ;
        RECT 6.155000 188.330000 6.475000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 188.735000 6.475000 189.055000 ;
      LAYER met4 ;
        RECT 6.155000 188.735000 6.475000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 189.140000 6.475000 189.460000 ;
      LAYER met4 ;
        RECT 6.155000 189.140000 6.475000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 189.545000 6.475000 189.865000 ;
      LAYER met4 ;
        RECT 6.155000 189.545000 6.475000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 189.950000 6.475000 190.270000 ;
      LAYER met4 ;
        RECT 6.155000 189.950000 6.475000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 190.355000 6.475000 190.675000 ;
      LAYER met4 ;
        RECT 6.155000 190.355000 6.475000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 190.760000 6.475000 191.080000 ;
      LAYER met4 ;
        RECT 6.155000 190.760000 6.475000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 191.165000 6.475000 191.485000 ;
      LAYER met4 ;
        RECT 6.155000 191.165000 6.475000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 191.570000 6.475000 191.890000 ;
      LAYER met4 ;
        RECT 6.155000 191.570000 6.475000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 191.975000 6.475000 192.295000 ;
      LAYER met4 ;
        RECT 6.155000 191.975000 6.475000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 192.380000 6.475000 192.700000 ;
      LAYER met4 ;
        RECT 6.155000 192.380000 6.475000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 192.785000 6.475000 193.105000 ;
      LAYER met4 ;
        RECT 6.155000 192.785000 6.475000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 193.190000 6.475000 193.510000 ;
      LAYER met4 ;
        RECT 6.155000 193.190000 6.475000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 193.595000 6.475000 193.915000 ;
      LAYER met4 ;
        RECT 6.155000 193.595000 6.475000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 194.000000 6.475000 194.320000 ;
      LAYER met4 ;
        RECT 6.155000 194.000000 6.475000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 194.405000 6.475000 194.725000 ;
      LAYER met4 ;
        RECT 6.155000 194.405000 6.475000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 194.810000 6.475000 195.130000 ;
      LAYER met4 ;
        RECT 6.155000 194.810000 6.475000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 195.215000 6.475000 195.535000 ;
      LAYER met4 ;
        RECT 6.155000 195.215000 6.475000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 195.620000 6.475000 195.940000 ;
      LAYER met4 ;
        RECT 6.155000 195.620000 6.475000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 196.025000 6.475000 196.345000 ;
      LAYER met4 ;
        RECT 6.155000 196.025000 6.475000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 196.430000 6.475000 196.750000 ;
      LAYER met4 ;
        RECT 6.155000 196.430000 6.475000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 196.835000 6.475000 197.155000 ;
      LAYER met4 ;
        RECT 6.155000 196.835000 6.475000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 197.240000 6.475000 197.560000 ;
      LAYER met4 ;
        RECT 6.155000 197.240000 6.475000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155000 197.645000 6.475000 197.965000 ;
      LAYER met4 ;
        RECT 6.155000 197.645000 6.475000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.215000 173.900000 6.415000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.215000 174.300000 6.415000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.215000 174.700000 6.415000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.215000 175.100000 6.415000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.215000 175.500000 6.415000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.215000 175.900000 6.415000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.215000 176.300000 6.415000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.215000 176.700000 6.415000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.215000 177.100000 6.415000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.215000 177.500000 6.415000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.215000 177.900000 6.415000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.215000 178.300000 6.415000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.215000 178.700000 6.415000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.215000 179.100000 6.415000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.215000 179.500000 6.415000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.215000 179.900000 6.415000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.215000 180.300000 6.415000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.215000 180.700000 6.415000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.215000 181.100000 6.415000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 23.850000 6.550000 24.170000 ;
      LAYER met4 ;
        RECT 6.230000 23.850000 6.550000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 24.280000 6.550000 24.600000 ;
      LAYER met4 ;
        RECT 6.230000 24.280000 6.550000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 24.710000 6.550000 25.030000 ;
      LAYER met4 ;
        RECT 6.230000 24.710000 6.550000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 25.140000 6.550000 25.460000 ;
      LAYER met4 ;
        RECT 6.230000 25.140000 6.550000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 25.570000 6.550000 25.890000 ;
      LAYER met4 ;
        RECT 6.230000 25.570000 6.550000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 26.000000 6.550000 26.320000 ;
      LAYER met4 ;
        RECT 6.230000 26.000000 6.550000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 26.430000 6.550000 26.750000 ;
      LAYER met4 ;
        RECT 6.230000 26.430000 6.550000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 26.860000 6.550000 27.180000 ;
      LAYER met4 ;
        RECT 6.230000 26.860000 6.550000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 27.290000 6.550000 27.610000 ;
      LAYER met4 ;
        RECT 6.230000 27.290000 6.550000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 27.720000 6.550000 28.040000 ;
      LAYER met4 ;
        RECT 6.230000 27.720000 6.550000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 28.150000 6.550000 28.470000 ;
      LAYER met4 ;
        RECT 6.230000 28.150000 6.550000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 181.445000 6.875000 181.765000 ;
      LAYER met4 ;
        RECT 6.555000 181.445000 6.875000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 181.850000 6.875000 182.170000 ;
      LAYER met4 ;
        RECT 6.555000 181.850000 6.875000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 182.255000 6.875000 182.575000 ;
      LAYER met4 ;
        RECT 6.555000 182.255000 6.875000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 182.660000 6.875000 182.980000 ;
      LAYER met4 ;
        RECT 6.555000 182.660000 6.875000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 183.065000 6.875000 183.385000 ;
      LAYER met4 ;
        RECT 6.555000 183.065000 6.875000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 183.470000 6.875000 183.790000 ;
      LAYER met4 ;
        RECT 6.555000 183.470000 6.875000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 183.875000 6.875000 184.195000 ;
      LAYER met4 ;
        RECT 6.555000 183.875000 6.875000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 184.280000 6.875000 184.600000 ;
      LAYER met4 ;
        RECT 6.555000 184.280000 6.875000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 184.685000 6.875000 185.005000 ;
      LAYER met4 ;
        RECT 6.555000 184.685000 6.875000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 185.090000 6.875000 185.410000 ;
      LAYER met4 ;
        RECT 6.555000 185.090000 6.875000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 185.495000 6.875000 185.815000 ;
      LAYER met4 ;
        RECT 6.555000 185.495000 6.875000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 185.900000 6.875000 186.220000 ;
      LAYER met4 ;
        RECT 6.555000 185.900000 6.875000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 186.305000 6.875000 186.625000 ;
      LAYER met4 ;
        RECT 6.555000 186.305000 6.875000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 186.710000 6.875000 187.030000 ;
      LAYER met4 ;
        RECT 6.555000 186.710000 6.875000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 187.115000 6.875000 187.435000 ;
      LAYER met4 ;
        RECT 6.555000 187.115000 6.875000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 187.520000 6.875000 187.840000 ;
      LAYER met4 ;
        RECT 6.555000 187.520000 6.875000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 187.925000 6.875000 188.245000 ;
      LAYER met4 ;
        RECT 6.555000 187.925000 6.875000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 188.330000 6.875000 188.650000 ;
      LAYER met4 ;
        RECT 6.555000 188.330000 6.875000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 188.735000 6.875000 189.055000 ;
      LAYER met4 ;
        RECT 6.555000 188.735000 6.875000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 189.140000 6.875000 189.460000 ;
      LAYER met4 ;
        RECT 6.555000 189.140000 6.875000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 189.545000 6.875000 189.865000 ;
      LAYER met4 ;
        RECT 6.555000 189.545000 6.875000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 189.950000 6.875000 190.270000 ;
      LAYER met4 ;
        RECT 6.555000 189.950000 6.875000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 190.355000 6.875000 190.675000 ;
      LAYER met4 ;
        RECT 6.555000 190.355000 6.875000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 190.760000 6.875000 191.080000 ;
      LAYER met4 ;
        RECT 6.555000 190.760000 6.875000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 191.165000 6.875000 191.485000 ;
      LAYER met4 ;
        RECT 6.555000 191.165000 6.875000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 191.570000 6.875000 191.890000 ;
      LAYER met4 ;
        RECT 6.555000 191.570000 6.875000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 191.975000 6.875000 192.295000 ;
      LAYER met4 ;
        RECT 6.555000 191.975000 6.875000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 192.380000 6.875000 192.700000 ;
      LAYER met4 ;
        RECT 6.555000 192.380000 6.875000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 192.785000 6.875000 193.105000 ;
      LAYER met4 ;
        RECT 6.555000 192.785000 6.875000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 193.190000 6.875000 193.510000 ;
      LAYER met4 ;
        RECT 6.555000 193.190000 6.875000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 193.595000 6.875000 193.915000 ;
      LAYER met4 ;
        RECT 6.555000 193.595000 6.875000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 194.000000 6.875000 194.320000 ;
      LAYER met4 ;
        RECT 6.555000 194.000000 6.875000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 194.405000 6.875000 194.725000 ;
      LAYER met4 ;
        RECT 6.555000 194.405000 6.875000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 194.810000 6.875000 195.130000 ;
      LAYER met4 ;
        RECT 6.555000 194.810000 6.875000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 195.215000 6.875000 195.535000 ;
      LAYER met4 ;
        RECT 6.555000 195.215000 6.875000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 195.620000 6.875000 195.940000 ;
      LAYER met4 ;
        RECT 6.555000 195.620000 6.875000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 196.025000 6.875000 196.345000 ;
      LAYER met4 ;
        RECT 6.555000 196.025000 6.875000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 196.430000 6.875000 196.750000 ;
      LAYER met4 ;
        RECT 6.555000 196.430000 6.875000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 196.835000 6.875000 197.155000 ;
      LAYER met4 ;
        RECT 6.555000 196.835000 6.875000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 197.240000 6.875000 197.560000 ;
      LAYER met4 ;
        RECT 6.555000 197.240000 6.875000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555000 197.645000 6.875000 197.965000 ;
      LAYER met4 ;
        RECT 6.555000 197.645000 6.875000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.615000 173.900000 6.815000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.615000 174.300000 6.815000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.615000 174.700000 6.815000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.615000 175.100000 6.815000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.615000 175.500000 6.815000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.615000 175.900000 6.815000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.615000 176.300000 6.815000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.615000 176.700000 6.815000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.615000 177.100000 6.815000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.615000 177.500000 6.815000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.615000 177.900000 6.815000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.615000 178.300000 6.815000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.615000 178.700000 6.815000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.615000 179.100000 6.815000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.615000 179.500000 6.815000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.615000 179.900000 6.815000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.615000 180.300000 6.815000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.615000 180.700000 6.815000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.615000 181.100000 6.815000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 23.850000 6.955000 24.170000 ;
      LAYER met4 ;
        RECT 6.635000 23.850000 6.955000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 24.280000 6.955000 24.600000 ;
      LAYER met4 ;
        RECT 6.635000 24.280000 6.955000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 24.710000 6.955000 25.030000 ;
      LAYER met4 ;
        RECT 6.635000 24.710000 6.955000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 25.140000 6.955000 25.460000 ;
      LAYER met4 ;
        RECT 6.635000 25.140000 6.955000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 25.570000 6.955000 25.890000 ;
      LAYER met4 ;
        RECT 6.635000 25.570000 6.955000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 26.000000 6.955000 26.320000 ;
      LAYER met4 ;
        RECT 6.635000 26.000000 6.955000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 26.430000 6.955000 26.750000 ;
      LAYER met4 ;
        RECT 6.635000 26.430000 6.955000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 26.860000 6.955000 27.180000 ;
      LAYER met4 ;
        RECT 6.635000 26.860000 6.955000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 27.290000 6.955000 27.610000 ;
      LAYER met4 ;
        RECT 6.635000 27.290000 6.955000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 27.720000 6.955000 28.040000 ;
      LAYER met4 ;
        RECT 6.635000 27.720000 6.955000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 28.150000 6.955000 28.470000 ;
      LAYER met4 ;
        RECT 6.635000 28.150000 6.955000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 181.445000 7.275000 181.765000 ;
      LAYER met4 ;
        RECT 6.955000 181.445000 7.275000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 181.850000 7.275000 182.170000 ;
      LAYER met4 ;
        RECT 6.955000 181.850000 7.275000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 182.255000 7.275000 182.575000 ;
      LAYER met4 ;
        RECT 6.955000 182.255000 7.275000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 182.660000 7.275000 182.980000 ;
      LAYER met4 ;
        RECT 6.955000 182.660000 7.275000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 183.065000 7.275000 183.385000 ;
      LAYER met4 ;
        RECT 6.955000 183.065000 7.275000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 183.470000 7.275000 183.790000 ;
      LAYER met4 ;
        RECT 6.955000 183.470000 7.275000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 183.875000 7.275000 184.195000 ;
      LAYER met4 ;
        RECT 6.955000 183.875000 7.275000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 184.280000 7.275000 184.600000 ;
      LAYER met4 ;
        RECT 6.955000 184.280000 7.275000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 184.685000 7.275000 185.005000 ;
      LAYER met4 ;
        RECT 6.955000 184.685000 7.275000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 185.090000 7.275000 185.410000 ;
      LAYER met4 ;
        RECT 6.955000 185.090000 7.275000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 185.495000 7.275000 185.815000 ;
      LAYER met4 ;
        RECT 6.955000 185.495000 7.275000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 185.900000 7.275000 186.220000 ;
      LAYER met4 ;
        RECT 6.955000 185.900000 7.275000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 186.305000 7.275000 186.625000 ;
      LAYER met4 ;
        RECT 6.955000 186.305000 7.275000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 186.710000 7.275000 187.030000 ;
      LAYER met4 ;
        RECT 6.955000 186.710000 7.275000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 187.115000 7.275000 187.435000 ;
      LAYER met4 ;
        RECT 6.955000 187.115000 7.275000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 187.520000 7.275000 187.840000 ;
      LAYER met4 ;
        RECT 6.955000 187.520000 7.275000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 187.925000 7.275000 188.245000 ;
      LAYER met4 ;
        RECT 6.955000 187.925000 7.275000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 188.330000 7.275000 188.650000 ;
      LAYER met4 ;
        RECT 6.955000 188.330000 7.275000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 188.735000 7.275000 189.055000 ;
      LAYER met4 ;
        RECT 6.955000 188.735000 7.275000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 189.140000 7.275000 189.460000 ;
      LAYER met4 ;
        RECT 6.955000 189.140000 7.275000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 189.545000 7.275000 189.865000 ;
      LAYER met4 ;
        RECT 6.955000 189.545000 7.275000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 189.950000 7.275000 190.270000 ;
      LAYER met4 ;
        RECT 6.955000 189.950000 7.275000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 190.355000 7.275000 190.675000 ;
      LAYER met4 ;
        RECT 6.955000 190.355000 7.275000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 190.760000 7.275000 191.080000 ;
      LAYER met4 ;
        RECT 6.955000 190.760000 7.275000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 191.165000 7.275000 191.485000 ;
      LAYER met4 ;
        RECT 6.955000 191.165000 7.275000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 191.570000 7.275000 191.890000 ;
      LAYER met4 ;
        RECT 6.955000 191.570000 7.275000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 191.975000 7.275000 192.295000 ;
      LAYER met4 ;
        RECT 6.955000 191.975000 7.275000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 192.380000 7.275000 192.700000 ;
      LAYER met4 ;
        RECT 6.955000 192.380000 7.275000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 192.785000 7.275000 193.105000 ;
      LAYER met4 ;
        RECT 6.955000 192.785000 7.275000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 193.190000 7.275000 193.510000 ;
      LAYER met4 ;
        RECT 6.955000 193.190000 7.275000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 193.595000 7.275000 193.915000 ;
      LAYER met4 ;
        RECT 6.955000 193.595000 7.275000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 194.000000 7.275000 194.320000 ;
      LAYER met4 ;
        RECT 6.955000 194.000000 7.275000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 194.405000 7.275000 194.725000 ;
      LAYER met4 ;
        RECT 6.955000 194.405000 7.275000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 194.810000 7.275000 195.130000 ;
      LAYER met4 ;
        RECT 6.955000 194.810000 7.275000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 195.215000 7.275000 195.535000 ;
      LAYER met4 ;
        RECT 6.955000 195.215000 7.275000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 195.620000 7.275000 195.940000 ;
      LAYER met4 ;
        RECT 6.955000 195.620000 7.275000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 196.025000 7.275000 196.345000 ;
      LAYER met4 ;
        RECT 6.955000 196.025000 7.275000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 196.430000 7.275000 196.750000 ;
      LAYER met4 ;
        RECT 6.955000 196.430000 7.275000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 196.835000 7.275000 197.155000 ;
      LAYER met4 ;
        RECT 6.955000 196.835000 7.275000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 197.240000 7.275000 197.560000 ;
      LAYER met4 ;
        RECT 6.955000 197.240000 7.275000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955000 197.645000 7.275000 197.965000 ;
      LAYER met4 ;
        RECT 6.955000 197.645000 7.275000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 23.850000 60.490000 24.170000 ;
      LAYER met4 ;
        RECT 60.170000 23.850000 60.490000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 24.280000 60.490000 24.600000 ;
      LAYER met4 ;
        RECT 60.170000 24.280000 60.490000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 24.710000 60.490000 25.030000 ;
      LAYER met4 ;
        RECT 60.170000 24.710000 60.490000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 25.140000 60.490000 25.460000 ;
      LAYER met4 ;
        RECT 60.170000 25.140000 60.490000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 25.570000 60.490000 25.890000 ;
      LAYER met4 ;
        RECT 60.170000 25.570000 60.490000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 26.000000 60.490000 26.320000 ;
      LAYER met4 ;
        RECT 60.170000 26.000000 60.490000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 26.430000 60.490000 26.750000 ;
      LAYER met4 ;
        RECT 60.170000 26.430000 60.490000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 26.860000 60.490000 27.180000 ;
      LAYER met4 ;
        RECT 60.170000 26.860000 60.490000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 27.290000 60.490000 27.610000 ;
      LAYER met4 ;
        RECT 60.170000 27.290000 60.490000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 27.720000 60.490000 28.040000 ;
      LAYER met4 ;
        RECT 60.170000 27.720000 60.490000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 28.150000 60.490000 28.470000 ;
      LAYER met4 ;
        RECT 60.170000 28.150000 60.490000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 23.850000 60.895000 24.170000 ;
      LAYER met4 ;
        RECT 60.575000 23.850000 60.895000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 24.280000 60.895000 24.600000 ;
      LAYER met4 ;
        RECT 60.575000 24.280000 60.895000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 24.710000 60.895000 25.030000 ;
      LAYER met4 ;
        RECT 60.575000 24.710000 60.895000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 25.140000 60.895000 25.460000 ;
      LAYER met4 ;
        RECT 60.575000 25.140000 60.895000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 25.570000 60.895000 25.890000 ;
      LAYER met4 ;
        RECT 60.575000 25.570000 60.895000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 26.000000 60.895000 26.320000 ;
      LAYER met4 ;
        RECT 60.575000 26.000000 60.895000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 26.430000 60.895000 26.750000 ;
      LAYER met4 ;
        RECT 60.575000 26.430000 60.895000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 26.860000 60.895000 27.180000 ;
      LAYER met4 ;
        RECT 60.575000 26.860000 60.895000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 27.290000 60.895000 27.610000 ;
      LAYER met4 ;
        RECT 60.575000 27.290000 60.895000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 27.720000 60.895000 28.040000 ;
      LAYER met4 ;
        RECT 60.575000 27.720000 60.895000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 28.150000 60.895000 28.470000 ;
      LAYER met4 ;
        RECT 60.575000 28.150000 60.895000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 23.850000 61.300000 24.170000 ;
      LAYER met4 ;
        RECT 60.980000 23.850000 61.300000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 24.280000 61.300000 24.600000 ;
      LAYER met4 ;
        RECT 60.980000 24.280000 61.300000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 24.710000 61.300000 25.030000 ;
      LAYER met4 ;
        RECT 60.980000 24.710000 61.300000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 25.140000 61.300000 25.460000 ;
      LAYER met4 ;
        RECT 60.980000 25.140000 61.300000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 25.570000 61.300000 25.890000 ;
      LAYER met4 ;
        RECT 60.980000 25.570000 61.300000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 26.000000 61.300000 26.320000 ;
      LAYER met4 ;
        RECT 60.980000 26.000000 61.300000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 26.430000 61.300000 26.750000 ;
      LAYER met4 ;
        RECT 60.980000 26.430000 61.300000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 26.860000 61.300000 27.180000 ;
      LAYER met4 ;
        RECT 60.980000 26.860000 61.300000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 27.290000 61.300000 27.610000 ;
      LAYER met4 ;
        RECT 60.980000 27.290000 61.300000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 27.720000 61.300000 28.040000 ;
      LAYER met4 ;
        RECT 60.980000 27.720000 61.300000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 28.150000 61.300000 28.470000 ;
      LAYER met4 ;
        RECT 60.980000 28.150000 61.300000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 23.850000 61.705000 24.170000 ;
      LAYER met4 ;
        RECT 61.385000 23.850000 61.705000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 24.280000 61.705000 24.600000 ;
      LAYER met4 ;
        RECT 61.385000 24.280000 61.705000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 24.710000 61.705000 25.030000 ;
      LAYER met4 ;
        RECT 61.385000 24.710000 61.705000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 25.140000 61.705000 25.460000 ;
      LAYER met4 ;
        RECT 61.385000 25.140000 61.705000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 25.570000 61.705000 25.890000 ;
      LAYER met4 ;
        RECT 61.385000 25.570000 61.705000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 26.000000 61.705000 26.320000 ;
      LAYER met4 ;
        RECT 61.385000 26.000000 61.705000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 26.430000 61.705000 26.750000 ;
      LAYER met4 ;
        RECT 61.385000 26.430000 61.705000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 26.860000 61.705000 27.180000 ;
      LAYER met4 ;
        RECT 61.385000 26.860000 61.705000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 27.290000 61.705000 27.610000 ;
      LAYER met4 ;
        RECT 61.385000 27.290000 61.705000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 27.720000 61.705000 28.040000 ;
      LAYER met4 ;
        RECT 61.385000 27.720000 61.705000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 28.150000 61.705000 28.470000 ;
      LAYER met4 ;
        RECT 61.385000 28.150000 61.705000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 23.850000 62.110000 24.170000 ;
      LAYER met4 ;
        RECT 61.790000 23.850000 62.110000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 24.280000 62.110000 24.600000 ;
      LAYER met4 ;
        RECT 61.790000 24.280000 62.110000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 24.710000 62.110000 25.030000 ;
      LAYER met4 ;
        RECT 61.790000 24.710000 62.110000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 25.140000 62.110000 25.460000 ;
      LAYER met4 ;
        RECT 61.790000 25.140000 62.110000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 25.570000 62.110000 25.890000 ;
      LAYER met4 ;
        RECT 61.790000 25.570000 62.110000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 26.000000 62.110000 26.320000 ;
      LAYER met4 ;
        RECT 61.790000 26.000000 62.110000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 26.430000 62.110000 26.750000 ;
      LAYER met4 ;
        RECT 61.790000 26.430000 62.110000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 26.860000 62.110000 27.180000 ;
      LAYER met4 ;
        RECT 61.790000 26.860000 62.110000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 27.290000 62.110000 27.610000 ;
      LAYER met4 ;
        RECT 61.790000 27.290000 62.110000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 27.720000 62.110000 28.040000 ;
      LAYER met4 ;
        RECT 61.790000 27.720000 62.110000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 28.150000 62.110000 28.470000 ;
      LAYER met4 ;
        RECT 61.790000 28.150000 62.110000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 173.840000 62.400000 174.160000 ;
      LAYER met4 ;
        RECT 62.080000 173.840000 62.400000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 174.240000 62.400000 174.560000 ;
      LAYER met4 ;
        RECT 62.080000 174.240000 62.400000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 174.640000 62.400000 174.960000 ;
      LAYER met4 ;
        RECT 62.080000 174.640000 62.400000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 175.040000 62.400000 175.360000 ;
      LAYER met4 ;
        RECT 62.080000 175.040000 62.400000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 175.440000 62.400000 175.760000 ;
      LAYER met4 ;
        RECT 62.080000 175.440000 62.400000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 175.840000 62.400000 176.160000 ;
      LAYER met4 ;
        RECT 62.080000 175.840000 62.400000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 176.240000 62.400000 176.560000 ;
      LAYER met4 ;
        RECT 62.080000 176.240000 62.400000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 176.640000 62.400000 176.960000 ;
      LAYER met4 ;
        RECT 62.080000 176.640000 62.400000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 177.040000 62.400000 177.360000 ;
      LAYER met4 ;
        RECT 62.080000 177.040000 62.400000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 177.440000 62.400000 177.760000 ;
      LAYER met4 ;
        RECT 62.080000 177.440000 62.400000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 177.840000 62.400000 178.160000 ;
      LAYER met4 ;
        RECT 62.080000 177.840000 62.400000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 178.240000 62.400000 178.560000 ;
      LAYER met4 ;
        RECT 62.080000 178.240000 62.400000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 178.640000 62.400000 178.960000 ;
      LAYER met4 ;
        RECT 62.080000 178.640000 62.400000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 179.040000 62.400000 179.360000 ;
      LAYER met4 ;
        RECT 62.080000 179.040000 62.400000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 179.440000 62.400000 179.760000 ;
      LAYER met4 ;
        RECT 62.080000 179.440000 62.400000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 179.840000 62.400000 180.160000 ;
      LAYER met4 ;
        RECT 62.080000 179.840000 62.400000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 180.240000 62.400000 180.560000 ;
      LAYER met4 ;
        RECT 62.080000 180.240000 62.400000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 180.640000 62.400000 180.960000 ;
      LAYER met4 ;
        RECT 62.080000 180.640000 62.400000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 181.040000 62.400000 181.360000 ;
      LAYER met4 ;
        RECT 62.080000 181.040000 62.400000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 181.445000 62.400000 181.765000 ;
      LAYER met4 ;
        RECT 62.080000 181.445000 62.400000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 181.850000 62.400000 182.170000 ;
      LAYER met4 ;
        RECT 62.080000 181.850000 62.400000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 182.255000 62.400000 182.575000 ;
      LAYER met4 ;
        RECT 62.080000 182.255000 62.400000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 182.660000 62.400000 182.980000 ;
      LAYER met4 ;
        RECT 62.080000 182.660000 62.400000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 183.065000 62.400000 183.385000 ;
      LAYER met4 ;
        RECT 62.080000 183.065000 62.400000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 183.470000 62.400000 183.790000 ;
      LAYER met4 ;
        RECT 62.080000 183.470000 62.400000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 183.875000 62.400000 184.195000 ;
      LAYER met4 ;
        RECT 62.080000 183.875000 62.400000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 184.280000 62.400000 184.600000 ;
      LAYER met4 ;
        RECT 62.080000 184.280000 62.400000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 184.685000 62.400000 185.005000 ;
      LAYER met4 ;
        RECT 62.080000 184.685000 62.400000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 185.090000 62.400000 185.410000 ;
      LAYER met4 ;
        RECT 62.080000 185.090000 62.400000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 185.495000 62.400000 185.815000 ;
      LAYER met4 ;
        RECT 62.080000 185.495000 62.400000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 185.900000 62.400000 186.220000 ;
      LAYER met4 ;
        RECT 62.080000 185.900000 62.400000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 186.305000 62.400000 186.625000 ;
      LAYER met4 ;
        RECT 62.080000 186.305000 62.400000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 186.710000 62.400000 187.030000 ;
      LAYER met4 ;
        RECT 62.080000 186.710000 62.400000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 187.115000 62.400000 187.435000 ;
      LAYER met4 ;
        RECT 62.080000 187.115000 62.400000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 187.520000 62.400000 187.840000 ;
      LAYER met4 ;
        RECT 62.080000 187.520000 62.400000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 187.925000 62.400000 188.245000 ;
      LAYER met4 ;
        RECT 62.080000 187.925000 62.400000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 188.330000 62.400000 188.650000 ;
      LAYER met4 ;
        RECT 62.080000 188.330000 62.400000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 188.735000 62.400000 189.055000 ;
      LAYER met4 ;
        RECT 62.080000 188.735000 62.400000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 189.140000 62.400000 189.460000 ;
      LAYER met4 ;
        RECT 62.080000 189.140000 62.400000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 189.545000 62.400000 189.865000 ;
      LAYER met4 ;
        RECT 62.080000 189.545000 62.400000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 189.950000 62.400000 190.270000 ;
      LAYER met4 ;
        RECT 62.080000 189.950000 62.400000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 190.355000 62.400000 190.675000 ;
      LAYER met4 ;
        RECT 62.080000 190.355000 62.400000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 190.760000 62.400000 191.080000 ;
      LAYER met4 ;
        RECT 62.080000 190.760000 62.400000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 191.165000 62.400000 191.485000 ;
      LAYER met4 ;
        RECT 62.080000 191.165000 62.400000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 191.570000 62.400000 191.890000 ;
      LAYER met4 ;
        RECT 62.080000 191.570000 62.400000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 191.975000 62.400000 192.295000 ;
      LAYER met4 ;
        RECT 62.080000 191.975000 62.400000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 192.380000 62.400000 192.700000 ;
      LAYER met4 ;
        RECT 62.080000 192.380000 62.400000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 192.785000 62.400000 193.105000 ;
      LAYER met4 ;
        RECT 62.080000 192.785000 62.400000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 193.190000 62.400000 193.510000 ;
      LAYER met4 ;
        RECT 62.080000 193.190000 62.400000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 193.595000 62.400000 193.915000 ;
      LAYER met4 ;
        RECT 62.080000 193.595000 62.400000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 194.000000 62.400000 194.320000 ;
      LAYER met4 ;
        RECT 62.080000 194.000000 62.400000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 194.405000 62.400000 194.725000 ;
      LAYER met4 ;
        RECT 62.080000 194.405000 62.400000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 194.810000 62.400000 195.130000 ;
      LAYER met4 ;
        RECT 62.080000 194.810000 62.400000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 195.215000 62.400000 195.535000 ;
      LAYER met4 ;
        RECT 62.080000 195.215000 62.400000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 195.620000 62.400000 195.940000 ;
      LAYER met4 ;
        RECT 62.080000 195.620000 62.400000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 196.025000 62.400000 196.345000 ;
      LAYER met4 ;
        RECT 62.080000 196.025000 62.400000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 196.430000 62.400000 196.750000 ;
      LAYER met4 ;
        RECT 62.080000 196.430000 62.400000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 196.835000 62.400000 197.155000 ;
      LAYER met4 ;
        RECT 62.080000 196.835000 62.400000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 197.240000 62.400000 197.560000 ;
      LAYER met4 ;
        RECT 62.080000 197.240000 62.400000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.080000 197.645000 62.400000 197.965000 ;
      LAYER met4 ;
        RECT 62.080000 197.645000 62.400000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 23.850000 62.515000 24.170000 ;
      LAYER met4 ;
        RECT 62.195000 23.850000 62.515000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 24.280000 62.515000 24.600000 ;
      LAYER met4 ;
        RECT 62.195000 24.280000 62.515000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 24.710000 62.515000 25.030000 ;
      LAYER met4 ;
        RECT 62.195000 24.710000 62.515000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 25.140000 62.515000 25.460000 ;
      LAYER met4 ;
        RECT 62.195000 25.140000 62.515000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 25.570000 62.515000 25.890000 ;
      LAYER met4 ;
        RECT 62.195000 25.570000 62.515000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 26.000000 62.515000 26.320000 ;
      LAYER met4 ;
        RECT 62.195000 26.000000 62.515000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 26.430000 62.515000 26.750000 ;
      LAYER met4 ;
        RECT 62.195000 26.430000 62.515000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 26.860000 62.515000 27.180000 ;
      LAYER met4 ;
        RECT 62.195000 26.860000 62.515000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 27.290000 62.515000 27.610000 ;
      LAYER met4 ;
        RECT 62.195000 27.290000 62.515000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 27.720000 62.515000 28.040000 ;
      LAYER met4 ;
        RECT 62.195000 27.720000 62.515000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 28.150000 62.515000 28.470000 ;
      LAYER met4 ;
        RECT 62.195000 28.150000 62.515000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 173.840000 62.810000 174.160000 ;
      LAYER met4 ;
        RECT 62.490000 173.840000 62.810000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 174.240000 62.810000 174.560000 ;
      LAYER met4 ;
        RECT 62.490000 174.240000 62.810000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 174.640000 62.810000 174.960000 ;
      LAYER met4 ;
        RECT 62.490000 174.640000 62.810000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 175.040000 62.810000 175.360000 ;
      LAYER met4 ;
        RECT 62.490000 175.040000 62.810000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 175.440000 62.810000 175.760000 ;
      LAYER met4 ;
        RECT 62.490000 175.440000 62.810000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 175.840000 62.810000 176.160000 ;
      LAYER met4 ;
        RECT 62.490000 175.840000 62.810000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 176.240000 62.810000 176.560000 ;
      LAYER met4 ;
        RECT 62.490000 176.240000 62.810000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 176.640000 62.810000 176.960000 ;
      LAYER met4 ;
        RECT 62.490000 176.640000 62.810000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 177.040000 62.810000 177.360000 ;
      LAYER met4 ;
        RECT 62.490000 177.040000 62.810000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 177.440000 62.810000 177.760000 ;
      LAYER met4 ;
        RECT 62.490000 177.440000 62.810000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 177.840000 62.810000 178.160000 ;
      LAYER met4 ;
        RECT 62.490000 177.840000 62.810000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 178.240000 62.810000 178.560000 ;
      LAYER met4 ;
        RECT 62.490000 178.240000 62.810000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 178.640000 62.810000 178.960000 ;
      LAYER met4 ;
        RECT 62.490000 178.640000 62.810000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 179.040000 62.810000 179.360000 ;
      LAYER met4 ;
        RECT 62.490000 179.040000 62.810000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 179.440000 62.810000 179.760000 ;
      LAYER met4 ;
        RECT 62.490000 179.440000 62.810000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 179.840000 62.810000 180.160000 ;
      LAYER met4 ;
        RECT 62.490000 179.840000 62.810000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 180.240000 62.810000 180.560000 ;
      LAYER met4 ;
        RECT 62.490000 180.240000 62.810000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 180.640000 62.810000 180.960000 ;
      LAYER met4 ;
        RECT 62.490000 180.640000 62.810000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 181.040000 62.810000 181.360000 ;
      LAYER met4 ;
        RECT 62.490000 181.040000 62.810000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 181.445000 62.810000 181.765000 ;
      LAYER met4 ;
        RECT 62.490000 181.445000 62.810000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 181.850000 62.810000 182.170000 ;
      LAYER met4 ;
        RECT 62.490000 181.850000 62.810000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 182.255000 62.810000 182.575000 ;
      LAYER met4 ;
        RECT 62.490000 182.255000 62.810000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 182.660000 62.810000 182.980000 ;
      LAYER met4 ;
        RECT 62.490000 182.660000 62.810000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 183.065000 62.810000 183.385000 ;
      LAYER met4 ;
        RECT 62.490000 183.065000 62.810000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 183.470000 62.810000 183.790000 ;
      LAYER met4 ;
        RECT 62.490000 183.470000 62.810000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 183.875000 62.810000 184.195000 ;
      LAYER met4 ;
        RECT 62.490000 183.875000 62.810000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 184.280000 62.810000 184.600000 ;
      LAYER met4 ;
        RECT 62.490000 184.280000 62.810000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 184.685000 62.810000 185.005000 ;
      LAYER met4 ;
        RECT 62.490000 184.685000 62.810000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 185.090000 62.810000 185.410000 ;
      LAYER met4 ;
        RECT 62.490000 185.090000 62.810000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 185.495000 62.810000 185.815000 ;
      LAYER met4 ;
        RECT 62.490000 185.495000 62.810000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 185.900000 62.810000 186.220000 ;
      LAYER met4 ;
        RECT 62.490000 185.900000 62.810000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 186.305000 62.810000 186.625000 ;
      LAYER met4 ;
        RECT 62.490000 186.305000 62.810000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 186.710000 62.810000 187.030000 ;
      LAYER met4 ;
        RECT 62.490000 186.710000 62.810000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 187.115000 62.810000 187.435000 ;
      LAYER met4 ;
        RECT 62.490000 187.115000 62.810000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 187.520000 62.810000 187.840000 ;
      LAYER met4 ;
        RECT 62.490000 187.520000 62.810000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 187.925000 62.810000 188.245000 ;
      LAYER met4 ;
        RECT 62.490000 187.925000 62.810000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 188.330000 62.810000 188.650000 ;
      LAYER met4 ;
        RECT 62.490000 188.330000 62.810000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 188.735000 62.810000 189.055000 ;
      LAYER met4 ;
        RECT 62.490000 188.735000 62.810000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 189.140000 62.810000 189.460000 ;
      LAYER met4 ;
        RECT 62.490000 189.140000 62.810000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 189.545000 62.810000 189.865000 ;
      LAYER met4 ;
        RECT 62.490000 189.545000 62.810000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 189.950000 62.810000 190.270000 ;
      LAYER met4 ;
        RECT 62.490000 189.950000 62.810000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 190.355000 62.810000 190.675000 ;
      LAYER met4 ;
        RECT 62.490000 190.355000 62.810000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 190.760000 62.810000 191.080000 ;
      LAYER met4 ;
        RECT 62.490000 190.760000 62.810000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 191.165000 62.810000 191.485000 ;
      LAYER met4 ;
        RECT 62.490000 191.165000 62.810000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 191.570000 62.810000 191.890000 ;
      LAYER met4 ;
        RECT 62.490000 191.570000 62.810000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 191.975000 62.810000 192.295000 ;
      LAYER met4 ;
        RECT 62.490000 191.975000 62.810000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 192.380000 62.810000 192.700000 ;
      LAYER met4 ;
        RECT 62.490000 192.380000 62.810000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 192.785000 62.810000 193.105000 ;
      LAYER met4 ;
        RECT 62.490000 192.785000 62.810000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 193.190000 62.810000 193.510000 ;
      LAYER met4 ;
        RECT 62.490000 193.190000 62.810000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 193.595000 62.810000 193.915000 ;
      LAYER met4 ;
        RECT 62.490000 193.595000 62.810000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 194.000000 62.810000 194.320000 ;
      LAYER met4 ;
        RECT 62.490000 194.000000 62.810000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 194.405000 62.810000 194.725000 ;
      LAYER met4 ;
        RECT 62.490000 194.405000 62.810000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 194.810000 62.810000 195.130000 ;
      LAYER met4 ;
        RECT 62.490000 194.810000 62.810000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 195.215000 62.810000 195.535000 ;
      LAYER met4 ;
        RECT 62.490000 195.215000 62.810000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 195.620000 62.810000 195.940000 ;
      LAYER met4 ;
        RECT 62.490000 195.620000 62.810000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 196.025000 62.810000 196.345000 ;
      LAYER met4 ;
        RECT 62.490000 196.025000 62.810000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 196.430000 62.810000 196.750000 ;
      LAYER met4 ;
        RECT 62.490000 196.430000 62.810000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 196.835000 62.810000 197.155000 ;
      LAYER met4 ;
        RECT 62.490000 196.835000 62.810000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 197.240000 62.810000 197.560000 ;
      LAYER met4 ;
        RECT 62.490000 197.240000 62.810000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.490000 197.645000 62.810000 197.965000 ;
      LAYER met4 ;
        RECT 62.490000 197.645000 62.810000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 23.850000 62.920000 24.170000 ;
      LAYER met4 ;
        RECT 62.600000 23.850000 62.920000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 24.280000 62.920000 24.600000 ;
      LAYER met4 ;
        RECT 62.600000 24.280000 62.920000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 24.710000 62.920000 25.030000 ;
      LAYER met4 ;
        RECT 62.600000 24.710000 62.920000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 25.140000 62.920000 25.460000 ;
      LAYER met4 ;
        RECT 62.600000 25.140000 62.920000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 25.570000 62.920000 25.890000 ;
      LAYER met4 ;
        RECT 62.600000 25.570000 62.920000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 26.000000 62.920000 26.320000 ;
      LAYER met4 ;
        RECT 62.600000 26.000000 62.920000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 26.430000 62.920000 26.750000 ;
      LAYER met4 ;
        RECT 62.600000 26.430000 62.920000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 26.860000 62.920000 27.180000 ;
      LAYER met4 ;
        RECT 62.600000 26.860000 62.920000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 27.290000 62.920000 27.610000 ;
      LAYER met4 ;
        RECT 62.600000 27.290000 62.920000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 27.720000 62.920000 28.040000 ;
      LAYER met4 ;
        RECT 62.600000 27.720000 62.920000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 28.150000 62.920000 28.470000 ;
      LAYER met4 ;
        RECT 62.600000 28.150000 62.920000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 173.840000 63.220000 174.160000 ;
      LAYER met4 ;
        RECT 62.900000 173.840000 63.220000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 174.240000 63.220000 174.560000 ;
      LAYER met4 ;
        RECT 62.900000 174.240000 63.220000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 174.640000 63.220000 174.960000 ;
      LAYER met4 ;
        RECT 62.900000 174.640000 63.220000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 175.040000 63.220000 175.360000 ;
      LAYER met4 ;
        RECT 62.900000 175.040000 63.220000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 175.440000 63.220000 175.760000 ;
      LAYER met4 ;
        RECT 62.900000 175.440000 63.220000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 175.840000 63.220000 176.160000 ;
      LAYER met4 ;
        RECT 62.900000 175.840000 63.220000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 176.240000 63.220000 176.560000 ;
      LAYER met4 ;
        RECT 62.900000 176.240000 63.220000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 176.640000 63.220000 176.960000 ;
      LAYER met4 ;
        RECT 62.900000 176.640000 63.220000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 177.040000 63.220000 177.360000 ;
      LAYER met4 ;
        RECT 62.900000 177.040000 63.220000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 177.440000 63.220000 177.760000 ;
      LAYER met4 ;
        RECT 62.900000 177.440000 63.220000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 177.840000 63.220000 178.160000 ;
      LAYER met4 ;
        RECT 62.900000 177.840000 63.220000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 178.240000 63.220000 178.560000 ;
      LAYER met4 ;
        RECT 62.900000 178.240000 63.220000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 178.640000 63.220000 178.960000 ;
      LAYER met4 ;
        RECT 62.900000 178.640000 63.220000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 179.040000 63.220000 179.360000 ;
      LAYER met4 ;
        RECT 62.900000 179.040000 63.220000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 179.440000 63.220000 179.760000 ;
      LAYER met4 ;
        RECT 62.900000 179.440000 63.220000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 179.840000 63.220000 180.160000 ;
      LAYER met4 ;
        RECT 62.900000 179.840000 63.220000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 180.240000 63.220000 180.560000 ;
      LAYER met4 ;
        RECT 62.900000 180.240000 63.220000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 180.640000 63.220000 180.960000 ;
      LAYER met4 ;
        RECT 62.900000 180.640000 63.220000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 181.040000 63.220000 181.360000 ;
      LAYER met4 ;
        RECT 62.900000 181.040000 63.220000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 181.445000 63.220000 181.765000 ;
      LAYER met4 ;
        RECT 62.900000 181.445000 63.220000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 181.850000 63.220000 182.170000 ;
      LAYER met4 ;
        RECT 62.900000 181.850000 63.220000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 182.255000 63.220000 182.575000 ;
      LAYER met4 ;
        RECT 62.900000 182.255000 63.220000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 182.660000 63.220000 182.980000 ;
      LAYER met4 ;
        RECT 62.900000 182.660000 63.220000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 183.065000 63.220000 183.385000 ;
      LAYER met4 ;
        RECT 62.900000 183.065000 63.220000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 183.470000 63.220000 183.790000 ;
      LAYER met4 ;
        RECT 62.900000 183.470000 63.220000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 183.875000 63.220000 184.195000 ;
      LAYER met4 ;
        RECT 62.900000 183.875000 63.220000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 184.280000 63.220000 184.600000 ;
      LAYER met4 ;
        RECT 62.900000 184.280000 63.220000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 184.685000 63.220000 185.005000 ;
      LAYER met4 ;
        RECT 62.900000 184.685000 63.220000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 185.090000 63.220000 185.410000 ;
      LAYER met4 ;
        RECT 62.900000 185.090000 63.220000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 185.495000 63.220000 185.815000 ;
      LAYER met4 ;
        RECT 62.900000 185.495000 63.220000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 185.900000 63.220000 186.220000 ;
      LAYER met4 ;
        RECT 62.900000 185.900000 63.220000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 186.305000 63.220000 186.625000 ;
      LAYER met4 ;
        RECT 62.900000 186.305000 63.220000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 186.710000 63.220000 187.030000 ;
      LAYER met4 ;
        RECT 62.900000 186.710000 63.220000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 187.115000 63.220000 187.435000 ;
      LAYER met4 ;
        RECT 62.900000 187.115000 63.220000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 187.520000 63.220000 187.840000 ;
      LAYER met4 ;
        RECT 62.900000 187.520000 63.220000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 187.925000 63.220000 188.245000 ;
      LAYER met4 ;
        RECT 62.900000 187.925000 63.220000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 188.330000 63.220000 188.650000 ;
      LAYER met4 ;
        RECT 62.900000 188.330000 63.220000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 188.735000 63.220000 189.055000 ;
      LAYER met4 ;
        RECT 62.900000 188.735000 63.220000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 189.140000 63.220000 189.460000 ;
      LAYER met4 ;
        RECT 62.900000 189.140000 63.220000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 189.545000 63.220000 189.865000 ;
      LAYER met4 ;
        RECT 62.900000 189.545000 63.220000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 189.950000 63.220000 190.270000 ;
      LAYER met4 ;
        RECT 62.900000 189.950000 63.220000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 190.355000 63.220000 190.675000 ;
      LAYER met4 ;
        RECT 62.900000 190.355000 63.220000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 190.760000 63.220000 191.080000 ;
      LAYER met4 ;
        RECT 62.900000 190.760000 63.220000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 191.165000 63.220000 191.485000 ;
      LAYER met4 ;
        RECT 62.900000 191.165000 63.220000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 191.570000 63.220000 191.890000 ;
      LAYER met4 ;
        RECT 62.900000 191.570000 63.220000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 191.975000 63.220000 192.295000 ;
      LAYER met4 ;
        RECT 62.900000 191.975000 63.220000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 192.380000 63.220000 192.700000 ;
      LAYER met4 ;
        RECT 62.900000 192.380000 63.220000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 192.785000 63.220000 193.105000 ;
      LAYER met4 ;
        RECT 62.900000 192.785000 63.220000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 193.190000 63.220000 193.510000 ;
      LAYER met4 ;
        RECT 62.900000 193.190000 63.220000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 193.595000 63.220000 193.915000 ;
      LAYER met4 ;
        RECT 62.900000 193.595000 63.220000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 194.000000 63.220000 194.320000 ;
      LAYER met4 ;
        RECT 62.900000 194.000000 63.220000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 194.405000 63.220000 194.725000 ;
      LAYER met4 ;
        RECT 62.900000 194.405000 63.220000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 194.810000 63.220000 195.130000 ;
      LAYER met4 ;
        RECT 62.900000 194.810000 63.220000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 195.215000 63.220000 195.535000 ;
      LAYER met4 ;
        RECT 62.900000 195.215000 63.220000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 195.620000 63.220000 195.940000 ;
      LAYER met4 ;
        RECT 62.900000 195.620000 63.220000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 196.025000 63.220000 196.345000 ;
      LAYER met4 ;
        RECT 62.900000 196.025000 63.220000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 196.430000 63.220000 196.750000 ;
      LAYER met4 ;
        RECT 62.900000 196.430000 63.220000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 196.835000 63.220000 197.155000 ;
      LAYER met4 ;
        RECT 62.900000 196.835000 63.220000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 197.240000 63.220000 197.560000 ;
      LAYER met4 ;
        RECT 62.900000 197.240000 63.220000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.900000 197.645000 63.220000 197.965000 ;
      LAYER met4 ;
        RECT 62.900000 197.645000 63.220000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 23.850000 63.325000 24.170000 ;
      LAYER met4 ;
        RECT 63.005000 23.850000 63.325000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 24.280000 63.325000 24.600000 ;
      LAYER met4 ;
        RECT 63.005000 24.280000 63.325000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 24.710000 63.325000 25.030000 ;
      LAYER met4 ;
        RECT 63.005000 24.710000 63.325000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 25.140000 63.325000 25.460000 ;
      LAYER met4 ;
        RECT 63.005000 25.140000 63.325000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 25.570000 63.325000 25.890000 ;
      LAYER met4 ;
        RECT 63.005000 25.570000 63.325000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 26.000000 63.325000 26.320000 ;
      LAYER met4 ;
        RECT 63.005000 26.000000 63.325000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 26.430000 63.325000 26.750000 ;
      LAYER met4 ;
        RECT 63.005000 26.430000 63.325000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 26.860000 63.325000 27.180000 ;
      LAYER met4 ;
        RECT 63.005000 26.860000 63.325000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 27.290000 63.325000 27.610000 ;
      LAYER met4 ;
        RECT 63.005000 27.290000 63.325000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 27.720000 63.325000 28.040000 ;
      LAYER met4 ;
        RECT 63.005000 27.720000 63.325000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 28.150000 63.325000 28.470000 ;
      LAYER met4 ;
        RECT 63.005000 28.150000 63.325000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 173.840000 63.630000 174.160000 ;
      LAYER met4 ;
        RECT 63.310000 173.840000 63.630000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 174.240000 63.630000 174.560000 ;
      LAYER met4 ;
        RECT 63.310000 174.240000 63.630000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 174.640000 63.630000 174.960000 ;
      LAYER met4 ;
        RECT 63.310000 174.640000 63.630000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 175.040000 63.630000 175.360000 ;
      LAYER met4 ;
        RECT 63.310000 175.040000 63.630000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 175.440000 63.630000 175.760000 ;
      LAYER met4 ;
        RECT 63.310000 175.440000 63.630000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 175.840000 63.630000 176.160000 ;
      LAYER met4 ;
        RECT 63.310000 175.840000 63.630000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 176.240000 63.630000 176.560000 ;
      LAYER met4 ;
        RECT 63.310000 176.240000 63.630000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 176.640000 63.630000 176.960000 ;
      LAYER met4 ;
        RECT 63.310000 176.640000 63.630000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 177.040000 63.630000 177.360000 ;
      LAYER met4 ;
        RECT 63.310000 177.040000 63.630000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 177.440000 63.630000 177.760000 ;
      LAYER met4 ;
        RECT 63.310000 177.440000 63.630000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 177.840000 63.630000 178.160000 ;
      LAYER met4 ;
        RECT 63.310000 177.840000 63.630000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 178.240000 63.630000 178.560000 ;
      LAYER met4 ;
        RECT 63.310000 178.240000 63.630000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 178.640000 63.630000 178.960000 ;
      LAYER met4 ;
        RECT 63.310000 178.640000 63.630000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 179.040000 63.630000 179.360000 ;
      LAYER met4 ;
        RECT 63.310000 179.040000 63.630000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 179.440000 63.630000 179.760000 ;
      LAYER met4 ;
        RECT 63.310000 179.440000 63.630000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 179.840000 63.630000 180.160000 ;
      LAYER met4 ;
        RECT 63.310000 179.840000 63.630000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 180.240000 63.630000 180.560000 ;
      LAYER met4 ;
        RECT 63.310000 180.240000 63.630000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 180.640000 63.630000 180.960000 ;
      LAYER met4 ;
        RECT 63.310000 180.640000 63.630000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 181.040000 63.630000 181.360000 ;
      LAYER met4 ;
        RECT 63.310000 181.040000 63.630000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 181.445000 63.630000 181.765000 ;
      LAYER met4 ;
        RECT 63.310000 181.445000 63.630000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 181.850000 63.630000 182.170000 ;
      LAYER met4 ;
        RECT 63.310000 181.850000 63.630000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 182.255000 63.630000 182.575000 ;
      LAYER met4 ;
        RECT 63.310000 182.255000 63.630000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 182.660000 63.630000 182.980000 ;
      LAYER met4 ;
        RECT 63.310000 182.660000 63.630000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 183.065000 63.630000 183.385000 ;
      LAYER met4 ;
        RECT 63.310000 183.065000 63.630000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 183.470000 63.630000 183.790000 ;
      LAYER met4 ;
        RECT 63.310000 183.470000 63.630000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 183.875000 63.630000 184.195000 ;
      LAYER met4 ;
        RECT 63.310000 183.875000 63.630000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 184.280000 63.630000 184.600000 ;
      LAYER met4 ;
        RECT 63.310000 184.280000 63.630000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 184.685000 63.630000 185.005000 ;
      LAYER met4 ;
        RECT 63.310000 184.685000 63.630000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 185.090000 63.630000 185.410000 ;
      LAYER met4 ;
        RECT 63.310000 185.090000 63.630000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 185.495000 63.630000 185.815000 ;
      LAYER met4 ;
        RECT 63.310000 185.495000 63.630000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 185.900000 63.630000 186.220000 ;
      LAYER met4 ;
        RECT 63.310000 185.900000 63.630000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 186.305000 63.630000 186.625000 ;
      LAYER met4 ;
        RECT 63.310000 186.305000 63.630000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 186.710000 63.630000 187.030000 ;
      LAYER met4 ;
        RECT 63.310000 186.710000 63.630000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 187.115000 63.630000 187.435000 ;
      LAYER met4 ;
        RECT 63.310000 187.115000 63.630000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 187.520000 63.630000 187.840000 ;
      LAYER met4 ;
        RECT 63.310000 187.520000 63.630000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 187.925000 63.630000 188.245000 ;
      LAYER met4 ;
        RECT 63.310000 187.925000 63.630000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 188.330000 63.630000 188.650000 ;
      LAYER met4 ;
        RECT 63.310000 188.330000 63.630000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 188.735000 63.630000 189.055000 ;
      LAYER met4 ;
        RECT 63.310000 188.735000 63.630000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 189.140000 63.630000 189.460000 ;
      LAYER met4 ;
        RECT 63.310000 189.140000 63.630000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 189.545000 63.630000 189.865000 ;
      LAYER met4 ;
        RECT 63.310000 189.545000 63.630000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 189.950000 63.630000 190.270000 ;
      LAYER met4 ;
        RECT 63.310000 189.950000 63.630000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 190.355000 63.630000 190.675000 ;
      LAYER met4 ;
        RECT 63.310000 190.355000 63.630000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 190.760000 63.630000 191.080000 ;
      LAYER met4 ;
        RECT 63.310000 190.760000 63.630000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 191.165000 63.630000 191.485000 ;
      LAYER met4 ;
        RECT 63.310000 191.165000 63.630000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 191.570000 63.630000 191.890000 ;
      LAYER met4 ;
        RECT 63.310000 191.570000 63.630000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 191.975000 63.630000 192.295000 ;
      LAYER met4 ;
        RECT 63.310000 191.975000 63.630000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 192.380000 63.630000 192.700000 ;
      LAYER met4 ;
        RECT 63.310000 192.380000 63.630000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 192.785000 63.630000 193.105000 ;
      LAYER met4 ;
        RECT 63.310000 192.785000 63.630000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 193.190000 63.630000 193.510000 ;
      LAYER met4 ;
        RECT 63.310000 193.190000 63.630000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 193.595000 63.630000 193.915000 ;
      LAYER met4 ;
        RECT 63.310000 193.595000 63.630000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 194.000000 63.630000 194.320000 ;
      LAYER met4 ;
        RECT 63.310000 194.000000 63.630000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 194.405000 63.630000 194.725000 ;
      LAYER met4 ;
        RECT 63.310000 194.405000 63.630000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 194.810000 63.630000 195.130000 ;
      LAYER met4 ;
        RECT 63.310000 194.810000 63.630000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 195.215000 63.630000 195.535000 ;
      LAYER met4 ;
        RECT 63.310000 195.215000 63.630000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 195.620000 63.630000 195.940000 ;
      LAYER met4 ;
        RECT 63.310000 195.620000 63.630000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 196.025000 63.630000 196.345000 ;
      LAYER met4 ;
        RECT 63.310000 196.025000 63.630000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 196.430000 63.630000 196.750000 ;
      LAYER met4 ;
        RECT 63.310000 196.430000 63.630000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 196.835000 63.630000 197.155000 ;
      LAYER met4 ;
        RECT 63.310000 196.835000 63.630000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 197.240000 63.630000 197.560000 ;
      LAYER met4 ;
        RECT 63.310000 197.240000 63.630000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.310000 197.645000 63.630000 197.965000 ;
      LAYER met4 ;
        RECT 63.310000 197.645000 63.630000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 23.850000 63.730000 24.170000 ;
      LAYER met4 ;
        RECT 63.410000 23.850000 63.730000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 24.280000 63.730000 24.600000 ;
      LAYER met4 ;
        RECT 63.410000 24.280000 63.730000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 24.710000 63.730000 25.030000 ;
      LAYER met4 ;
        RECT 63.410000 24.710000 63.730000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 25.140000 63.730000 25.460000 ;
      LAYER met4 ;
        RECT 63.410000 25.140000 63.730000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 25.570000 63.730000 25.890000 ;
      LAYER met4 ;
        RECT 63.410000 25.570000 63.730000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 26.000000 63.730000 26.320000 ;
      LAYER met4 ;
        RECT 63.410000 26.000000 63.730000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 26.430000 63.730000 26.750000 ;
      LAYER met4 ;
        RECT 63.410000 26.430000 63.730000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 26.860000 63.730000 27.180000 ;
      LAYER met4 ;
        RECT 63.410000 26.860000 63.730000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 27.290000 63.730000 27.610000 ;
      LAYER met4 ;
        RECT 63.410000 27.290000 63.730000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 27.720000 63.730000 28.040000 ;
      LAYER met4 ;
        RECT 63.410000 27.720000 63.730000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 28.150000 63.730000 28.470000 ;
      LAYER met4 ;
        RECT 63.410000 28.150000 63.730000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 173.840000 64.040000 174.160000 ;
      LAYER met4 ;
        RECT 63.720000 173.840000 64.040000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 174.240000 64.040000 174.560000 ;
      LAYER met4 ;
        RECT 63.720000 174.240000 64.040000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 174.640000 64.040000 174.960000 ;
      LAYER met4 ;
        RECT 63.720000 174.640000 64.040000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 175.040000 64.040000 175.360000 ;
      LAYER met4 ;
        RECT 63.720000 175.040000 64.040000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 175.440000 64.040000 175.760000 ;
      LAYER met4 ;
        RECT 63.720000 175.440000 64.040000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 175.840000 64.040000 176.160000 ;
      LAYER met4 ;
        RECT 63.720000 175.840000 64.040000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 176.240000 64.040000 176.560000 ;
      LAYER met4 ;
        RECT 63.720000 176.240000 64.040000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 176.640000 64.040000 176.960000 ;
      LAYER met4 ;
        RECT 63.720000 176.640000 64.040000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 177.040000 64.040000 177.360000 ;
      LAYER met4 ;
        RECT 63.720000 177.040000 64.040000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 177.440000 64.040000 177.760000 ;
      LAYER met4 ;
        RECT 63.720000 177.440000 64.040000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 177.840000 64.040000 178.160000 ;
      LAYER met4 ;
        RECT 63.720000 177.840000 64.040000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 178.240000 64.040000 178.560000 ;
      LAYER met4 ;
        RECT 63.720000 178.240000 64.040000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 178.640000 64.040000 178.960000 ;
      LAYER met4 ;
        RECT 63.720000 178.640000 64.040000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 179.040000 64.040000 179.360000 ;
      LAYER met4 ;
        RECT 63.720000 179.040000 64.040000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 179.440000 64.040000 179.760000 ;
      LAYER met4 ;
        RECT 63.720000 179.440000 64.040000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 179.840000 64.040000 180.160000 ;
      LAYER met4 ;
        RECT 63.720000 179.840000 64.040000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 180.240000 64.040000 180.560000 ;
      LAYER met4 ;
        RECT 63.720000 180.240000 64.040000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 180.640000 64.040000 180.960000 ;
      LAYER met4 ;
        RECT 63.720000 180.640000 64.040000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 181.040000 64.040000 181.360000 ;
      LAYER met4 ;
        RECT 63.720000 181.040000 64.040000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 181.445000 64.040000 181.765000 ;
      LAYER met4 ;
        RECT 63.720000 181.445000 64.040000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 181.850000 64.040000 182.170000 ;
      LAYER met4 ;
        RECT 63.720000 181.850000 64.040000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 182.255000 64.040000 182.575000 ;
      LAYER met4 ;
        RECT 63.720000 182.255000 64.040000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 182.660000 64.040000 182.980000 ;
      LAYER met4 ;
        RECT 63.720000 182.660000 64.040000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 183.065000 64.040000 183.385000 ;
      LAYER met4 ;
        RECT 63.720000 183.065000 64.040000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 183.470000 64.040000 183.790000 ;
      LAYER met4 ;
        RECT 63.720000 183.470000 64.040000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 183.875000 64.040000 184.195000 ;
      LAYER met4 ;
        RECT 63.720000 183.875000 64.040000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 184.280000 64.040000 184.600000 ;
      LAYER met4 ;
        RECT 63.720000 184.280000 64.040000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 184.685000 64.040000 185.005000 ;
      LAYER met4 ;
        RECT 63.720000 184.685000 64.040000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 185.090000 64.040000 185.410000 ;
      LAYER met4 ;
        RECT 63.720000 185.090000 64.040000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 185.495000 64.040000 185.815000 ;
      LAYER met4 ;
        RECT 63.720000 185.495000 64.040000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 185.900000 64.040000 186.220000 ;
      LAYER met4 ;
        RECT 63.720000 185.900000 64.040000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 186.305000 64.040000 186.625000 ;
      LAYER met4 ;
        RECT 63.720000 186.305000 64.040000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 186.710000 64.040000 187.030000 ;
      LAYER met4 ;
        RECT 63.720000 186.710000 64.040000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 187.115000 64.040000 187.435000 ;
      LAYER met4 ;
        RECT 63.720000 187.115000 64.040000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 187.520000 64.040000 187.840000 ;
      LAYER met4 ;
        RECT 63.720000 187.520000 64.040000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 187.925000 64.040000 188.245000 ;
      LAYER met4 ;
        RECT 63.720000 187.925000 64.040000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 188.330000 64.040000 188.650000 ;
      LAYER met4 ;
        RECT 63.720000 188.330000 64.040000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 188.735000 64.040000 189.055000 ;
      LAYER met4 ;
        RECT 63.720000 188.735000 64.040000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 189.140000 64.040000 189.460000 ;
      LAYER met4 ;
        RECT 63.720000 189.140000 64.040000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 189.545000 64.040000 189.865000 ;
      LAYER met4 ;
        RECT 63.720000 189.545000 64.040000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 189.950000 64.040000 190.270000 ;
      LAYER met4 ;
        RECT 63.720000 189.950000 64.040000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 190.355000 64.040000 190.675000 ;
      LAYER met4 ;
        RECT 63.720000 190.355000 64.040000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 190.760000 64.040000 191.080000 ;
      LAYER met4 ;
        RECT 63.720000 190.760000 64.040000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 191.165000 64.040000 191.485000 ;
      LAYER met4 ;
        RECT 63.720000 191.165000 64.040000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 191.570000 64.040000 191.890000 ;
      LAYER met4 ;
        RECT 63.720000 191.570000 64.040000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 191.975000 64.040000 192.295000 ;
      LAYER met4 ;
        RECT 63.720000 191.975000 64.040000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 192.380000 64.040000 192.700000 ;
      LAYER met4 ;
        RECT 63.720000 192.380000 64.040000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 192.785000 64.040000 193.105000 ;
      LAYER met4 ;
        RECT 63.720000 192.785000 64.040000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 193.190000 64.040000 193.510000 ;
      LAYER met4 ;
        RECT 63.720000 193.190000 64.040000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 193.595000 64.040000 193.915000 ;
      LAYER met4 ;
        RECT 63.720000 193.595000 64.040000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 194.000000 64.040000 194.320000 ;
      LAYER met4 ;
        RECT 63.720000 194.000000 64.040000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 194.405000 64.040000 194.725000 ;
      LAYER met4 ;
        RECT 63.720000 194.405000 64.040000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 194.810000 64.040000 195.130000 ;
      LAYER met4 ;
        RECT 63.720000 194.810000 64.040000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 195.215000 64.040000 195.535000 ;
      LAYER met4 ;
        RECT 63.720000 195.215000 64.040000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 195.620000 64.040000 195.940000 ;
      LAYER met4 ;
        RECT 63.720000 195.620000 64.040000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 196.025000 64.040000 196.345000 ;
      LAYER met4 ;
        RECT 63.720000 196.025000 64.040000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 196.430000 64.040000 196.750000 ;
      LAYER met4 ;
        RECT 63.720000 196.430000 64.040000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 196.835000 64.040000 197.155000 ;
      LAYER met4 ;
        RECT 63.720000 196.835000 64.040000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 197.240000 64.040000 197.560000 ;
      LAYER met4 ;
        RECT 63.720000 197.240000 64.040000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.720000 197.645000 64.040000 197.965000 ;
      LAYER met4 ;
        RECT 63.720000 197.645000 64.040000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 23.850000 64.135000 24.170000 ;
      LAYER met4 ;
        RECT 63.815000 23.850000 64.135000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 24.280000 64.135000 24.600000 ;
      LAYER met4 ;
        RECT 63.815000 24.280000 64.135000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 24.710000 64.135000 25.030000 ;
      LAYER met4 ;
        RECT 63.815000 24.710000 64.135000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 25.140000 64.135000 25.460000 ;
      LAYER met4 ;
        RECT 63.815000 25.140000 64.135000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 25.570000 64.135000 25.890000 ;
      LAYER met4 ;
        RECT 63.815000 25.570000 64.135000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 26.000000 64.135000 26.320000 ;
      LAYER met4 ;
        RECT 63.815000 26.000000 64.135000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 26.430000 64.135000 26.750000 ;
      LAYER met4 ;
        RECT 63.815000 26.430000 64.135000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 26.860000 64.135000 27.180000 ;
      LAYER met4 ;
        RECT 63.815000 26.860000 64.135000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 27.290000 64.135000 27.610000 ;
      LAYER met4 ;
        RECT 63.815000 27.290000 64.135000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 27.720000 64.135000 28.040000 ;
      LAYER met4 ;
        RECT 63.815000 27.720000 64.135000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 28.150000 64.135000 28.470000 ;
      LAYER met4 ;
        RECT 63.815000 28.150000 64.135000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 173.840000 64.450000 174.160000 ;
      LAYER met4 ;
        RECT 64.130000 173.840000 64.450000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 174.240000 64.450000 174.560000 ;
      LAYER met4 ;
        RECT 64.130000 174.240000 64.450000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 174.640000 64.450000 174.960000 ;
      LAYER met4 ;
        RECT 64.130000 174.640000 64.450000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 175.040000 64.450000 175.360000 ;
      LAYER met4 ;
        RECT 64.130000 175.040000 64.450000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 175.440000 64.450000 175.760000 ;
      LAYER met4 ;
        RECT 64.130000 175.440000 64.450000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 175.840000 64.450000 176.160000 ;
      LAYER met4 ;
        RECT 64.130000 175.840000 64.450000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 176.240000 64.450000 176.560000 ;
      LAYER met4 ;
        RECT 64.130000 176.240000 64.450000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 176.640000 64.450000 176.960000 ;
      LAYER met4 ;
        RECT 64.130000 176.640000 64.450000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 177.040000 64.450000 177.360000 ;
      LAYER met4 ;
        RECT 64.130000 177.040000 64.450000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 177.440000 64.450000 177.760000 ;
      LAYER met4 ;
        RECT 64.130000 177.440000 64.450000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 177.840000 64.450000 178.160000 ;
      LAYER met4 ;
        RECT 64.130000 177.840000 64.450000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 178.240000 64.450000 178.560000 ;
      LAYER met4 ;
        RECT 64.130000 178.240000 64.450000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 178.640000 64.450000 178.960000 ;
      LAYER met4 ;
        RECT 64.130000 178.640000 64.450000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 179.040000 64.450000 179.360000 ;
      LAYER met4 ;
        RECT 64.130000 179.040000 64.450000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 179.440000 64.450000 179.760000 ;
      LAYER met4 ;
        RECT 64.130000 179.440000 64.450000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 179.840000 64.450000 180.160000 ;
      LAYER met4 ;
        RECT 64.130000 179.840000 64.450000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 180.240000 64.450000 180.560000 ;
      LAYER met4 ;
        RECT 64.130000 180.240000 64.450000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 180.640000 64.450000 180.960000 ;
      LAYER met4 ;
        RECT 64.130000 180.640000 64.450000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 181.040000 64.450000 181.360000 ;
      LAYER met4 ;
        RECT 64.130000 181.040000 64.450000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 181.445000 64.450000 181.765000 ;
      LAYER met4 ;
        RECT 64.130000 181.445000 64.450000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 181.850000 64.450000 182.170000 ;
      LAYER met4 ;
        RECT 64.130000 181.850000 64.450000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 182.255000 64.450000 182.575000 ;
      LAYER met4 ;
        RECT 64.130000 182.255000 64.450000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 182.660000 64.450000 182.980000 ;
      LAYER met4 ;
        RECT 64.130000 182.660000 64.450000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 183.065000 64.450000 183.385000 ;
      LAYER met4 ;
        RECT 64.130000 183.065000 64.450000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 183.470000 64.450000 183.790000 ;
      LAYER met4 ;
        RECT 64.130000 183.470000 64.450000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 183.875000 64.450000 184.195000 ;
      LAYER met4 ;
        RECT 64.130000 183.875000 64.450000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 184.280000 64.450000 184.600000 ;
      LAYER met4 ;
        RECT 64.130000 184.280000 64.450000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 184.685000 64.450000 185.005000 ;
      LAYER met4 ;
        RECT 64.130000 184.685000 64.450000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 185.090000 64.450000 185.410000 ;
      LAYER met4 ;
        RECT 64.130000 185.090000 64.450000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 185.495000 64.450000 185.815000 ;
      LAYER met4 ;
        RECT 64.130000 185.495000 64.450000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 185.900000 64.450000 186.220000 ;
      LAYER met4 ;
        RECT 64.130000 185.900000 64.450000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 186.305000 64.450000 186.625000 ;
      LAYER met4 ;
        RECT 64.130000 186.305000 64.450000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 186.710000 64.450000 187.030000 ;
      LAYER met4 ;
        RECT 64.130000 186.710000 64.450000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 187.115000 64.450000 187.435000 ;
      LAYER met4 ;
        RECT 64.130000 187.115000 64.450000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 187.520000 64.450000 187.840000 ;
      LAYER met4 ;
        RECT 64.130000 187.520000 64.450000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 187.925000 64.450000 188.245000 ;
      LAYER met4 ;
        RECT 64.130000 187.925000 64.450000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 188.330000 64.450000 188.650000 ;
      LAYER met4 ;
        RECT 64.130000 188.330000 64.450000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 188.735000 64.450000 189.055000 ;
      LAYER met4 ;
        RECT 64.130000 188.735000 64.450000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 189.140000 64.450000 189.460000 ;
      LAYER met4 ;
        RECT 64.130000 189.140000 64.450000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 189.545000 64.450000 189.865000 ;
      LAYER met4 ;
        RECT 64.130000 189.545000 64.450000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 189.950000 64.450000 190.270000 ;
      LAYER met4 ;
        RECT 64.130000 189.950000 64.450000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 190.355000 64.450000 190.675000 ;
      LAYER met4 ;
        RECT 64.130000 190.355000 64.450000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 190.760000 64.450000 191.080000 ;
      LAYER met4 ;
        RECT 64.130000 190.760000 64.450000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 191.165000 64.450000 191.485000 ;
      LAYER met4 ;
        RECT 64.130000 191.165000 64.450000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 191.570000 64.450000 191.890000 ;
      LAYER met4 ;
        RECT 64.130000 191.570000 64.450000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 191.975000 64.450000 192.295000 ;
      LAYER met4 ;
        RECT 64.130000 191.975000 64.450000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 192.380000 64.450000 192.700000 ;
      LAYER met4 ;
        RECT 64.130000 192.380000 64.450000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 192.785000 64.450000 193.105000 ;
      LAYER met4 ;
        RECT 64.130000 192.785000 64.450000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 193.190000 64.450000 193.510000 ;
      LAYER met4 ;
        RECT 64.130000 193.190000 64.450000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 193.595000 64.450000 193.915000 ;
      LAYER met4 ;
        RECT 64.130000 193.595000 64.450000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 194.000000 64.450000 194.320000 ;
      LAYER met4 ;
        RECT 64.130000 194.000000 64.450000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 194.405000 64.450000 194.725000 ;
      LAYER met4 ;
        RECT 64.130000 194.405000 64.450000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 194.810000 64.450000 195.130000 ;
      LAYER met4 ;
        RECT 64.130000 194.810000 64.450000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 195.215000 64.450000 195.535000 ;
      LAYER met4 ;
        RECT 64.130000 195.215000 64.450000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 195.620000 64.450000 195.940000 ;
      LAYER met4 ;
        RECT 64.130000 195.620000 64.450000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 196.025000 64.450000 196.345000 ;
      LAYER met4 ;
        RECT 64.130000 196.025000 64.450000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 196.430000 64.450000 196.750000 ;
      LAYER met4 ;
        RECT 64.130000 196.430000 64.450000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 196.835000 64.450000 197.155000 ;
      LAYER met4 ;
        RECT 64.130000 196.835000 64.450000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 197.240000 64.450000 197.560000 ;
      LAYER met4 ;
        RECT 64.130000 197.240000 64.450000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.130000 197.645000 64.450000 197.965000 ;
      LAYER met4 ;
        RECT 64.130000 197.645000 64.450000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 23.850000 64.540000 24.170000 ;
      LAYER met4 ;
        RECT 64.220000 23.850000 64.540000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 24.280000 64.540000 24.600000 ;
      LAYER met4 ;
        RECT 64.220000 24.280000 64.540000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 24.710000 64.540000 25.030000 ;
      LAYER met4 ;
        RECT 64.220000 24.710000 64.540000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 25.140000 64.540000 25.460000 ;
      LAYER met4 ;
        RECT 64.220000 25.140000 64.540000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 25.570000 64.540000 25.890000 ;
      LAYER met4 ;
        RECT 64.220000 25.570000 64.540000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 26.000000 64.540000 26.320000 ;
      LAYER met4 ;
        RECT 64.220000 26.000000 64.540000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 26.430000 64.540000 26.750000 ;
      LAYER met4 ;
        RECT 64.220000 26.430000 64.540000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 26.860000 64.540000 27.180000 ;
      LAYER met4 ;
        RECT 64.220000 26.860000 64.540000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 27.290000 64.540000 27.610000 ;
      LAYER met4 ;
        RECT 64.220000 27.290000 64.540000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 27.720000 64.540000 28.040000 ;
      LAYER met4 ;
        RECT 64.220000 27.720000 64.540000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 28.150000 64.540000 28.470000 ;
      LAYER met4 ;
        RECT 64.220000 28.150000 64.540000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 173.840000 64.860000 174.160000 ;
      LAYER met4 ;
        RECT 64.540000 173.840000 64.860000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 174.240000 64.860000 174.560000 ;
      LAYER met4 ;
        RECT 64.540000 174.240000 64.860000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 174.640000 64.860000 174.960000 ;
      LAYER met4 ;
        RECT 64.540000 174.640000 64.860000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 175.040000 64.860000 175.360000 ;
      LAYER met4 ;
        RECT 64.540000 175.040000 64.860000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 175.440000 64.860000 175.760000 ;
      LAYER met4 ;
        RECT 64.540000 175.440000 64.860000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 175.840000 64.860000 176.160000 ;
      LAYER met4 ;
        RECT 64.540000 175.840000 64.860000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 176.240000 64.860000 176.560000 ;
      LAYER met4 ;
        RECT 64.540000 176.240000 64.860000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 176.640000 64.860000 176.960000 ;
      LAYER met4 ;
        RECT 64.540000 176.640000 64.860000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 177.040000 64.860000 177.360000 ;
      LAYER met4 ;
        RECT 64.540000 177.040000 64.860000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 177.440000 64.860000 177.760000 ;
      LAYER met4 ;
        RECT 64.540000 177.440000 64.860000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 177.840000 64.860000 178.160000 ;
      LAYER met4 ;
        RECT 64.540000 177.840000 64.860000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 178.240000 64.860000 178.560000 ;
      LAYER met4 ;
        RECT 64.540000 178.240000 64.860000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 178.640000 64.860000 178.960000 ;
      LAYER met4 ;
        RECT 64.540000 178.640000 64.860000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 179.040000 64.860000 179.360000 ;
      LAYER met4 ;
        RECT 64.540000 179.040000 64.860000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 179.440000 64.860000 179.760000 ;
      LAYER met4 ;
        RECT 64.540000 179.440000 64.860000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 179.840000 64.860000 180.160000 ;
      LAYER met4 ;
        RECT 64.540000 179.840000 64.860000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 180.240000 64.860000 180.560000 ;
      LAYER met4 ;
        RECT 64.540000 180.240000 64.860000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 180.640000 64.860000 180.960000 ;
      LAYER met4 ;
        RECT 64.540000 180.640000 64.860000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 181.040000 64.860000 181.360000 ;
      LAYER met4 ;
        RECT 64.540000 181.040000 64.860000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 181.445000 64.860000 181.765000 ;
      LAYER met4 ;
        RECT 64.540000 181.445000 64.860000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 181.850000 64.860000 182.170000 ;
      LAYER met4 ;
        RECT 64.540000 181.850000 64.860000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 182.255000 64.860000 182.575000 ;
      LAYER met4 ;
        RECT 64.540000 182.255000 64.860000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 182.660000 64.860000 182.980000 ;
      LAYER met4 ;
        RECT 64.540000 182.660000 64.860000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 183.065000 64.860000 183.385000 ;
      LAYER met4 ;
        RECT 64.540000 183.065000 64.860000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 183.470000 64.860000 183.790000 ;
      LAYER met4 ;
        RECT 64.540000 183.470000 64.860000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 183.875000 64.860000 184.195000 ;
      LAYER met4 ;
        RECT 64.540000 183.875000 64.860000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 184.280000 64.860000 184.600000 ;
      LAYER met4 ;
        RECT 64.540000 184.280000 64.860000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 184.685000 64.860000 185.005000 ;
      LAYER met4 ;
        RECT 64.540000 184.685000 64.860000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 185.090000 64.860000 185.410000 ;
      LAYER met4 ;
        RECT 64.540000 185.090000 64.860000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 185.495000 64.860000 185.815000 ;
      LAYER met4 ;
        RECT 64.540000 185.495000 64.860000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 185.900000 64.860000 186.220000 ;
      LAYER met4 ;
        RECT 64.540000 185.900000 64.860000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 186.305000 64.860000 186.625000 ;
      LAYER met4 ;
        RECT 64.540000 186.305000 64.860000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 186.710000 64.860000 187.030000 ;
      LAYER met4 ;
        RECT 64.540000 186.710000 64.860000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 187.115000 64.860000 187.435000 ;
      LAYER met4 ;
        RECT 64.540000 187.115000 64.860000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 187.520000 64.860000 187.840000 ;
      LAYER met4 ;
        RECT 64.540000 187.520000 64.860000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 187.925000 64.860000 188.245000 ;
      LAYER met4 ;
        RECT 64.540000 187.925000 64.860000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 188.330000 64.860000 188.650000 ;
      LAYER met4 ;
        RECT 64.540000 188.330000 64.860000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 188.735000 64.860000 189.055000 ;
      LAYER met4 ;
        RECT 64.540000 188.735000 64.860000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 189.140000 64.860000 189.460000 ;
      LAYER met4 ;
        RECT 64.540000 189.140000 64.860000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 189.545000 64.860000 189.865000 ;
      LAYER met4 ;
        RECT 64.540000 189.545000 64.860000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 189.950000 64.860000 190.270000 ;
      LAYER met4 ;
        RECT 64.540000 189.950000 64.860000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 190.355000 64.860000 190.675000 ;
      LAYER met4 ;
        RECT 64.540000 190.355000 64.860000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 190.760000 64.860000 191.080000 ;
      LAYER met4 ;
        RECT 64.540000 190.760000 64.860000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 191.165000 64.860000 191.485000 ;
      LAYER met4 ;
        RECT 64.540000 191.165000 64.860000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 191.570000 64.860000 191.890000 ;
      LAYER met4 ;
        RECT 64.540000 191.570000 64.860000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 191.975000 64.860000 192.295000 ;
      LAYER met4 ;
        RECT 64.540000 191.975000 64.860000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 192.380000 64.860000 192.700000 ;
      LAYER met4 ;
        RECT 64.540000 192.380000 64.860000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 192.785000 64.860000 193.105000 ;
      LAYER met4 ;
        RECT 64.540000 192.785000 64.860000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 193.190000 64.860000 193.510000 ;
      LAYER met4 ;
        RECT 64.540000 193.190000 64.860000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 193.595000 64.860000 193.915000 ;
      LAYER met4 ;
        RECT 64.540000 193.595000 64.860000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 194.000000 64.860000 194.320000 ;
      LAYER met4 ;
        RECT 64.540000 194.000000 64.860000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 194.405000 64.860000 194.725000 ;
      LAYER met4 ;
        RECT 64.540000 194.405000 64.860000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 194.810000 64.860000 195.130000 ;
      LAYER met4 ;
        RECT 64.540000 194.810000 64.860000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 195.215000 64.860000 195.535000 ;
      LAYER met4 ;
        RECT 64.540000 195.215000 64.860000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 195.620000 64.860000 195.940000 ;
      LAYER met4 ;
        RECT 64.540000 195.620000 64.860000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 196.025000 64.860000 196.345000 ;
      LAYER met4 ;
        RECT 64.540000 196.025000 64.860000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 196.430000 64.860000 196.750000 ;
      LAYER met4 ;
        RECT 64.540000 196.430000 64.860000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 196.835000 64.860000 197.155000 ;
      LAYER met4 ;
        RECT 64.540000 196.835000 64.860000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 197.240000 64.860000 197.560000 ;
      LAYER met4 ;
        RECT 64.540000 197.240000 64.860000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.540000 197.645000 64.860000 197.965000 ;
      LAYER met4 ;
        RECT 64.540000 197.645000 64.860000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 23.850000 64.945000 24.170000 ;
      LAYER met4 ;
        RECT 64.625000 23.850000 64.945000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 24.280000 64.945000 24.600000 ;
      LAYER met4 ;
        RECT 64.625000 24.280000 64.945000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 24.710000 64.945000 25.030000 ;
      LAYER met4 ;
        RECT 64.625000 24.710000 64.945000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 25.140000 64.945000 25.460000 ;
      LAYER met4 ;
        RECT 64.625000 25.140000 64.945000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 25.570000 64.945000 25.890000 ;
      LAYER met4 ;
        RECT 64.625000 25.570000 64.945000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 26.000000 64.945000 26.320000 ;
      LAYER met4 ;
        RECT 64.625000 26.000000 64.945000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 26.430000 64.945000 26.750000 ;
      LAYER met4 ;
        RECT 64.625000 26.430000 64.945000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 26.860000 64.945000 27.180000 ;
      LAYER met4 ;
        RECT 64.625000 26.860000 64.945000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 27.290000 64.945000 27.610000 ;
      LAYER met4 ;
        RECT 64.625000 27.290000 64.945000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 27.720000 64.945000 28.040000 ;
      LAYER met4 ;
        RECT 64.625000 27.720000 64.945000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 28.150000 64.945000 28.470000 ;
      LAYER met4 ;
        RECT 64.625000 28.150000 64.945000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 173.840000 65.270000 174.160000 ;
      LAYER met4 ;
        RECT 64.950000 173.840000 65.270000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 174.240000 65.270000 174.560000 ;
      LAYER met4 ;
        RECT 64.950000 174.240000 65.270000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 174.640000 65.270000 174.960000 ;
      LAYER met4 ;
        RECT 64.950000 174.640000 65.270000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 175.040000 65.270000 175.360000 ;
      LAYER met4 ;
        RECT 64.950000 175.040000 65.270000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 175.440000 65.270000 175.760000 ;
      LAYER met4 ;
        RECT 64.950000 175.440000 65.270000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 175.840000 65.270000 176.160000 ;
      LAYER met4 ;
        RECT 64.950000 175.840000 65.270000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 176.240000 65.270000 176.560000 ;
      LAYER met4 ;
        RECT 64.950000 176.240000 65.270000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 176.640000 65.270000 176.960000 ;
      LAYER met4 ;
        RECT 64.950000 176.640000 65.270000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 177.040000 65.270000 177.360000 ;
      LAYER met4 ;
        RECT 64.950000 177.040000 65.270000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 177.440000 65.270000 177.760000 ;
      LAYER met4 ;
        RECT 64.950000 177.440000 65.270000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 177.840000 65.270000 178.160000 ;
      LAYER met4 ;
        RECT 64.950000 177.840000 65.270000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 178.240000 65.270000 178.560000 ;
      LAYER met4 ;
        RECT 64.950000 178.240000 65.270000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 178.640000 65.270000 178.960000 ;
      LAYER met4 ;
        RECT 64.950000 178.640000 65.270000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 179.040000 65.270000 179.360000 ;
      LAYER met4 ;
        RECT 64.950000 179.040000 65.270000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 179.440000 65.270000 179.760000 ;
      LAYER met4 ;
        RECT 64.950000 179.440000 65.270000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 179.840000 65.270000 180.160000 ;
      LAYER met4 ;
        RECT 64.950000 179.840000 65.270000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 180.240000 65.270000 180.560000 ;
      LAYER met4 ;
        RECT 64.950000 180.240000 65.270000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 180.640000 65.270000 180.960000 ;
      LAYER met4 ;
        RECT 64.950000 180.640000 65.270000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 181.040000 65.270000 181.360000 ;
      LAYER met4 ;
        RECT 64.950000 181.040000 65.270000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 181.445000 65.270000 181.765000 ;
      LAYER met4 ;
        RECT 64.950000 181.445000 65.270000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 181.850000 65.270000 182.170000 ;
      LAYER met4 ;
        RECT 64.950000 181.850000 65.270000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 182.255000 65.270000 182.575000 ;
      LAYER met4 ;
        RECT 64.950000 182.255000 65.270000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 182.660000 65.270000 182.980000 ;
      LAYER met4 ;
        RECT 64.950000 182.660000 65.270000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 183.065000 65.270000 183.385000 ;
      LAYER met4 ;
        RECT 64.950000 183.065000 65.270000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 183.470000 65.270000 183.790000 ;
      LAYER met4 ;
        RECT 64.950000 183.470000 65.270000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 183.875000 65.270000 184.195000 ;
      LAYER met4 ;
        RECT 64.950000 183.875000 65.270000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 184.280000 65.270000 184.600000 ;
      LAYER met4 ;
        RECT 64.950000 184.280000 65.270000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 184.685000 65.270000 185.005000 ;
      LAYER met4 ;
        RECT 64.950000 184.685000 65.270000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 185.090000 65.270000 185.410000 ;
      LAYER met4 ;
        RECT 64.950000 185.090000 65.270000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 185.495000 65.270000 185.815000 ;
      LAYER met4 ;
        RECT 64.950000 185.495000 65.270000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 185.900000 65.270000 186.220000 ;
      LAYER met4 ;
        RECT 64.950000 185.900000 65.270000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 186.305000 65.270000 186.625000 ;
      LAYER met4 ;
        RECT 64.950000 186.305000 65.270000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 186.710000 65.270000 187.030000 ;
      LAYER met4 ;
        RECT 64.950000 186.710000 65.270000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 187.115000 65.270000 187.435000 ;
      LAYER met4 ;
        RECT 64.950000 187.115000 65.270000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 187.520000 65.270000 187.840000 ;
      LAYER met4 ;
        RECT 64.950000 187.520000 65.270000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 187.925000 65.270000 188.245000 ;
      LAYER met4 ;
        RECT 64.950000 187.925000 65.270000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 188.330000 65.270000 188.650000 ;
      LAYER met4 ;
        RECT 64.950000 188.330000 65.270000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 188.735000 65.270000 189.055000 ;
      LAYER met4 ;
        RECT 64.950000 188.735000 65.270000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 189.140000 65.270000 189.460000 ;
      LAYER met4 ;
        RECT 64.950000 189.140000 65.270000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 189.545000 65.270000 189.865000 ;
      LAYER met4 ;
        RECT 64.950000 189.545000 65.270000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 189.950000 65.270000 190.270000 ;
      LAYER met4 ;
        RECT 64.950000 189.950000 65.270000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 190.355000 65.270000 190.675000 ;
      LAYER met4 ;
        RECT 64.950000 190.355000 65.270000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 190.760000 65.270000 191.080000 ;
      LAYER met4 ;
        RECT 64.950000 190.760000 65.270000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 191.165000 65.270000 191.485000 ;
      LAYER met4 ;
        RECT 64.950000 191.165000 65.270000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 191.570000 65.270000 191.890000 ;
      LAYER met4 ;
        RECT 64.950000 191.570000 65.270000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 191.975000 65.270000 192.295000 ;
      LAYER met4 ;
        RECT 64.950000 191.975000 65.270000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 192.380000 65.270000 192.700000 ;
      LAYER met4 ;
        RECT 64.950000 192.380000 65.270000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 192.785000 65.270000 193.105000 ;
      LAYER met4 ;
        RECT 64.950000 192.785000 65.270000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 193.190000 65.270000 193.510000 ;
      LAYER met4 ;
        RECT 64.950000 193.190000 65.270000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 193.595000 65.270000 193.915000 ;
      LAYER met4 ;
        RECT 64.950000 193.595000 65.270000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 194.000000 65.270000 194.320000 ;
      LAYER met4 ;
        RECT 64.950000 194.000000 65.270000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 194.405000 65.270000 194.725000 ;
      LAYER met4 ;
        RECT 64.950000 194.405000 65.270000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 194.810000 65.270000 195.130000 ;
      LAYER met4 ;
        RECT 64.950000 194.810000 65.270000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 195.215000 65.270000 195.535000 ;
      LAYER met4 ;
        RECT 64.950000 195.215000 65.270000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 195.620000 65.270000 195.940000 ;
      LAYER met4 ;
        RECT 64.950000 195.620000 65.270000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 196.025000 65.270000 196.345000 ;
      LAYER met4 ;
        RECT 64.950000 196.025000 65.270000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 196.430000 65.270000 196.750000 ;
      LAYER met4 ;
        RECT 64.950000 196.430000 65.270000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 196.835000 65.270000 197.155000 ;
      LAYER met4 ;
        RECT 64.950000 196.835000 65.270000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 197.240000 65.270000 197.560000 ;
      LAYER met4 ;
        RECT 64.950000 197.240000 65.270000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 197.645000 65.270000 197.965000 ;
      LAYER met4 ;
        RECT 64.950000 197.645000 65.270000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 23.850000 65.350000 24.170000 ;
      LAYER met4 ;
        RECT 65.030000 23.850000 65.350000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 24.280000 65.350000 24.600000 ;
      LAYER met4 ;
        RECT 65.030000 24.280000 65.350000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 24.710000 65.350000 25.030000 ;
      LAYER met4 ;
        RECT 65.030000 24.710000 65.350000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 25.140000 65.350000 25.460000 ;
      LAYER met4 ;
        RECT 65.030000 25.140000 65.350000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 25.570000 65.350000 25.890000 ;
      LAYER met4 ;
        RECT 65.030000 25.570000 65.350000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 26.000000 65.350000 26.320000 ;
      LAYER met4 ;
        RECT 65.030000 26.000000 65.350000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 26.430000 65.350000 26.750000 ;
      LAYER met4 ;
        RECT 65.030000 26.430000 65.350000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 26.860000 65.350000 27.180000 ;
      LAYER met4 ;
        RECT 65.030000 26.860000 65.350000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 27.290000 65.350000 27.610000 ;
      LAYER met4 ;
        RECT 65.030000 27.290000 65.350000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 27.720000 65.350000 28.040000 ;
      LAYER met4 ;
        RECT 65.030000 27.720000 65.350000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 28.150000 65.350000 28.470000 ;
      LAYER met4 ;
        RECT 65.030000 28.150000 65.350000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 173.840000 65.680000 174.160000 ;
      LAYER met4 ;
        RECT 65.360000 173.840000 65.680000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 174.240000 65.680000 174.560000 ;
      LAYER met4 ;
        RECT 65.360000 174.240000 65.680000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 174.640000 65.680000 174.960000 ;
      LAYER met4 ;
        RECT 65.360000 174.640000 65.680000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 175.040000 65.680000 175.360000 ;
      LAYER met4 ;
        RECT 65.360000 175.040000 65.680000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 175.440000 65.680000 175.760000 ;
      LAYER met4 ;
        RECT 65.360000 175.440000 65.680000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 175.840000 65.680000 176.160000 ;
      LAYER met4 ;
        RECT 65.360000 175.840000 65.680000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 176.240000 65.680000 176.560000 ;
      LAYER met4 ;
        RECT 65.360000 176.240000 65.680000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 176.640000 65.680000 176.960000 ;
      LAYER met4 ;
        RECT 65.360000 176.640000 65.680000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 177.040000 65.680000 177.360000 ;
      LAYER met4 ;
        RECT 65.360000 177.040000 65.680000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 177.440000 65.680000 177.760000 ;
      LAYER met4 ;
        RECT 65.360000 177.440000 65.680000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 177.840000 65.680000 178.160000 ;
      LAYER met4 ;
        RECT 65.360000 177.840000 65.680000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 178.240000 65.680000 178.560000 ;
      LAYER met4 ;
        RECT 65.360000 178.240000 65.680000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 178.640000 65.680000 178.960000 ;
      LAYER met4 ;
        RECT 65.360000 178.640000 65.680000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 179.040000 65.680000 179.360000 ;
      LAYER met4 ;
        RECT 65.360000 179.040000 65.680000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 179.440000 65.680000 179.760000 ;
      LAYER met4 ;
        RECT 65.360000 179.440000 65.680000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 179.840000 65.680000 180.160000 ;
      LAYER met4 ;
        RECT 65.360000 179.840000 65.680000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 180.240000 65.680000 180.560000 ;
      LAYER met4 ;
        RECT 65.360000 180.240000 65.680000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 180.640000 65.680000 180.960000 ;
      LAYER met4 ;
        RECT 65.360000 180.640000 65.680000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 181.040000 65.680000 181.360000 ;
      LAYER met4 ;
        RECT 65.360000 181.040000 65.680000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 181.445000 65.680000 181.765000 ;
      LAYER met4 ;
        RECT 65.360000 181.445000 65.680000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 181.850000 65.680000 182.170000 ;
      LAYER met4 ;
        RECT 65.360000 181.850000 65.680000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 182.255000 65.680000 182.575000 ;
      LAYER met4 ;
        RECT 65.360000 182.255000 65.680000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 182.660000 65.680000 182.980000 ;
      LAYER met4 ;
        RECT 65.360000 182.660000 65.680000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 183.065000 65.680000 183.385000 ;
      LAYER met4 ;
        RECT 65.360000 183.065000 65.680000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 183.470000 65.680000 183.790000 ;
      LAYER met4 ;
        RECT 65.360000 183.470000 65.680000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 183.875000 65.680000 184.195000 ;
      LAYER met4 ;
        RECT 65.360000 183.875000 65.680000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 184.280000 65.680000 184.600000 ;
      LAYER met4 ;
        RECT 65.360000 184.280000 65.680000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 184.685000 65.680000 185.005000 ;
      LAYER met4 ;
        RECT 65.360000 184.685000 65.680000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 185.090000 65.680000 185.410000 ;
      LAYER met4 ;
        RECT 65.360000 185.090000 65.680000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 185.495000 65.680000 185.815000 ;
      LAYER met4 ;
        RECT 65.360000 185.495000 65.680000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 185.900000 65.680000 186.220000 ;
      LAYER met4 ;
        RECT 65.360000 185.900000 65.680000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 186.305000 65.680000 186.625000 ;
      LAYER met4 ;
        RECT 65.360000 186.305000 65.680000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 186.710000 65.680000 187.030000 ;
      LAYER met4 ;
        RECT 65.360000 186.710000 65.680000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 187.115000 65.680000 187.435000 ;
      LAYER met4 ;
        RECT 65.360000 187.115000 65.680000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 187.520000 65.680000 187.840000 ;
      LAYER met4 ;
        RECT 65.360000 187.520000 65.680000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 187.925000 65.680000 188.245000 ;
      LAYER met4 ;
        RECT 65.360000 187.925000 65.680000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 188.330000 65.680000 188.650000 ;
      LAYER met4 ;
        RECT 65.360000 188.330000 65.680000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 188.735000 65.680000 189.055000 ;
      LAYER met4 ;
        RECT 65.360000 188.735000 65.680000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 189.140000 65.680000 189.460000 ;
      LAYER met4 ;
        RECT 65.360000 189.140000 65.680000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 189.545000 65.680000 189.865000 ;
      LAYER met4 ;
        RECT 65.360000 189.545000 65.680000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 189.950000 65.680000 190.270000 ;
      LAYER met4 ;
        RECT 65.360000 189.950000 65.680000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 190.355000 65.680000 190.675000 ;
      LAYER met4 ;
        RECT 65.360000 190.355000 65.680000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 190.760000 65.680000 191.080000 ;
      LAYER met4 ;
        RECT 65.360000 190.760000 65.680000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 191.165000 65.680000 191.485000 ;
      LAYER met4 ;
        RECT 65.360000 191.165000 65.680000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 191.570000 65.680000 191.890000 ;
      LAYER met4 ;
        RECT 65.360000 191.570000 65.680000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 191.975000 65.680000 192.295000 ;
      LAYER met4 ;
        RECT 65.360000 191.975000 65.680000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 192.380000 65.680000 192.700000 ;
      LAYER met4 ;
        RECT 65.360000 192.380000 65.680000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 192.785000 65.680000 193.105000 ;
      LAYER met4 ;
        RECT 65.360000 192.785000 65.680000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 193.190000 65.680000 193.510000 ;
      LAYER met4 ;
        RECT 65.360000 193.190000 65.680000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 193.595000 65.680000 193.915000 ;
      LAYER met4 ;
        RECT 65.360000 193.595000 65.680000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 194.000000 65.680000 194.320000 ;
      LAYER met4 ;
        RECT 65.360000 194.000000 65.680000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 194.405000 65.680000 194.725000 ;
      LAYER met4 ;
        RECT 65.360000 194.405000 65.680000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 194.810000 65.680000 195.130000 ;
      LAYER met4 ;
        RECT 65.360000 194.810000 65.680000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 195.215000 65.680000 195.535000 ;
      LAYER met4 ;
        RECT 65.360000 195.215000 65.680000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 195.620000 65.680000 195.940000 ;
      LAYER met4 ;
        RECT 65.360000 195.620000 65.680000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 196.025000 65.680000 196.345000 ;
      LAYER met4 ;
        RECT 65.360000 196.025000 65.680000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 196.430000 65.680000 196.750000 ;
      LAYER met4 ;
        RECT 65.360000 196.430000 65.680000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 196.835000 65.680000 197.155000 ;
      LAYER met4 ;
        RECT 65.360000 196.835000 65.680000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 197.240000 65.680000 197.560000 ;
      LAYER met4 ;
        RECT 65.360000 197.240000 65.680000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.360000 197.645000 65.680000 197.965000 ;
      LAYER met4 ;
        RECT 65.360000 197.645000 65.680000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 23.850000 65.755000 24.170000 ;
      LAYER met4 ;
        RECT 65.435000 23.850000 65.755000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 24.280000 65.755000 24.600000 ;
      LAYER met4 ;
        RECT 65.435000 24.280000 65.755000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 24.710000 65.755000 25.030000 ;
      LAYER met4 ;
        RECT 65.435000 24.710000 65.755000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 25.140000 65.755000 25.460000 ;
      LAYER met4 ;
        RECT 65.435000 25.140000 65.755000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 25.570000 65.755000 25.890000 ;
      LAYER met4 ;
        RECT 65.435000 25.570000 65.755000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 26.000000 65.755000 26.320000 ;
      LAYER met4 ;
        RECT 65.435000 26.000000 65.755000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 26.430000 65.755000 26.750000 ;
      LAYER met4 ;
        RECT 65.435000 26.430000 65.755000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 26.860000 65.755000 27.180000 ;
      LAYER met4 ;
        RECT 65.435000 26.860000 65.755000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 27.290000 65.755000 27.610000 ;
      LAYER met4 ;
        RECT 65.435000 27.290000 65.755000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 27.720000 65.755000 28.040000 ;
      LAYER met4 ;
        RECT 65.435000 27.720000 65.755000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 28.150000 65.755000 28.470000 ;
      LAYER met4 ;
        RECT 65.435000 28.150000 65.755000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 173.840000 66.090000 174.160000 ;
      LAYER met4 ;
        RECT 65.770000 173.840000 66.090000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 174.240000 66.090000 174.560000 ;
      LAYER met4 ;
        RECT 65.770000 174.240000 66.090000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 174.640000 66.090000 174.960000 ;
      LAYER met4 ;
        RECT 65.770000 174.640000 66.090000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 175.040000 66.090000 175.360000 ;
      LAYER met4 ;
        RECT 65.770000 175.040000 66.090000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 175.440000 66.090000 175.760000 ;
      LAYER met4 ;
        RECT 65.770000 175.440000 66.090000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 175.840000 66.090000 176.160000 ;
      LAYER met4 ;
        RECT 65.770000 175.840000 66.090000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 176.240000 66.090000 176.560000 ;
      LAYER met4 ;
        RECT 65.770000 176.240000 66.090000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 176.640000 66.090000 176.960000 ;
      LAYER met4 ;
        RECT 65.770000 176.640000 66.090000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 177.040000 66.090000 177.360000 ;
      LAYER met4 ;
        RECT 65.770000 177.040000 66.090000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 177.440000 66.090000 177.760000 ;
      LAYER met4 ;
        RECT 65.770000 177.440000 66.090000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 177.840000 66.090000 178.160000 ;
      LAYER met4 ;
        RECT 65.770000 177.840000 66.090000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 178.240000 66.090000 178.560000 ;
      LAYER met4 ;
        RECT 65.770000 178.240000 66.090000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 178.640000 66.090000 178.960000 ;
      LAYER met4 ;
        RECT 65.770000 178.640000 66.090000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 179.040000 66.090000 179.360000 ;
      LAYER met4 ;
        RECT 65.770000 179.040000 66.090000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 179.440000 66.090000 179.760000 ;
      LAYER met4 ;
        RECT 65.770000 179.440000 66.090000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 179.840000 66.090000 180.160000 ;
      LAYER met4 ;
        RECT 65.770000 179.840000 66.090000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 180.240000 66.090000 180.560000 ;
      LAYER met4 ;
        RECT 65.770000 180.240000 66.090000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 180.640000 66.090000 180.960000 ;
      LAYER met4 ;
        RECT 65.770000 180.640000 66.090000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 181.040000 66.090000 181.360000 ;
      LAYER met4 ;
        RECT 65.770000 181.040000 66.090000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 181.445000 66.090000 181.765000 ;
      LAYER met4 ;
        RECT 65.770000 181.445000 66.090000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 181.850000 66.090000 182.170000 ;
      LAYER met4 ;
        RECT 65.770000 181.850000 66.090000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 182.255000 66.090000 182.575000 ;
      LAYER met4 ;
        RECT 65.770000 182.255000 66.090000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 182.660000 66.090000 182.980000 ;
      LAYER met4 ;
        RECT 65.770000 182.660000 66.090000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 183.065000 66.090000 183.385000 ;
      LAYER met4 ;
        RECT 65.770000 183.065000 66.090000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 183.470000 66.090000 183.790000 ;
      LAYER met4 ;
        RECT 65.770000 183.470000 66.090000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 183.875000 66.090000 184.195000 ;
      LAYER met4 ;
        RECT 65.770000 183.875000 66.090000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 184.280000 66.090000 184.600000 ;
      LAYER met4 ;
        RECT 65.770000 184.280000 66.090000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 184.685000 66.090000 185.005000 ;
      LAYER met4 ;
        RECT 65.770000 184.685000 66.090000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 185.090000 66.090000 185.410000 ;
      LAYER met4 ;
        RECT 65.770000 185.090000 66.090000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 185.495000 66.090000 185.815000 ;
      LAYER met4 ;
        RECT 65.770000 185.495000 66.090000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 185.900000 66.090000 186.220000 ;
      LAYER met4 ;
        RECT 65.770000 185.900000 66.090000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 186.305000 66.090000 186.625000 ;
      LAYER met4 ;
        RECT 65.770000 186.305000 66.090000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 186.710000 66.090000 187.030000 ;
      LAYER met4 ;
        RECT 65.770000 186.710000 66.090000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 187.115000 66.090000 187.435000 ;
      LAYER met4 ;
        RECT 65.770000 187.115000 66.090000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 187.520000 66.090000 187.840000 ;
      LAYER met4 ;
        RECT 65.770000 187.520000 66.090000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 187.925000 66.090000 188.245000 ;
      LAYER met4 ;
        RECT 65.770000 187.925000 66.090000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 188.330000 66.090000 188.650000 ;
      LAYER met4 ;
        RECT 65.770000 188.330000 66.090000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 188.735000 66.090000 189.055000 ;
      LAYER met4 ;
        RECT 65.770000 188.735000 66.090000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 189.140000 66.090000 189.460000 ;
      LAYER met4 ;
        RECT 65.770000 189.140000 66.090000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 189.545000 66.090000 189.865000 ;
      LAYER met4 ;
        RECT 65.770000 189.545000 66.090000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 189.950000 66.090000 190.270000 ;
      LAYER met4 ;
        RECT 65.770000 189.950000 66.090000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 190.355000 66.090000 190.675000 ;
      LAYER met4 ;
        RECT 65.770000 190.355000 66.090000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 190.760000 66.090000 191.080000 ;
      LAYER met4 ;
        RECT 65.770000 190.760000 66.090000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 191.165000 66.090000 191.485000 ;
      LAYER met4 ;
        RECT 65.770000 191.165000 66.090000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 191.570000 66.090000 191.890000 ;
      LAYER met4 ;
        RECT 65.770000 191.570000 66.090000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 191.975000 66.090000 192.295000 ;
      LAYER met4 ;
        RECT 65.770000 191.975000 66.090000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 192.380000 66.090000 192.700000 ;
      LAYER met4 ;
        RECT 65.770000 192.380000 66.090000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 192.785000 66.090000 193.105000 ;
      LAYER met4 ;
        RECT 65.770000 192.785000 66.090000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 193.190000 66.090000 193.510000 ;
      LAYER met4 ;
        RECT 65.770000 193.190000 66.090000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 193.595000 66.090000 193.915000 ;
      LAYER met4 ;
        RECT 65.770000 193.595000 66.090000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 194.000000 66.090000 194.320000 ;
      LAYER met4 ;
        RECT 65.770000 194.000000 66.090000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 194.405000 66.090000 194.725000 ;
      LAYER met4 ;
        RECT 65.770000 194.405000 66.090000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 194.810000 66.090000 195.130000 ;
      LAYER met4 ;
        RECT 65.770000 194.810000 66.090000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 195.215000 66.090000 195.535000 ;
      LAYER met4 ;
        RECT 65.770000 195.215000 66.090000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 195.620000 66.090000 195.940000 ;
      LAYER met4 ;
        RECT 65.770000 195.620000 66.090000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 196.025000 66.090000 196.345000 ;
      LAYER met4 ;
        RECT 65.770000 196.025000 66.090000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 196.430000 66.090000 196.750000 ;
      LAYER met4 ;
        RECT 65.770000 196.430000 66.090000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 196.835000 66.090000 197.155000 ;
      LAYER met4 ;
        RECT 65.770000 196.835000 66.090000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 197.240000 66.090000 197.560000 ;
      LAYER met4 ;
        RECT 65.770000 197.240000 66.090000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 197.645000 66.090000 197.965000 ;
      LAYER met4 ;
        RECT 65.770000 197.645000 66.090000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 23.850000 66.160000 24.170000 ;
      LAYER met4 ;
        RECT 65.840000 23.850000 66.160000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 24.280000 66.160000 24.600000 ;
      LAYER met4 ;
        RECT 65.840000 24.280000 66.160000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 24.710000 66.160000 25.030000 ;
      LAYER met4 ;
        RECT 65.840000 24.710000 66.160000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 25.140000 66.160000 25.460000 ;
      LAYER met4 ;
        RECT 65.840000 25.140000 66.160000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 25.570000 66.160000 25.890000 ;
      LAYER met4 ;
        RECT 65.840000 25.570000 66.160000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 26.000000 66.160000 26.320000 ;
      LAYER met4 ;
        RECT 65.840000 26.000000 66.160000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 26.430000 66.160000 26.750000 ;
      LAYER met4 ;
        RECT 65.840000 26.430000 66.160000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 26.860000 66.160000 27.180000 ;
      LAYER met4 ;
        RECT 65.840000 26.860000 66.160000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 27.290000 66.160000 27.610000 ;
      LAYER met4 ;
        RECT 65.840000 27.290000 66.160000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 27.720000 66.160000 28.040000 ;
      LAYER met4 ;
        RECT 65.840000 27.720000 66.160000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 28.150000 66.160000 28.470000 ;
      LAYER met4 ;
        RECT 65.840000 28.150000 66.160000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 173.840000 66.500000 174.160000 ;
      LAYER met4 ;
        RECT 66.180000 173.840000 66.500000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 174.240000 66.500000 174.560000 ;
      LAYER met4 ;
        RECT 66.180000 174.240000 66.500000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 174.640000 66.500000 174.960000 ;
      LAYER met4 ;
        RECT 66.180000 174.640000 66.500000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 175.040000 66.500000 175.360000 ;
      LAYER met4 ;
        RECT 66.180000 175.040000 66.500000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 175.440000 66.500000 175.760000 ;
      LAYER met4 ;
        RECT 66.180000 175.440000 66.500000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 175.840000 66.500000 176.160000 ;
      LAYER met4 ;
        RECT 66.180000 175.840000 66.500000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 176.240000 66.500000 176.560000 ;
      LAYER met4 ;
        RECT 66.180000 176.240000 66.500000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 176.640000 66.500000 176.960000 ;
      LAYER met4 ;
        RECT 66.180000 176.640000 66.500000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 177.040000 66.500000 177.360000 ;
      LAYER met4 ;
        RECT 66.180000 177.040000 66.500000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 177.440000 66.500000 177.760000 ;
      LAYER met4 ;
        RECT 66.180000 177.440000 66.500000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 177.840000 66.500000 178.160000 ;
      LAYER met4 ;
        RECT 66.180000 177.840000 66.500000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 178.240000 66.500000 178.560000 ;
      LAYER met4 ;
        RECT 66.180000 178.240000 66.500000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 178.640000 66.500000 178.960000 ;
      LAYER met4 ;
        RECT 66.180000 178.640000 66.500000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 179.040000 66.500000 179.360000 ;
      LAYER met4 ;
        RECT 66.180000 179.040000 66.500000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 179.440000 66.500000 179.760000 ;
      LAYER met4 ;
        RECT 66.180000 179.440000 66.500000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 179.840000 66.500000 180.160000 ;
      LAYER met4 ;
        RECT 66.180000 179.840000 66.500000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 180.240000 66.500000 180.560000 ;
      LAYER met4 ;
        RECT 66.180000 180.240000 66.500000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 180.640000 66.500000 180.960000 ;
      LAYER met4 ;
        RECT 66.180000 180.640000 66.500000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 181.040000 66.500000 181.360000 ;
      LAYER met4 ;
        RECT 66.180000 181.040000 66.500000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 181.445000 66.500000 181.765000 ;
      LAYER met4 ;
        RECT 66.180000 181.445000 66.500000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 181.850000 66.500000 182.170000 ;
      LAYER met4 ;
        RECT 66.180000 181.850000 66.500000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 182.255000 66.500000 182.575000 ;
      LAYER met4 ;
        RECT 66.180000 182.255000 66.500000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 182.660000 66.500000 182.980000 ;
      LAYER met4 ;
        RECT 66.180000 182.660000 66.500000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 183.065000 66.500000 183.385000 ;
      LAYER met4 ;
        RECT 66.180000 183.065000 66.500000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 183.470000 66.500000 183.790000 ;
      LAYER met4 ;
        RECT 66.180000 183.470000 66.500000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 183.875000 66.500000 184.195000 ;
      LAYER met4 ;
        RECT 66.180000 183.875000 66.500000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 184.280000 66.500000 184.600000 ;
      LAYER met4 ;
        RECT 66.180000 184.280000 66.500000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 184.685000 66.500000 185.005000 ;
      LAYER met4 ;
        RECT 66.180000 184.685000 66.500000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 185.090000 66.500000 185.410000 ;
      LAYER met4 ;
        RECT 66.180000 185.090000 66.500000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 185.495000 66.500000 185.815000 ;
      LAYER met4 ;
        RECT 66.180000 185.495000 66.500000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 185.900000 66.500000 186.220000 ;
      LAYER met4 ;
        RECT 66.180000 185.900000 66.500000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 186.305000 66.500000 186.625000 ;
      LAYER met4 ;
        RECT 66.180000 186.305000 66.500000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 186.710000 66.500000 187.030000 ;
      LAYER met4 ;
        RECT 66.180000 186.710000 66.500000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 187.115000 66.500000 187.435000 ;
      LAYER met4 ;
        RECT 66.180000 187.115000 66.500000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 187.520000 66.500000 187.840000 ;
      LAYER met4 ;
        RECT 66.180000 187.520000 66.500000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 187.925000 66.500000 188.245000 ;
      LAYER met4 ;
        RECT 66.180000 187.925000 66.500000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 188.330000 66.500000 188.650000 ;
      LAYER met4 ;
        RECT 66.180000 188.330000 66.500000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 188.735000 66.500000 189.055000 ;
      LAYER met4 ;
        RECT 66.180000 188.735000 66.500000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 189.140000 66.500000 189.460000 ;
      LAYER met4 ;
        RECT 66.180000 189.140000 66.500000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 189.545000 66.500000 189.865000 ;
      LAYER met4 ;
        RECT 66.180000 189.545000 66.500000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 189.950000 66.500000 190.270000 ;
      LAYER met4 ;
        RECT 66.180000 189.950000 66.500000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 190.355000 66.500000 190.675000 ;
      LAYER met4 ;
        RECT 66.180000 190.355000 66.500000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 190.760000 66.500000 191.080000 ;
      LAYER met4 ;
        RECT 66.180000 190.760000 66.500000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 191.165000 66.500000 191.485000 ;
      LAYER met4 ;
        RECT 66.180000 191.165000 66.500000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 191.570000 66.500000 191.890000 ;
      LAYER met4 ;
        RECT 66.180000 191.570000 66.500000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 191.975000 66.500000 192.295000 ;
      LAYER met4 ;
        RECT 66.180000 191.975000 66.500000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 192.380000 66.500000 192.700000 ;
      LAYER met4 ;
        RECT 66.180000 192.380000 66.500000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 192.785000 66.500000 193.105000 ;
      LAYER met4 ;
        RECT 66.180000 192.785000 66.500000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 193.190000 66.500000 193.510000 ;
      LAYER met4 ;
        RECT 66.180000 193.190000 66.500000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 193.595000 66.500000 193.915000 ;
      LAYER met4 ;
        RECT 66.180000 193.595000 66.500000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 194.000000 66.500000 194.320000 ;
      LAYER met4 ;
        RECT 66.180000 194.000000 66.500000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 194.405000 66.500000 194.725000 ;
      LAYER met4 ;
        RECT 66.180000 194.405000 66.500000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 194.810000 66.500000 195.130000 ;
      LAYER met4 ;
        RECT 66.180000 194.810000 66.500000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 195.215000 66.500000 195.535000 ;
      LAYER met4 ;
        RECT 66.180000 195.215000 66.500000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 195.620000 66.500000 195.940000 ;
      LAYER met4 ;
        RECT 66.180000 195.620000 66.500000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 196.025000 66.500000 196.345000 ;
      LAYER met4 ;
        RECT 66.180000 196.025000 66.500000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 196.430000 66.500000 196.750000 ;
      LAYER met4 ;
        RECT 66.180000 196.430000 66.500000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 196.835000 66.500000 197.155000 ;
      LAYER met4 ;
        RECT 66.180000 196.835000 66.500000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 197.240000 66.500000 197.560000 ;
      LAYER met4 ;
        RECT 66.180000 197.240000 66.500000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 197.645000 66.500000 197.965000 ;
      LAYER met4 ;
        RECT 66.180000 197.645000 66.500000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 23.850000 66.565000 24.170000 ;
      LAYER met4 ;
        RECT 66.245000 23.850000 66.565000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 24.280000 66.565000 24.600000 ;
      LAYER met4 ;
        RECT 66.245000 24.280000 66.565000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 24.710000 66.565000 25.030000 ;
      LAYER met4 ;
        RECT 66.245000 24.710000 66.565000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 25.140000 66.565000 25.460000 ;
      LAYER met4 ;
        RECT 66.245000 25.140000 66.565000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 25.570000 66.565000 25.890000 ;
      LAYER met4 ;
        RECT 66.245000 25.570000 66.565000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 26.000000 66.565000 26.320000 ;
      LAYER met4 ;
        RECT 66.245000 26.000000 66.565000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 26.430000 66.565000 26.750000 ;
      LAYER met4 ;
        RECT 66.245000 26.430000 66.565000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 26.860000 66.565000 27.180000 ;
      LAYER met4 ;
        RECT 66.245000 26.860000 66.565000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 27.290000 66.565000 27.610000 ;
      LAYER met4 ;
        RECT 66.245000 27.290000 66.565000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 27.720000 66.565000 28.040000 ;
      LAYER met4 ;
        RECT 66.245000 27.720000 66.565000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 28.150000 66.565000 28.470000 ;
      LAYER met4 ;
        RECT 66.245000 28.150000 66.565000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 173.840000 66.910000 174.160000 ;
      LAYER met4 ;
        RECT 66.590000 173.840000 66.910000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 174.240000 66.910000 174.560000 ;
      LAYER met4 ;
        RECT 66.590000 174.240000 66.910000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 174.640000 66.910000 174.960000 ;
      LAYER met4 ;
        RECT 66.590000 174.640000 66.910000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 175.040000 66.910000 175.360000 ;
      LAYER met4 ;
        RECT 66.590000 175.040000 66.910000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 175.440000 66.910000 175.760000 ;
      LAYER met4 ;
        RECT 66.590000 175.440000 66.910000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 175.840000 66.910000 176.160000 ;
      LAYER met4 ;
        RECT 66.590000 175.840000 66.910000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 176.240000 66.910000 176.560000 ;
      LAYER met4 ;
        RECT 66.590000 176.240000 66.910000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 176.640000 66.910000 176.960000 ;
      LAYER met4 ;
        RECT 66.590000 176.640000 66.910000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 177.040000 66.910000 177.360000 ;
      LAYER met4 ;
        RECT 66.590000 177.040000 66.910000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 177.440000 66.910000 177.760000 ;
      LAYER met4 ;
        RECT 66.590000 177.440000 66.910000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 177.840000 66.910000 178.160000 ;
      LAYER met4 ;
        RECT 66.590000 177.840000 66.910000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 178.240000 66.910000 178.560000 ;
      LAYER met4 ;
        RECT 66.590000 178.240000 66.910000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 178.640000 66.910000 178.960000 ;
      LAYER met4 ;
        RECT 66.590000 178.640000 66.910000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 179.040000 66.910000 179.360000 ;
      LAYER met4 ;
        RECT 66.590000 179.040000 66.910000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 179.440000 66.910000 179.760000 ;
      LAYER met4 ;
        RECT 66.590000 179.440000 66.910000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 179.840000 66.910000 180.160000 ;
      LAYER met4 ;
        RECT 66.590000 179.840000 66.910000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 180.240000 66.910000 180.560000 ;
      LAYER met4 ;
        RECT 66.590000 180.240000 66.910000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 180.640000 66.910000 180.960000 ;
      LAYER met4 ;
        RECT 66.590000 180.640000 66.910000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 181.040000 66.910000 181.360000 ;
      LAYER met4 ;
        RECT 66.590000 181.040000 66.910000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 181.445000 66.910000 181.765000 ;
      LAYER met4 ;
        RECT 66.590000 181.445000 66.910000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 181.850000 66.910000 182.170000 ;
      LAYER met4 ;
        RECT 66.590000 181.850000 66.910000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 182.255000 66.910000 182.575000 ;
      LAYER met4 ;
        RECT 66.590000 182.255000 66.910000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 182.660000 66.910000 182.980000 ;
      LAYER met4 ;
        RECT 66.590000 182.660000 66.910000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 183.065000 66.910000 183.385000 ;
      LAYER met4 ;
        RECT 66.590000 183.065000 66.910000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 183.470000 66.910000 183.790000 ;
      LAYER met4 ;
        RECT 66.590000 183.470000 66.910000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 183.875000 66.910000 184.195000 ;
      LAYER met4 ;
        RECT 66.590000 183.875000 66.910000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 184.280000 66.910000 184.600000 ;
      LAYER met4 ;
        RECT 66.590000 184.280000 66.910000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 184.685000 66.910000 185.005000 ;
      LAYER met4 ;
        RECT 66.590000 184.685000 66.910000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 185.090000 66.910000 185.410000 ;
      LAYER met4 ;
        RECT 66.590000 185.090000 66.910000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 185.495000 66.910000 185.815000 ;
      LAYER met4 ;
        RECT 66.590000 185.495000 66.910000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 185.900000 66.910000 186.220000 ;
      LAYER met4 ;
        RECT 66.590000 185.900000 66.910000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 186.305000 66.910000 186.625000 ;
      LAYER met4 ;
        RECT 66.590000 186.305000 66.910000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 186.710000 66.910000 187.030000 ;
      LAYER met4 ;
        RECT 66.590000 186.710000 66.910000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 187.115000 66.910000 187.435000 ;
      LAYER met4 ;
        RECT 66.590000 187.115000 66.910000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 187.520000 66.910000 187.840000 ;
      LAYER met4 ;
        RECT 66.590000 187.520000 66.910000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 187.925000 66.910000 188.245000 ;
      LAYER met4 ;
        RECT 66.590000 187.925000 66.910000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 188.330000 66.910000 188.650000 ;
      LAYER met4 ;
        RECT 66.590000 188.330000 66.910000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 188.735000 66.910000 189.055000 ;
      LAYER met4 ;
        RECT 66.590000 188.735000 66.910000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 189.140000 66.910000 189.460000 ;
      LAYER met4 ;
        RECT 66.590000 189.140000 66.910000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 189.545000 66.910000 189.865000 ;
      LAYER met4 ;
        RECT 66.590000 189.545000 66.910000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 189.950000 66.910000 190.270000 ;
      LAYER met4 ;
        RECT 66.590000 189.950000 66.910000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 190.355000 66.910000 190.675000 ;
      LAYER met4 ;
        RECT 66.590000 190.355000 66.910000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 190.760000 66.910000 191.080000 ;
      LAYER met4 ;
        RECT 66.590000 190.760000 66.910000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 191.165000 66.910000 191.485000 ;
      LAYER met4 ;
        RECT 66.590000 191.165000 66.910000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 191.570000 66.910000 191.890000 ;
      LAYER met4 ;
        RECT 66.590000 191.570000 66.910000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 191.975000 66.910000 192.295000 ;
      LAYER met4 ;
        RECT 66.590000 191.975000 66.910000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 192.380000 66.910000 192.700000 ;
      LAYER met4 ;
        RECT 66.590000 192.380000 66.910000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 192.785000 66.910000 193.105000 ;
      LAYER met4 ;
        RECT 66.590000 192.785000 66.910000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 193.190000 66.910000 193.510000 ;
      LAYER met4 ;
        RECT 66.590000 193.190000 66.910000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 193.595000 66.910000 193.915000 ;
      LAYER met4 ;
        RECT 66.590000 193.595000 66.910000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 194.000000 66.910000 194.320000 ;
      LAYER met4 ;
        RECT 66.590000 194.000000 66.910000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 194.405000 66.910000 194.725000 ;
      LAYER met4 ;
        RECT 66.590000 194.405000 66.910000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 194.810000 66.910000 195.130000 ;
      LAYER met4 ;
        RECT 66.590000 194.810000 66.910000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 195.215000 66.910000 195.535000 ;
      LAYER met4 ;
        RECT 66.590000 195.215000 66.910000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 195.620000 66.910000 195.940000 ;
      LAYER met4 ;
        RECT 66.590000 195.620000 66.910000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 196.025000 66.910000 196.345000 ;
      LAYER met4 ;
        RECT 66.590000 196.025000 66.910000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 196.430000 66.910000 196.750000 ;
      LAYER met4 ;
        RECT 66.590000 196.430000 66.910000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 196.835000 66.910000 197.155000 ;
      LAYER met4 ;
        RECT 66.590000 196.835000 66.910000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 197.240000 66.910000 197.560000 ;
      LAYER met4 ;
        RECT 66.590000 197.240000 66.910000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.590000 197.645000 66.910000 197.965000 ;
      LAYER met4 ;
        RECT 66.590000 197.645000 66.910000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 23.850000 66.970000 24.170000 ;
      LAYER met4 ;
        RECT 66.650000 23.850000 66.970000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 24.280000 66.970000 24.600000 ;
      LAYER met4 ;
        RECT 66.650000 24.280000 66.970000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 24.710000 66.970000 25.030000 ;
      LAYER met4 ;
        RECT 66.650000 24.710000 66.970000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 25.140000 66.970000 25.460000 ;
      LAYER met4 ;
        RECT 66.650000 25.140000 66.970000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 25.570000 66.970000 25.890000 ;
      LAYER met4 ;
        RECT 66.650000 25.570000 66.970000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 26.000000 66.970000 26.320000 ;
      LAYER met4 ;
        RECT 66.650000 26.000000 66.970000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 26.430000 66.970000 26.750000 ;
      LAYER met4 ;
        RECT 66.650000 26.430000 66.970000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 26.860000 66.970000 27.180000 ;
      LAYER met4 ;
        RECT 66.650000 26.860000 66.970000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 27.290000 66.970000 27.610000 ;
      LAYER met4 ;
        RECT 66.650000 27.290000 66.970000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 27.720000 66.970000 28.040000 ;
      LAYER met4 ;
        RECT 66.650000 27.720000 66.970000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 28.150000 66.970000 28.470000 ;
      LAYER met4 ;
        RECT 66.650000 28.150000 66.970000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 173.840000 67.320000 174.160000 ;
      LAYER met4 ;
        RECT 67.000000 173.840000 67.320000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 174.240000 67.320000 174.560000 ;
      LAYER met4 ;
        RECT 67.000000 174.240000 67.320000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 174.640000 67.320000 174.960000 ;
      LAYER met4 ;
        RECT 67.000000 174.640000 67.320000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 175.040000 67.320000 175.360000 ;
      LAYER met4 ;
        RECT 67.000000 175.040000 67.320000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 175.440000 67.320000 175.760000 ;
      LAYER met4 ;
        RECT 67.000000 175.440000 67.320000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 175.840000 67.320000 176.160000 ;
      LAYER met4 ;
        RECT 67.000000 175.840000 67.320000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 176.240000 67.320000 176.560000 ;
      LAYER met4 ;
        RECT 67.000000 176.240000 67.320000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 176.640000 67.320000 176.960000 ;
      LAYER met4 ;
        RECT 67.000000 176.640000 67.320000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 177.040000 67.320000 177.360000 ;
      LAYER met4 ;
        RECT 67.000000 177.040000 67.320000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 177.440000 67.320000 177.760000 ;
      LAYER met4 ;
        RECT 67.000000 177.440000 67.320000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 177.840000 67.320000 178.160000 ;
      LAYER met4 ;
        RECT 67.000000 177.840000 67.320000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 178.240000 67.320000 178.560000 ;
      LAYER met4 ;
        RECT 67.000000 178.240000 67.320000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 178.640000 67.320000 178.960000 ;
      LAYER met4 ;
        RECT 67.000000 178.640000 67.320000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 179.040000 67.320000 179.360000 ;
      LAYER met4 ;
        RECT 67.000000 179.040000 67.320000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 179.440000 67.320000 179.760000 ;
      LAYER met4 ;
        RECT 67.000000 179.440000 67.320000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 179.840000 67.320000 180.160000 ;
      LAYER met4 ;
        RECT 67.000000 179.840000 67.320000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 180.240000 67.320000 180.560000 ;
      LAYER met4 ;
        RECT 67.000000 180.240000 67.320000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 180.640000 67.320000 180.960000 ;
      LAYER met4 ;
        RECT 67.000000 180.640000 67.320000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 181.040000 67.320000 181.360000 ;
      LAYER met4 ;
        RECT 67.000000 181.040000 67.320000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 181.445000 67.320000 181.765000 ;
      LAYER met4 ;
        RECT 67.000000 181.445000 67.320000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 181.850000 67.320000 182.170000 ;
      LAYER met4 ;
        RECT 67.000000 181.850000 67.320000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 182.255000 67.320000 182.575000 ;
      LAYER met4 ;
        RECT 67.000000 182.255000 67.320000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 182.660000 67.320000 182.980000 ;
      LAYER met4 ;
        RECT 67.000000 182.660000 67.320000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 183.065000 67.320000 183.385000 ;
      LAYER met4 ;
        RECT 67.000000 183.065000 67.320000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 183.470000 67.320000 183.790000 ;
      LAYER met4 ;
        RECT 67.000000 183.470000 67.320000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 183.875000 67.320000 184.195000 ;
      LAYER met4 ;
        RECT 67.000000 183.875000 67.320000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 184.280000 67.320000 184.600000 ;
      LAYER met4 ;
        RECT 67.000000 184.280000 67.320000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 184.685000 67.320000 185.005000 ;
      LAYER met4 ;
        RECT 67.000000 184.685000 67.320000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 185.090000 67.320000 185.410000 ;
      LAYER met4 ;
        RECT 67.000000 185.090000 67.320000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 185.495000 67.320000 185.815000 ;
      LAYER met4 ;
        RECT 67.000000 185.495000 67.320000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 185.900000 67.320000 186.220000 ;
      LAYER met4 ;
        RECT 67.000000 185.900000 67.320000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 186.305000 67.320000 186.625000 ;
      LAYER met4 ;
        RECT 67.000000 186.305000 67.320000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 186.710000 67.320000 187.030000 ;
      LAYER met4 ;
        RECT 67.000000 186.710000 67.320000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 187.115000 67.320000 187.435000 ;
      LAYER met4 ;
        RECT 67.000000 187.115000 67.320000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 187.520000 67.320000 187.840000 ;
      LAYER met4 ;
        RECT 67.000000 187.520000 67.320000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 187.925000 67.320000 188.245000 ;
      LAYER met4 ;
        RECT 67.000000 187.925000 67.320000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 188.330000 67.320000 188.650000 ;
      LAYER met4 ;
        RECT 67.000000 188.330000 67.320000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 188.735000 67.320000 189.055000 ;
      LAYER met4 ;
        RECT 67.000000 188.735000 67.320000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 189.140000 67.320000 189.460000 ;
      LAYER met4 ;
        RECT 67.000000 189.140000 67.320000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 189.545000 67.320000 189.865000 ;
      LAYER met4 ;
        RECT 67.000000 189.545000 67.320000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 189.950000 67.320000 190.270000 ;
      LAYER met4 ;
        RECT 67.000000 189.950000 67.320000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 190.355000 67.320000 190.675000 ;
      LAYER met4 ;
        RECT 67.000000 190.355000 67.320000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 190.760000 67.320000 191.080000 ;
      LAYER met4 ;
        RECT 67.000000 190.760000 67.320000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 191.165000 67.320000 191.485000 ;
      LAYER met4 ;
        RECT 67.000000 191.165000 67.320000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 191.570000 67.320000 191.890000 ;
      LAYER met4 ;
        RECT 67.000000 191.570000 67.320000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 191.975000 67.320000 192.295000 ;
      LAYER met4 ;
        RECT 67.000000 191.975000 67.320000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 192.380000 67.320000 192.700000 ;
      LAYER met4 ;
        RECT 67.000000 192.380000 67.320000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 192.785000 67.320000 193.105000 ;
      LAYER met4 ;
        RECT 67.000000 192.785000 67.320000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 193.190000 67.320000 193.510000 ;
      LAYER met4 ;
        RECT 67.000000 193.190000 67.320000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 193.595000 67.320000 193.915000 ;
      LAYER met4 ;
        RECT 67.000000 193.595000 67.320000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 194.000000 67.320000 194.320000 ;
      LAYER met4 ;
        RECT 67.000000 194.000000 67.320000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 194.405000 67.320000 194.725000 ;
      LAYER met4 ;
        RECT 67.000000 194.405000 67.320000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 194.810000 67.320000 195.130000 ;
      LAYER met4 ;
        RECT 67.000000 194.810000 67.320000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 195.215000 67.320000 195.535000 ;
      LAYER met4 ;
        RECT 67.000000 195.215000 67.320000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 195.620000 67.320000 195.940000 ;
      LAYER met4 ;
        RECT 67.000000 195.620000 67.320000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 196.025000 67.320000 196.345000 ;
      LAYER met4 ;
        RECT 67.000000 196.025000 67.320000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 196.430000 67.320000 196.750000 ;
      LAYER met4 ;
        RECT 67.000000 196.430000 67.320000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 196.835000 67.320000 197.155000 ;
      LAYER met4 ;
        RECT 67.000000 196.835000 67.320000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 197.240000 67.320000 197.560000 ;
      LAYER met4 ;
        RECT 67.000000 197.240000 67.320000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.000000 197.645000 67.320000 197.965000 ;
      LAYER met4 ;
        RECT 67.000000 197.645000 67.320000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 23.850000 67.375000 24.170000 ;
      LAYER met4 ;
        RECT 67.055000 23.850000 67.375000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 24.280000 67.375000 24.600000 ;
      LAYER met4 ;
        RECT 67.055000 24.280000 67.375000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 24.710000 67.375000 25.030000 ;
      LAYER met4 ;
        RECT 67.055000 24.710000 67.375000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 25.140000 67.375000 25.460000 ;
      LAYER met4 ;
        RECT 67.055000 25.140000 67.375000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 25.570000 67.375000 25.890000 ;
      LAYER met4 ;
        RECT 67.055000 25.570000 67.375000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 26.000000 67.375000 26.320000 ;
      LAYER met4 ;
        RECT 67.055000 26.000000 67.375000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 26.430000 67.375000 26.750000 ;
      LAYER met4 ;
        RECT 67.055000 26.430000 67.375000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 26.860000 67.375000 27.180000 ;
      LAYER met4 ;
        RECT 67.055000 26.860000 67.375000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 27.290000 67.375000 27.610000 ;
      LAYER met4 ;
        RECT 67.055000 27.290000 67.375000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 27.720000 67.375000 28.040000 ;
      LAYER met4 ;
        RECT 67.055000 27.720000 67.375000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 28.150000 67.375000 28.470000 ;
      LAYER met4 ;
        RECT 67.055000 28.150000 67.375000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 173.840000 67.730000 174.160000 ;
      LAYER met4 ;
        RECT 67.410000 173.840000 67.730000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 174.240000 67.730000 174.560000 ;
      LAYER met4 ;
        RECT 67.410000 174.240000 67.730000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 174.640000 67.730000 174.960000 ;
      LAYER met4 ;
        RECT 67.410000 174.640000 67.730000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 175.040000 67.730000 175.360000 ;
      LAYER met4 ;
        RECT 67.410000 175.040000 67.730000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 175.440000 67.730000 175.760000 ;
      LAYER met4 ;
        RECT 67.410000 175.440000 67.730000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 175.840000 67.730000 176.160000 ;
      LAYER met4 ;
        RECT 67.410000 175.840000 67.730000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 176.240000 67.730000 176.560000 ;
      LAYER met4 ;
        RECT 67.410000 176.240000 67.730000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 176.640000 67.730000 176.960000 ;
      LAYER met4 ;
        RECT 67.410000 176.640000 67.730000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 177.040000 67.730000 177.360000 ;
      LAYER met4 ;
        RECT 67.410000 177.040000 67.730000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 177.440000 67.730000 177.760000 ;
      LAYER met4 ;
        RECT 67.410000 177.440000 67.730000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 177.840000 67.730000 178.160000 ;
      LAYER met4 ;
        RECT 67.410000 177.840000 67.730000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 178.240000 67.730000 178.560000 ;
      LAYER met4 ;
        RECT 67.410000 178.240000 67.730000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 178.640000 67.730000 178.960000 ;
      LAYER met4 ;
        RECT 67.410000 178.640000 67.730000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 179.040000 67.730000 179.360000 ;
      LAYER met4 ;
        RECT 67.410000 179.040000 67.730000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 179.440000 67.730000 179.760000 ;
      LAYER met4 ;
        RECT 67.410000 179.440000 67.730000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 179.840000 67.730000 180.160000 ;
      LAYER met4 ;
        RECT 67.410000 179.840000 67.730000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 180.240000 67.730000 180.560000 ;
      LAYER met4 ;
        RECT 67.410000 180.240000 67.730000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 180.640000 67.730000 180.960000 ;
      LAYER met4 ;
        RECT 67.410000 180.640000 67.730000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 181.040000 67.730000 181.360000 ;
      LAYER met4 ;
        RECT 67.410000 181.040000 67.730000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 181.445000 67.730000 181.765000 ;
      LAYER met4 ;
        RECT 67.410000 181.445000 67.730000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 181.850000 67.730000 182.170000 ;
      LAYER met4 ;
        RECT 67.410000 181.850000 67.730000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 182.255000 67.730000 182.575000 ;
      LAYER met4 ;
        RECT 67.410000 182.255000 67.730000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 182.660000 67.730000 182.980000 ;
      LAYER met4 ;
        RECT 67.410000 182.660000 67.730000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 183.065000 67.730000 183.385000 ;
      LAYER met4 ;
        RECT 67.410000 183.065000 67.730000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 183.470000 67.730000 183.790000 ;
      LAYER met4 ;
        RECT 67.410000 183.470000 67.730000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 183.875000 67.730000 184.195000 ;
      LAYER met4 ;
        RECT 67.410000 183.875000 67.730000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 184.280000 67.730000 184.600000 ;
      LAYER met4 ;
        RECT 67.410000 184.280000 67.730000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 184.685000 67.730000 185.005000 ;
      LAYER met4 ;
        RECT 67.410000 184.685000 67.730000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 185.090000 67.730000 185.410000 ;
      LAYER met4 ;
        RECT 67.410000 185.090000 67.730000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 185.495000 67.730000 185.815000 ;
      LAYER met4 ;
        RECT 67.410000 185.495000 67.730000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 185.900000 67.730000 186.220000 ;
      LAYER met4 ;
        RECT 67.410000 185.900000 67.730000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 186.305000 67.730000 186.625000 ;
      LAYER met4 ;
        RECT 67.410000 186.305000 67.730000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 186.710000 67.730000 187.030000 ;
      LAYER met4 ;
        RECT 67.410000 186.710000 67.730000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 187.115000 67.730000 187.435000 ;
      LAYER met4 ;
        RECT 67.410000 187.115000 67.730000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 187.520000 67.730000 187.840000 ;
      LAYER met4 ;
        RECT 67.410000 187.520000 67.730000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 187.925000 67.730000 188.245000 ;
      LAYER met4 ;
        RECT 67.410000 187.925000 67.730000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 188.330000 67.730000 188.650000 ;
      LAYER met4 ;
        RECT 67.410000 188.330000 67.730000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 188.735000 67.730000 189.055000 ;
      LAYER met4 ;
        RECT 67.410000 188.735000 67.730000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 189.140000 67.730000 189.460000 ;
      LAYER met4 ;
        RECT 67.410000 189.140000 67.730000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 189.545000 67.730000 189.865000 ;
      LAYER met4 ;
        RECT 67.410000 189.545000 67.730000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 189.950000 67.730000 190.270000 ;
      LAYER met4 ;
        RECT 67.410000 189.950000 67.730000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 190.355000 67.730000 190.675000 ;
      LAYER met4 ;
        RECT 67.410000 190.355000 67.730000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 190.760000 67.730000 191.080000 ;
      LAYER met4 ;
        RECT 67.410000 190.760000 67.730000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 191.165000 67.730000 191.485000 ;
      LAYER met4 ;
        RECT 67.410000 191.165000 67.730000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 191.570000 67.730000 191.890000 ;
      LAYER met4 ;
        RECT 67.410000 191.570000 67.730000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 191.975000 67.730000 192.295000 ;
      LAYER met4 ;
        RECT 67.410000 191.975000 67.730000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 192.380000 67.730000 192.700000 ;
      LAYER met4 ;
        RECT 67.410000 192.380000 67.730000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 192.785000 67.730000 193.105000 ;
      LAYER met4 ;
        RECT 67.410000 192.785000 67.730000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 193.190000 67.730000 193.510000 ;
      LAYER met4 ;
        RECT 67.410000 193.190000 67.730000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 193.595000 67.730000 193.915000 ;
      LAYER met4 ;
        RECT 67.410000 193.595000 67.730000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 194.000000 67.730000 194.320000 ;
      LAYER met4 ;
        RECT 67.410000 194.000000 67.730000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 194.405000 67.730000 194.725000 ;
      LAYER met4 ;
        RECT 67.410000 194.405000 67.730000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 194.810000 67.730000 195.130000 ;
      LAYER met4 ;
        RECT 67.410000 194.810000 67.730000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 195.215000 67.730000 195.535000 ;
      LAYER met4 ;
        RECT 67.410000 195.215000 67.730000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 195.620000 67.730000 195.940000 ;
      LAYER met4 ;
        RECT 67.410000 195.620000 67.730000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 196.025000 67.730000 196.345000 ;
      LAYER met4 ;
        RECT 67.410000 196.025000 67.730000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 196.430000 67.730000 196.750000 ;
      LAYER met4 ;
        RECT 67.410000 196.430000 67.730000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 196.835000 67.730000 197.155000 ;
      LAYER met4 ;
        RECT 67.410000 196.835000 67.730000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 197.240000 67.730000 197.560000 ;
      LAYER met4 ;
        RECT 67.410000 197.240000 67.730000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410000 197.645000 67.730000 197.965000 ;
      LAYER met4 ;
        RECT 67.410000 197.645000 67.730000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 23.850000 67.780000 24.170000 ;
      LAYER met4 ;
        RECT 67.460000 23.850000 67.780000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 24.280000 67.780000 24.600000 ;
      LAYER met4 ;
        RECT 67.460000 24.280000 67.780000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 24.710000 67.780000 25.030000 ;
      LAYER met4 ;
        RECT 67.460000 24.710000 67.780000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 25.140000 67.780000 25.460000 ;
      LAYER met4 ;
        RECT 67.460000 25.140000 67.780000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 25.570000 67.780000 25.890000 ;
      LAYER met4 ;
        RECT 67.460000 25.570000 67.780000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 26.000000 67.780000 26.320000 ;
      LAYER met4 ;
        RECT 67.460000 26.000000 67.780000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 26.430000 67.780000 26.750000 ;
      LAYER met4 ;
        RECT 67.460000 26.430000 67.780000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 26.860000 67.780000 27.180000 ;
      LAYER met4 ;
        RECT 67.460000 26.860000 67.780000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 27.290000 67.780000 27.610000 ;
      LAYER met4 ;
        RECT 67.460000 27.290000 67.780000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 27.720000 67.780000 28.040000 ;
      LAYER met4 ;
        RECT 67.460000 27.720000 67.780000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 28.150000 67.780000 28.470000 ;
      LAYER met4 ;
        RECT 67.460000 28.150000 67.780000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 173.840000 68.140000 174.160000 ;
      LAYER met4 ;
        RECT 67.820000 173.840000 68.140000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 174.240000 68.140000 174.560000 ;
      LAYER met4 ;
        RECT 67.820000 174.240000 68.140000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 174.640000 68.140000 174.960000 ;
      LAYER met4 ;
        RECT 67.820000 174.640000 68.140000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 175.040000 68.140000 175.360000 ;
      LAYER met4 ;
        RECT 67.820000 175.040000 68.140000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 175.440000 68.140000 175.760000 ;
      LAYER met4 ;
        RECT 67.820000 175.440000 68.140000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 175.840000 68.140000 176.160000 ;
      LAYER met4 ;
        RECT 67.820000 175.840000 68.140000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 176.240000 68.140000 176.560000 ;
      LAYER met4 ;
        RECT 67.820000 176.240000 68.140000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 176.640000 68.140000 176.960000 ;
      LAYER met4 ;
        RECT 67.820000 176.640000 68.140000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 177.040000 68.140000 177.360000 ;
      LAYER met4 ;
        RECT 67.820000 177.040000 68.140000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 177.440000 68.140000 177.760000 ;
      LAYER met4 ;
        RECT 67.820000 177.440000 68.140000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 177.840000 68.140000 178.160000 ;
      LAYER met4 ;
        RECT 67.820000 177.840000 68.140000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 178.240000 68.140000 178.560000 ;
      LAYER met4 ;
        RECT 67.820000 178.240000 68.140000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 178.640000 68.140000 178.960000 ;
      LAYER met4 ;
        RECT 67.820000 178.640000 68.140000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 179.040000 68.140000 179.360000 ;
      LAYER met4 ;
        RECT 67.820000 179.040000 68.140000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 179.440000 68.140000 179.760000 ;
      LAYER met4 ;
        RECT 67.820000 179.440000 68.140000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 179.840000 68.140000 180.160000 ;
      LAYER met4 ;
        RECT 67.820000 179.840000 68.140000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 180.240000 68.140000 180.560000 ;
      LAYER met4 ;
        RECT 67.820000 180.240000 68.140000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 180.640000 68.140000 180.960000 ;
      LAYER met4 ;
        RECT 67.820000 180.640000 68.140000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 181.040000 68.140000 181.360000 ;
      LAYER met4 ;
        RECT 67.820000 181.040000 68.140000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 181.445000 68.140000 181.765000 ;
      LAYER met4 ;
        RECT 67.820000 181.445000 68.140000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 181.850000 68.140000 182.170000 ;
      LAYER met4 ;
        RECT 67.820000 181.850000 68.140000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 182.255000 68.140000 182.575000 ;
      LAYER met4 ;
        RECT 67.820000 182.255000 68.140000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 182.660000 68.140000 182.980000 ;
      LAYER met4 ;
        RECT 67.820000 182.660000 68.140000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 183.065000 68.140000 183.385000 ;
      LAYER met4 ;
        RECT 67.820000 183.065000 68.140000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 183.470000 68.140000 183.790000 ;
      LAYER met4 ;
        RECT 67.820000 183.470000 68.140000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 183.875000 68.140000 184.195000 ;
      LAYER met4 ;
        RECT 67.820000 183.875000 68.140000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 184.280000 68.140000 184.600000 ;
      LAYER met4 ;
        RECT 67.820000 184.280000 68.140000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 184.685000 68.140000 185.005000 ;
      LAYER met4 ;
        RECT 67.820000 184.685000 68.140000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 185.090000 68.140000 185.410000 ;
      LAYER met4 ;
        RECT 67.820000 185.090000 68.140000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 185.495000 68.140000 185.815000 ;
      LAYER met4 ;
        RECT 67.820000 185.495000 68.140000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 185.900000 68.140000 186.220000 ;
      LAYER met4 ;
        RECT 67.820000 185.900000 68.140000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 186.305000 68.140000 186.625000 ;
      LAYER met4 ;
        RECT 67.820000 186.305000 68.140000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 186.710000 68.140000 187.030000 ;
      LAYER met4 ;
        RECT 67.820000 186.710000 68.140000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 187.115000 68.140000 187.435000 ;
      LAYER met4 ;
        RECT 67.820000 187.115000 68.140000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 187.520000 68.140000 187.840000 ;
      LAYER met4 ;
        RECT 67.820000 187.520000 68.140000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 187.925000 68.140000 188.245000 ;
      LAYER met4 ;
        RECT 67.820000 187.925000 68.140000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 188.330000 68.140000 188.650000 ;
      LAYER met4 ;
        RECT 67.820000 188.330000 68.140000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 188.735000 68.140000 189.055000 ;
      LAYER met4 ;
        RECT 67.820000 188.735000 68.140000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 189.140000 68.140000 189.460000 ;
      LAYER met4 ;
        RECT 67.820000 189.140000 68.140000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 189.545000 68.140000 189.865000 ;
      LAYER met4 ;
        RECT 67.820000 189.545000 68.140000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 189.950000 68.140000 190.270000 ;
      LAYER met4 ;
        RECT 67.820000 189.950000 68.140000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 190.355000 68.140000 190.675000 ;
      LAYER met4 ;
        RECT 67.820000 190.355000 68.140000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 190.760000 68.140000 191.080000 ;
      LAYER met4 ;
        RECT 67.820000 190.760000 68.140000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 191.165000 68.140000 191.485000 ;
      LAYER met4 ;
        RECT 67.820000 191.165000 68.140000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 191.570000 68.140000 191.890000 ;
      LAYER met4 ;
        RECT 67.820000 191.570000 68.140000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 191.975000 68.140000 192.295000 ;
      LAYER met4 ;
        RECT 67.820000 191.975000 68.140000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 192.380000 68.140000 192.700000 ;
      LAYER met4 ;
        RECT 67.820000 192.380000 68.140000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 192.785000 68.140000 193.105000 ;
      LAYER met4 ;
        RECT 67.820000 192.785000 68.140000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 193.190000 68.140000 193.510000 ;
      LAYER met4 ;
        RECT 67.820000 193.190000 68.140000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 193.595000 68.140000 193.915000 ;
      LAYER met4 ;
        RECT 67.820000 193.595000 68.140000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 194.000000 68.140000 194.320000 ;
      LAYER met4 ;
        RECT 67.820000 194.000000 68.140000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 194.405000 68.140000 194.725000 ;
      LAYER met4 ;
        RECT 67.820000 194.405000 68.140000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 194.810000 68.140000 195.130000 ;
      LAYER met4 ;
        RECT 67.820000 194.810000 68.140000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 195.215000 68.140000 195.535000 ;
      LAYER met4 ;
        RECT 67.820000 195.215000 68.140000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 195.620000 68.140000 195.940000 ;
      LAYER met4 ;
        RECT 67.820000 195.620000 68.140000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 196.025000 68.140000 196.345000 ;
      LAYER met4 ;
        RECT 67.820000 196.025000 68.140000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 196.430000 68.140000 196.750000 ;
      LAYER met4 ;
        RECT 67.820000 196.430000 68.140000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 196.835000 68.140000 197.155000 ;
      LAYER met4 ;
        RECT 67.820000 196.835000 68.140000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 197.240000 68.140000 197.560000 ;
      LAYER met4 ;
        RECT 67.820000 197.240000 68.140000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.820000 197.645000 68.140000 197.965000 ;
      LAYER met4 ;
        RECT 67.820000 197.645000 68.140000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 23.850000 68.185000 24.170000 ;
      LAYER met4 ;
        RECT 67.865000 23.850000 68.185000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 24.280000 68.185000 24.600000 ;
      LAYER met4 ;
        RECT 67.865000 24.280000 68.185000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 24.710000 68.185000 25.030000 ;
      LAYER met4 ;
        RECT 67.865000 24.710000 68.185000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 25.140000 68.185000 25.460000 ;
      LAYER met4 ;
        RECT 67.865000 25.140000 68.185000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 25.570000 68.185000 25.890000 ;
      LAYER met4 ;
        RECT 67.865000 25.570000 68.185000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 26.000000 68.185000 26.320000 ;
      LAYER met4 ;
        RECT 67.865000 26.000000 68.185000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 26.430000 68.185000 26.750000 ;
      LAYER met4 ;
        RECT 67.865000 26.430000 68.185000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 26.860000 68.185000 27.180000 ;
      LAYER met4 ;
        RECT 67.865000 26.860000 68.185000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 27.290000 68.185000 27.610000 ;
      LAYER met4 ;
        RECT 67.865000 27.290000 68.185000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 27.720000 68.185000 28.040000 ;
      LAYER met4 ;
        RECT 67.865000 27.720000 68.185000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 28.150000 68.185000 28.470000 ;
      LAYER met4 ;
        RECT 67.865000 28.150000 68.185000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 173.840000 68.550000 174.160000 ;
      LAYER met4 ;
        RECT 68.230000 173.840000 68.550000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 174.240000 68.550000 174.560000 ;
      LAYER met4 ;
        RECT 68.230000 174.240000 68.550000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 174.640000 68.550000 174.960000 ;
      LAYER met4 ;
        RECT 68.230000 174.640000 68.550000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 175.040000 68.550000 175.360000 ;
      LAYER met4 ;
        RECT 68.230000 175.040000 68.550000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 175.440000 68.550000 175.760000 ;
      LAYER met4 ;
        RECT 68.230000 175.440000 68.550000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 175.840000 68.550000 176.160000 ;
      LAYER met4 ;
        RECT 68.230000 175.840000 68.550000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 176.240000 68.550000 176.560000 ;
      LAYER met4 ;
        RECT 68.230000 176.240000 68.550000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 176.640000 68.550000 176.960000 ;
      LAYER met4 ;
        RECT 68.230000 176.640000 68.550000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 177.040000 68.550000 177.360000 ;
      LAYER met4 ;
        RECT 68.230000 177.040000 68.550000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 177.440000 68.550000 177.760000 ;
      LAYER met4 ;
        RECT 68.230000 177.440000 68.550000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 177.840000 68.550000 178.160000 ;
      LAYER met4 ;
        RECT 68.230000 177.840000 68.550000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 178.240000 68.550000 178.560000 ;
      LAYER met4 ;
        RECT 68.230000 178.240000 68.550000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 178.640000 68.550000 178.960000 ;
      LAYER met4 ;
        RECT 68.230000 178.640000 68.550000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 179.040000 68.550000 179.360000 ;
      LAYER met4 ;
        RECT 68.230000 179.040000 68.550000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 179.440000 68.550000 179.760000 ;
      LAYER met4 ;
        RECT 68.230000 179.440000 68.550000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 179.840000 68.550000 180.160000 ;
      LAYER met4 ;
        RECT 68.230000 179.840000 68.550000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 180.240000 68.550000 180.560000 ;
      LAYER met4 ;
        RECT 68.230000 180.240000 68.550000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 180.640000 68.550000 180.960000 ;
      LAYER met4 ;
        RECT 68.230000 180.640000 68.550000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 181.040000 68.550000 181.360000 ;
      LAYER met4 ;
        RECT 68.230000 181.040000 68.550000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 181.445000 68.550000 181.765000 ;
      LAYER met4 ;
        RECT 68.230000 181.445000 68.550000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 181.850000 68.550000 182.170000 ;
      LAYER met4 ;
        RECT 68.230000 181.850000 68.550000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 182.255000 68.550000 182.575000 ;
      LAYER met4 ;
        RECT 68.230000 182.255000 68.550000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 182.660000 68.550000 182.980000 ;
      LAYER met4 ;
        RECT 68.230000 182.660000 68.550000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 183.065000 68.550000 183.385000 ;
      LAYER met4 ;
        RECT 68.230000 183.065000 68.550000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 183.470000 68.550000 183.790000 ;
      LAYER met4 ;
        RECT 68.230000 183.470000 68.550000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 183.875000 68.550000 184.195000 ;
      LAYER met4 ;
        RECT 68.230000 183.875000 68.550000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 184.280000 68.550000 184.600000 ;
      LAYER met4 ;
        RECT 68.230000 184.280000 68.550000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 184.685000 68.550000 185.005000 ;
      LAYER met4 ;
        RECT 68.230000 184.685000 68.550000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 185.090000 68.550000 185.410000 ;
      LAYER met4 ;
        RECT 68.230000 185.090000 68.550000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 185.495000 68.550000 185.815000 ;
      LAYER met4 ;
        RECT 68.230000 185.495000 68.550000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 185.900000 68.550000 186.220000 ;
      LAYER met4 ;
        RECT 68.230000 185.900000 68.550000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 186.305000 68.550000 186.625000 ;
      LAYER met4 ;
        RECT 68.230000 186.305000 68.550000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 186.710000 68.550000 187.030000 ;
      LAYER met4 ;
        RECT 68.230000 186.710000 68.550000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 187.115000 68.550000 187.435000 ;
      LAYER met4 ;
        RECT 68.230000 187.115000 68.550000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 187.520000 68.550000 187.840000 ;
      LAYER met4 ;
        RECT 68.230000 187.520000 68.550000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 187.925000 68.550000 188.245000 ;
      LAYER met4 ;
        RECT 68.230000 187.925000 68.550000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 188.330000 68.550000 188.650000 ;
      LAYER met4 ;
        RECT 68.230000 188.330000 68.550000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 188.735000 68.550000 189.055000 ;
      LAYER met4 ;
        RECT 68.230000 188.735000 68.550000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 189.140000 68.550000 189.460000 ;
      LAYER met4 ;
        RECT 68.230000 189.140000 68.550000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 189.545000 68.550000 189.865000 ;
      LAYER met4 ;
        RECT 68.230000 189.545000 68.550000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 189.950000 68.550000 190.270000 ;
      LAYER met4 ;
        RECT 68.230000 189.950000 68.550000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 190.355000 68.550000 190.675000 ;
      LAYER met4 ;
        RECT 68.230000 190.355000 68.550000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 190.760000 68.550000 191.080000 ;
      LAYER met4 ;
        RECT 68.230000 190.760000 68.550000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 191.165000 68.550000 191.485000 ;
      LAYER met4 ;
        RECT 68.230000 191.165000 68.550000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 191.570000 68.550000 191.890000 ;
      LAYER met4 ;
        RECT 68.230000 191.570000 68.550000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 191.975000 68.550000 192.295000 ;
      LAYER met4 ;
        RECT 68.230000 191.975000 68.550000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 192.380000 68.550000 192.700000 ;
      LAYER met4 ;
        RECT 68.230000 192.380000 68.550000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 192.785000 68.550000 193.105000 ;
      LAYER met4 ;
        RECT 68.230000 192.785000 68.550000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 193.190000 68.550000 193.510000 ;
      LAYER met4 ;
        RECT 68.230000 193.190000 68.550000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 193.595000 68.550000 193.915000 ;
      LAYER met4 ;
        RECT 68.230000 193.595000 68.550000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 194.000000 68.550000 194.320000 ;
      LAYER met4 ;
        RECT 68.230000 194.000000 68.550000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 194.405000 68.550000 194.725000 ;
      LAYER met4 ;
        RECT 68.230000 194.405000 68.550000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 194.810000 68.550000 195.130000 ;
      LAYER met4 ;
        RECT 68.230000 194.810000 68.550000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 195.215000 68.550000 195.535000 ;
      LAYER met4 ;
        RECT 68.230000 195.215000 68.550000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 195.620000 68.550000 195.940000 ;
      LAYER met4 ;
        RECT 68.230000 195.620000 68.550000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 196.025000 68.550000 196.345000 ;
      LAYER met4 ;
        RECT 68.230000 196.025000 68.550000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 196.430000 68.550000 196.750000 ;
      LAYER met4 ;
        RECT 68.230000 196.430000 68.550000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 196.835000 68.550000 197.155000 ;
      LAYER met4 ;
        RECT 68.230000 196.835000 68.550000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 197.240000 68.550000 197.560000 ;
      LAYER met4 ;
        RECT 68.230000 197.240000 68.550000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 197.645000 68.550000 197.965000 ;
      LAYER met4 ;
        RECT 68.230000 197.645000 68.550000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 23.850000 68.590000 24.170000 ;
      LAYER met4 ;
        RECT 68.270000 23.850000 68.590000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 24.280000 68.590000 24.600000 ;
      LAYER met4 ;
        RECT 68.270000 24.280000 68.590000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 24.710000 68.590000 25.030000 ;
      LAYER met4 ;
        RECT 68.270000 24.710000 68.590000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 25.140000 68.590000 25.460000 ;
      LAYER met4 ;
        RECT 68.270000 25.140000 68.590000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 25.570000 68.590000 25.890000 ;
      LAYER met4 ;
        RECT 68.270000 25.570000 68.590000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 26.000000 68.590000 26.320000 ;
      LAYER met4 ;
        RECT 68.270000 26.000000 68.590000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 26.430000 68.590000 26.750000 ;
      LAYER met4 ;
        RECT 68.270000 26.430000 68.590000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 26.860000 68.590000 27.180000 ;
      LAYER met4 ;
        RECT 68.270000 26.860000 68.590000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 27.290000 68.590000 27.610000 ;
      LAYER met4 ;
        RECT 68.270000 27.290000 68.590000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 27.720000 68.590000 28.040000 ;
      LAYER met4 ;
        RECT 68.270000 27.720000 68.590000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 28.150000 68.590000 28.470000 ;
      LAYER met4 ;
        RECT 68.270000 28.150000 68.590000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 173.840000 68.960000 174.160000 ;
      LAYER met4 ;
        RECT 68.640000 173.840000 68.960000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 174.240000 68.960000 174.560000 ;
      LAYER met4 ;
        RECT 68.640000 174.240000 68.960000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 174.640000 68.960000 174.960000 ;
      LAYER met4 ;
        RECT 68.640000 174.640000 68.960000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 175.040000 68.960000 175.360000 ;
      LAYER met4 ;
        RECT 68.640000 175.040000 68.960000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 175.440000 68.960000 175.760000 ;
      LAYER met4 ;
        RECT 68.640000 175.440000 68.960000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 175.840000 68.960000 176.160000 ;
      LAYER met4 ;
        RECT 68.640000 175.840000 68.960000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 176.240000 68.960000 176.560000 ;
      LAYER met4 ;
        RECT 68.640000 176.240000 68.960000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 176.640000 68.960000 176.960000 ;
      LAYER met4 ;
        RECT 68.640000 176.640000 68.960000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 177.040000 68.960000 177.360000 ;
      LAYER met4 ;
        RECT 68.640000 177.040000 68.960000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 177.440000 68.960000 177.760000 ;
      LAYER met4 ;
        RECT 68.640000 177.440000 68.960000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 177.840000 68.960000 178.160000 ;
      LAYER met4 ;
        RECT 68.640000 177.840000 68.960000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 178.240000 68.960000 178.560000 ;
      LAYER met4 ;
        RECT 68.640000 178.240000 68.960000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 178.640000 68.960000 178.960000 ;
      LAYER met4 ;
        RECT 68.640000 178.640000 68.960000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 179.040000 68.960000 179.360000 ;
      LAYER met4 ;
        RECT 68.640000 179.040000 68.960000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 179.440000 68.960000 179.760000 ;
      LAYER met4 ;
        RECT 68.640000 179.440000 68.960000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 179.840000 68.960000 180.160000 ;
      LAYER met4 ;
        RECT 68.640000 179.840000 68.960000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 180.240000 68.960000 180.560000 ;
      LAYER met4 ;
        RECT 68.640000 180.240000 68.960000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 180.640000 68.960000 180.960000 ;
      LAYER met4 ;
        RECT 68.640000 180.640000 68.960000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 181.040000 68.960000 181.360000 ;
      LAYER met4 ;
        RECT 68.640000 181.040000 68.960000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 181.445000 68.960000 181.765000 ;
      LAYER met4 ;
        RECT 68.640000 181.445000 68.960000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 181.850000 68.960000 182.170000 ;
      LAYER met4 ;
        RECT 68.640000 181.850000 68.960000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 182.255000 68.960000 182.575000 ;
      LAYER met4 ;
        RECT 68.640000 182.255000 68.960000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 182.660000 68.960000 182.980000 ;
      LAYER met4 ;
        RECT 68.640000 182.660000 68.960000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 183.065000 68.960000 183.385000 ;
      LAYER met4 ;
        RECT 68.640000 183.065000 68.960000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 183.470000 68.960000 183.790000 ;
      LAYER met4 ;
        RECT 68.640000 183.470000 68.960000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 183.875000 68.960000 184.195000 ;
      LAYER met4 ;
        RECT 68.640000 183.875000 68.960000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 184.280000 68.960000 184.600000 ;
      LAYER met4 ;
        RECT 68.640000 184.280000 68.960000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 184.685000 68.960000 185.005000 ;
      LAYER met4 ;
        RECT 68.640000 184.685000 68.960000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 185.090000 68.960000 185.410000 ;
      LAYER met4 ;
        RECT 68.640000 185.090000 68.960000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 185.495000 68.960000 185.815000 ;
      LAYER met4 ;
        RECT 68.640000 185.495000 68.960000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 185.900000 68.960000 186.220000 ;
      LAYER met4 ;
        RECT 68.640000 185.900000 68.960000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 186.305000 68.960000 186.625000 ;
      LAYER met4 ;
        RECT 68.640000 186.305000 68.960000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 186.710000 68.960000 187.030000 ;
      LAYER met4 ;
        RECT 68.640000 186.710000 68.960000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 187.115000 68.960000 187.435000 ;
      LAYER met4 ;
        RECT 68.640000 187.115000 68.960000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 187.520000 68.960000 187.840000 ;
      LAYER met4 ;
        RECT 68.640000 187.520000 68.960000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 187.925000 68.960000 188.245000 ;
      LAYER met4 ;
        RECT 68.640000 187.925000 68.960000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 188.330000 68.960000 188.650000 ;
      LAYER met4 ;
        RECT 68.640000 188.330000 68.960000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 188.735000 68.960000 189.055000 ;
      LAYER met4 ;
        RECT 68.640000 188.735000 68.960000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 189.140000 68.960000 189.460000 ;
      LAYER met4 ;
        RECT 68.640000 189.140000 68.960000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 189.545000 68.960000 189.865000 ;
      LAYER met4 ;
        RECT 68.640000 189.545000 68.960000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 189.950000 68.960000 190.270000 ;
      LAYER met4 ;
        RECT 68.640000 189.950000 68.960000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 190.355000 68.960000 190.675000 ;
      LAYER met4 ;
        RECT 68.640000 190.355000 68.960000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 190.760000 68.960000 191.080000 ;
      LAYER met4 ;
        RECT 68.640000 190.760000 68.960000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 191.165000 68.960000 191.485000 ;
      LAYER met4 ;
        RECT 68.640000 191.165000 68.960000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 191.570000 68.960000 191.890000 ;
      LAYER met4 ;
        RECT 68.640000 191.570000 68.960000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 191.975000 68.960000 192.295000 ;
      LAYER met4 ;
        RECT 68.640000 191.975000 68.960000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 192.380000 68.960000 192.700000 ;
      LAYER met4 ;
        RECT 68.640000 192.380000 68.960000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 192.785000 68.960000 193.105000 ;
      LAYER met4 ;
        RECT 68.640000 192.785000 68.960000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 193.190000 68.960000 193.510000 ;
      LAYER met4 ;
        RECT 68.640000 193.190000 68.960000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 193.595000 68.960000 193.915000 ;
      LAYER met4 ;
        RECT 68.640000 193.595000 68.960000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 194.000000 68.960000 194.320000 ;
      LAYER met4 ;
        RECT 68.640000 194.000000 68.960000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 194.405000 68.960000 194.725000 ;
      LAYER met4 ;
        RECT 68.640000 194.405000 68.960000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 194.810000 68.960000 195.130000 ;
      LAYER met4 ;
        RECT 68.640000 194.810000 68.960000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 195.215000 68.960000 195.535000 ;
      LAYER met4 ;
        RECT 68.640000 195.215000 68.960000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 195.620000 68.960000 195.940000 ;
      LAYER met4 ;
        RECT 68.640000 195.620000 68.960000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 196.025000 68.960000 196.345000 ;
      LAYER met4 ;
        RECT 68.640000 196.025000 68.960000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 196.430000 68.960000 196.750000 ;
      LAYER met4 ;
        RECT 68.640000 196.430000 68.960000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 196.835000 68.960000 197.155000 ;
      LAYER met4 ;
        RECT 68.640000 196.835000 68.960000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 197.240000 68.960000 197.560000 ;
      LAYER met4 ;
        RECT 68.640000 197.240000 68.960000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.640000 197.645000 68.960000 197.965000 ;
      LAYER met4 ;
        RECT 68.640000 197.645000 68.960000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 23.850000 68.995000 24.170000 ;
      LAYER met4 ;
        RECT 68.675000 23.850000 68.995000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 24.280000 68.995000 24.600000 ;
      LAYER met4 ;
        RECT 68.675000 24.280000 68.995000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 24.710000 68.995000 25.030000 ;
      LAYER met4 ;
        RECT 68.675000 24.710000 68.995000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 25.140000 68.995000 25.460000 ;
      LAYER met4 ;
        RECT 68.675000 25.140000 68.995000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 25.570000 68.995000 25.890000 ;
      LAYER met4 ;
        RECT 68.675000 25.570000 68.995000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 26.000000 68.995000 26.320000 ;
      LAYER met4 ;
        RECT 68.675000 26.000000 68.995000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 26.430000 68.995000 26.750000 ;
      LAYER met4 ;
        RECT 68.675000 26.430000 68.995000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 26.860000 68.995000 27.180000 ;
      LAYER met4 ;
        RECT 68.675000 26.860000 68.995000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 27.290000 68.995000 27.610000 ;
      LAYER met4 ;
        RECT 68.675000 27.290000 68.995000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 27.720000 68.995000 28.040000 ;
      LAYER met4 ;
        RECT 68.675000 27.720000 68.995000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 28.150000 68.995000 28.470000 ;
      LAYER met4 ;
        RECT 68.675000 28.150000 68.995000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 173.840000 69.370000 174.160000 ;
      LAYER met4 ;
        RECT 69.050000 173.840000 69.370000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 174.240000 69.370000 174.560000 ;
      LAYER met4 ;
        RECT 69.050000 174.240000 69.370000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 174.640000 69.370000 174.960000 ;
      LAYER met4 ;
        RECT 69.050000 174.640000 69.370000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 175.040000 69.370000 175.360000 ;
      LAYER met4 ;
        RECT 69.050000 175.040000 69.370000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 175.440000 69.370000 175.760000 ;
      LAYER met4 ;
        RECT 69.050000 175.440000 69.370000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 175.840000 69.370000 176.160000 ;
      LAYER met4 ;
        RECT 69.050000 175.840000 69.370000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 176.240000 69.370000 176.560000 ;
      LAYER met4 ;
        RECT 69.050000 176.240000 69.370000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 176.640000 69.370000 176.960000 ;
      LAYER met4 ;
        RECT 69.050000 176.640000 69.370000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 177.040000 69.370000 177.360000 ;
      LAYER met4 ;
        RECT 69.050000 177.040000 69.370000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 177.440000 69.370000 177.760000 ;
      LAYER met4 ;
        RECT 69.050000 177.440000 69.370000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 177.840000 69.370000 178.160000 ;
      LAYER met4 ;
        RECT 69.050000 177.840000 69.370000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 178.240000 69.370000 178.560000 ;
      LAYER met4 ;
        RECT 69.050000 178.240000 69.370000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 178.640000 69.370000 178.960000 ;
      LAYER met4 ;
        RECT 69.050000 178.640000 69.370000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 179.040000 69.370000 179.360000 ;
      LAYER met4 ;
        RECT 69.050000 179.040000 69.370000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 179.440000 69.370000 179.760000 ;
      LAYER met4 ;
        RECT 69.050000 179.440000 69.370000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 179.840000 69.370000 180.160000 ;
      LAYER met4 ;
        RECT 69.050000 179.840000 69.370000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 180.240000 69.370000 180.560000 ;
      LAYER met4 ;
        RECT 69.050000 180.240000 69.370000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 180.640000 69.370000 180.960000 ;
      LAYER met4 ;
        RECT 69.050000 180.640000 69.370000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 181.040000 69.370000 181.360000 ;
      LAYER met4 ;
        RECT 69.050000 181.040000 69.370000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 181.445000 69.370000 181.765000 ;
      LAYER met4 ;
        RECT 69.050000 181.445000 69.370000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 181.850000 69.370000 182.170000 ;
      LAYER met4 ;
        RECT 69.050000 181.850000 69.370000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 182.255000 69.370000 182.575000 ;
      LAYER met4 ;
        RECT 69.050000 182.255000 69.370000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 182.660000 69.370000 182.980000 ;
      LAYER met4 ;
        RECT 69.050000 182.660000 69.370000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 183.065000 69.370000 183.385000 ;
      LAYER met4 ;
        RECT 69.050000 183.065000 69.370000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 183.470000 69.370000 183.790000 ;
      LAYER met4 ;
        RECT 69.050000 183.470000 69.370000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 183.875000 69.370000 184.195000 ;
      LAYER met4 ;
        RECT 69.050000 183.875000 69.370000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 184.280000 69.370000 184.600000 ;
      LAYER met4 ;
        RECT 69.050000 184.280000 69.370000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 184.685000 69.370000 185.005000 ;
      LAYER met4 ;
        RECT 69.050000 184.685000 69.370000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 185.090000 69.370000 185.410000 ;
      LAYER met4 ;
        RECT 69.050000 185.090000 69.370000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 185.495000 69.370000 185.815000 ;
      LAYER met4 ;
        RECT 69.050000 185.495000 69.370000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 185.900000 69.370000 186.220000 ;
      LAYER met4 ;
        RECT 69.050000 185.900000 69.370000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 186.305000 69.370000 186.625000 ;
      LAYER met4 ;
        RECT 69.050000 186.305000 69.370000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 186.710000 69.370000 187.030000 ;
      LAYER met4 ;
        RECT 69.050000 186.710000 69.370000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 187.115000 69.370000 187.435000 ;
      LAYER met4 ;
        RECT 69.050000 187.115000 69.370000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 187.520000 69.370000 187.840000 ;
      LAYER met4 ;
        RECT 69.050000 187.520000 69.370000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 187.925000 69.370000 188.245000 ;
      LAYER met4 ;
        RECT 69.050000 187.925000 69.370000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 188.330000 69.370000 188.650000 ;
      LAYER met4 ;
        RECT 69.050000 188.330000 69.370000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 188.735000 69.370000 189.055000 ;
      LAYER met4 ;
        RECT 69.050000 188.735000 69.370000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 189.140000 69.370000 189.460000 ;
      LAYER met4 ;
        RECT 69.050000 189.140000 69.370000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 189.545000 69.370000 189.865000 ;
      LAYER met4 ;
        RECT 69.050000 189.545000 69.370000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 189.950000 69.370000 190.270000 ;
      LAYER met4 ;
        RECT 69.050000 189.950000 69.370000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 190.355000 69.370000 190.675000 ;
      LAYER met4 ;
        RECT 69.050000 190.355000 69.370000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 190.760000 69.370000 191.080000 ;
      LAYER met4 ;
        RECT 69.050000 190.760000 69.370000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 191.165000 69.370000 191.485000 ;
      LAYER met4 ;
        RECT 69.050000 191.165000 69.370000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 191.570000 69.370000 191.890000 ;
      LAYER met4 ;
        RECT 69.050000 191.570000 69.370000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 191.975000 69.370000 192.295000 ;
      LAYER met4 ;
        RECT 69.050000 191.975000 69.370000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 192.380000 69.370000 192.700000 ;
      LAYER met4 ;
        RECT 69.050000 192.380000 69.370000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 192.785000 69.370000 193.105000 ;
      LAYER met4 ;
        RECT 69.050000 192.785000 69.370000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 193.190000 69.370000 193.510000 ;
      LAYER met4 ;
        RECT 69.050000 193.190000 69.370000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 193.595000 69.370000 193.915000 ;
      LAYER met4 ;
        RECT 69.050000 193.595000 69.370000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 194.000000 69.370000 194.320000 ;
      LAYER met4 ;
        RECT 69.050000 194.000000 69.370000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 194.405000 69.370000 194.725000 ;
      LAYER met4 ;
        RECT 69.050000 194.405000 69.370000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 194.810000 69.370000 195.130000 ;
      LAYER met4 ;
        RECT 69.050000 194.810000 69.370000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 195.215000 69.370000 195.535000 ;
      LAYER met4 ;
        RECT 69.050000 195.215000 69.370000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 195.620000 69.370000 195.940000 ;
      LAYER met4 ;
        RECT 69.050000 195.620000 69.370000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 196.025000 69.370000 196.345000 ;
      LAYER met4 ;
        RECT 69.050000 196.025000 69.370000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 196.430000 69.370000 196.750000 ;
      LAYER met4 ;
        RECT 69.050000 196.430000 69.370000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 196.835000 69.370000 197.155000 ;
      LAYER met4 ;
        RECT 69.050000 196.835000 69.370000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 197.240000 69.370000 197.560000 ;
      LAYER met4 ;
        RECT 69.050000 197.240000 69.370000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 197.645000 69.370000 197.965000 ;
      LAYER met4 ;
        RECT 69.050000 197.645000 69.370000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 23.850000 69.400000 24.170000 ;
      LAYER met4 ;
        RECT 69.080000 23.850000 69.400000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 24.280000 69.400000 24.600000 ;
      LAYER met4 ;
        RECT 69.080000 24.280000 69.400000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 24.710000 69.400000 25.030000 ;
      LAYER met4 ;
        RECT 69.080000 24.710000 69.400000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 25.140000 69.400000 25.460000 ;
      LAYER met4 ;
        RECT 69.080000 25.140000 69.400000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 25.570000 69.400000 25.890000 ;
      LAYER met4 ;
        RECT 69.080000 25.570000 69.400000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 26.000000 69.400000 26.320000 ;
      LAYER met4 ;
        RECT 69.080000 26.000000 69.400000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 26.430000 69.400000 26.750000 ;
      LAYER met4 ;
        RECT 69.080000 26.430000 69.400000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 26.860000 69.400000 27.180000 ;
      LAYER met4 ;
        RECT 69.080000 26.860000 69.400000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 27.290000 69.400000 27.610000 ;
      LAYER met4 ;
        RECT 69.080000 27.290000 69.400000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 27.720000 69.400000 28.040000 ;
      LAYER met4 ;
        RECT 69.080000 27.720000 69.400000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 28.150000 69.400000 28.470000 ;
      LAYER met4 ;
        RECT 69.080000 28.150000 69.400000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 173.840000 69.780000 174.160000 ;
      LAYER met4 ;
        RECT 69.460000 173.840000 69.780000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 174.240000 69.780000 174.560000 ;
      LAYER met4 ;
        RECT 69.460000 174.240000 69.780000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 174.640000 69.780000 174.960000 ;
      LAYER met4 ;
        RECT 69.460000 174.640000 69.780000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 175.040000 69.780000 175.360000 ;
      LAYER met4 ;
        RECT 69.460000 175.040000 69.780000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 175.440000 69.780000 175.760000 ;
      LAYER met4 ;
        RECT 69.460000 175.440000 69.780000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 175.840000 69.780000 176.160000 ;
      LAYER met4 ;
        RECT 69.460000 175.840000 69.780000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 176.240000 69.780000 176.560000 ;
      LAYER met4 ;
        RECT 69.460000 176.240000 69.780000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 176.640000 69.780000 176.960000 ;
      LAYER met4 ;
        RECT 69.460000 176.640000 69.780000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 177.040000 69.780000 177.360000 ;
      LAYER met4 ;
        RECT 69.460000 177.040000 69.780000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 177.440000 69.780000 177.760000 ;
      LAYER met4 ;
        RECT 69.460000 177.440000 69.780000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 177.840000 69.780000 178.160000 ;
      LAYER met4 ;
        RECT 69.460000 177.840000 69.780000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 178.240000 69.780000 178.560000 ;
      LAYER met4 ;
        RECT 69.460000 178.240000 69.780000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 178.640000 69.780000 178.960000 ;
      LAYER met4 ;
        RECT 69.460000 178.640000 69.780000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 179.040000 69.780000 179.360000 ;
      LAYER met4 ;
        RECT 69.460000 179.040000 69.780000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 179.440000 69.780000 179.760000 ;
      LAYER met4 ;
        RECT 69.460000 179.440000 69.780000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 179.840000 69.780000 180.160000 ;
      LAYER met4 ;
        RECT 69.460000 179.840000 69.780000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 180.240000 69.780000 180.560000 ;
      LAYER met4 ;
        RECT 69.460000 180.240000 69.780000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 180.640000 69.780000 180.960000 ;
      LAYER met4 ;
        RECT 69.460000 180.640000 69.780000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 181.040000 69.780000 181.360000 ;
      LAYER met4 ;
        RECT 69.460000 181.040000 69.780000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 181.445000 69.780000 181.765000 ;
      LAYER met4 ;
        RECT 69.460000 181.445000 69.780000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 181.850000 69.780000 182.170000 ;
      LAYER met4 ;
        RECT 69.460000 181.850000 69.780000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 182.255000 69.780000 182.575000 ;
      LAYER met4 ;
        RECT 69.460000 182.255000 69.780000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 182.660000 69.780000 182.980000 ;
      LAYER met4 ;
        RECT 69.460000 182.660000 69.780000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 183.065000 69.780000 183.385000 ;
      LAYER met4 ;
        RECT 69.460000 183.065000 69.780000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 183.470000 69.780000 183.790000 ;
      LAYER met4 ;
        RECT 69.460000 183.470000 69.780000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 183.875000 69.780000 184.195000 ;
      LAYER met4 ;
        RECT 69.460000 183.875000 69.780000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 184.280000 69.780000 184.600000 ;
      LAYER met4 ;
        RECT 69.460000 184.280000 69.780000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 184.685000 69.780000 185.005000 ;
      LAYER met4 ;
        RECT 69.460000 184.685000 69.780000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 185.090000 69.780000 185.410000 ;
      LAYER met4 ;
        RECT 69.460000 185.090000 69.780000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 185.495000 69.780000 185.815000 ;
      LAYER met4 ;
        RECT 69.460000 185.495000 69.780000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 185.900000 69.780000 186.220000 ;
      LAYER met4 ;
        RECT 69.460000 185.900000 69.780000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 186.305000 69.780000 186.625000 ;
      LAYER met4 ;
        RECT 69.460000 186.305000 69.780000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 186.710000 69.780000 187.030000 ;
      LAYER met4 ;
        RECT 69.460000 186.710000 69.780000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 187.115000 69.780000 187.435000 ;
      LAYER met4 ;
        RECT 69.460000 187.115000 69.780000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 187.520000 69.780000 187.840000 ;
      LAYER met4 ;
        RECT 69.460000 187.520000 69.780000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 187.925000 69.780000 188.245000 ;
      LAYER met4 ;
        RECT 69.460000 187.925000 69.780000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 188.330000 69.780000 188.650000 ;
      LAYER met4 ;
        RECT 69.460000 188.330000 69.780000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 188.735000 69.780000 189.055000 ;
      LAYER met4 ;
        RECT 69.460000 188.735000 69.780000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 189.140000 69.780000 189.460000 ;
      LAYER met4 ;
        RECT 69.460000 189.140000 69.780000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 189.545000 69.780000 189.865000 ;
      LAYER met4 ;
        RECT 69.460000 189.545000 69.780000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 189.950000 69.780000 190.270000 ;
      LAYER met4 ;
        RECT 69.460000 189.950000 69.780000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 190.355000 69.780000 190.675000 ;
      LAYER met4 ;
        RECT 69.460000 190.355000 69.780000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 190.760000 69.780000 191.080000 ;
      LAYER met4 ;
        RECT 69.460000 190.760000 69.780000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 191.165000 69.780000 191.485000 ;
      LAYER met4 ;
        RECT 69.460000 191.165000 69.780000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 191.570000 69.780000 191.890000 ;
      LAYER met4 ;
        RECT 69.460000 191.570000 69.780000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 191.975000 69.780000 192.295000 ;
      LAYER met4 ;
        RECT 69.460000 191.975000 69.780000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 192.380000 69.780000 192.700000 ;
      LAYER met4 ;
        RECT 69.460000 192.380000 69.780000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 192.785000 69.780000 193.105000 ;
      LAYER met4 ;
        RECT 69.460000 192.785000 69.780000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 193.190000 69.780000 193.510000 ;
      LAYER met4 ;
        RECT 69.460000 193.190000 69.780000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 193.595000 69.780000 193.915000 ;
      LAYER met4 ;
        RECT 69.460000 193.595000 69.780000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 194.000000 69.780000 194.320000 ;
      LAYER met4 ;
        RECT 69.460000 194.000000 69.780000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 194.405000 69.780000 194.725000 ;
      LAYER met4 ;
        RECT 69.460000 194.405000 69.780000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 194.810000 69.780000 195.130000 ;
      LAYER met4 ;
        RECT 69.460000 194.810000 69.780000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 195.215000 69.780000 195.535000 ;
      LAYER met4 ;
        RECT 69.460000 195.215000 69.780000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 195.620000 69.780000 195.940000 ;
      LAYER met4 ;
        RECT 69.460000 195.620000 69.780000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 196.025000 69.780000 196.345000 ;
      LAYER met4 ;
        RECT 69.460000 196.025000 69.780000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 196.430000 69.780000 196.750000 ;
      LAYER met4 ;
        RECT 69.460000 196.430000 69.780000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 196.835000 69.780000 197.155000 ;
      LAYER met4 ;
        RECT 69.460000 196.835000 69.780000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 197.240000 69.780000 197.560000 ;
      LAYER met4 ;
        RECT 69.460000 197.240000 69.780000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.460000 197.645000 69.780000 197.965000 ;
      LAYER met4 ;
        RECT 69.460000 197.645000 69.780000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 23.850000 69.805000 24.170000 ;
      LAYER met4 ;
        RECT 69.485000 23.850000 69.805000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 24.280000 69.805000 24.600000 ;
      LAYER met4 ;
        RECT 69.485000 24.280000 69.805000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 24.710000 69.805000 25.030000 ;
      LAYER met4 ;
        RECT 69.485000 24.710000 69.805000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 25.140000 69.805000 25.460000 ;
      LAYER met4 ;
        RECT 69.485000 25.140000 69.805000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 25.570000 69.805000 25.890000 ;
      LAYER met4 ;
        RECT 69.485000 25.570000 69.805000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 26.000000 69.805000 26.320000 ;
      LAYER met4 ;
        RECT 69.485000 26.000000 69.805000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 26.430000 69.805000 26.750000 ;
      LAYER met4 ;
        RECT 69.485000 26.430000 69.805000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 26.860000 69.805000 27.180000 ;
      LAYER met4 ;
        RECT 69.485000 26.860000 69.805000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 27.290000 69.805000 27.610000 ;
      LAYER met4 ;
        RECT 69.485000 27.290000 69.805000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 27.720000 69.805000 28.040000 ;
      LAYER met4 ;
        RECT 69.485000 27.720000 69.805000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 28.150000 69.805000 28.470000 ;
      LAYER met4 ;
        RECT 69.485000 28.150000 69.805000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 173.840000 70.190000 174.160000 ;
      LAYER met4 ;
        RECT 69.870000 173.840000 70.190000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 174.240000 70.190000 174.560000 ;
      LAYER met4 ;
        RECT 69.870000 174.240000 70.190000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 174.640000 70.190000 174.960000 ;
      LAYER met4 ;
        RECT 69.870000 174.640000 70.190000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 175.040000 70.190000 175.360000 ;
      LAYER met4 ;
        RECT 69.870000 175.040000 70.190000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 175.440000 70.190000 175.760000 ;
      LAYER met4 ;
        RECT 69.870000 175.440000 70.190000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 175.840000 70.190000 176.160000 ;
      LAYER met4 ;
        RECT 69.870000 175.840000 70.190000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 176.240000 70.190000 176.560000 ;
      LAYER met4 ;
        RECT 69.870000 176.240000 70.190000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 176.640000 70.190000 176.960000 ;
      LAYER met4 ;
        RECT 69.870000 176.640000 70.190000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 177.040000 70.190000 177.360000 ;
      LAYER met4 ;
        RECT 69.870000 177.040000 70.190000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 177.440000 70.190000 177.760000 ;
      LAYER met4 ;
        RECT 69.870000 177.440000 70.190000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 177.840000 70.190000 178.160000 ;
      LAYER met4 ;
        RECT 69.870000 177.840000 70.190000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 178.240000 70.190000 178.560000 ;
      LAYER met4 ;
        RECT 69.870000 178.240000 70.190000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 178.640000 70.190000 178.960000 ;
      LAYER met4 ;
        RECT 69.870000 178.640000 70.190000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 179.040000 70.190000 179.360000 ;
      LAYER met4 ;
        RECT 69.870000 179.040000 70.190000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 179.440000 70.190000 179.760000 ;
      LAYER met4 ;
        RECT 69.870000 179.440000 70.190000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 179.840000 70.190000 180.160000 ;
      LAYER met4 ;
        RECT 69.870000 179.840000 70.190000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 180.240000 70.190000 180.560000 ;
      LAYER met4 ;
        RECT 69.870000 180.240000 70.190000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 180.640000 70.190000 180.960000 ;
      LAYER met4 ;
        RECT 69.870000 180.640000 70.190000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 181.040000 70.190000 181.360000 ;
      LAYER met4 ;
        RECT 69.870000 181.040000 70.190000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 181.445000 70.190000 181.765000 ;
      LAYER met4 ;
        RECT 69.870000 181.445000 70.190000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 181.850000 70.190000 182.170000 ;
      LAYER met4 ;
        RECT 69.870000 181.850000 70.190000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 182.255000 70.190000 182.575000 ;
      LAYER met4 ;
        RECT 69.870000 182.255000 70.190000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 182.660000 70.190000 182.980000 ;
      LAYER met4 ;
        RECT 69.870000 182.660000 70.190000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 183.065000 70.190000 183.385000 ;
      LAYER met4 ;
        RECT 69.870000 183.065000 70.190000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 183.470000 70.190000 183.790000 ;
      LAYER met4 ;
        RECT 69.870000 183.470000 70.190000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 183.875000 70.190000 184.195000 ;
      LAYER met4 ;
        RECT 69.870000 183.875000 70.190000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 184.280000 70.190000 184.600000 ;
      LAYER met4 ;
        RECT 69.870000 184.280000 70.190000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 184.685000 70.190000 185.005000 ;
      LAYER met4 ;
        RECT 69.870000 184.685000 70.190000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 185.090000 70.190000 185.410000 ;
      LAYER met4 ;
        RECT 69.870000 185.090000 70.190000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 185.495000 70.190000 185.815000 ;
      LAYER met4 ;
        RECT 69.870000 185.495000 70.190000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 185.900000 70.190000 186.220000 ;
      LAYER met4 ;
        RECT 69.870000 185.900000 70.190000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 186.305000 70.190000 186.625000 ;
      LAYER met4 ;
        RECT 69.870000 186.305000 70.190000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 186.710000 70.190000 187.030000 ;
      LAYER met4 ;
        RECT 69.870000 186.710000 70.190000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 187.115000 70.190000 187.435000 ;
      LAYER met4 ;
        RECT 69.870000 187.115000 70.190000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 187.520000 70.190000 187.840000 ;
      LAYER met4 ;
        RECT 69.870000 187.520000 70.190000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 187.925000 70.190000 188.245000 ;
      LAYER met4 ;
        RECT 69.870000 187.925000 70.190000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 188.330000 70.190000 188.650000 ;
      LAYER met4 ;
        RECT 69.870000 188.330000 70.190000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 188.735000 70.190000 189.055000 ;
      LAYER met4 ;
        RECT 69.870000 188.735000 70.190000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 189.140000 70.190000 189.460000 ;
      LAYER met4 ;
        RECT 69.870000 189.140000 70.190000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 189.545000 70.190000 189.865000 ;
      LAYER met4 ;
        RECT 69.870000 189.545000 70.190000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 189.950000 70.190000 190.270000 ;
      LAYER met4 ;
        RECT 69.870000 189.950000 70.190000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 190.355000 70.190000 190.675000 ;
      LAYER met4 ;
        RECT 69.870000 190.355000 70.190000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 190.760000 70.190000 191.080000 ;
      LAYER met4 ;
        RECT 69.870000 190.760000 70.190000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 191.165000 70.190000 191.485000 ;
      LAYER met4 ;
        RECT 69.870000 191.165000 70.190000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 191.570000 70.190000 191.890000 ;
      LAYER met4 ;
        RECT 69.870000 191.570000 70.190000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 191.975000 70.190000 192.295000 ;
      LAYER met4 ;
        RECT 69.870000 191.975000 70.190000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 192.380000 70.190000 192.700000 ;
      LAYER met4 ;
        RECT 69.870000 192.380000 70.190000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 192.785000 70.190000 193.105000 ;
      LAYER met4 ;
        RECT 69.870000 192.785000 70.190000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 193.190000 70.190000 193.510000 ;
      LAYER met4 ;
        RECT 69.870000 193.190000 70.190000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 193.595000 70.190000 193.915000 ;
      LAYER met4 ;
        RECT 69.870000 193.595000 70.190000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 194.000000 70.190000 194.320000 ;
      LAYER met4 ;
        RECT 69.870000 194.000000 70.190000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 194.405000 70.190000 194.725000 ;
      LAYER met4 ;
        RECT 69.870000 194.405000 70.190000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 194.810000 70.190000 195.130000 ;
      LAYER met4 ;
        RECT 69.870000 194.810000 70.190000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 195.215000 70.190000 195.535000 ;
      LAYER met4 ;
        RECT 69.870000 195.215000 70.190000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 195.620000 70.190000 195.940000 ;
      LAYER met4 ;
        RECT 69.870000 195.620000 70.190000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 196.025000 70.190000 196.345000 ;
      LAYER met4 ;
        RECT 69.870000 196.025000 70.190000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 196.430000 70.190000 196.750000 ;
      LAYER met4 ;
        RECT 69.870000 196.430000 70.190000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 196.835000 70.190000 197.155000 ;
      LAYER met4 ;
        RECT 69.870000 196.835000 70.190000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 197.240000 70.190000 197.560000 ;
      LAYER met4 ;
        RECT 69.870000 197.240000 70.190000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.870000 197.645000 70.190000 197.965000 ;
      LAYER met4 ;
        RECT 69.870000 197.645000 70.190000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 23.850000 70.210000 24.170000 ;
      LAYER met4 ;
        RECT 69.890000 23.850000 70.210000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 24.280000 70.210000 24.600000 ;
      LAYER met4 ;
        RECT 69.890000 24.280000 70.210000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 24.710000 70.210000 25.030000 ;
      LAYER met4 ;
        RECT 69.890000 24.710000 70.210000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 25.140000 70.210000 25.460000 ;
      LAYER met4 ;
        RECT 69.890000 25.140000 70.210000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 25.570000 70.210000 25.890000 ;
      LAYER met4 ;
        RECT 69.890000 25.570000 70.210000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 26.000000 70.210000 26.320000 ;
      LAYER met4 ;
        RECT 69.890000 26.000000 70.210000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 26.430000 70.210000 26.750000 ;
      LAYER met4 ;
        RECT 69.890000 26.430000 70.210000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 26.860000 70.210000 27.180000 ;
      LAYER met4 ;
        RECT 69.890000 26.860000 70.210000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 27.290000 70.210000 27.610000 ;
      LAYER met4 ;
        RECT 69.890000 27.290000 70.210000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 27.720000 70.210000 28.040000 ;
      LAYER met4 ;
        RECT 69.890000 27.720000 70.210000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 28.150000 70.210000 28.470000 ;
      LAYER met4 ;
        RECT 69.890000 28.150000 70.210000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.015000 173.900000 7.215000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.015000 174.300000 7.215000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.015000 174.700000 7.215000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.015000 175.100000 7.215000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.015000 175.500000 7.215000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.015000 175.900000 7.215000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.015000 176.300000 7.215000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.015000 176.700000 7.215000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.015000 177.100000 7.215000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.015000 177.500000 7.215000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.015000 177.900000 7.215000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.015000 178.300000 7.215000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.015000 178.700000 7.215000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.015000 179.100000 7.215000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.015000 179.500000 7.215000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.015000 179.900000 7.215000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.015000 180.300000 7.215000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.015000 180.700000 7.215000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.015000 181.100000 7.215000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 23.850000 7.360000 24.170000 ;
      LAYER met4 ;
        RECT 7.040000 23.850000 7.360000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 24.280000 7.360000 24.600000 ;
      LAYER met4 ;
        RECT 7.040000 24.280000 7.360000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 24.710000 7.360000 25.030000 ;
      LAYER met4 ;
        RECT 7.040000 24.710000 7.360000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 25.140000 7.360000 25.460000 ;
      LAYER met4 ;
        RECT 7.040000 25.140000 7.360000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 25.570000 7.360000 25.890000 ;
      LAYER met4 ;
        RECT 7.040000 25.570000 7.360000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 26.000000 7.360000 26.320000 ;
      LAYER met4 ;
        RECT 7.040000 26.000000 7.360000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 26.430000 7.360000 26.750000 ;
      LAYER met4 ;
        RECT 7.040000 26.430000 7.360000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 26.860000 7.360000 27.180000 ;
      LAYER met4 ;
        RECT 7.040000 26.860000 7.360000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 27.290000 7.360000 27.610000 ;
      LAYER met4 ;
        RECT 7.040000 27.290000 7.360000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 27.720000 7.360000 28.040000 ;
      LAYER met4 ;
        RECT 7.040000 27.720000 7.360000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 28.150000 7.360000 28.470000 ;
      LAYER met4 ;
        RECT 7.040000 28.150000 7.360000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 181.445000 7.675000 181.765000 ;
      LAYER met4 ;
        RECT 7.355000 181.445000 7.675000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 181.850000 7.675000 182.170000 ;
      LAYER met4 ;
        RECT 7.355000 181.850000 7.675000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 182.255000 7.675000 182.575000 ;
      LAYER met4 ;
        RECT 7.355000 182.255000 7.675000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 182.660000 7.675000 182.980000 ;
      LAYER met4 ;
        RECT 7.355000 182.660000 7.675000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 183.065000 7.675000 183.385000 ;
      LAYER met4 ;
        RECT 7.355000 183.065000 7.675000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 183.470000 7.675000 183.790000 ;
      LAYER met4 ;
        RECT 7.355000 183.470000 7.675000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 183.875000 7.675000 184.195000 ;
      LAYER met4 ;
        RECT 7.355000 183.875000 7.675000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 184.280000 7.675000 184.600000 ;
      LAYER met4 ;
        RECT 7.355000 184.280000 7.675000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 184.685000 7.675000 185.005000 ;
      LAYER met4 ;
        RECT 7.355000 184.685000 7.675000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 185.090000 7.675000 185.410000 ;
      LAYER met4 ;
        RECT 7.355000 185.090000 7.675000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 185.495000 7.675000 185.815000 ;
      LAYER met4 ;
        RECT 7.355000 185.495000 7.675000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 185.900000 7.675000 186.220000 ;
      LAYER met4 ;
        RECT 7.355000 185.900000 7.675000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 186.305000 7.675000 186.625000 ;
      LAYER met4 ;
        RECT 7.355000 186.305000 7.675000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 186.710000 7.675000 187.030000 ;
      LAYER met4 ;
        RECT 7.355000 186.710000 7.675000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 187.115000 7.675000 187.435000 ;
      LAYER met4 ;
        RECT 7.355000 187.115000 7.675000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 187.520000 7.675000 187.840000 ;
      LAYER met4 ;
        RECT 7.355000 187.520000 7.675000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 187.925000 7.675000 188.245000 ;
      LAYER met4 ;
        RECT 7.355000 187.925000 7.675000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 188.330000 7.675000 188.650000 ;
      LAYER met4 ;
        RECT 7.355000 188.330000 7.675000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 188.735000 7.675000 189.055000 ;
      LAYER met4 ;
        RECT 7.355000 188.735000 7.675000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 189.140000 7.675000 189.460000 ;
      LAYER met4 ;
        RECT 7.355000 189.140000 7.675000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 189.545000 7.675000 189.865000 ;
      LAYER met4 ;
        RECT 7.355000 189.545000 7.675000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 189.950000 7.675000 190.270000 ;
      LAYER met4 ;
        RECT 7.355000 189.950000 7.675000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 190.355000 7.675000 190.675000 ;
      LAYER met4 ;
        RECT 7.355000 190.355000 7.675000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 190.760000 7.675000 191.080000 ;
      LAYER met4 ;
        RECT 7.355000 190.760000 7.675000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 191.165000 7.675000 191.485000 ;
      LAYER met4 ;
        RECT 7.355000 191.165000 7.675000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 191.570000 7.675000 191.890000 ;
      LAYER met4 ;
        RECT 7.355000 191.570000 7.675000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 191.975000 7.675000 192.295000 ;
      LAYER met4 ;
        RECT 7.355000 191.975000 7.675000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 192.380000 7.675000 192.700000 ;
      LAYER met4 ;
        RECT 7.355000 192.380000 7.675000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 192.785000 7.675000 193.105000 ;
      LAYER met4 ;
        RECT 7.355000 192.785000 7.675000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 193.190000 7.675000 193.510000 ;
      LAYER met4 ;
        RECT 7.355000 193.190000 7.675000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 193.595000 7.675000 193.915000 ;
      LAYER met4 ;
        RECT 7.355000 193.595000 7.675000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 194.000000 7.675000 194.320000 ;
      LAYER met4 ;
        RECT 7.355000 194.000000 7.675000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 194.405000 7.675000 194.725000 ;
      LAYER met4 ;
        RECT 7.355000 194.405000 7.675000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 194.810000 7.675000 195.130000 ;
      LAYER met4 ;
        RECT 7.355000 194.810000 7.675000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 195.215000 7.675000 195.535000 ;
      LAYER met4 ;
        RECT 7.355000 195.215000 7.675000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 195.620000 7.675000 195.940000 ;
      LAYER met4 ;
        RECT 7.355000 195.620000 7.675000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 196.025000 7.675000 196.345000 ;
      LAYER met4 ;
        RECT 7.355000 196.025000 7.675000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 196.430000 7.675000 196.750000 ;
      LAYER met4 ;
        RECT 7.355000 196.430000 7.675000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 196.835000 7.675000 197.155000 ;
      LAYER met4 ;
        RECT 7.355000 196.835000 7.675000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 197.240000 7.675000 197.560000 ;
      LAYER met4 ;
        RECT 7.355000 197.240000 7.675000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355000 197.645000 7.675000 197.965000 ;
      LAYER met4 ;
        RECT 7.355000 197.645000 7.675000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.415000 173.900000 7.615000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.415000 174.300000 7.615000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.415000 174.700000 7.615000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.415000 175.100000 7.615000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.415000 175.500000 7.615000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.415000 175.900000 7.615000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.415000 176.300000 7.615000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.415000 176.700000 7.615000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.415000 177.100000 7.615000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.415000 177.500000 7.615000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.415000 177.900000 7.615000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.415000 178.300000 7.615000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.415000 178.700000 7.615000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.415000 179.100000 7.615000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.415000 179.500000 7.615000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.415000 179.900000 7.615000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.415000 180.300000 7.615000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.415000 180.700000 7.615000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.415000 181.100000 7.615000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 23.850000 7.765000 24.170000 ;
      LAYER met4 ;
        RECT 7.445000 23.850000 7.765000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 24.280000 7.765000 24.600000 ;
      LAYER met4 ;
        RECT 7.445000 24.280000 7.765000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 24.710000 7.765000 25.030000 ;
      LAYER met4 ;
        RECT 7.445000 24.710000 7.765000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 25.140000 7.765000 25.460000 ;
      LAYER met4 ;
        RECT 7.445000 25.140000 7.765000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 25.570000 7.765000 25.890000 ;
      LAYER met4 ;
        RECT 7.445000 25.570000 7.765000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 26.000000 7.765000 26.320000 ;
      LAYER met4 ;
        RECT 7.445000 26.000000 7.765000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 26.430000 7.765000 26.750000 ;
      LAYER met4 ;
        RECT 7.445000 26.430000 7.765000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 26.860000 7.765000 27.180000 ;
      LAYER met4 ;
        RECT 7.445000 26.860000 7.765000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 27.290000 7.765000 27.610000 ;
      LAYER met4 ;
        RECT 7.445000 27.290000 7.765000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 27.720000 7.765000 28.040000 ;
      LAYER met4 ;
        RECT 7.445000 27.720000 7.765000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 28.150000 7.765000 28.470000 ;
      LAYER met4 ;
        RECT 7.445000 28.150000 7.765000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 181.445000 8.075000 181.765000 ;
      LAYER met4 ;
        RECT 7.755000 181.445000 8.075000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 181.850000 8.075000 182.170000 ;
      LAYER met4 ;
        RECT 7.755000 181.850000 8.075000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 182.255000 8.075000 182.575000 ;
      LAYER met4 ;
        RECT 7.755000 182.255000 8.075000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 182.660000 8.075000 182.980000 ;
      LAYER met4 ;
        RECT 7.755000 182.660000 8.075000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 183.065000 8.075000 183.385000 ;
      LAYER met4 ;
        RECT 7.755000 183.065000 8.075000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 183.470000 8.075000 183.790000 ;
      LAYER met4 ;
        RECT 7.755000 183.470000 8.075000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 183.875000 8.075000 184.195000 ;
      LAYER met4 ;
        RECT 7.755000 183.875000 8.075000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 184.280000 8.075000 184.600000 ;
      LAYER met4 ;
        RECT 7.755000 184.280000 8.075000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 184.685000 8.075000 185.005000 ;
      LAYER met4 ;
        RECT 7.755000 184.685000 8.075000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 185.090000 8.075000 185.410000 ;
      LAYER met4 ;
        RECT 7.755000 185.090000 8.075000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 185.495000 8.075000 185.815000 ;
      LAYER met4 ;
        RECT 7.755000 185.495000 8.075000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 185.900000 8.075000 186.220000 ;
      LAYER met4 ;
        RECT 7.755000 185.900000 8.075000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 186.305000 8.075000 186.625000 ;
      LAYER met4 ;
        RECT 7.755000 186.305000 8.075000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 186.710000 8.075000 187.030000 ;
      LAYER met4 ;
        RECT 7.755000 186.710000 8.075000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 187.115000 8.075000 187.435000 ;
      LAYER met4 ;
        RECT 7.755000 187.115000 8.075000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 187.520000 8.075000 187.840000 ;
      LAYER met4 ;
        RECT 7.755000 187.520000 8.075000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 187.925000 8.075000 188.245000 ;
      LAYER met4 ;
        RECT 7.755000 187.925000 8.075000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 188.330000 8.075000 188.650000 ;
      LAYER met4 ;
        RECT 7.755000 188.330000 8.075000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 188.735000 8.075000 189.055000 ;
      LAYER met4 ;
        RECT 7.755000 188.735000 8.075000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 189.140000 8.075000 189.460000 ;
      LAYER met4 ;
        RECT 7.755000 189.140000 8.075000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 189.545000 8.075000 189.865000 ;
      LAYER met4 ;
        RECT 7.755000 189.545000 8.075000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 189.950000 8.075000 190.270000 ;
      LAYER met4 ;
        RECT 7.755000 189.950000 8.075000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 190.355000 8.075000 190.675000 ;
      LAYER met4 ;
        RECT 7.755000 190.355000 8.075000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 190.760000 8.075000 191.080000 ;
      LAYER met4 ;
        RECT 7.755000 190.760000 8.075000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 191.165000 8.075000 191.485000 ;
      LAYER met4 ;
        RECT 7.755000 191.165000 8.075000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 191.570000 8.075000 191.890000 ;
      LAYER met4 ;
        RECT 7.755000 191.570000 8.075000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 191.975000 8.075000 192.295000 ;
      LAYER met4 ;
        RECT 7.755000 191.975000 8.075000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 192.380000 8.075000 192.700000 ;
      LAYER met4 ;
        RECT 7.755000 192.380000 8.075000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 192.785000 8.075000 193.105000 ;
      LAYER met4 ;
        RECT 7.755000 192.785000 8.075000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 193.190000 8.075000 193.510000 ;
      LAYER met4 ;
        RECT 7.755000 193.190000 8.075000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 193.595000 8.075000 193.915000 ;
      LAYER met4 ;
        RECT 7.755000 193.595000 8.075000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 194.000000 8.075000 194.320000 ;
      LAYER met4 ;
        RECT 7.755000 194.000000 8.075000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 194.405000 8.075000 194.725000 ;
      LAYER met4 ;
        RECT 7.755000 194.405000 8.075000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 194.810000 8.075000 195.130000 ;
      LAYER met4 ;
        RECT 7.755000 194.810000 8.075000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 195.215000 8.075000 195.535000 ;
      LAYER met4 ;
        RECT 7.755000 195.215000 8.075000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 195.620000 8.075000 195.940000 ;
      LAYER met4 ;
        RECT 7.755000 195.620000 8.075000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 196.025000 8.075000 196.345000 ;
      LAYER met4 ;
        RECT 7.755000 196.025000 8.075000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 196.430000 8.075000 196.750000 ;
      LAYER met4 ;
        RECT 7.755000 196.430000 8.075000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 196.835000 8.075000 197.155000 ;
      LAYER met4 ;
        RECT 7.755000 196.835000 8.075000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 197.240000 8.075000 197.560000 ;
      LAYER met4 ;
        RECT 7.755000 197.240000 8.075000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755000 197.645000 8.075000 197.965000 ;
      LAYER met4 ;
        RECT 7.755000 197.645000 8.075000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.815000 173.900000 8.015000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.815000 174.300000 8.015000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.815000 174.700000 8.015000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.815000 175.100000 8.015000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.815000 175.500000 8.015000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.815000 175.900000 8.015000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.815000 176.300000 8.015000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.815000 176.700000 8.015000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.815000 177.100000 8.015000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.815000 177.500000 8.015000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.815000 177.900000 8.015000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.815000 178.300000 8.015000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.815000 178.700000 8.015000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.815000 179.100000 8.015000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.815000 179.500000 8.015000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.815000 179.900000 8.015000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.815000 180.300000 8.015000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.815000 180.700000 8.015000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.815000 181.100000 8.015000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 23.850000 8.170000 24.170000 ;
      LAYER met4 ;
        RECT 7.850000 23.850000 8.170000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 24.280000 8.170000 24.600000 ;
      LAYER met4 ;
        RECT 7.850000 24.280000 8.170000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 24.710000 8.170000 25.030000 ;
      LAYER met4 ;
        RECT 7.850000 24.710000 8.170000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 25.140000 8.170000 25.460000 ;
      LAYER met4 ;
        RECT 7.850000 25.140000 8.170000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 25.570000 8.170000 25.890000 ;
      LAYER met4 ;
        RECT 7.850000 25.570000 8.170000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 26.000000 8.170000 26.320000 ;
      LAYER met4 ;
        RECT 7.850000 26.000000 8.170000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 26.430000 8.170000 26.750000 ;
      LAYER met4 ;
        RECT 7.850000 26.430000 8.170000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 26.860000 8.170000 27.180000 ;
      LAYER met4 ;
        RECT 7.850000 26.860000 8.170000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 27.290000 8.170000 27.610000 ;
      LAYER met4 ;
        RECT 7.850000 27.290000 8.170000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 27.720000 8.170000 28.040000 ;
      LAYER met4 ;
        RECT 7.850000 27.720000 8.170000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 28.150000 8.170000 28.470000 ;
      LAYER met4 ;
        RECT 7.850000 28.150000 8.170000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 173.840000 70.600000 174.160000 ;
      LAYER met4 ;
        RECT 70.280000 173.840000 70.600000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 174.240000 70.600000 174.560000 ;
      LAYER met4 ;
        RECT 70.280000 174.240000 70.600000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 174.640000 70.600000 174.960000 ;
      LAYER met4 ;
        RECT 70.280000 174.640000 70.600000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 175.040000 70.600000 175.360000 ;
      LAYER met4 ;
        RECT 70.280000 175.040000 70.600000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 175.440000 70.600000 175.760000 ;
      LAYER met4 ;
        RECT 70.280000 175.440000 70.600000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 175.840000 70.600000 176.160000 ;
      LAYER met4 ;
        RECT 70.280000 175.840000 70.600000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 176.240000 70.600000 176.560000 ;
      LAYER met4 ;
        RECT 70.280000 176.240000 70.600000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 176.640000 70.600000 176.960000 ;
      LAYER met4 ;
        RECT 70.280000 176.640000 70.600000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 177.040000 70.600000 177.360000 ;
      LAYER met4 ;
        RECT 70.280000 177.040000 70.600000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 177.440000 70.600000 177.760000 ;
      LAYER met4 ;
        RECT 70.280000 177.440000 70.600000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 177.840000 70.600000 178.160000 ;
      LAYER met4 ;
        RECT 70.280000 177.840000 70.600000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 178.240000 70.600000 178.560000 ;
      LAYER met4 ;
        RECT 70.280000 178.240000 70.600000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 178.640000 70.600000 178.960000 ;
      LAYER met4 ;
        RECT 70.280000 178.640000 70.600000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 179.040000 70.600000 179.360000 ;
      LAYER met4 ;
        RECT 70.280000 179.040000 70.600000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 179.440000 70.600000 179.760000 ;
      LAYER met4 ;
        RECT 70.280000 179.440000 70.600000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 179.840000 70.600000 180.160000 ;
      LAYER met4 ;
        RECT 70.280000 179.840000 70.600000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 180.240000 70.600000 180.560000 ;
      LAYER met4 ;
        RECT 70.280000 180.240000 70.600000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 180.640000 70.600000 180.960000 ;
      LAYER met4 ;
        RECT 70.280000 180.640000 70.600000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 181.040000 70.600000 181.360000 ;
      LAYER met4 ;
        RECT 70.280000 181.040000 70.600000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 181.445000 70.600000 181.765000 ;
      LAYER met4 ;
        RECT 70.280000 181.445000 70.600000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 181.850000 70.600000 182.170000 ;
      LAYER met4 ;
        RECT 70.280000 181.850000 70.600000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 182.255000 70.600000 182.575000 ;
      LAYER met4 ;
        RECT 70.280000 182.255000 70.600000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 182.660000 70.600000 182.980000 ;
      LAYER met4 ;
        RECT 70.280000 182.660000 70.600000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 183.065000 70.600000 183.385000 ;
      LAYER met4 ;
        RECT 70.280000 183.065000 70.600000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 183.470000 70.600000 183.790000 ;
      LAYER met4 ;
        RECT 70.280000 183.470000 70.600000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 183.875000 70.600000 184.195000 ;
      LAYER met4 ;
        RECT 70.280000 183.875000 70.600000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 184.280000 70.600000 184.600000 ;
      LAYER met4 ;
        RECT 70.280000 184.280000 70.600000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 184.685000 70.600000 185.005000 ;
      LAYER met4 ;
        RECT 70.280000 184.685000 70.600000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 185.090000 70.600000 185.410000 ;
      LAYER met4 ;
        RECT 70.280000 185.090000 70.600000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 185.495000 70.600000 185.815000 ;
      LAYER met4 ;
        RECT 70.280000 185.495000 70.600000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 185.900000 70.600000 186.220000 ;
      LAYER met4 ;
        RECT 70.280000 185.900000 70.600000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 186.305000 70.600000 186.625000 ;
      LAYER met4 ;
        RECT 70.280000 186.305000 70.600000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 186.710000 70.600000 187.030000 ;
      LAYER met4 ;
        RECT 70.280000 186.710000 70.600000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 187.115000 70.600000 187.435000 ;
      LAYER met4 ;
        RECT 70.280000 187.115000 70.600000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 187.520000 70.600000 187.840000 ;
      LAYER met4 ;
        RECT 70.280000 187.520000 70.600000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 187.925000 70.600000 188.245000 ;
      LAYER met4 ;
        RECT 70.280000 187.925000 70.600000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 188.330000 70.600000 188.650000 ;
      LAYER met4 ;
        RECT 70.280000 188.330000 70.600000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 188.735000 70.600000 189.055000 ;
      LAYER met4 ;
        RECT 70.280000 188.735000 70.600000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 189.140000 70.600000 189.460000 ;
      LAYER met4 ;
        RECT 70.280000 189.140000 70.600000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 189.545000 70.600000 189.865000 ;
      LAYER met4 ;
        RECT 70.280000 189.545000 70.600000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 189.950000 70.600000 190.270000 ;
      LAYER met4 ;
        RECT 70.280000 189.950000 70.600000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 190.355000 70.600000 190.675000 ;
      LAYER met4 ;
        RECT 70.280000 190.355000 70.600000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 190.760000 70.600000 191.080000 ;
      LAYER met4 ;
        RECT 70.280000 190.760000 70.600000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 191.165000 70.600000 191.485000 ;
      LAYER met4 ;
        RECT 70.280000 191.165000 70.600000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 191.570000 70.600000 191.890000 ;
      LAYER met4 ;
        RECT 70.280000 191.570000 70.600000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 191.975000 70.600000 192.295000 ;
      LAYER met4 ;
        RECT 70.280000 191.975000 70.600000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 192.380000 70.600000 192.700000 ;
      LAYER met4 ;
        RECT 70.280000 192.380000 70.600000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 192.785000 70.600000 193.105000 ;
      LAYER met4 ;
        RECT 70.280000 192.785000 70.600000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 193.190000 70.600000 193.510000 ;
      LAYER met4 ;
        RECT 70.280000 193.190000 70.600000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 193.595000 70.600000 193.915000 ;
      LAYER met4 ;
        RECT 70.280000 193.595000 70.600000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 194.000000 70.600000 194.320000 ;
      LAYER met4 ;
        RECT 70.280000 194.000000 70.600000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 194.405000 70.600000 194.725000 ;
      LAYER met4 ;
        RECT 70.280000 194.405000 70.600000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 194.810000 70.600000 195.130000 ;
      LAYER met4 ;
        RECT 70.280000 194.810000 70.600000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 195.215000 70.600000 195.535000 ;
      LAYER met4 ;
        RECT 70.280000 195.215000 70.600000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 195.620000 70.600000 195.940000 ;
      LAYER met4 ;
        RECT 70.280000 195.620000 70.600000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 196.025000 70.600000 196.345000 ;
      LAYER met4 ;
        RECT 70.280000 196.025000 70.600000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 196.430000 70.600000 196.750000 ;
      LAYER met4 ;
        RECT 70.280000 196.430000 70.600000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 196.835000 70.600000 197.155000 ;
      LAYER met4 ;
        RECT 70.280000 196.835000 70.600000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 197.240000 70.600000 197.560000 ;
      LAYER met4 ;
        RECT 70.280000 197.240000 70.600000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.280000 197.645000 70.600000 197.965000 ;
      LAYER met4 ;
        RECT 70.280000 197.645000 70.600000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 23.850000 70.615000 24.170000 ;
      LAYER met4 ;
        RECT 70.295000 23.850000 70.615000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 24.280000 70.615000 24.600000 ;
      LAYER met4 ;
        RECT 70.295000 24.280000 70.615000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 24.710000 70.615000 25.030000 ;
      LAYER met4 ;
        RECT 70.295000 24.710000 70.615000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 25.140000 70.615000 25.460000 ;
      LAYER met4 ;
        RECT 70.295000 25.140000 70.615000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 25.570000 70.615000 25.890000 ;
      LAYER met4 ;
        RECT 70.295000 25.570000 70.615000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 26.000000 70.615000 26.320000 ;
      LAYER met4 ;
        RECT 70.295000 26.000000 70.615000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 26.430000 70.615000 26.750000 ;
      LAYER met4 ;
        RECT 70.295000 26.430000 70.615000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 26.860000 70.615000 27.180000 ;
      LAYER met4 ;
        RECT 70.295000 26.860000 70.615000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 27.290000 70.615000 27.610000 ;
      LAYER met4 ;
        RECT 70.295000 27.290000 70.615000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 27.720000 70.615000 28.040000 ;
      LAYER met4 ;
        RECT 70.295000 27.720000 70.615000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 28.150000 70.615000 28.470000 ;
      LAYER met4 ;
        RECT 70.295000 28.150000 70.615000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 173.840000 71.010000 174.160000 ;
      LAYER met4 ;
        RECT 70.690000 173.840000 71.010000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 174.240000 71.010000 174.560000 ;
      LAYER met4 ;
        RECT 70.690000 174.240000 71.010000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 174.640000 71.010000 174.960000 ;
      LAYER met4 ;
        RECT 70.690000 174.640000 71.010000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 175.040000 71.010000 175.360000 ;
      LAYER met4 ;
        RECT 70.690000 175.040000 71.010000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 175.440000 71.010000 175.760000 ;
      LAYER met4 ;
        RECT 70.690000 175.440000 71.010000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 175.840000 71.010000 176.160000 ;
      LAYER met4 ;
        RECT 70.690000 175.840000 71.010000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 176.240000 71.010000 176.560000 ;
      LAYER met4 ;
        RECT 70.690000 176.240000 71.010000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 176.640000 71.010000 176.960000 ;
      LAYER met4 ;
        RECT 70.690000 176.640000 71.010000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 177.040000 71.010000 177.360000 ;
      LAYER met4 ;
        RECT 70.690000 177.040000 71.010000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 177.440000 71.010000 177.760000 ;
      LAYER met4 ;
        RECT 70.690000 177.440000 71.010000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 177.840000 71.010000 178.160000 ;
      LAYER met4 ;
        RECT 70.690000 177.840000 71.010000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 178.240000 71.010000 178.560000 ;
      LAYER met4 ;
        RECT 70.690000 178.240000 71.010000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 178.640000 71.010000 178.960000 ;
      LAYER met4 ;
        RECT 70.690000 178.640000 71.010000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 179.040000 71.010000 179.360000 ;
      LAYER met4 ;
        RECT 70.690000 179.040000 71.010000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 179.440000 71.010000 179.760000 ;
      LAYER met4 ;
        RECT 70.690000 179.440000 71.010000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 179.840000 71.010000 180.160000 ;
      LAYER met4 ;
        RECT 70.690000 179.840000 71.010000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 180.240000 71.010000 180.560000 ;
      LAYER met4 ;
        RECT 70.690000 180.240000 71.010000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 180.640000 71.010000 180.960000 ;
      LAYER met4 ;
        RECT 70.690000 180.640000 71.010000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 181.040000 71.010000 181.360000 ;
      LAYER met4 ;
        RECT 70.690000 181.040000 71.010000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 181.445000 71.010000 181.765000 ;
      LAYER met4 ;
        RECT 70.690000 181.445000 71.010000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 181.850000 71.010000 182.170000 ;
      LAYER met4 ;
        RECT 70.690000 181.850000 71.010000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 182.255000 71.010000 182.575000 ;
      LAYER met4 ;
        RECT 70.690000 182.255000 71.010000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 182.660000 71.010000 182.980000 ;
      LAYER met4 ;
        RECT 70.690000 182.660000 71.010000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 183.065000 71.010000 183.385000 ;
      LAYER met4 ;
        RECT 70.690000 183.065000 71.010000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 183.470000 71.010000 183.790000 ;
      LAYER met4 ;
        RECT 70.690000 183.470000 71.010000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 183.875000 71.010000 184.195000 ;
      LAYER met4 ;
        RECT 70.690000 183.875000 71.010000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 184.280000 71.010000 184.600000 ;
      LAYER met4 ;
        RECT 70.690000 184.280000 71.010000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 184.685000 71.010000 185.005000 ;
      LAYER met4 ;
        RECT 70.690000 184.685000 71.010000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 185.090000 71.010000 185.410000 ;
      LAYER met4 ;
        RECT 70.690000 185.090000 71.010000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 185.495000 71.010000 185.815000 ;
      LAYER met4 ;
        RECT 70.690000 185.495000 71.010000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 185.900000 71.010000 186.220000 ;
      LAYER met4 ;
        RECT 70.690000 185.900000 71.010000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 186.305000 71.010000 186.625000 ;
      LAYER met4 ;
        RECT 70.690000 186.305000 71.010000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 186.710000 71.010000 187.030000 ;
      LAYER met4 ;
        RECT 70.690000 186.710000 71.010000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 187.115000 71.010000 187.435000 ;
      LAYER met4 ;
        RECT 70.690000 187.115000 71.010000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 187.520000 71.010000 187.840000 ;
      LAYER met4 ;
        RECT 70.690000 187.520000 71.010000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 187.925000 71.010000 188.245000 ;
      LAYER met4 ;
        RECT 70.690000 187.925000 71.010000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 188.330000 71.010000 188.650000 ;
      LAYER met4 ;
        RECT 70.690000 188.330000 71.010000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 188.735000 71.010000 189.055000 ;
      LAYER met4 ;
        RECT 70.690000 188.735000 71.010000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 189.140000 71.010000 189.460000 ;
      LAYER met4 ;
        RECT 70.690000 189.140000 71.010000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 189.545000 71.010000 189.865000 ;
      LAYER met4 ;
        RECT 70.690000 189.545000 71.010000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 189.950000 71.010000 190.270000 ;
      LAYER met4 ;
        RECT 70.690000 189.950000 71.010000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 190.355000 71.010000 190.675000 ;
      LAYER met4 ;
        RECT 70.690000 190.355000 71.010000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 190.760000 71.010000 191.080000 ;
      LAYER met4 ;
        RECT 70.690000 190.760000 71.010000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 191.165000 71.010000 191.485000 ;
      LAYER met4 ;
        RECT 70.690000 191.165000 71.010000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 191.570000 71.010000 191.890000 ;
      LAYER met4 ;
        RECT 70.690000 191.570000 71.010000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 191.975000 71.010000 192.295000 ;
      LAYER met4 ;
        RECT 70.690000 191.975000 71.010000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 192.380000 71.010000 192.700000 ;
      LAYER met4 ;
        RECT 70.690000 192.380000 71.010000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 192.785000 71.010000 193.105000 ;
      LAYER met4 ;
        RECT 70.690000 192.785000 71.010000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 193.190000 71.010000 193.510000 ;
      LAYER met4 ;
        RECT 70.690000 193.190000 71.010000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 193.595000 71.010000 193.915000 ;
      LAYER met4 ;
        RECT 70.690000 193.595000 71.010000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 194.000000 71.010000 194.320000 ;
      LAYER met4 ;
        RECT 70.690000 194.000000 71.010000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 194.405000 71.010000 194.725000 ;
      LAYER met4 ;
        RECT 70.690000 194.405000 71.010000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 194.810000 71.010000 195.130000 ;
      LAYER met4 ;
        RECT 70.690000 194.810000 71.010000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 195.215000 71.010000 195.535000 ;
      LAYER met4 ;
        RECT 70.690000 195.215000 71.010000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 195.620000 71.010000 195.940000 ;
      LAYER met4 ;
        RECT 70.690000 195.620000 71.010000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 196.025000 71.010000 196.345000 ;
      LAYER met4 ;
        RECT 70.690000 196.025000 71.010000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 196.430000 71.010000 196.750000 ;
      LAYER met4 ;
        RECT 70.690000 196.430000 71.010000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 196.835000 71.010000 197.155000 ;
      LAYER met4 ;
        RECT 70.690000 196.835000 71.010000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 197.240000 71.010000 197.560000 ;
      LAYER met4 ;
        RECT 70.690000 197.240000 71.010000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690000 197.645000 71.010000 197.965000 ;
      LAYER met4 ;
        RECT 70.690000 197.645000 71.010000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 23.850000 71.020000 24.170000 ;
      LAYER met4 ;
        RECT 70.700000 23.850000 71.020000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 24.280000 71.020000 24.600000 ;
      LAYER met4 ;
        RECT 70.700000 24.280000 71.020000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 24.710000 71.020000 25.030000 ;
      LAYER met4 ;
        RECT 70.700000 24.710000 71.020000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 25.140000 71.020000 25.460000 ;
      LAYER met4 ;
        RECT 70.700000 25.140000 71.020000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 25.570000 71.020000 25.890000 ;
      LAYER met4 ;
        RECT 70.700000 25.570000 71.020000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 26.000000 71.020000 26.320000 ;
      LAYER met4 ;
        RECT 70.700000 26.000000 71.020000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 26.430000 71.020000 26.750000 ;
      LAYER met4 ;
        RECT 70.700000 26.430000 71.020000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 26.860000 71.020000 27.180000 ;
      LAYER met4 ;
        RECT 70.700000 26.860000 71.020000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 27.290000 71.020000 27.610000 ;
      LAYER met4 ;
        RECT 70.700000 27.290000 71.020000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 27.720000 71.020000 28.040000 ;
      LAYER met4 ;
        RECT 70.700000 27.720000 71.020000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 28.150000 71.020000 28.470000 ;
      LAYER met4 ;
        RECT 70.700000 28.150000 71.020000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 173.840000 71.420000 174.160000 ;
      LAYER met4 ;
        RECT 71.100000 173.840000 71.420000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 174.240000 71.420000 174.560000 ;
      LAYER met4 ;
        RECT 71.100000 174.240000 71.420000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 174.640000 71.420000 174.960000 ;
      LAYER met4 ;
        RECT 71.100000 174.640000 71.420000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 175.040000 71.420000 175.360000 ;
      LAYER met4 ;
        RECT 71.100000 175.040000 71.420000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 175.440000 71.420000 175.760000 ;
      LAYER met4 ;
        RECT 71.100000 175.440000 71.420000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 175.840000 71.420000 176.160000 ;
      LAYER met4 ;
        RECT 71.100000 175.840000 71.420000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 176.240000 71.420000 176.560000 ;
      LAYER met4 ;
        RECT 71.100000 176.240000 71.420000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 176.640000 71.420000 176.960000 ;
      LAYER met4 ;
        RECT 71.100000 176.640000 71.420000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 177.040000 71.420000 177.360000 ;
      LAYER met4 ;
        RECT 71.100000 177.040000 71.420000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 177.440000 71.420000 177.760000 ;
      LAYER met4 ;
        RECT 71.100000 177.440000 71.420000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 177.840000 71.420000 178.160000 ;
      LAYER met4 ;
        RECT 71.100000 177.840000 71.420000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 178.240000 71.420000 178.560000 ;
      LAYER met4 ;
        RECT 71.100000 178.240000 71.420000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 178.640000 71.420000 178.960000 ;
      LAYER met4 ;
        RECT 71.100000 178.640000 71.420000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 179.040000 71.420000 179.360000 ;
      LAYER met4 ;
        RECT 71.100000 179.040000 71.420000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 179.440000 71.420000 179.760000 ;
      LAYER met4 ;
        RECT 71.100000 179.440000 71.420000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 179.840000 71.420000 180.160000 ;
      LAYER met4 ;
        RECT 71.100000 179.840000 71.420000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 180.240000 71.420000 180.560000 ;
      LAYER met4 ;
        RECT 71.100000 180.240000 71.420000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 180.640000 71.420000 180.960000 ;
      LAYER met4 ;
        RECT 71.100000 180.640000 71.420000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 181.040000 71.420000 181.360000 ;
      LAYER met4 ;
        RECT 71.100000 181.040000 71.420000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 181.445000 71.420000 181.765000 ;
      LAYER met4 ;
        RECT 71.100000 181.445000 71.420000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 181.850000 71.420000 182.170000 ;
      LAYER met4 ;
        RECT 71.100000 181.850000 71.420000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 182.255000 71.420000 182.575000 ;
      LAYER met4 ;
        RECT 71.100000 182.255000 71.420000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 182.660000 71.420000 182.980000 ;
      LAYER met4 ;
        RECT 71.100000 182.660000 71.420000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 183.065000 71.420000 183.385000 ;
      LAYER met4 ;
        RECT 71.100000 183.065000 71.420000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 183.470000 71.420000 183.790000 ;
      LAYER met4 ;
        RECT 71.100000 183.470000 71.420000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 183.875000 71.420000 184.195000 ;
      LAYER met4 ;
        RECT 71.100000 183.875000 71.420000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 184.280000 71.420000 184.600000 ;
      LAYER met4 ;
        RECT 71.100000 184.280000 71.420000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 184.685000 71.420000 185.005000 ;
      LAYER met4 ;
        RECT 71.100000 184.685000 71.420000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 185.090000 71.420000 185.410000 ;
      LAYER met4 ;
        RECT 71.100000 185.090000 71.420000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 185.495000 71.420000 185.815000 ;
      LAYER met4 ;
        RECT 71.100000 185.495000 71.420000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 185.900000 71.420000 186.220000 ;
      LAYER met4 ;
        RECT 71.100000 185.900000 71.420000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 186.305000 71.420000 186.625000 ;
      LAYER met4 ;
        RECT 71.100000 186.305000 71.420000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 186.710000 71.420000 187.030000 ;
      LAYER met4 ;
        RECT 71.100000 186.710000 71.420000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 187.115000 71.420000 187.435000 ;
      LAYER met4 ;
        RECT 71.100000 187.115000 71.420000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 187.520000 71.420000 187.840000 ;
      LAYER met4 ;
        RECT 71.100000 187.520000 71.420000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 187.925000 71.420000 188.245000 ;
      LAYER met4 ;
        RECT 71.100000 187.925000 71.420000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 188.330000 71.420000 188.650000 ;
      LAYER met4 ;
        RECT 71.100000 188.330000 71.420000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 188.735000 71.420000 189.055000 ;
      LAYER met4 ;
        RECT 71.100000 188.735000 71.420000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 189.140000 71.420000 189.460000 ;
      LAYER met4 ;
        RECT 71.100000 189.140000 71.420000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 189.545000 71.420000 189.865000 ;
      LAYER met4 ;
        RECT 71.100000 189.545000 71.420000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 189.950000 71.420000 190.270000 ;
      LAYER met4 ;
        RECT 71.100000 189.950000 71.420000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 190.355000 71.420000 190.675000 ;
      LAYER met4 ;
        RECT 71.100000 190.355000 71.420000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 190.760000 71.420000 191.080000 ;
      LAYER met4 ;
        RECT 71.100000 190.760000 71.420000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 191.165000 71.420000 191.485000 ;
      LAYER met4 ;
        RECT 71.100000 191.165000 71.420000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 191.570000 71.420000 191.890000 ;
      LAYER met4 ;
        RECT 71.100000 191.570000 71.420000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 191.975000 71.420000 192.295000 ;
      LAYER met4 ;
        RECT 71.100000 191.975000 71.420000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 192.380000 71.420000 192.700000 ;
      LAYER met4 ;
        RECT 71.100000 192.380000 71.420000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 192.785000 71.420000 193.105000 ;
      LAYER met4 ;
        RECT 71.100000 192.785000 71.420000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 193.190000 71.420000 193.510000 ;
      LAYER met4 ;
        RECT 71.100000 193.190000 71.420000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 193.595000 71.420000 193.915000 ;
      LAYER met4 ;
        RECT 71.100000 193.595000 71.420000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 194.000000 71.420000 194.320000 ;
      LAYER met4 ;
        RECT 71.100000 194.000000 71.420000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 194.405000 71.420000 194.725000 ;
      LAYER met4 ;
        RECT 71.100000 194.405000 71.420000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 194.810000 71.420000 195.130000 ;
      LAYER met4 ;
        RECT 71.100000 194.810000 71.420000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 195.215000 71.420000 195.535000 ;
      LAYER met4 ;
        RECT 71.100000 195.215000 71.420000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 195.620000 71.420000 195.940000 ;
      LAYER met4 ;
        RECT 71.100000 195.620000 71.420000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 196.025000 71.420000 196.345000 ;
      LAYER met4 ;
        RECT 71.100000 196.025000 71.420000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 196.430000 71.420000 196.750000 ;
      LAYER met4 ;
        RECT 71.100000 196.430000 71.420000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 196.835000 71.420000 197.155000 ;
      LAYER met4 ;
        RECT 71.100000 196.835000 71.420000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 197.240000 71.420000 197.560000 ;
      LAYER met4 ;
        RECT 71.100000 197.240000 71.420000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.100000 197.645000 71.420000 197.965000 ;
      LAYER met4 ;
        RECT 71.100000 197.645000 71.420000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 23.850000 71.425000 24.170000 ;
      LAYER met4 ;
        RECT 71.105000 23.850000 71.425000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 24.280000 71.425000 24.600000 ;
      LAYER met4 ;
        RECT 71.105000 24.280000 71.425000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 24.710000 71.425000 25.030000 ;
      LAYER met4 ;
        RECT 71.105000 24.710000 71.425000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 25.140000 71.425000 25.460000 ;
      LAYER met4 ;
        RECT 71.105000 25.140000 71.425000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 25.570000 71.425000 25.890000 ;
      LAYER met4 ;
        RECT 71.105000 25.570000 71.425000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 26.000000 71.425000 26.320000 ;
      LAYER met4 ;
        RECT 71.105000 26.000000 71.425000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 26.430000 71.425000 26.750000 ;
      LAYER met4 ;
        RECT 71.105000 26.430000 71.425000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 26.860000 71.425000 27.180000 ;
      LAYER met4 ;
        RECT 71.105000 26.860000 71.425000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 27.290000 71.425000 27.610000 ;
      LAYER met4 ;
        RECT 71.105000 27.290000 71.425000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 27.720000 71.425000 28.040000 ;
      LAYER met4 ;
        RECT 71.105000 27.720000 71.425000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 28.150000 71.425000 28.470000 ;
      LAYER met4 ;
        RECT 71.105000 28.150000 71.425000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 173.840000 71.830000 174.160000 ;
      LAYER met4 ;
        RECT 71.510000 173.840000 71.830000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 174.240000 71.830000 174.560000 ;
      LAYER met4 ;
        RECT 71.510000 174.240000 71.830000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 174.640000 71.830000 174.960000 ;
      LAYER met4 ;
        RECT 71.510000 174.640000 71.830000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 175.040000 71.830000 175.360000 ;
      LAYER met4 ;
        RECT 71.510000 175.040000 71.830000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 175.440000 71.830000 175.760000 ;
      LAYER met4 ;
        RECT 71.510000 175.440000 71.830000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 175.840000 71.830000 176.160000 ;
      LAYER met4 ;
        RECT 71.510000 175.840000 71.830000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 176.240000 71.830000 176.560000 ;
      LAYER met4 ;
        RECT 71.510000 176.240000 71.830000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 176.640000 71.830000 176.960000 ;
      LAYER met4 ;
        RECT 71.510000 176.640000 71.830000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 177.040000 71.830000 177.360000 ;
      LAYER met4 ;
        RECT 71.510000 177.040000 71.830000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 177.440000 71.830000 177.760000 ;
      LAYER met4 ;
        RECT 71.510000 177.440000 71.830000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 177.840000 71.830000 178.160000 ;
      LAYER met4 ;
        RECT 71.510000 177.840000 71.830000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 178.240000 71.830000 178.560000 ;
      LAYER met4 ;
        RECT 71.510000 178.240000 71.830000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 178.640000 71.830000 178.960000 ;
      LAYER met4 ;
        RECT 71.510000 178.640000 71.830000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 179.040000 71.830000 179.360000 ;
      LAYER met4 ;
        RECT 71.510000 179.040000 71.830000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 179.440000 71.830000 179.760000 ;
      LAYER met4 ;
        RECT 71.510000 179.440000 71.830000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 179.840000 71.830000 180.160000 ;
      LAYER met4 ;
        RECT 71.510000 179.840000 71.830000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 180.240000 71.830000 180.560000 ;
      LAYER met4 ;
        RECT 71.510000 180.240000 71.830000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 180.640000 71.830000 180.960000 ;
      LAYER met4 ;
        RECT 71.510000 180.640000 71.830000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 181.040000 71.830000 181.360000 ;
      LAYER met4 ;
        RECT 71.510000 181.040000 71.830000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 181.445000 71.830000 181.765000 ;
      LAYER met4 ;
        RECT 71.510000 181.445000 71.830000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 181.850000 71.830000 182.170000 ;
      LAYER met4 ;
        RECT 71.510000 181.850000 71.830000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 182.255000 71.830000 182.575000 ;
      LAYER met4 ;
        RECT 71.510000 182.255000 71.830000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 182.660000 71.830000 182.980000 ;
      LAYER met4 ;
        RECT 71.510000 182.660000 71.830000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 183.065000 71.830000 183.385000 ;
      LAYER met4 ;
        RECT 71.510000 183.065000 71.830000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 183.470000 71.830000 183.790000 ;
      LAYER met4 ;
        RECT 71.510000 183.470000 71.830000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 183.875000 71.830000 184.195000 ;
      LAYER met4 ;
        RECT 71.510000 183.875000 71.830000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 184.280000 71.830000 184.600000 ;
      LAYER met4 ;
        RECT 71.510000 184.280000 71.830000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 184.685000 71.830000 185.005000 ;
      LAYER met4 ;
        RECT 71.510000 184.685000 71.830000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 185.090000 71.830000 185.410000 ;
      LAYER met4 ;
        RECT 71.510000 185.090000 71.830000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 185.495000 71.830000 185.815000 ;
      LAYER met4 ;
        RECT 71.510000 185.495000 71.830000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 185.900000 71.830000 186.220000 ;
      LAYER met4 ;
        RECT 71.510000 185.900000 71.830000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 186.305000 71.830000 186.625000 ;
      LAYER met4 ;
        RECT 71.510000 186.305000 71.830000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 186.710000 71.830000 187.030000 ;
      LAYER met4 ;
        RECT 71.510000 186.710000 71.830000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 187.115000 71.830000 187.435000 ;
      LAYER met4 ;
        RECT 71.510000 187.115000 71.830000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 187.520000 71.830000 187.840000 ;
      LAYER met4 ;
        RECT 71.510000 187.520000 71.830000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 187.925000 71.830000 188.245000 ;
      LAYER met4 ;
        RECT 71.510000 187.925000 71.830000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 188.330000 71.830000 188.650000 ;
      LAYER met4 ;
        RECT 71.510000 188.330000 71.830000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 188.735000 71.830000 189.055000 ;
      LAYER met4 ;
        RECT 71.510000 188.735000 71.830000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 189.140000 71.830000 189.460000 ;
      LAYER met4 ;
        RECT 71.510000 189.140000 71.830000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 189.545000 71.830000 189.865000 ;
      LAYER met4 ;
        RECT 71.510000 189.545000 71.830000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 189.950000 71.830000 190.270000 ;
      LAYER met4 ;
        RECT 71.510000 189.950000 71.830000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 190.355000 71.830000 190.675000 ;
      LAYER met4 ;
        RECT 71.510000 190.355000 71.830000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 190.760000 71.830000 191.080000 ;
      LAYER met4 ;
        RECT 71.510000 190.760000 71.830000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 191.165000 71.830000 191.485000 ;
      LAYER met4 ;
        RECT 71.510000 191.165000 71.830000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 191.570000 71.830000 191.890000 ;
      LAYER met4 ;
        RECT 71.510000 191.570000 71.830000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 191.975000 71.830000 192.295000 ;
      LAYER met4 ;
        RECT 71.510000 191.975000 71.830000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 192.380000 71.830000 192.700000 ;
      LAYER met4 ;
        RECT 71.510000 192.380000 71.830000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 192.785000 71.830000 193.105000 ;
      LAYER met4 ;
        RECT 71.510000 192.785000 71.830000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 193.190000 71.830000 193.510000 ;
      LAYER met4 ;
        RECT 71.510000 193.190000 71.830000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 193.595000 71.830000 193.915000 ;
      LAYER met4 ;
        RECT 71.510000 193.595000 71.830000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 194.000000 71.830000 194.320000 ;
      LAYER met4 ;
        RECT 71.510000 194.000000 71.830000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 194.405000 71.830000 194.725000 ;
      LAYER met4 ;
        RECT 71.510000 194.405000 71.830000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 194.810000 71.830000 195.130000 ;
      LAYER met4 ;
        RECT 71.510000 194.810000 71.830000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 195.215000 71.830000 195.535000 ;
      LAYER met4 ;
        RECT 71.510000 195.215000 71.830000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 195.620000 71.830000 195.940000 ;
      LAYER met4 ;
        RECT 71.510000 195.620000 71.830000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 196.025000 71.830000 196.345000 ;
      LAYER met4 ;
        RECT 71.510000 196.025000 71.830000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 196.430000 71.830000 196.750000 ;
      LAYER met4 ;
        RECT 71.510000 196.430000 71.830000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 196.835000 71.830000 197.155000 ;
      LAYER met4 ;
        RECT 71.510000 196.835000 71.830000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 197.240000 71.830000 197.560000 ;
      LAYER met4 ;
        RECT 71.510000 197.240000 71.830000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 197.645000 71.830000 197.965000 ;
      LAYER met4 ;
        RECT 71.510000 197.645000 71.830000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 23.850000 71.830000 24.170000 ;
      LAYER met4 ;
        RECT 71.510000 23.850000 71.830000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 24.280000 71.830000 24.600000 ;
      LAYER met4 ;
        RECT 71.510000 24.280000 71.830000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 24.710000 71.830000 25.030000 ;
      LAYER met4 ;
        RECT 71.510000 24.710000 71.830000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 25.140000 71.830000 25.460000 ;
      LAYER met4 ;
        RECT 71.510000 25.140000 71.830000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 25.570000 71.830000 25.890000 ;
      LAYER met4 ;
        RECT 71.510000 25.570000 71.830000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 26.000000 71.830000 26.320000 ;
      LAYER met4 ;
        RECT 71.510000 26.000000 71.830000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 26.430000 71.830000 26.750000 ;
      LAYER met4 ;
        RECT 71.510000 26.430000 71.830000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 26.860000 71.830000 27.180000 ;
      LAYER met4 ;
        RECT 71.510000 26.860000 71.830000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 27.290000 71.830000 27.610000 ;
      LAYER met4 ;
        RECT 71.510000 27.290000 71.830000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 27.720000 71.830000 28.040000 ;
      LAYER met4 ;
        RECT 71.510000 27.720000 71.830000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 28.150000 71.830000 28.470000 ;
      LAYER met4 ;
        RECT 71.510000 28.150000 71.830000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 23.850000 72.235000 24.170000 ;
      LAYER met4 ;
        RECT 71.915000 23.850000 72.235000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 24.280000 72.235000 24.600000 ;
      LAYER met4 ;
        RECT 71.915000 24.280000 72.235000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 24.710000 72.235000 25.030000 ;
      LAYER met4 ;
        RECT 71.915000 24.710000 72.235000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 25.140000 72.235000 25.460000 ;
      LAYER met4 ;
        RECT 71.915000 25.140000 72.235000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 25.570000 72.235000 25.890000 ;
      LAYER met4 ;
        RECT 71.915000 25.570000 72.235000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 26.000000 72.235000 26.320000 ;
      LAYER met4 ;
        RECT 71.915000 26.000000 72.235000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 26.430000 72.235000 26.750000 ;
      LAYER met4 ;
        RECT 71.915000 26.430000 72.235000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 26.860000 72.235000 27.180000 ;
      LAYER met4 ;
        RECT 71.915000 26.860000 72.235000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 27.290000 72.235000 27.610000 ;
      LAYER met4 ;
        RECT 71.915000 27.290000 72.235000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 27.720000 72.235000 28.040000 ;
      LAYER met4 ;
        RECT 71.915000 27.720000 72.235000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 28.150000 72.235000 28.470000 ;
      LAYER met4 ;
        RECT 71.915000 28.150000 72.235000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 173.840000 72.240000 174.160000 ;
      LAYER met4 ;
        RECT 71.920000 173.840000 72.240000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 174.240000 72.240000 174.560000 ;
      LAYER met4 ;
        RECT 71.920000 174.240000 72.240000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 174.640000 72.240000 174.960000 ;
      LAYER met4 ;
        RECT 71.920000 174.640000 72.240000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 175.040000 72.240000 175.360000 ;
      LAYER met4 ;
        RECT 71.920000 175.040000 72.240000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 175.440000 72.240000 175.760000 ;
      LAYER met4 ;
        RECT 71.920000 175.440000 72.240000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 175.840000 72.240000 176.160000 ;
      LAYER met4 ;
        RECT 71.920000 175.840000 72.240000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 176.240000 72.240000 176.560000 ;
      LAYER met4 ;
        RECT 71.920000 176.240000 72.240000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 176.640000 72.240000 176.960000 ;
      LAYER met4 ;
        RECT 71.920000 176.640000 72.240000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 177.040000 72.240000 177.360000 ;
      LAYER met4 ;
        RECT 71.920000 177.040000 72.240000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 177.440000 72.240000 177.760000 ;
      LAYER met4 ;
        RECT 71.920000 177.440000 72.240000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 177.840000 72.240000 178.160000 ;
      LAYER met4 ;
        RECT 71.920000 177.840000 72.240000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 178.240000 72.240000 178.560000 ;
      LAYER met4 ;
        RECT 71.920000 178.240000 72.240000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 178.640000 72.240000 178.960000 ;
      LAYER met4 ;
        RECT 71.920000 178.640000 72.240000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 179.040000 72.240000 179.360000 ;
      LAYER met4 ;
        RECT 71.920000 179.040000 72.240000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 179.440000 72.240000 179.760000 ;
      LAYER met4 ;
        RECT 71.920000 179.440000 72.240000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 179.840000 72.240000 180.160000 ;
      LAYER met4 ;
        RECT 71.920000 179.840000 72.240000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 180.240000 72.240000 180.560000 ;
      LAYER met4 ;
        RECT 71.920000 180.240000 72.240000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 180.640000 72.240000 180.960000 ;
      LAYER met4 ;
        RECT 71.920000 180.640000 72.240000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 181.040000 72.240000 181.360000 ;
      LAYER met4 ;
        RECT 71.920000 181.040000 72.240000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 181.445000 72.240000 181.765000 ;
      LAYER met4 ;
        RECT 71.920000 181.445000 72.240000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 181.850000 72.240000 182.170000 ;
      LAYER met4 ;
        RECT 71.920000 181.850000 72.240000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 182.255000 72.240000 182.575000 ;
      LAYER met4 ;
        RECT 71.920000 182.255000 72.240000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 182.660000 72.240000 182.980000 ;
      LAYER met4 ;
        RECT 71.920000 182.660000 72.240000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 183.065000 72.240000 183.385000 ;
      LAYER met4 ;
        RECT 71.920000 183.065000 72.240000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 183.470000 72.240000 183.790000 ;
      LAYER met4 ;
        RECT 71.920000 183.470000 72.240000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 183.875000 72.240000 184.195000 ;
      LAYER met4 ;
        RECT 71.920000 183.875000 72.240000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 184.280000 72.240000 184.600000 ;
      LAYER met4 ;
        RECT 71.920000 184.280000 72.240000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 184.685000 72.240000 185.005000 ;
      LAYER met4 ;
        RECT 71.920000 184.685000 72.240000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 185.090000 72.240000 185.410000 ;
      LAYER met4 ;
        RECT 71.920000 185.090000 72.240000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 185.495000 72.240000 185.815000 ;
      LAYER met4 ;
        RECT 71.920000 185.495000 72.240000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 185.900000 72.240000 186.220000 ;
      LAYER met4 ;
        RECT 71.920000 185.900000 72.240000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 186.305000 72.240000 186.625000 ;
      LAYER met4 ;
        RECT 71.920000 186.305000 72.240000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 186.710000 72.240000 187.030000 ;
      LAYER met4 ;
        RECT 71.920000 186.710000 72.240000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 187.115000 72.240000 187.435000 ;
      LAYER met4 ;
        RECT 71.920000 187.115000 72.240000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 187.520000 72.240000 187.840000 ;
      LAYER met4 ;
        RECT 71.920000 187.520000 72.240000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 187.925000 72.240000 188.245000 ;
      LAYER met4 ;
        RECT 71.920000 187.925000 72.240000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 188.330000 72.240000 188.650000 ;
      LAYER met4 ;
        RECT 71.920000 188.330000 72.240000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 188.735000 72.240000 189.055000 ;
      LAYER met4 ;
        RECT 71.920000 188.735000 72.240000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 189.140000 72.240000 189.460000 ;
      LAYER met4 ;
        RECT 71.920000 189.140000 72.240000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 189.545000 72.240000 189.865000 ;
      LAYER met4 ;
        RECT 71.920000 189.545000 72.240000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 189.950000 72.240000 190.270000 ;
      LAYER met4 ;
        RECT 71.920000 189.950000 72.240000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 190.355000 72.240000 190.675000 ;
      LAYER met4 ;
        RECT 71.920000 190.355000 72.240000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 190.760000 72.240000 191.080000 ;
      LAYER met4 ;
        RECT 71.920000 190.760000 72.240000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 191.165000 72.240000 191.485000 ;
      LAYER met4 ;
        RECT 71.920000 191.165000 72.240000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 191.570000 72.240000 191.890000 ;
      LAYER met4 ;
        RECT 71.920000 191.570000 72.240000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 191.975000 72.240000 192.295000 ;
      LAYER met4 ;
        RECT 71.920000 191.975000 72.240000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 192.380000 72.240000 192.700000 ;
      LAYER met4 ;
        RECT 71.920000 192.380000 72.240000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 192.785000 72.240000 193.105000 ;
      LAYER met4 ;
        RECT 71.920000 192.785000 72.240000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 193.190000 72.240000 193.510000 ;
      LAYER met4 ;
        RECT 71.920000 193.190000 72.240000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 193.595000 72.240000 193.915000 ;
      LAYER met4 ;
        RECT 71.920000 193.595000 72.240000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 194.000000 72.240000 194.320000 ;
      LAYER met4 ;
        RECT 71.920000 194.000000 72.240000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 194.405000 72.240000 194.725000 ;
      LAYER met4 ;
        RECT 71.920000 194.405000 72.240000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 194.810000 72.240000 195.130000 ;
      LAYER met4 ;
        RECT 71.920000 194.810000 72.240000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 195.215000 72.240000 195.535000 ;
      LAYER met4 ;
        RECT 71.920000 195.215000 72.240000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 195.620000 72.240000 195.940000 ;
      LAYER met4 ;
        RECT 71.920000 195.620000 72.240000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 196.025000 72.240000 196.345000 ;
      LAYER met4 ;
        RECT 71.920000 196.025000 72.240000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 196.430000 72.240000 196.750000 ;
      LAYER met4 ;
        RECT 71.920000 196.430000 72.240000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 196.835000 72.240000 197.155000 ;
      LAYER met4 ;
        RECT 71.920000 196.835000 72.240000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 197.240000 72.240000 197.560000 ;
      LAYER met4 ;
        RECT 71.920000 197.240000 72.240000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.920000 197.645000 72.240000 197.965000 ;
      LAYER met4 ;
        RECT 71.920000 197.645000 72.240000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 23.850000 72.640000 24.170000 ;
      LAYER met4 ;
        RECT 72.320000 23.850000 72.640000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 24.280000 72.640000 24.600000 ;
      LAYER met4 ;
        RECT 72.320000 24.280000 72.640000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 24.710000 72.640000 25.030000 ;
      LAYER met4 ;
        RECT 72.320000 24.710000 72.640000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 25.140000 72.640000 25.460000 ;
      LAYER met4 ;
        RECT 72.320000 25.140000 72.640000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 25.570000 72.640000 25.890000 ;
      LAYER met4 ;
        RECT 72.320000 25.570000 72.640000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 26.000000 72.640000 26.320000 ;
      LAYER met4 ;
        RECT 72.320000 26.000000 72.640000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 26.430000 72.640000 26.750000 ;
      LAYER met4 ;
        RECT 72.320000 26.430000 72.640000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 26.860000 72.640000 27.180000 ;
      LAYER met4 ;
        RECT 72.320000 26.860000 72.640000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 27.290000 72.640000 27.610000 ;
      LAYER met4 ;
        RECT 72.320000 27.290000 72.640000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 27.720000 72.640000 28.040000 ;
      LAYER met4 ;
        RECT 72.320000 27.720000 72.640000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 28.150000 72.640000 28.470000 ;
      LAYER met4 ;
        RECT 72.320000 28.150000 72.640000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 173.840000 72.650000 174.160000 ;
      LAYER met4 ;
        RECT 72.330000 173.840000 72.650000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 174.240000 72.650000 174.560000 ;
      LAYER met4 ;
        RECT 72.330000 174.240000 72.650000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 174.640000 72.650000 174.960000 ;
      LAYER met4 ;
        RECT 72.330000 174.640000 72.650000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 175.040000 72.650000 175.360000 ;
      LAYER met4 ;
        RECT 72.330000 175.040000 72.650000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 175.440000 72.650000 175.760000 ;
      LAYER met4 ;
        RECT 72.330000 175.440000 72.650000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 175.840000 72.650000 176.160000 ;
      LAYER met4 ;
        RECT 72.330000 175.840000 72.650000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 176.240000 72.650000 176.560000 ;
      LAYER met4 ;
        RECT 72.330000 176.240000 72.650000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 176.640000 72.650000 176.960000 ;
      LAYER met4 ;
        RECT 72.330000 176.640000 72.650000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 177.040000 72.650000 177.360000 ;
      LAYER met4 ;
        RECT 72.330000 177.040000 72.650000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 177.440000 72.650000 177.760000 ;
      LAYER met4 ;
        RECT 72.330000 177.440000 72.650000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 177.840000 72.650000 178.160000 ;
      LAYER met4 ;
        RECT 72.330000 177.840000 72.650000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 178.240000 72.650000 178.560000 ;
      LAYER met4 ;
        RECT 72.330000 178.240000 72.650000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 178.640000 72.650000 178.960000 ;
      LAYER met4 ;
        RECT 72.330000 178.640000 72.650000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 179.040000 72.650000 179.360000 ;
      LAYER met4 ;
        RECT 72.330000 179.040000 72.650000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 179.440000 72.650000 179.760000 ;
      LAYER met4 ;
        RECT 72.330000 179.440000 72.650000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 179.840000 72.650000 180.160000 ;
      LAYER met4 ;
        RECT 72.330000 179.840000 72.650000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 180.240000 72.650000 180.560000 ;
      LAYER met4 ;
        RECT 72.330000 180.240000 72.650000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 180.640000 72.650000 180.960000 ;
      LAYER met4 ;
        RECT 72.330000 180.640000 72.650000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 181.040000 72.650000 181.360000 ;
      LAYER met4 ;
        RECT 72.330000 181.040000 72.650000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 181.445000 72.650000 181.765000 ;
      LAYER met4 ;
        RECT 72.330000 181.445000 72.650000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 181.850000 72.650000 182.170000 ;
      LAYER met4 ;
        RECT 72.330000 181.850000 72.650000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 182.255000 72.650000 182.575000 ;
      LAYER met4 ;
        RECT 72.330000 182.255000 72.650000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 182.660000 72.650000 182.980000 ;
      LAYER met4 ;
        RECT 72.330000 182.660000 72.650000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 183.065000 72.650000 183.385000 ;
      LAYER met4 ;
        RECT 72.330000 183.065000 72.650000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 183.470000 72.650000 183.790000 ;
      LAYER met4 ;
        RECT 72.330000 183.470000 72.650000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 183.875000 72.650000 184.195000 ;
      LAYER met4 ;
        RECT 72.330000 183.875000 72.650000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 184.280000 72.650000 184.600000 ;
      LAYER met4 ;
        RECT 72.330000 184.280000 72.650000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 184.685000 72.650000 185.005000 ;
      LAYER met4 ;
        RECT 72.330000 184.685000 72.650000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 185.090000 72.650000 185.410000 ;
      LAYER met4 ;
        RECT 72.330000 185.090000 72.650000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 185.495000 72.650000 185.815000 ;
      LAYER met4 ;
        RECT 72.330000 185.495000 72.650000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 185.900000 72.650000 186.220000 ;
      LAYER met4 ;
        RECT 72.330000 185.900000 72.650000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 186.305000 72.650000 186.625000 ;
      LAYER met4 ;
        RECT 72.330000 186.305000 72.650000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 186.710000 72.650000 187.030000 ;
      LAYER met4 ;
        RECT 72.330000 186.710000 72.650000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 187.115000 72.650000 187.435000 ;
      LAYER met4 ;
        RECT 72.330000 187.115000 72.650000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 187.520000 72.650000 187.840000 ;
      LAYER met4 ;
        RECT 72.330000 187.520000 72.650000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 187.925000 72.650000 188.245000 ;
      LAYER met4 ;
        RECT 72.330000 187.925000 72.650000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 188.330000 72.650000 188.650000 ;
      LAYER met4 ;
        RECT 72.330000 188.330000 72.650000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 188.735000 72.650000 189.055000 ;
      LAYER met4 ;
        RECT 72.330000 188.735000 72.650000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 189.140000 72.650000 189.460000 ;
      LAYER met4 ;
        RECT 72.330000 189.140000 72.650000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 189.545000 72.650000 189.865000 ;
      LAYER met4 ;
        RECT 72.330000 189.545000 72.650000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 189.950000 72.650000 190.270000 ;
      LAYER met4 ;
        RECT 72.330000 189.950000 72.650000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 190.355000 72.650000 190.675000 ;
      LAYER met4 ;
        RECT 72.330000 190.355000 72.650000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 190.760000 72.650000 191.080000 ;
      LAYER met4 ;
        RECT 72.330000 190.760000 72.650000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 191.165000 72.650000 191.485000 ;
      LAYER met4 ;
        RECT 72.330000 191.165000 72.650000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 191.570000 72.650000 191.890000 ;
      LAYER met4 ;
        RECT 72.330000 191.570000 72.650000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 191.975000 72.650000 192.295000 ;
      LAYER met4 ;
        RECT 72.330000 191.975000 72.650000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 192.380000 72.650000 192.700000 ;
      LAYER met4 ;
        RECT 72.330000 192.380000 72.650000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 192.785000 72.650000 193.105000 ;
      LAYER met4 ;
        RECT 72.330000 192.785000 72.650000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 193.190000 72.650000 193.510000 ;
      LAYER met4 ;
        RECT 72.330000 193.190000 72.650000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 193.595000 72.650000 193.915000 ;
      LAYER met4 ;
        RECT 72.330000 193.595000 72.650000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 194.000000 72.650000 194.320000 ;
      LAYER met4 ;
        RECT 72.330000 194.000000 72.650000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 194.405000 72.650000 194.725000 ;
      LAYER met4 ;
        RECT 72.330000 194.405000 72.650000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 194.810000 72.650000 195.130000 ;
      LAYER met4 ;
        RECT 72.330000 194.810000 72.650000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 195.215000 72.650000 195.535000 ;
      LAYER met4 ;
        RECT 72.330000 195.215000 72.650000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 195.620000 72.650000 195.940000 ;
      LAYER met4 ;
        RECT 72.330000 195.620000 72.650000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 196.025000 72.650000 196.345000 ;
      LAYER met4 ;
        RECT 72.330000 196.025000 72.650000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 196.430000 72.650000 196.750000 ;
      LAYER met4 ;
        RECT 72.330000 196.430000 72.650000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 196.835000 72.650000 197.155000 ;
      LAYER met4 ;
        RECT 72.330000 196.835000 72.650000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 197.240000 72.650000 197.560000 ;
      LAYER met4 ;
        RECT 72.330000 197.240000 72.650000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330000 197.645000 72.650000 197.965000 ;
      LAYER met4 ;
        RECT 72.330000 197.645000 72.650000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 23.850000 73.045000 24.170000 ;
      LAYER met4 ;
        RECT 72.725000 23.850000 73.045000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 24.280000 73.045000 24.600000 ;
      LAYER met4 ;
        RECT 72.725000 24.280000 73.045000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 24.710000 73.045000 25.030000 ;
      LAYER met4 ;
        RECT 72.725000 24.710000 73.045000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 25.140000 73.045000 25.460000 ;
      LAYER met4 ;
        RECT 72.725000 25.140000 73.045000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 25.570000 73.045000 25.890000 ;
      LAYER met4 ;
        RECT 72.725000 25.570000 73.045000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 26.000000 73.045000 26.320000 ;
      LAYER met4 ;
        RECT 72.725000 26.000000 73.045000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 26.430000 73.045000 26.750000 ;
      LAYER met4 ;
        RECT 72.725000 26.430000 73.045000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 26.860000 73.045000 27.180000 ;
      LAYER met4 ;
        RECT 72.725000 26.860000 73.045000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 27.290000 73.045000 27.610000 ;
      LAYER met4 ;
        RECT 72.725000 27.290000 73.045000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 27.720000 73.045000 28.040000 ;
      LAYER met4 ;
        RECT 72.725000 27.720000 73.045000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 28.150000 73.045000 28.470000 ;
      LAYER met4 ;
        RECT 72.725000 28.150000 73.045000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 173.840000 73.060000 174.160000 ;
      LAYER met4 ;
        RECT 72.740000 173.840000 73.060000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 174.240000 73.060000 174.560000 ;
      LAYER met4 ;
        RECT 72.740000 174.240000 73.060000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 174.640000 73.060000 174.960000 ;
      LAYER met4 ;
        RECT 72.740000 174.640000 73.060000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 175.040000 73.060000 175.360000 ;
      LAYER met4 ;
        RECT 72.740000 175.040000 73.060000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 175.440000 73.060000 175.760000 ;
      LAYER met4 ;
        RECT 72.740000 175.440000 73.060000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 175.840000 73.060000 176.160000 ;
      LAYER met4 ;
        RECT 72.740000 175.840000 73.060000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 176.240000 73.060000 176.560000 ;
      LAYER met4 ;
        RECT 72.740000 176.240000 73.060000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 176.640000 73.060000 176.960000 ;
      LAYER met4 ;
        RECT 72.740000 176.640000 73.060000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 177.040000 73.060000 177.360000 ;
      LAYER met4 ;
        RECT 72.740000 177.040000 73.060000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 177.440000 73.060000 177.760000 ;
      LAYER met4 ;
        RECT 72.740000 177.440000 73.060000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 177.840000 73.060000 178.160000 ;
      LAYER met4 ;
        RECT 72.740000 177.840000 73.060000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 178.240000 73.060000 178.560000 ;
      LAYER met4 ;
        RECT 72.740000 178.240000 73.060000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 178.640000 73.060000 178.960000 ;
      LAYER met4 ;
        RECT 72.740000 178.640000 73.060000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 179.040000 73.060000 179.360000 ;
      LAYER met4 ;
        RECT 72.740000 179.040000 73.060000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 179.440000 73.060000 179.760000 ;
      LAYER met4 ;
        RECT 72.740000 179.440000 73.060000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 179.840000 73.060000 180.160000 ;
      LAYER met4 ;
        RECT 72.740000 179.840000 73.060000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 180.240000 73.060000 180.560000 ;
      LAYER met4 ;
        RECT 72.740000 180.240000 73.060000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 180.640000 73.060000 180.960000 ;
      LAYER met4 ;
        RECT 72.740000 180.640000 73.060000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 181.040000 73.060000 181.360000 ;
      LAYER met4 ;
        RECT 72.740000 181.040000 73.060000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 181.445000 73.060000 181.765000 ;
      LAYER met4 ;
        RECT 72.740000 181.445000 73.060000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 181.850000 73.060000 182.170000 ;
      LAYER met4 ;
        RECT 72.740000 181.850000 73.060000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 182.255000 73.060000 182.575000 ;
      LAYER met4 ;
        RECT 72.740000 182.255000 73.060000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 182.660000 73.060000 182.980000 ;
      LAYER met4 ;
        RECT 72.740000 182.660000 73.060000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 183.065000 73.060000 183.385000 ;
      LAYER met4 ;
        RECT 72.740000 183.065000 73.060000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 183.470000 73.060000 183.790000 ;
      LAYER met4 ;
        RECT 72.740000 183.470000 73.060000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 183.875000 73.060000 184.195000 ;
      LAYER met4 ;
        RECT 72.740000 183.875000 73.060000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 184.280000 73.060000 184.600000 ;
      LAYER met4 ;
        RECT 72.740000 184.280000 73.060000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 184.685000 73.060000 185.005000 ;
      LAYER met4 ;
        RECT 72.740000 184.685000 73.060000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 185.090000 73.060000 185.410000 ;
      LAYER met4 ;
        RECT 72.740000 185.090000 73.060000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 185.495000 73.060000 185.815000 ;
      LAYER met4 ;
        RECT 72.740000 185.495000 73.060000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 185.900000 73.060000 186.220000 ;
      LAYER met4 ;
        RECT 72.740000 185.900000 73.060000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 186.305000 73.060000 186.625000 ;
      LAYER met4 ;
        RECT 72.740000 186.305000 73.060000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 186.710000 73.060000 187.030000 ;
      LAYER met4 ;
        RECT 72.740000 186.710000 73.060000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 187.115000 73.060000 187.435000 ;
      LAYER met4 ;
        RECT 72.740000 187.115000 73.060000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 187.520000 73.060000 187.840000 ;
      LAYER met4 ;
        RECT 72.740000 187.520000 73.060000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 187.925000 73.060000 188.245000 ;
      LAYER met4 ;
        RECT 72.740000 187.925000 73.060000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 188.330000 73.060000 188.650000 ;
      LAYER met4 ;
        RECT 72.740000 188.330000 73.060000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 188.735000 73.060000 189.055000 ;
      LAYER met4 ;
        RECT 72.740000 188.735000 73.060000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 189.140000 73.060000 189.460000 ;
      LAYER met4 ;
        RECT 72.740000 189.140000 73.060000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 189.545000 73.060000 189.865000 ;
      LAYER met4 ;
        RECT 72.740000 189.545000 73.060000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 189.950000 73.060000 190.270000 ;
      LAYER met4 ;
        RECT 72.740000 189.950000 73.060000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 190.355000 73.060000 190.675000 ;
      LAYER met4 ;
        RECT 72.740000 190.355000 73.060000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 190.760000 73.060000 191.080000 ;
      LAYER met4 ;
        RECT 72.740000 190.760000 73.060000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 191.165000 73.060000 191.485000 ;
      LAYER met4 ;
        RECT 72.740000 191.165000 73.060000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 191.570000 73.060000 191.890000 ;
      LAYER met4 ;
        RECT 72.740000 191.570000 73.060000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 191.975000 73.060000 192.295000 ;
      LAYER met4 ;
        RECT 72.740000 191.975000 73.060000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 192.380000 73.060000 192.700000 ;
      LAYER met4 ;
        RECT 72.740000 192.380000 73.060000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 192.785000 73.060000 193.105000 ;
      LAYER met4 ;
        RECT 72.740000 192.785000 73.060000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 193.190000 73.060000 193.510000 ;
      LAYER met4 ;
        RECT 72.740000 193.190000 73.060000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 193.595000 73.060000 193.915000 ;
      LAYER met4 ;
        RECT 72.740000 193.595000 73.060000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 194.000000 73.060000 194.320000 ;
      LAYER met4 ;
        RECT 72.740000 194.000000 73.060000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 194.405000 73.060000 194.725000 ;
      LAYER met4 ;
        RECT 72.740000 194.405000 73.060000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 194.810000 73.060000 195.130000 ;
      LAYER met4 ;
        RECT 72.740000 194.810000 73.060000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 195.215000 73.060000 195.535000 ;
      LAYER met4 ;
        RECT 72.740000 195.215000 73.060000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 195.620000 73.060000 195.940000 ;
      LAYER met4 ;
        RECT 72.740000 195.620000 73.060000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 196.025000 73.060000 196.345000 ;
      LAYER met4 ;
        RECT 72.740000 196.025000 73.060000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 196.430000 73.060000 196.750000 ;
      LAYER met4 ;
        RECT 72.740000 196.430000 73.060000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 196.835000 73.060000 197.155000 ;
      LAYER met4 ;
        RECT 72.740000 196.835000 73.060000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 197.240000 73.060000 197.560000 ;
      LAYER met4 ;
        RECT 72.740000 197.240000 73.060000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.740000 197.645000 73.060000 197.965000 ;
      LAYER met4 ;
        RECT 72.740000 197.645000 73.060000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 23.850000 73.450000 24.170000 ;
      LAYER met4 ;
        RECT 73.130000 23.850000 73.450000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 24.280000 73.450000 24.600000 ;
      LAYER met4 ;
        RECT 73.130000 24.280000 73.450000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 24.710000 73.450000 25.030000 ;
      LAYER met4 ;
        RECT 73.130000 24.710000 73.450000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 25.140000 73.450000 25.460000 ;
      LAYER met4 ;
        RECT 73.130000 25.140000 73.450000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 25.570000 73.450000 25.890000 ;
      LAYER met4 ;
        RECT 73.130000 25.570000 73.450000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 26.000000 73.450000 26.320000 ;
      LAYER met4 ;
        RECT 73.130000 26.000000 73.450000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 26.430000 73.450000 26.750000 ;
      LAYER met4 ;
        RECT 73.130000 26.430000 73.450000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 26.860000 73.450000 27.180000 ;
      LAYER met4 ;
        RECT 73.130000 26.860000 73.450000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 27.290000 73.450000 27.610000 ;
      LAYER met4 ;
        RECT 73.130000 27.290000 73.450000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 27.720000 73.450000 28.040000 ;
      LAYER met4 ;
        RECT 73.130000 27.720000 73.450000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 28.150000 73.450000 28.470000 ;
      LAYER met4 ;
        RECT 73.130000 28.150000 73.450000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 173.840000 73.470000 174.160000 ;
      LAYER met4 ;
        RECT 73.150000 173.840000 73.470000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 174.240000 73.470000 174.560000 ;
      LAYER met4 ;
        RECT 73.150000 174.240000 73.470000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 174.640000 73.470000 174.960000 ;
      LAYER met4 ;
        RECT 73.150000 174.640000 73.470000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 175.040000 73.470000 175.360000 ;
      LAYER met4 ;
        RECT 73.150000 175.040000 73.470000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 175.440000 73.470000 175.760000 ;
      LAYER met4 ;
        RECT 73.150000 175.440000 73.470000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 175.840000 73.470000 176.160000 ;
      LAYER met4 ;
        RECT 73.150000 175.840000 73.470000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 176.240000 73.470000 176.560000 ;
      LAYER met4 ;
        RECT 73.150000 176.240000 73.470000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 176.640000 73.470000 176.960000 ;
      LAYER met4 ;
        RECT 73.150000 176.640000 73.470000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 177.040000 73.470000 177.360000 ;
      LAYER met4 ;
        RECT 73.150000 177.040000 73.470000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 177.440000 73.470000 177.760000 ;
      LAYER met4 ;
        RECT 73.150000 177.440000 73.470000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 177.840000 73.470000 178.160000 ;
      LAYER met4 ;
        RECT 73.150000 177.840000 73.470000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 178.240000 73.470000 178.560000 ;
      LAYER met4 ;
        RECT 73.150000 178.240000 73.470000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 178.640000 73.470000 178.960000 ;
      LAYER met4 ;
        RECT 73.150000 178.640000 73.470000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 179.040000 73.470000 179.360000 ;
      LAYER met4 ;
        RECT 73.150000 179.040000 73.470000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 179.440000 73.470000 179.760000 ;
      LAYER met4 ;
        RECT 73.150000 179.440000 73.470000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 179.840000 73.470000 180.160000 ;
      LAYER met4 ;
        RECT 73.150000 179.840000 73.470000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 180.240000 73.470000 180.560000 ;
      LAYER met4 ;
        RECT 73.150000 180.240000 73.470000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 180.640000 73.470000 180.960000 ;
      LAYER met4 ;
        RECT 73.150000 180.640000 73.470000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 181.040000 73.470000 181.360000 ;
      LAYER met4 ;
        RECT 73.150000 181.040000 73.470000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 181.445000 73.470000 181.765000 ;
      LAYER met4 ;
        RECT 73.150000 181.445000 73.470000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 181.850000 73.470000 182.170000 ;
      LAYER met4 ;
        RECT 73.150000 181.850000 73.470000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 182.255000 73.470000 182.575000 ;
      LAYER met4 ;
        RECT 73.150000 182.255000 73.470000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 182.660000 73.470000 182.980000 ;
      LAYER met4 ;
        RECT 73.150000 182.660000 73.470000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 183.065000 73.470000 183.385000 ;
      LAYER met4 ;
        RECT 73.150000 183.065000 73.470000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 183.470000 73.470000 183.790000 ;
      LAYER met4 ;
        RECT 73.150000 183.470000 73.470000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 183.875000 73.470000 184.195000 ;
      LAYER met4 ;
        RECT 73.150000 183.875000 73.470000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 184.280000 73.470000 184.600000 ;
      LAYER met4 ;
        RECT 73.150000 184.280000 73.470000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 184.685000 73.470000 185.005000 ;
      LAYER met4 ;
        RECT 73.150000 184.685000 73.470000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 185.090000 73.470000 185.410000 ;
      LAYER met4 ;
        RECT 73.150000 185.090000 73.470000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 185.495000 73.470000 185.815000 ;
      LAYER met4 ;
        RECT 73.150000 185.495000 73.470000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 185.900000 73.470000 186.220000 ;
      LAYER met4 ;
        RECT 73.150000 185.900000 73.470000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 186.305000 73.470000 186.625000 ;
      LAYER met4 ;
        RECT 73.150000 186.305000 73.470000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 186.710000 73.470000 187.030000 ;
      LAYER met4 ;
        RECT 73.150000 186.710000 73.470000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 187.115000 73.470000 187.435000 ;
      LAYER met4 ;
        RECT 73.150000 187.115000 73.470000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 187.520000 73.470000 187.840000 ;
      LAYER met4 ;
        RECT 73.150000 187.520000 73.470000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 187.925000 73.470000 188.245000 ;
      LAYER met4 ;
        RECT 73.150000 187.925000 73.470000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 188.330000 73.470000 188.650000 ;
      LAYER met4 ;
        RECT 73.150000 188.330000 73.470000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 188.735000 73.470000 189.055000 ;
      LAYER met4 ;
        RECT 73.150000 188.735000 73.470000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 189.140000 73.470000 189.460000 ;
      LAYER met4 ;
        RECT 73.150000 189.140000 73.470000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 189.545000 73.470000 189.865000 ;
      LAYER met4 ;
        RECT 73.150000 189.545000 73.470000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 189.950000 73.470000 190.270000 ;
      LAYER met4 ;
        RECT 73.150000 189.950000 73.470000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 190.355000 73.470000 190.675000 ;
      LAYER met4 ;
        RECT 73.150000 190.355000 73.470000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 190.760000 73.470000 191.080000 ;
      LAYER met4 ;
        RECT 73.150000 190.760000 73.470000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 191.165000 73.470000 191.485000 ;
      LAYER met4 ;
        RECT 73.150000 191.165000 73.470000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 191.570000 73.470000 191.890000 ;
      LAYER met4 ;
        RECT 73.150000 191.570000 73.470000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 191.975000 73.470000 192.295000 ;
      LAYER met4 ;
        RECT 73.150000 191.975000 73.470000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 192.380000 73.470000 192.700000 ;
      LAYER met4 ;
        RECT 73.150000 192.380000 73.470000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 192.785000 73.470000 193.105000 ;
      LAYER met4 ;
        RECT 73.150000 192.785000 73.470000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 193.190000 73.470000 193.510000 ;
      LAYER met4 ;
        RECT 73.150000 193.190000 73.470000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 193.595000 73.470000 193.915000 ;
      LAYER met4 ;
        RECT 73.150000 193.595000 73.470000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 194.000000 73.470000 194.320000 ;
      LAYER met4 ;
        RECT 73.150000 194.000000 73.470000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 194.405000 73.470000 194.725000 ;
      LAYER met4 ;
        RECT 73.150000 194.405000 73.470000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 194.810000 73.470000 195.130000 ;
      LAYER met4 ;
        RECT 73.150000 194.810000 73.470000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 195.215000 73.470000 195.535000 ;
      LAYER met4 ;
        RECT 73.150000 195.215000 73.470000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 195.620000 73.470000 195.940000 ;
      LAYER met4 ;
        RECT 73.150000 195.620000 73.470000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 196.025000 73.470000 196.345000 ;
      LAYER met4 ;
        RECT 73.150000 196.025000 73.470000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 196.430000 73.470000 196.750000 ;
      LAYER met4 ;
        RECT 73.150000 196.430000 73.470000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 196.835000 73.470000 197.155000 ;
      LAYER met4 ;
        RECT 73.150000 196.835000 73.470000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 197.240000 73.470000 197.560000 ;
      LAYER met4 ;
        RECT 73.150000 197.240000 73.470000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150000 197.645000 73.470000 197.965000 ;
      LAYER met4 ;
        RECT 73.150000 197.645000 73.470000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 23.850000 73.855000 24.170000 ;
      LAYER met4 ;
        RECT 73.535000 23.850000 73.855000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 24.280000 73.855000 24.600000 ;
      LAYER met4 ;
        RECT 73.535000 24.280000 73.855000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 24.710000 73.855000 25.030000 ;
      LAYER met4 ;
        RECT 73.535000 24.710000 73.855000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 25.140000 73.855000 25.460000 ;
      LAYER met4 ;
        RECT 73.535000 25.140000 73.855000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 25.570000 73.855000 25.890000 ;
      LAYER met4 ;
        RECT 73.535000 25.570000 73.855000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 26.000000 73.855000 26.320000 ;
      LAYER met4 ;
        RECT 73.535000 26.000000 73.855000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 26.430000 73.855000 26.750000 ;
      LAYER met4 ;
        RECT 73.535000 26.430000 73.855000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 26.860000 73.855000 27.180000 ;
      LAYER met4 ;
        RECT 73.535000 26.860000 73.855000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 27.290000 73.855000 27.610000 ;
      LAYER met4 ;
        RECT 73.535000 27.290000 73.855000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 27.720000 73.855000 28.040000 ;
      LAYER met4 ;
        RECT 73.535000 27.720000 73.855000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 28.150000 73.855000 28.470000 ;
      LAYER met4 ;
        RECT 73.535000 28.150000 73.855000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 173.840000 73.880000 174.160000 ;
      LAYER met4 ;
        RECT 73.560000 173.840000 73.880000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 174.240000 73.880000 174.560000 ;
      LAYER met4 ;
        RECT 73.560000 174.240000 73.880000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 174.640000 73.880000 174.960000 ;
      LAYER met4 ;
        RECT 73.560000 174.640000 73.880000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 175.040000 73.880000 175.360000 ;
      LAYER met4 ;
        RECT 73.560000 175.040000 73.880000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 175.440000 73.880000 175.760000 ;
      LAYER met4 ;
        RECT 73.560000 175.440000 73.880000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 175.840000 73.880000 176.160000 ;
      LAYER met4 ;
        RECT 73.560000 175.840000 73.880000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 176.240000 73.880000 176.560000 ;
      LAYER met4 ;
        RECT 73.560000 176.240000 73.880000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 176.640000 73.880000 176.960000 ;
      LAYER met4 ;
        RECT 73.560000 176.640000 73.880000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 177.040000 73.880000 177.360000 ;
      LAYER met4 ;
        RECT 73.560000 177.040000 73.880000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 177.440000 73.880000 177.760000 ;
      LAYER met4 ;
        RECT 73.560000 177.440000 73.880000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 177.840000 73.880000 178.160000 ;
      LAYER met4 ;
        RECT 73.560000 177.840000 73.880000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 178.240000 73.880000 178.560000 ;
      LAYER met4 ;
        RECT 73.560000 178.240000 73.880000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 178.640000 73.880000 178.960000 ;
      LAYER met4 ;
        RECT 73.560000 178.640000 73.880000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 179.040000 73.880000 179.360000 ;
      LAYER met4 ;
        RECT 73.560000 179.040000 73.880000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 179.440000 73.880000 179.760000 ;
      LAYER met4 ;
        RECT 73.560000 179.440000 73.880000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 179.840000 73.880000 180.160000 ;
      LAYER met4 ;
        RECT 73.560000 179.840000 73.880000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 180.240000 73.880000 180.560000 ;
      LAYER met4 ;
        RECT 73.560000 180.240000 73.880000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 180.640000 73.880000 180.960000 ;
      LAYER met4 ;
        RECT 73.560000 180.640000 73.880000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 181.040000 73.880000 181.360000 ;
      LAYER met4 ;
        RECT 73.560000 181.040000 73.880000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 181.445000 73.880000 181.765000 ;
      LAYER met4 ;
        RECT 73.560000 181.445000 73.880000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 181.850000 73.880000 182.170000 ;
      LAYER met4 ;
        RECT 73.560000 181.850000 73.880000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 182.255000 73.880000 182.575000 ;
      LAYER met4 ;
        RECT 73.560000 182.255000 73.880000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 182.660000 73.880000 182.980000 ;
      LAYER met4 ;
        RECT 73.560000 182.660000 73.880000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 183.065000 73.880000 183.385000 ;
      LAYER met4 ;
        RECT 73.560000 183.065000 73.880000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 183.470000 73.880000 183.790000 ;
      LAYER met4 ;
        RECT 73.560000 183.470000 73.880000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 183.875000 73.880000 184.195000 ;
      LAYER met4 ;
        RECT 73.560000 183.875000 73.880000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 184.280000 73.880000 184.600000 ;
      LAYER met4 ;
        RECT 73.560000 184.280000 73.880000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 184.685000 73.880000 185.005000 ;
      LAYER met4 ;
        RECT 73.560000 184.685000 73.880000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 185.090000 73.880000 185.410000 ;
      LAYER met4 ;
        RECT 73.560000 185.090000 73.880000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 185.495000 73.880000 185.815000 ;
      LAYER met4 ;
        RECT 73.560000 185.495000 73.880000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 185.900000 73.880000 186.220000 ;
      LAYER met4 ;
        RECT 73.560000 185.900000 73.880000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 186.305000 73.880000 186.625000 ;
      LAYER met4 ;
        RECT 73.560000 186.305000 73.880000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 186.710000 73.880000 187.030000 ;
      LAYER met4 ;
        RECT 73.560000 186.710000 73.880000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 187.115000 73.880000 187.435000 ;
      LAYER met4 ;
        RECT 73.560000 187.115000 73.880000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 187.520000 73.880000 187.840000 ;
      LAYER met4 ;
        RECT 73.560000 187.520000 73.880000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 187.925000 73.880000 188.245000 ;
      LAYER met4 ;
        RECT 73.560000 187.925000 73.880000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 188.330000 73.880000 188.650000 ;
      LAYER met4 ;
        RECT 73.560000 188.330000 73.880000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 188.735000 73.880000 189.055000 ;
      LAYER met4 ;
        RECT 73.560000 188.735000 73.880000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 189.140000 73.880000 189.460000 ;
      LAYER met4 ;
        RECT 73.560000 189.140000 73.880000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 189.545000 73.880000 189.865000 ;
      LAYER met4 ;
        RECT 73.560000 189.545000 73.880000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 189.950000 73.880000 190.270000 ;
      LAYER met4 ;
        RECT 73.560000 189.950000 73.880000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 190.355000 73.880000 190.675000 ;
      LAYER met4 ;
        RECT 73.560000 190.355000 73.880000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 190.760000 73.880000 191.080000 ;
      LAYER met4 ;
        RECT 73.560000 190.760000 73.880000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 191.165000 73.880000 191.485000 ;
      LAYER met4 ;
        RECT 73.560000 191.165000 73.880000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 191.570000 73.880000 191.890000 ;
      LAYER met4 ;
        RECT 73.560000 191.570000 73.880000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 191.975000 73.880000 192.295000 ;
      LAYER met4 ;
        RECT 73.560000 191.975000 73.880000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 192.380000 73.880000 192.700000 ;
      LAYER met4 ;
        RECT 73.560000 192.380000 73.880000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 192.785000 73.880000 193.105000 ;
      LAYER met4 ;
        RECT 73.560000 192.785000 73.880000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 193.190000 73.880000 193.510000 ;
      LAYER met4 ;
        RECT 73.560000 193.190000 73.880000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 193.595000 73.880000 193.915000 ;
      LAYER met4 ;
        RECT 73.560000 193.595000 73.880000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 194.000000 73.880000 194.320000 ;
      LAYER met4 ;
        RECT 73.560000 194.000000 73.880000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 194.405000 73.880000 194.725000 ;
      LAYER met4 ;
        RECT 73.560000 194.405000 73.880000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 194.810000 73.880000 195.130000 ;
      LAYER met4 ;
        RECT 73.560000 194.810000 73.880000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 195.215000 73.880000 195.535000 ;
      LAYER met4 ;
        RECT 73.560000 195.215000 73.880000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 195.620000 73.880000 195.940000 ;
      LAYER met4 ;
        RECT 73.560000 195.620000 73.880000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 196.025000 73.880000 196.345000 ;
      LAYER met4 ;
        RECT 73.560000 196.025000 73.880000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 196.430000 73.880000 196.750000 ;
      LAYER met4 ;
        RECT 73.560000 196.430000 73.880000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 196.835000 73.880000 197.155000 ;
      LAYER met4 ;
        RECT 73.560000 196.835000 73.880000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 197.240000 73.880000 197.560000 ;
      LAYER met4 ;
        RECT 73.560000 197.240000 73.880000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.560000 197.645000 73.880000 197.965000 ;
      LAYER met4 ;
        RECT 73.560000 197.645000 73.880000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 23.850000 74.260000 24.170000 ;
      LAYER met4 ;
        RECT 73.940000 23.850000 74.260000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 24.280000 74.260000 24.600000 ;
      LAYER met4 ;
        RECT 73.940000 24.280000 74.260000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 24.710000 74.260000 25.030000 ;
      LAYER met4 ;
        RECT 73.940000 24.710000 74.260000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 25.140000 74.260000 25.460000 ;
      LAYER met4 ;
        RECT 73.940000 25.140000 74.260000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 25.570000 74.260000 25.890000 ;
      LAYER met4 ;
        RECT 73.940000 25.570000 74.260000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 26.000000 74.260000 26.320000 ;
      LAYER met4 ;
        RECT 73.940000 26.000000 74.260000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 26.430000 74.260000 26.750000 ;
      LAYER met4 ;
        RECT 73.940000 26.430000 74.260000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 26.860000 74.260000 27.180000 ;
      LAYER met4 ;
        RECT 73.940000 26.860000 74.260000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 27.290000 74.260000 27.610000 ;
      LAYER met4 ;
        RECT 73.940000 27.290000 74.260000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 27.720000 74.260000 28.040000 ;
      LAYER met4 ;
        RECT 73.940000 27.720000 74.260000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 28.150000 74.260000 28.470000 ;
      LAYER met4 ;
        RECT 73.940000 28.150000 74.260000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 173.840000 74.290000 174.160000 ;
      LAYER met4 ;
        RECT 73.970000 173.840000 74.290000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 174.240000 74.290000 174.560000 ;
      LAYER met4 ;
        RECT 73.970000 174.240000 74.290000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 174.640000 74.290000 174.960000 ;
      LAYER met4 ;
        RECT 73.970000 174.640000 74.290000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 175.040000 74.290000 175.360000 ;
      LAYER met4 ;
        RECT 73.970000 175.040000 74.290000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 175.440000 74.290000 175.760000 ;
      LAYER met4 ;
        RECT 73.970000 175.440000 74.290000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 175.840000 74.290000 176.160000 ;
      LAYER met4 ;
        RECT 73.970000 175.840000 74.290000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 176.240000 74.290000 176.560000 ;
      LAYER met4 ;
        RECT 73.970000 176.240000 74.290000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 176.640000 74.290000 176.960000 ;
      LAYER met4 ;
        RECT 73.970000 176.640000 74.290000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 177.040000 74.290000 177.360000 ;
      LAYER met4 ;
        RECT 73.970000 177.040000 74.290000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 177.440000 74.290000 177.760000 ;
      LAYER met4 ;
        RECT 73.970000 177.440000 74.290000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 177.840000 74.290000 178.160000 ;
      LAYER met4 ;
        RECT 73.970000 177.840000 74.290000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 178.240000 74.290000 178.560000 ;
      LAYER met4 ;
        RECT 73.970000 178.240000 74.290000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 178.640000 74.290000 178.960000 ;
      LAYER met4 ;
        RECT 73.970000 178.640000 74.290000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 179.040000 74.290000 179.360000 ;
      LAYER met4 ;
        RECT 73.970000 179.040000 74.290000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 179.440000 74.290000 179.760000 ;
      LAYER met4 ;
        RECT 73.970000 179.440000 74.290000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 179.840000 74.290000 180.160000 ;
      LAYER met4 ;
        RECT 73.970000 179.840000 74.290000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 180.240000 74.290000 180.560000 ;
      LAYER met4 ;
        RECT 73.970000 180.240000 74.290000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 180.640000 74.290000 180.960000 ;
      LAYER met4 ;
        RECT 73.970000 180.640000 74.290000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 181.040000 74.290000 181.360000 ;
      LAYER met4 ;
        RECT 73.970000 181.040000 74.290000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 181.445000 74.290000 181.765000 ;
      LAYER met4 ;
        RECT 73.970000 181.445000 74.290000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 181.850000 74.290000 182.170000 ;
      LAYER met4 ;
        RECT 73.970000 181.850000 74.290000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 182.255000 74.290000 182.575000 ;
      LAYER met4 ;
        RECT 73.970000 182.255000 74.290000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 182.660000 74.290000 182.980000 ;
      LAYER met4 ;
        RECT 73.970000 182.660000 74.290000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 183.065000 74.290000 183.385000 ;
      LAYER met4 ;
        RECT 73.970000 183.065000 74.290000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 183.470000 74.290000 183.790000 ;
      LAYER met4 ;
        RECT 73.970000 183.470000 74.290000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 183.875000 74.290000 184.195000 ;
      LAYER met4 ;
        RECT 73.970000 183.875000 74.290000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 184.280000 74.290000 184.600000 ;
      LAYER met4 ;
        RECT 73.970000 184.280000 74.290000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 184.685000 74.290000 185.005000 ;
      LAYER met4 ;
        RECT 73.970000 184.685000 74.290000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 185.090000 74.290000 185.410000 ;
      LAYER met4 ;
        RECT 73.970000 185.090000 74.290000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 185.495000 74.290000 185.815000 ;
      LAYER met4 ;
        RECT 73.970000 185.495000 74.290000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 185.900000 74.290000 186.220000 ;
      LAYER met4 ;
        RECT 73.970000 185.900000 74.290000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 186.305000 74.290000 186.625000 ;
      LAYER met4 ;
        RECT 73.970000 186.305000 74.290000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 186.710000 74.290000 187.030000 ;
      LAYER met4 ;
        RECT 73.970000 186.710000 74.290000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 187.115000 74.290000 187.435000 ;
      LAYER met4 ;
        RECT 73.970000 187.115000 74.290000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 187.520000 74.290000 187.840000 ;
      LAYER met4 ;
        RECT 73.970000 187.520000 74.290000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 187.925000 74.290000 188.245000 ;
      LAYER met4 ;
        RECT 73.970000 187.925000 74.290000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 188.330000 74.290000 188.650000 ;
      LAYER met4 ;
        RECT 73.970000 188.330000 74.290000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 188.735000 74.290000 189.055000 ;
      LAYER met4 ;
        RECT 73.970000 188.735000 74.290000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 189.140000 74.290000 189.460000 ;
      LAYER met4 ;
        RECT 73.970000 189.140000 74.290000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 189.545000 74.290000 189.865000 ;
      LAYER met4 ;
        RECT 73.970000 189.545000 74.290000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 189.950000 74.290000 190.270000 ;
      LAYER met4 ;
        RECT 73.970000 189.950000 74.290000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 190.355000 74.290000 190.675000 ;
      LAYER met4 ;
        RECT 73.970000 190.355000 74.290000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 190.760000 74.290000 191.080000 ;
      LAYER met4 ;
        RECT 73.970000 190.760000 74.290000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 191.165000 74.290000 191.485000 ;
      LAYER met4 ;
        RECT 73.970000 191.165000 74.290000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 191.570000 74.290000 191.890000 ;
      LAYER met4 ;
        RECT 73.970000 191.570000 74.290000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 191.975000 74.290000 192.295000 ;
      LAYER met4 ;
        RECT 73.970000 191.975000 74.290000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 192.380000 74.290000 192.700000 ;
      LAYER met4 ;
        RECT 73.970000 192.380000 74.290000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 192.785000 74.290000 193.105000 ;
      LAYER met4 ;
        RECT 73.970000 192.785000 74.290000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 193.190000 74.290000 193.510000 ;
      LAYER met4 ;
        RECT 73.970000 193.190000 74.290000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 193.595000 74.290000 193.915000 ;
      LAYER met4 ;
        RECT 73.970000 193.595000 74.290000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 194.000000 74.290000 194.320000 ;
      LAYER met4 ;
        RECT 73.970000 194.000000 74.290000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 194.405000 74.290000 194.725000 ;
      LAYER met4 ;
        RECT 73.970000 194.405000 74.290000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 194.810000 74.290000 195.130000 ;
      LAYER met4 ;
        RECT 73.970000 194.810000 74.290000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 195.215000 74.290000 195.535000 ;
      LAYER met4 ;
        RECT 73.970000 195.215000 74.290000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 195.620000 74.290000 195.940000 ;
      LAYER met4 ;
        RECT 73.970000 195.620000 74.290000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 196.025000 74.290000 196.345000 ;
      LAYER met4 ;
        RECT 73.970000 196.025000 74.290000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 196.430000 74.290000 196.750000 ;
      LAYER met4 ;
        RECT 73.970000 196.430000 74.290000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 196.835000 74.290000 197.155000 ;
      LAYER met4 ;
        RECT 73.970000 196.835000 74.290000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 197.240000 74.290000 197.560000 ;
      LAYER met4 ;
        RECT 73.970000 197.240000 74.290000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.970000 197.645000 74.290000 197.965000 ;
      LAYER met4 ;
        RECT 73.970000 197.645000 74.290000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 173.840000 74.700000 174.160000 ;
      LAYER met4 ;
        RECT 74.380000 173.840000 74.700000 174.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 174.240000 74.700000 174.560000 ;
      LAYER met4 ;
        RECT 74.380000 174.240000 74.700000 174.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 174.640000 74.700000 174.960000 ;
      LAYER met4 ;
        RECT 74.380000 174.640000 74.700000 174.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 175.040000 74.700000 175.360000 ;
      LAYER met4 ;
        RECT 74.380000 175.040000 74.700000 175.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 175.440000 74.700000 175.760000 ;
      LAYER met4 ;
        RECT 74.380000 175.440000 74.700000 175.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 175.840000 74.700000 176.160000 ;
      LAYER met4 ;
        RECT 74.380000 175.840000 74.700000 176.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 176.240000 74.700000 176.560000 ;
      LAYER met4 ;
        RECT 74.380000 176.240000 74.700000 176.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 176.640000 74.700000 176.960000 ;
      LAYER met4 ;
        RECT 74.380000 176.640000 74.700000 176.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 177.040000 74.700000 177.360000 ;
      LAYER met4 ;
        RECT 74.380000 177.040000 74.700000 177.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 177.440000 74.700000 177.760000 ;
      LAYER met4 ;
        RECT 74.380000 177.440000 74.700000 177.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 177.840000 74.700000 178.160000 ;
      LAYER met4 ;
        RECT 74.380000 177.840000 74.700000 178.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 178.240000 74.700000 178.560000 ;
      LAYER met4 ;
        RECT 74.380000 178.240000 74.700000 178.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 178.640000 74.700000 178.960000 ;
      LAYER met4 ;
        RECT 74.380000 178.640000 74.700000 178.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 179.040000 74.700000 179.360000 ;
      LAYER met4 ;
        RECT 74.380000 179.040000 74.700000 179.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 179.440000 74.700000 179.760000 ;
      LAYER met4 ;
        RECT 74.380000 179.440000 74.700000 179.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 179.840000 74.700000 180.160000 ;
      LAYER met4 ;
        RECT 74.380000 179.840000 74.700000 180.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 180.240000 74.700000 180.560000 ;
      LAYER met4 ;
        RECT 74.380000 180.240000 74.700000 180.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 180.640000 74.700000 180.960000 ;
      LAYER met4 ;
        RECT 74.380000 180.640000 74.700000 180.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 181.040000 74.700000 181.360000 ;
      LAYER met4 ;
        RECT 74.380000 181.040000 74.700000 181.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 181.445000 74.700000 181.765000 ;
      LAYER met4 ;
        RECT 74.380000 181.445000 74.700000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 181.850000 74.700000 182.170000 ;
      LAYER met4 ;
        RECT 74.380000 181.850000 74.700000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 182.255000 74.700000 182.575000 ;
      LAYER met4 ;
        RECT 74.380000 182.255000 74.700000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 182.660000 74.700000 182.980000 ;
      LAYER met4 ;
        RECT 74.380000 182.660000 74.700000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 183.065000 74.700000 183.385000 ;
      LAYER met4 ;
        RECT 74.380000 183.065000 74.700000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 183.470000 74.700000 183.790000 ;
      LAYER met4 ;
        RECT 74.380000 183.470000 74.700000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 183.875000 74.700000 184.195000 ;
      LAYER met4 ;
        RECT 74.380000 183.875000 74.700000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 184.280000 74.700000 184.600000 ;
      LAYER met4 ;
        RECT 74.380000 184.280000 74.700000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 184.685000 74.700000 185.005000 ;
      LAYER met4 ;
        RECT 74.380000 184.685000 74.700000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 185.090000 74.700000 185.410000 ;
      LAYER met4 ;
        RECT 74.380000 185.090000 74.700000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 185.495000 74.700000 185.815000 ;
      LAYER met4 ;
        RECT 74.380000 185.495000 74.700000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 185.900000 74.700000 186.220000 ;
      LAYER met4 ;
        RECT 74.380000 185.900000 74.700000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 186.305000 74.700000 186.625000 ;
      LAYER met4 ;
        RECT 74.380000 186.305000 74.700000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 186.710000 74.700000 187.030000 ;
      LAYER met4 ;
        RECT 74.380000 186.710000 74.700000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 187.115000 74.700000 187.435000 ;
      LAYER met4 ;
        RECT 74.380000 187.115000 74.700000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 187.520000 74.700000 187.840000 ;
      LAYER met4 ;
        RECT 74.380000 187.520000 74.700000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 187.925000 74.700000 188.245000 ;
      LAYER met4 ;
        RECT 74.380000 187.925000 74.700000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 188.330000 74.700000 188.650000 ;
      LAYER met4 ;
        RECT 74.380000 188.330000 74.700000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 188.735000 74.700000 189.055000 ;
      LAYER met4 ;
        RECT 74.380000 188.735000 74.700000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 189.140000 74.700000 189.460000 ;
      LAYER met4 ;
        RECT 74.380000 189.140000 74.700000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 189.545000 74.700000 189.865000 ;
      LAYER met4 ;
        RECT 74.380000 189.545000 74.700000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 189.950000 74.700000 190.270000 ;
      LAYER met4 ;
        RECT 74.380000 189.950000 74.700000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 190.355000 74.700000 190.675000 ;
      LAYER met4 ;
        RECT 74.380000 190.355000 74.700000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 190.760000 74.700000 191.080000 ;
      LAYER met4 ;
        RECT 74.380000 190.760000 74.700000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 191.165000 74.700000 191.485000 ;
      LAYER met4 ;
        RECT 74.380000 191.165000 74.700000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 191.570000 74.700000 191.890000 ;
      LAYER met4 ;
        RECT 74.380000 191.570000 74.700000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 191.975000 74.700000 192.295000 ;
      LAYER met4 ;
        RECT 74.380000 191.975000 74.700000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 192.380000 74.700000 192.700000 ;
      LAYER met4 ;
        RECT 74.380000 192.380000 74.700000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 192.785000 74.700000 193.105000 ;
      LAYER met4 ;
        RECT 74.380000 192.785000 74.700000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 193.190000 74.700000 193.510000 ;
      LAYER met4 ;
        RECT 74.380000 193.190000 74.700000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 193.595000 74.700000 193.915000 ;
      LAYER met4 ;
        RECT 74.380000 193.595000 74.700000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 194.000000 74.700000 194.320000 ;
      LAYER met4 ;
        RECT 74.380000 194.000000 74.700000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 194.405000 74.700000 194.725000 ;
      LAYER met4 ;
        RECT 74.380000 194.405000 74.700000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 194.810000 74.700000 195.130000 ;
      LAYER met4 ;
        RECT 74.380000 194.810000 74.700000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 195.215000 74.700000 195.535000 ;
      LAYER met4 ;
        RECT 74.380000 195.215000 74.700000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 195.620000 74.700000 195.940000 ;
      LAYER met4 ;
        RECT 74.380000 195.620000 74.700000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 196.025000 74.700000 196.345000 ;
      LAYER met4 ;
        RECT 74.380000 196.025000 74.700000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 196.430000 74.700000 196.750000 ;
      LAYER met4 ;
        RECT 74.380000 196.430000 74.700000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 196.835000 74.700000 197.155000 ;
      LAYER met4 ;
        RECT 74.380000 196.835000 74.700000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 197.240000 74.700000 197.560000 ;
      LAYER met4 ;
        RECT 74.380000 197.240000 74.700000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.380000 197.645000 74.700000 197.965000 ;
      LAYER met4 ;
        RECT 74.380000 197.645000 74.700000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 181.445000 8.475000 181.765000 ;
      LAYER met4 ;
        RECT 8.155000 181.445000 8.475000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 181.850000 8.475000 182.170000 ;
      LAYER met4 ;
        RECT 8.155000 181.850000 8.475000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 182.255000 8.475000 182.575000 ;
      LAYER met4 ;
        RECT 8.155000 182.255000 8.475000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 182.660000 8.475000 182.980000 ;
      LAYER met4 ;
        RECT 8.155000 182.660000 8.475000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 183.065000 8.475000 183.385000 ;
      LAYER met4 ;
        RECT 8.155000 183.065000 8.475000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 183.470000 8.475000 183.790000 ;
      LAYER met4 ;
        RECT 8.155000 183.470000 8.475000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 183.875000 8.475000 184.195000 ;
      LAYER met4 ;
        RECT 8.155000 183.875000 8.475000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 184.280000 8.475000 184.600000 ;
      LAYER met4 ;
        RECT 8.155000 184.280000 8.475000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 184.685000 8.475000 185.005000 ;
      LAYER met4 ;
        RECT 8.155000 184.685000 8.475000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 185.090000 8.475000 185.410000 ;
      LAYER met4 ;
        RECT 8.155000 185.090000 8.475000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 185.495000 8.475000 185.815000 ;
      LAYER met4 ;
        RECT 8.155000 185.495000 8.475000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 185.900000 8.475000 186.220000 ;
      LAYER met4 ;
        RECT 8.155000 185.900000 8.475000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 186.305000 8.475000 186.625000 ;
      LAYER met4 ;
        RECT 8.155000 186.305000 8.475000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 186.710000 8.475000 187.030000 ;
      LAYER met4 ;
        RECT 8.155000 186.710000 8.475000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 187.115000 8.475000 187.435000 ;
      LAYER met4 ;
        RECT 8.155000 187.115000 8.475000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 187.520000 8.475000 187.840000 ;
      LAYER met4 ;
        RECT 8.155000 187.520000 8.475000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 187.925000 8.475000 188.245000 ;
      LAYER met4 ;
        RECT 8.155000 187.925000 8.475000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 188.330000 8.475000 188.650000 ;
      LAYER met4 ;
        RECT 8.155000 188.330000 8.475000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 188.735000 8.475000 189.055000 ;
      LAYER met4 ;
        RECT 8.155000 188.735000 8.475000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 189.140000 8.475000 189.460000 ;
      LAYER met4 ;
        RECT 8.155000 189.140000 8.475000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 189.545000 8.475000 189.865000 ;
      LAYER met4 ;
        RECT 8.155000 189.545000 8.475000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 189.950000 8.475000 190.270000 ;
      LAYER met4 ;
        RECT 8.155000 189.950000 8.475000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 190.355000 8.475000 190.675000 ;
      LAYER met4 ;
        RECT 8.155000 190.355000 8.475000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 190.760000 8.475000 191.080000 ;
      LAYER met4 ;
        RECT 8.155000 190.760000 8.475000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 191.165000 8.475000 191.485000 ;
      LAYER met4 ;
        RECT 8.155000 191.165000 8.475000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 191.570000 8.475000 191.890000 ;
      LAYER met4 ;
        RECT 8.155000 191.570000 8.475000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 191.975000 8.475000 192.295000 ;
      LAYER met4 ;
        RECT 8.155000 191.975000 8.475000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 192.380000 8.475000 192.700000 ;
      LAYER met4 ;
        RECT 8.155000 192.380000 8.475000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 192.785000 8.475000 193.105000 ;
      LAYER met4 ;
        RECT 8.155000 192.785000 8.475000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 193.190000 8.475000 193.510000 ;
      LAYER met4 ;
        RECT 8.155000 193.190000 8.475000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 193.595000 8.475000 193.915000 ;
      LAYER met4 ;
        RECT 8.155000 193.595000 8.475000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 194.000000 8.475000 194.320000 ;
      LAYER met4 ;
        RECT 8.155000 194.000000 8.475000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 194.405000 8.475000 194.725000 ;
      LAYER met4 ;
        RECT 8.155000 194.405000 8.475000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 194.810000 8.475000 195.130000 ;
      LAYER met4 ;
        RECT 8.155000 194.810000 8.475000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 195.215000 8.475000 195.535000 ;
      LAYER met4 ;
        RECT 8.155000 195.215000 8.475000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 195.620000 8.475000 195.940000 ;
      LAYER met4 ;
        RECT 8.155000 195.620000 8.475000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 196.025000 8.475000 196.345000 ;
      LAYER met4 ;
        RECT 8.155000 196.025000 8.475000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 196.430000 8.475000 196.750000 ;
      LAYER met4 ;
        RECT 8.155000 196.430000 8.475000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 196.835000 8.475000 197.155000 ;
      LAYER met4 ;
        RECT 8.155000 196.835000 8.475000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 197.240000 8.475000 197.560000 ;
      LAYER met4 ;
        RECT 8.155000 197.240000 8.475000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155000 197.645000 8.475000 197.965000 ;
      LAYER met4 ;
        RECT 8.155000 197.645000 8.475000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.215000 173.900000 8.415000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.215000 174.300000 8.415000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.215000 174.700000 8.415000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.215000 175.100000 8.415000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.215000 175.500000 8.415000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.215000 175.900000 8.415000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.215000 176.300000 8.415000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.215000 176.700000 8.415000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.215000 177.100000 8.415000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.215000 177.500000 8.415000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.215000 177.900000 8.415000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.215000 178.300000 8.415000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.215000 178.700000 8.415000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.215000 179.100000 8.415000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.215000 179.500000 8.415000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.215000 179.900000 8.415000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.215000 180.300000 8.415000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.215000 180.700000 8.415000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.215000 181.100000 8.415000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 23.850000 8.575000 24.170000 ;
      LAYER met4 ;
        RECT 8.255000 23.850000 8.575000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 24.280000 8.575000 24.600000 ;
      LAYER met4 ;
        RECT 8.255000 24.280000 8.575000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 24.710000 8.575000 25.030000 ;
      LAYER met4 ;
        RECT 8.255000 24.710000 8.575000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 25.140000 8.575000 25.460000 ;
      LAYER met4 ;
        RECT 8.255000 25.140000 8.575000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 25.570000 8.575000 25.890000 ;
      LAYER met4 ;
        RECT 8.255000 25.570000 8.575000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 26.000000 8.575000 26.320000 ;
      LAYER met4 ;
        RECT 8.255000 26.000000 8.575000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 26.430000 8.575000 26.750000 ;
      LAYER met4 ;
        RECT 8.255000 26.430000 8.575000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 26.860000 8.575000 27.180000 ;
      LAYER met4 ;
        RECT 8.255000 26.860000 8.575000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 27.290000 8.575000 27.610000 ;
      LAYER met4 ;
        RECT 8.255000 27.290000 8.575000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 27.720000 8.575000 28.040000 ;
      LAYER met4 ;
        RECT 8.255000 27.720000 8.575000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 28.150000 8.575000 28.470000 ;
      LAYER met4 ;
        RECT 8.255000 28.150000 8.575000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 181.445000 8.875000 181.765000 ;
      LAYER met4 ;
        RECT 8.555000 181.445000 8.875000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 181.850000 8.875000 182.170000 ;
      LAYER met4 ;
        RECT 8.555000 181.850000 8.875000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 182.255000 8.875000 182.575000 ;
      LAYER met4 ;
        RECT 8.555000 182.255000 8.875000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 182.660000 8.875000 182.980000 ;
      LAYER met4 ;
        RECT 8.555000 182.660000 8.875000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 183.065000 8.875000 183.385000 ;
      LAYER met4 ;
        RECT 8.555000 183.065000 8.875000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 183.470000 8.875000 183.790000 ;
      LAYER met4 ;
        RECT 8.555000 183.470000 8.875000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 183.875000 8.875000 184.195000 ;
      LAYER met4 ;
        RECT 8.555000 183.875000 8.875000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 184.280000 8.875000 184.600000 ;
      LAYER met4 ;
        RECT 8.555000 184.280000 8.875000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 184.685000 8.875000 185.005000 ;
      LAYER met4 ;
        RECT 8.555000 184.685000 8.875000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 185.090000 8.875000 185.410000 ;
      LAYER met4 ;
        RECT 8.555000 185.090000 8.875000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 185.495000 8.875000 185.815000 ;
      LAYER met4 ;
        RECT 8.555000 185.495000 8.875000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 185.900000 8.875000 186.220000 ;
      LAYER met4 ;
        RECT 8.555000 185.900000 8.875000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 186.305000 8.875000 186.625000 ;
      LAYER met4 ;
        RECT 8.555000 186.305000 8.875000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 186.710000 8.875000 187.030000 ;
      LAYER met4 ;
        RECT 8.555000 186.710000 8.875000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 187.115000 8.875000 187.435000 ;
      LAYER met4 ;
        RECT 8.555000 187.115000 8.875000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 187.520000 8.875000 187.840000 ;
      LAYER met4 ;
        RECT 8.555000 187.520000 8.875000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 187.925000 8.875000 188.245000 ;
      LAYER met4 ;
        RECT 8.555000 187.925000 8.875000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 188.330000 8.875000 188.650000 ;
      LAYER met4 ;
        RECT 8.555000 188.330000 8.875000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 188.735000 8.875000 189.055000 ;
      LAYER met4 ;
        RECT 8.555000 188.735000 8.875000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 189.140000 8.875000 189.460000 ;
      LAYER met4 ;
        RECT 8.555000 189.140000 8.875000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 189.545000 8.875000 189.865000 ;
      LAYER met4 ;
        RECT 8.555000 189.545000 8.875000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 189.950000 8.875000 190.270000 ;
      LAYER met4 ;
        RECT 8.555000 189.950000 8.875000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 190.355000 8.875000 190.675000 ;
      LAYER met4 ;
        RECT 8.555000 190.355000 8.875000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 190.760000 8.875000 191.080000 ;
      LAYER met4 ;
        RECT 8.555000 190.760000 8.875000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 191.165000 8.875000 191.485000 ;
      LAYER met4 ;
        RECT 8.555000 191.165000 8.875000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 191.570000 8.875000 191.890000 ;
      LAYER met4 ;
        RECT 8.555000 191.570000 8.875000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 191.975000 8.875000 192.295000 ;
      LAYER met4 ;
        RECT 8.555000 191.975000 8.875000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 192.380000 8.875000 192.700000 ;
      LAYER met4 ;
        RECT 8.555000 192.380000 8.875000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 192.785000 8.875000 193.105000 ;
      LAYER met4 ;
        RECT 8.555000 192.785000 8.875000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 193.190000 8.875000 193.510000 ;
      LAYER met4 ;
        RECT 8.555000 193.190000 8.875000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 193.595000 8.875000 193.915000 ;
      LAYER met4 ;
        RECT 8.555000 193.595000 8.875000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 194.000000 8.875000 194.320000 ;
      LAYER met4 ;
        RECT 8.555000 194.000000 8.875000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 194.405000 8.875000 194.725000 ;
      LAYER met4 ;
        RECT 8.555000 194.405000 8.875000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 194.810000 8.875000 195.130000 ;
      LAYER met4 ;
        RECT 8.555000 194.810000 8.875000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 195.215000 8.875000 195.535000 ;
      LAYER met4 ;
        RECT 8.555000 195.215000 8.875000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 195.620000 8.875000 195.940000 ;
      LAYER met4 ;
        RECT 8.555000 195.620000 8.875000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 196.025000 8.875000 196.345000 ;
      LAYER met4 ;
        RECT 8.555000 196.025000 8.875000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 196.430000 8.875000 196.750000 ;
      LAYER met4 ;
        RECT 8.555000 196.430000 8.875000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 196.835000 8.875000 197.155000 ;
      LAYER met4 ;
        RECT 8.555000 196.835000 8.875000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 197.240000 8.875000 197.560000 ;
      LAYER met4 ;
        RECT 8.555000 197.240000 8.875000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555000 197.645000 8.875000 197.965000 ;
      LAYER met4 ;
        RECT 8.555000 197.645000 8.875000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.615000 173.900000 8.815000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.615000 174.300000 8.815000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.615000 174.700000 8.815000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.615000 175.100000 8.815000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.615000 175.500000 8.815000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.615000 175.900000 8.815000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.615000 176.300000 8.815000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.615000 176.700000 8.815000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.615000 177.100000 8.815000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.615000 177.500000 8.815000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.615000 177.900000 8.815000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.615000 178.300000 8.815000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.615000 178.700000 8.815000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.615000 179.100000 8.815000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.615000 179.500000 8.815000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.615000 179.900000 8.815000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.615000 180.300000 8.815000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.615000 180.700000 8.815000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.615000 181.100000 8.815000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 23.850000 8.980000 24.170000 ;
      LAYER met4 ;
        RECT 8.660000 23.850000 8.980000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 24.280000 8.980000 24.600000 ;
      LAYER met4 ;
        RECT 8.660000 24.280000 8.980000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 24.710000 8.980000 25.030000 ;
      LAYER met4 ;
        RECT 8.660000 24.710000 8.980000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 25.140000 8.980000 25.460000 ;
      LAYER met4 ;
        RECT 8.660000 25.140000 8.980000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 25.570000 8.980000 25.890000 ;
      LAYER met4 ;
        RECT 8.660000 25.570000 8.980000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 26.000000 8.980000 26.320000 ;
      LAYER met4 ;
        RECT 8.660000 26.000000 8.980000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 26.430000 8.980000 26.750000 ;
      LAYER met4 ;
        RECT 8.660000 26.430000 8.980000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 26.860000 8.980000 27.180000 ;
      LAYER met4 ;
        RECT 8.660000 26.860000 8.980000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 27.290000 8.980000 27.610000 ;
      LAYER met4 ;
        RECT 8.660000 27.290000 8.980000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 27.720000 8.980000 28.040000 ;
      LAYER met4 ;
        RECT 8.660000 27.720000 8.980000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 28.150000 8.980000 28.470000 ;
      LAYER met4 ;
        RECT 8.660000 28.150000 8.980000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 181.445000 9.275000 181.765000 ;
      LAYER met4 ;
        RECT 8.955000 181.445000 9.275000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 181.850000 9.275000 182.170000 ;
      LAYER met4 ;
        RECT 8.955000 181.850000 9.275000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 182.255000 9.275000 182.575000 ;
      LAYER met4 ;
        RECT 8.955000 182.255000 9.275000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 182.660000 9.275000 182.980000 ;
      LAYER met4 ;
        RECT 8.955000 182.660000 9.275000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 183.065000 9.275000 183.385000 ;
      LAYER met4 ;
        RECT 8.955000 183.065000 9.275000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 183.470000 9.275000 183.790000 ;
      LAYER met4 ;
        RECT 8.955000 183.470000 9.275000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 183.875000 9.275000 184.195000 ;
      LAYER met4 ;
        RECT 8.955000 183.875000 9.275000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 184.280000 9.275000 184.600000 ;
      LAYER met4 ;
        RECT 8.955000 184.280000 9.275000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 184.685000 9.275000 185.005000 ;
      LAYER met4 ;
        RECT 8.955000 184.685000 9.275000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 185.090000 9.275000 185.410000 ;
      LAYER met4 ;
        RECT 8.955000 185.090000 9.275000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 185.495000 9.275000 185.815000 ;
      LAYER met4 ;
        RECT 8.955000 185.495000 9.275000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 185.900000 9.275000 186.220000 ;
      LAYER met4 ;
        RECT 8.955000 185.900000 9.275000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 186.305000 9.275000 186.625000 ;
      LAYER met4 ;
        RECT 8.955000 186.305000 9.275000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 186.710000 9.275000 187.030000 ;
      LAYER met4 ;
        RECT 8.955000 186.710000 9.275000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 187.115000 9.275000 187.435000 ;
      LAYER met4 ;
        RECT 8.955000 187.115000 9.275000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 187.520000 9.275000 187.840000 ;
      LAYER met4 ;
        RECT 8.955000 187.520000 9.275000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 187.925000 9.275000 188.245000 ;
      LAYER met4 ;
        RECT 8.955000 187.925000 9.275000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 188.330000 9.275000 188.650000 ;
      LAYER met4 ;
        RECT 8.955000 188.330000 9.275000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 188.735000 9.275000 189.055000 ;
      LAYER met4 ;
        RECT 8.955000 188.735000 9.275000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 189.140000 9.275000 189.460000 ;
      LAYER met4 ;
        RECT 8.955000 189.140000 9.275000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 189.545000 9.275000 189.865000 ;
      LAYER met4 ;
        RECT 8.955000 189.545000 9.275000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 189.950000 9.275000 190.270000 ;
      LAYER met4 ;
        RECT 8.955000 189.950000 9.275000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 190.355000 9.275000 190.675000 ;
      LAYER met4 ;
        RECT 8.955000 190.355000 9.275000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 190.760000 9.275000 191.080000 ;
      LAYER met4 ;
        RECT 8.955000 190.760000 9.275000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 191.165000 9.275000 191.485000 ;
      LAYER met4 ;
        RECT 8.955000 191.165000 9.275000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 191.570000 9.275000 191.890000 ;
      LAYER met4 ;
        RECT 8.955000 191.570000 9.275000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 191.975000 9.275000 192.295000 ;
      LAYER met4 ;
        RECT 8.955000 191.975000 9.275000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 192.380000 9.275000 192.700000 ;
      LAYER met4 ;
        RECT 8.955000 192.380000 9.275000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 192.785000 9.275000 193.105000 ;
      LAYER met4 ;
        RECT 8.955000 192.785000 9.275000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 193.190000 9.275000 193.510000 ;
      LAYER met4 ;
        RECT 8.955000 193.190000 9.275000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 193.595000 9.275000 193.915000 ;
      LAYER met4 ;
        RECT 8.955000 193.595000 9.275000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 194.000000 9.275000 194.320000 ;
      LAYER met4 ;
        RECT 8.955000 194.000000 9.275000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 194.405000 9.275000 194.725000 ;
      LAYER met4 ;
        RECT 8.955000 194.405000 9.275000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 194.810000 9.275000 195.130000 ;
      LAYER met4 ;
        RECT 8.955000 194.810000 9.275000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 195.215000 9.275000 195.535000 ;
      LAYER met4 ;
        RECT 8.955000 195.215000 9.275000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 195.620000 9.275000 195.940000 ;
      LAYER met4 ;
        RECT 8.955000 195.620000 9.275000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 196.025000 9.275000 196.345000 ;
      LAYER met4 ;
        RECT 8.955000 196.025000 9.275000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 196.430000 9.275000 196.750000 ;
      LAYER met4 ;
        RECT 8.955000 196.430000 9.275000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 196.835000 9.275000 197.155000 ;
      LAYER met4 ;
        RECT 8.955000 196.835000 9.275000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 197.240000 9.275000 197.560000 ;
      LAYER met4 ;
        RECT 8.955000 197.240000 9.275000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955000 197.645000 9.275000 197.965000 ;
      LAYER met4 ;
        RECT 8.955000 197.645000 9.275000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.015000 173.900000 9.215000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.015000 174.300000 9.215000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.015000 174.700000 9.215000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.015000 175.100000 9.215000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.015000 175.500000 9.215000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.015000 175.900000 9.215000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.015000 176.300000 9.215000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.015000 176.700000 9.215000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.015000 177.100000 9.215000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.015000 177.500000 9.215000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.015000 177.900000 9.215000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.015000 178.300000 9.215000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.015000 178.700000 9.215000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.015000 179.100000 9.215000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.015000 179.500000 9.215000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.015000 179.900000 9.215000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.015000 180.300000 9.215000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.015000 180.700000 9.215000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.015000 181.100000 9.215000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 23.850000 9.385000 24.170000 ;
      LAYER met4 ;
        RECT 9.065000 23.850000 9.385000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 24.280000 9.385000 24.600000 ;
      LAYER met4 ;
        RECT 9.065000 24.280000 9.385000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 24.710000 9.385000 25.030000 ;
      LAYER met4 ;
        RECT 9.065000 24.710000 9.385000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 25.140000 9.385000 25.460000 ;
      LAYER met4 ;
        RECT 9.065000 25.140000 9.385000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 25.570000 9.385000 25.890000 ;
      LAYER met4 ;
        RECT 9.065000 25.570000 9.385000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 26.000000 9.385000 26.320000 ;
      LAYER met4 ;
        RECT 9.065000 26.000000 9.385000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 26.430000 9.385000 26.750000 ;
      LAYER met4 ;
        RECT 9.065000 26.430000 9.385000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 26.860000 9.385000 27.180000 ;
      LAYER met4 ;
        RECT 9.065000 26.860000 9.385000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 27.290000 9.385000 27.610000 ;
      LAYER met4 ;
        RECT 9.065000 27.290000 9.385000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 27.720000 9.385000 28.040000 ;
      LAYER met4 ;
        RECT 9.065000 27.720000 9.385000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 28.150000 9.385000 28.470000 ;
      LAYER met4 ;
        RECT 9.065000 28.150000 9.385000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 181.445000 9.675000 181.765000 ;
      LAYER met4 ;
        RECT 9.355000 181.445000 9.675000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 181.850000 9.675000 182.170000 ;
      LAYER met4 ;
        RECT 9.355000 181.850000 9.675000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 182.255000 9.675000 182.575000 ;
      LAYER met4 ;
        RECT 9.355000 182.255000 9.675000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 182.660000 9.675000 182.980000 ;
      LAYER met4 ;
        RECT 9.355000 182.660000 9.675000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 183.065000 9.675000 183.385000 ;
      LAYER met4 ;
        RECT 9.355000 183.065000 9.675000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 183.470000 9.675000 183.790000 ;
      LAYER met4 ;
        RECT 9.355000 183.470000 9.675000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 183.875000 9.675000 184.195000 ;
      LAYER met4 ;
        RECT 9.355000 183.875000 9.675000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 184.280000 9.675000 184.600000 ;
      LAYER met4 ;
        RECT 9.355000 184.280000 9.675000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 184.685000 9.675000 185.005000 ;
      LAYER met4 ;
        RECT 9.355000 184.685000 9.675000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 185.090000 9.675000 185.410000 ;
      LAYER met4 ;
        RECT 9.355000 185.090000 9.675000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 185.495000 9.675000 185.815000 ;
      LAYER met4 ;
        RECT 9.355000 185.495000 9.675000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 185.900000 9.675000 186.220000 ;
      LAYER met4 ;
        RECT 9.355000 185.900000 9.675000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 186.305000 9.675000 186.625000 ;
      LAYER met4 ;
        RECT 9.355000 186.305000 9.675000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 186.710000 9.675000 187.030000 ;
      LAYER met4 ;
        RECT 9.355000 186.710000 9.675000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 187.115000 9.675000 187.435000 ;
      LAYER met4 ;
        RECT 9.355000 187.115000 9.675000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 187.520000 9.675000 187.840000 ;
      LAYER met4 ;
        RECT 9.355000 187.520000 9.675000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 187.925000 9.675000 188.245000 ;
      LAYER met4 ;
        RECT 9.355000 187.925000 9.675000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 188.330000 9.675000 188.650000 ;
      LAYER met4 ;
        RECT 9.355000 188.330000 9.675000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 188.735000 9.675000 189.055000 ;
      LAYER met4 ;
        RECT 9.355000 188.735000 9.675000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 189.140000 9.675000 189.460000 ;
      LAYER met4 ;
        RECT 9.355000 189.140000 9.675000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 189.545000 9.675000 189.865000 ;
      LAYER met4 ;
        RECT 9.355000 189.545000 9.675000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 189.950000 9.675000 190.270000 ;
      LAYER met4 ;
        RECT 9.355000 189.950000 9.675000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 190.355000 9.675000 190.675000 ;
      LAYER met4 ;
        RECT 9.355000 190.355000 9.675000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 190.760000 9.675000 191.080000 ;
      LAYER met4 ;
        RECT 9.355000 190.760000 9.675000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 191.165000 9.675000 191.485000 ;
      LAYER met4 ;
        RECT 9.355000 191.165000 9.675000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 191.570000 9.675000 191.890000 ;
      LAYER met4 ;
        RECT 9.355000 191.570000 9.675000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 191.975000 9.675000 192.295000 ;
      LAYER met4 ;
        RECT 9.355000 191.975000 9.675000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 192.380000 9.675000 192.700000 ;
      LAYER met4 ;
        RECT 9.355000 192.380000 9.675000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 192.785000 9.675000 193.105000 ;
      LAYER met4 ;
        RECT 9.355000 192.785000 9.675000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 193.190000 9.675000 193.510000 ;
      LAYER met4 ;
        RECT 9.355000 193.190000 9.675000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 193.595000 9.675000 193.915000 ;
      LAYER met4 ;
        RECT 9.355000 193.595000 9.675000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 194.000000 9.675000 194.320000 ;
      LAYER met4 ;
        RECT 9.355000 194.000000 9.675000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 194.405000 9.675000 194.725000 ;
      LAYER met4 ;
        RECT 9.355000 194.405000 9.675000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 194.810000 9.675000 195.130000 ;
      LAYER met4 ;
        RECT 9.355000 194.810000 9.675000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 195.215000 9.675000 195.535000 ;
      LAYER met4 ;
        RECT 9.355000 195.215000 9.675000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 195.620000 9.675000 195.940000 ;
      LAYER met4 ;
        RECT 9.355000 195.620000 9.675000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 196.025000 9.675000 196.345000 ;
      LAYER met4 ;
        RECT 9.355000 196.025000 9.675000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 196.430000 9.675000 196.750000 ;
      LAYER met4 ;
        RECT 9.355000 196.430000 9.675000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 196.835000 9.675000 197.155000 ;
      LAYER met4 ;
        RECT 9.355000 196.835000 9.675000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 197.240000 9.675000 197.560000 ;
      LAYER met4 ;
        RECT 9.355000 197.240000 9.675000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355000 197.645000 9.675000 197.965000 ;
      LAYER met4 ;
        RECT 9.355000 197.645000 9.675000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.415000 173.900000 9.615000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.415000 174.300000 9.615000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.415000 174.700000 9.615000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.415000 175.100000 9.615000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.415000 175.500000 9.615000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.415000 175.900000 9.615000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.415000 176.300000 9.615000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.415000 176.700000 9.615000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.415000 177.100000 9.615000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.415000 177.500000 9.615000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.415000 177.900000 9.615000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.415000 178.300000 9.615000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.415000 178.700000 9.615000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.415000 179.100000 9.615000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.415000 179.500000 9.615000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.415000 179.900000 9.615000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.415000 180.300000 9.615000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.415000 180.700000 9.615000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.415000 181.100000 9.615000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 23.850000 9.790000 24.170000 ;
      LAYER met4 ;
        RECT 9.470000 23.850000 9.790000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 24.280000 9.790000 24.600000 ;
      LAYER met4 ;
        RECT 9.470000 24.280000 9.790000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 24.710000 9.790000 25.030000 ;
      LAYER met4 ;
        RECT 9.470000 24.710000 9.790000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 25.140000 9.790000 25.460000 ;
      LAYER met4 ;
        RECT 9.470000 25.140000 9.790000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 25.570000 9.790000 25.890000 ;
      LAYER met4 ;
        RECT 9.470000 25.570000 9.790000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 26.000000 9.790000 26.320000 ;
      LAYER met4 ;
        RECT 9.470000 26.000000 9.790000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 26.430000 9.790000 26.750000 ;
      LAYER met4 ;
        RECT 9.470000 26.430000 9.790000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 26.860000 9.790000 27.180000 ;
      LAYER met4 ;
        RECT 9.470000 26.860000 9.790000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 27.290000 9.790000 27.610000 ;
      LAYER met4 ;
        RECT 9.470000 27.290000 9.790000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 27.720000 9.790000 28.040000 ;
      LAYER met4 ;
        RECT 9.470000 27.720000 9.790000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 28.150000 9.790000 28.470000 ;
      LAYER met4 ;
        RECT 9.470000 28.150000 9.790000 28.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 181.445000 10.075000 181.765000 ;
      LAYER met4 ;
        RECT 9.755000 181.445000 10.075000 181.765000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 181.850000 10.075000 182.170000 ;
      LAYER met4 ;
        RECT 9.755000 181.850000 10.075000 182.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 182.255000 10.075000 182.575000 ;
      LAYER met4 ;
        RECT 9.755000 182.255000 10.075000 182.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 182.660000 10.075000 182.980000 ;
      LAYER met4 ;
        RECT 9.755000 182.660000 10.075000 182.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 183.065000 10.075000 183.385000 ;
      LAYER met4 ;
        RECT 9.755000 183.065000 10.075000 183.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 183.470000 10.075000 183.790000 ;
      LAYER met4 ;
        RECT 9.755000 183.470000 10.075000 183.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 183.875000 10.075000 184.195000 ;
      LAYER met4 ;
        RECT 9.755000 183.875000 10.075000 184.195000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 184.280000 10.075000 184.600000 ;
      LAYER met4 ;
        RECT 9.755000 184.280000 10.075000 184.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 184.685000 10.075000 185.005000 ;
      LAYER met4 ;
        RECT 9.755000 184.685000 10.075000 185.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 185.090000 10.075000 185.410000 ;
      LAYER met4 ;
        RECT 9.755000 185.090000 10.075000 185.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 185.495000 10.075000 185.815000 ;
      LAYER met4 ;
        RECT 9.755000 185.495000 10.075000 185.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 185.900000 10.075000 186.220000 ;
      LAYER met4 ;
        RECT 9.755000 185.900000 10.075000 186.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 186.305000 10.075000 186.625000 ;
      LAYER met4 ;
        RECT 9.755000 186.305000 10.075000 186.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 186.710000 10.075000 187.030000 ;
      LAYER met4 ;
        RECT 9.755000 186.710000 10.075000 187.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 187.115000 10.075000 187.435000 ;
      LAYER met4 ;
        RECT 9.755000 187.115000 10.075000 187.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 187.520000 10.075000 187.840000 ;
      LAYER met4 ;
        RECT 9.755000 187.520000 10.075000 187.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 187.925000 10.075000 188.245000 ;
      LAYER met4 ;
        RECT 9.755000 187.925000 10.075000 188.245000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 188.330000 10.075000 188.650000 ;
      LAYER met4 ;
        RECT 9.755000 188.330000 10.075000 188.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 188.735000 10.075000 189.055000 ;
      LAYER met4 ;
        RECT 9.755000 188.735000 10.075000 189.055000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 189.140000 10.075000 189.460000 ;
      LAYER met4 ;
        RECT 9.755000 189.140000 10.075000 189.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 189.545000 10.075000 189.865000 ;
      LAYER met4 ;
        RECT 9.755000 189.545000 10.075000 189.865000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 189.950000 10.075000 190.270000 ;
      LAYER met4 ;
        RECT 9.755000 189.950000 10.075000 190.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 190.355000 10.075000 190.675000 ;
      LAYER met4 ;
        RECT 9.755000 190.355000 10.075000 190.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 190.760000 10.075000 191.080000 ;
      LAYER met4 ;
        RECT 9.755000 190.760000 10.075000 191.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 191.165000 10.075000 191.485000 ;
      LAYER met4 ;
        RECT 9.755000 191.165000 10.075000 191.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 191.570000 10.075000 191.890000 ;
      LAYER met4 ;
        RECT 9.755000 191.570000 10.075000 191.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 191.975000 10.075000 192.295000 ;
      LAYER met4 ;
        RECT 9.755000 191.975000 10.075000 192.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 192.380000 10.075000 192.700000 ;
      LAYER met4 ;
        RECT 9.755000 192.380000 10.075000 192.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 192.785000 10.075000 193.105000 ;
      LAYER met4 ;
        RECT 9.755000 192.785000 10.075000 193.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 193.190000 10.075000 193.510000 ;
      LAYER met4 ;
        RECT 9.755000 193.190000 10.075000 193.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 193.595000 10.075000 193.915000 ;
      LAYER met4 ;
        RECT 9.755000 193.595000 10.075000 193.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 194.000000 10.075000 194.320000 ;
      LAYER met4 ;
        RECT 9.755000 194.000000 10.075000 194.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 194.405000 10.075000 194.725000 ;
      LAYER met4 ;
        RECT 9.755000 194.405000 10.075000 194.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 194.810000 10.075000 195.130000 ;
      LAYER met4 ;
        RECT 9.755000 194.810000 10.075000 195.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 195.215000 10.075000 195.535000 ;
      LAYER met4 ;
        RECT 9.755000 195.215000 10.075000 195.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 195.620000 10.075000 195.940000 ;
      LAYER met4 ;
        RECT 9.755000 195.620000 10.075000 195.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 196.025000 10.075000 196.345000 ;
      LAYER met4 ;
        RECT 9.755000 196.025000 10.075000 196.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 196.430000 10.075000 196.750000 ;
      LAYER met4 ;
        RECT 9.755000 196.430000 10.075000 196.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 196.835000 10.075000 197.155000 ;
      LAYER met4 ;
        RECT 9.755000 196.835000 10.075000 197.155000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 197.240000 10.075000 197.560000 ;
      LAYER met4 ;
        RECT 9.755000 197.240000 10.075000 197.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755000 197.645000 10.075000 197.965000 ;
      LAYER met4 ;
        RECT 9.755000 197.645000 10.075000 197.965000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.815000 173.900000 10.015000 174.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.815000 174.300000 10.015000 174.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.815000 174.700000 10.015000 174.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.815000 175.100000 10.015000 175.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.815000 175.500000 10.015000 175.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.815000 175.900000 10.015000 176.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.815000 176.300000 10.015000 176.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.815000 176.700000 10.015000 176.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.815000 177.100000 10.015000 177.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.815000 177.500000 10.015000 177.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.815000 177.900000 10.015000 178.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.815000 178.300000 10.015000 178.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.815000 178.700000 10.015000 178.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.815000 179.100000 10.015000 179.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.815000 179.500000 10.015000 179.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.815000 179.900000 10.015000 180.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.815000 180.300000 10.015000 180.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.815000 180.700000 10.015000 180.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.815000 181.100000 10.015000 181.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 23.850000 10.195000 24.170000 ;
      LAYER met4 ;
        RECT 9.875000 23.850000 10.195000 24.170000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 24.280000 10.195000 24.600000 ;
      LAYER met4 ;
        RECT 9.875000 24.280000 10.195000 24.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 24.710000 10.195000 25.030000 ;
      LAYER met4 ;
        RECT 9.875000 24.710000 10.195000 25.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 25.140000 10.195000 25.460000 ;
      LAYER met4 ;
        RECT 9.875000 25.140000 10.195000 25.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 25.570000 10.195000 25.890000 ;
      LAYER met4 ;
        RECT 9.875000 25.570000 10.195000 25.890000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 26.000000 10.195000 26.320000 ;
      LAYER met4 ;
        RECT 9.875000 26.000000 10.195000 26.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 26.430000 10.195000 26.750000 ;
      LAYER met4 ;
        RECT 9.875000 26.430000 10.195000 26.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 26.860000 10.195000 27.180000 ;
      LAYER met4 ;
        RECT 9.875000 26.860000 10.195000 27.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 27.290000 10.195000 27.610000 ;
      LAYER met4 ;
        RECT 9.875000 27.290000 10.195000 27.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 27.720000 10.195000 28.040000 ;
      LAYER met4 ;
        RECT 9.875000 27.720000 10.195000 28.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 28.150000 10.195000 28.470000 ;
      LAYER met4 ;
        RECT 9.875000 28.150000 10.195000 28.470000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.530000 56.250000 0.850000 56.570000 ;
      LAYER met4 ;
        RECT 0.530000 56.250000 0.850000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 56.660000 0.850000 56.980000 ;
      LAYER met4 ;
        RECT 0.530000 56.660000 0.850000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 57.070000 0.850000 57.390000 ;
      LAYER met4 ;
        RECT 0.530000 57.070000 0.850000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 57.480000 0.850000 57.800000 ;
      LAYER met4 ;
        RECT 0.530000 57.480000 0.850000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 57.890000 0.850000 58.210000 ;
      LAYER met4 ;
        RECT 0.530000 57.890000 0.850000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 58.300000 0.850000 58.620000 ;
      LAYER met4 ;
        RECT 0.530000 58.300000 0.850000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 58.710000 0.850000 59.030000 ;
      LAYER met4 ;
        RECT 0.530000 58.710000 0.850000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 59.120000 0.850000 59.440000 ;
      LAYER met4 ;
        RECT 0.530000 59.120000 0.850000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 59.530000 0.850000 59.850000 ;
      LAYER met4 ;
        RECT 0.530000 59.530000 0.850000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 59.940000 0.850000 60.260000 ;
      LAYER met4 ;
        RECT 0.530000 59.940000 0.850000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 60.350000 0.850000 60.670000 ;
      LAYER met4 ;
        RECT 0.530000 60.350000 0.850000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 56.250000 1.260000 56.570000 ;
      LAYER met4 ;
        RECT 0.940000 56.250000 1.260000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 56.660000 1.260000 56.980000 ;
      LAYER met4 ;
        RECT 0.940000 56.660000 1.260000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 57.070000 1.260000 57.390000 ;
      LAYER met4 ;
        RECT 0.940000 57.070000 1.260000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 57.480000 1.260000 57.800000 ;
      LAYER met4 ;
        RECT 0.940000 57.480000 1.260000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 57.890000 1.260000 58.210000 ;
      LAYER met4 ;
        RECT 0.940000 57.890000 1.260000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 58.300000 1.260000 58.620000 ;
      LAYER met4 ;
        RECT 0.940000 58.300000 1.260000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 58.710000 1.260000 59.030000 ;
      LAYER met4 ;
        RECT 0.940000 58.710000 1.260000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 59.120000 1.260000 59.440000 ;
      LAYER met4 ;
        RECT 0.940000 59.120000 1.260000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 59.530000 1.260000 59.850000 ;
      LAYER met4 ;
        RECT 0.940000 59.530000 1.260000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 59.940000 1.260000 60.260000 ;
      LAYER met4 ;
        RECT 0.940000 59.940000 1.260000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 60.350000 1.260000 60.670000 ;
      LAYER met4 ;
        RECT 0.940000 60.350000 1.260000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 56.250000 1.670000 56.570000 ;
      LAYER met4 ;
        RECT 1.350000 56.250000 1.670000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 56.660000 1.670000 56.980000 ;
      LAYER met4 ;
        RECT 1.350000 56.660000 1.670000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 57.070000 1.670000 57.390000 ;
      LAYER met4 ;
        RECT 1.350000 57.070000 1.670000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 57.480000 1.670000 57.800000 ;
      LAYER met4 ;
        RECT 1.350000 57.480000 1.670000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 57.890000 1.670000 58.210000 ;
      LAYER met4 ;
        RECT 1.350000 57.890000 1.670000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 58.300000 1.670000 58.620000 ;
      LAYER met4 ;
        RECT 1.350000 58.300000 1.670000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 58.710000 1.670000 59.030000 ;
      LAYER met4 ;
        RECT 1.350000 58.710000 1.670000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 59.120000 1.670000 59.440000 ;
      LAYER met4 ;
        RECT 1.350000 59.120000 1.670000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 59.530000 1.670000 59.850000 ;
      LAYER met4 ;
        RECT 1.350000 59.530000 1.670000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 59.940000 1.670000 60.260000 ;
      LAYER met4 ;
        RECT 1.350000 59.940000 1.670000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 60.350000 1.670000 60.670000 ;
      LAYER met4 ;
        RECT 1.350000 60.350000 1.670000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 56.250000 2.080000 56.570000 ;
      LAYER met4 ;
        RECT 1.760000 56.250000 2.080000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 56.660000 2.080000 56.980000 ;
      LAYER met4 ;
        RECT 1.760000 56.660000 2.080000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 57.070000 2.080000 57.390000 ;
      LAYER met4 ;
        RECT 1.760000 57.070000 2.080000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 57.480000 2.080000 57.800000 ;
      LAYER met4 ;
        RECT 1.760000 57.480000 2.080000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 57.890000 2.080000 58.210000 ;
      LAYER met4 ;
        RECT 1.760000 57.890000 2.080000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 58.300000 2.080000 58.620000 ;
      LAYER met4 ;
        RECT 1.760000 58.300000 2.080000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 58.710000 2.080000 59.030000 ;
      LAYER met4 ;
        RECT 1.760000 58.710000 2.080000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 59.120000 2.080000 59.440000 ;
      LAYER met4 ;
        RECT 1.760000 59.120000 2.080000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 59.530000 2.080000 59.850000 ;
      LAYER met4 ;
        RECT 1.760000 59.530000 2.080000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 59.940000 2.080000 60.260000 ;
      LAYER met4 ;
        RECT 1.760000 59.940000 2.080000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 60.350000 2.080000 60.670000 ;
      LAYER met4 ;
        RECT 1.760000 60.350000 2.080000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 56.250000 10.600000 56.570000 ;
      LAYER met4 ;
        RECT 10.280000 56.250000 10.600000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 56.660000 10.600000 56.980000 ;
      LAYER met4 ;
        RECT 10.280000 56.660000 10.600000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 57.070000 10.600000 57.390000 ;
      LAYER met4 ;
        RECT 10.280000 57.070000 10.600000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 57.480000 10.600000 57.800000 ;
      LAYER met4 ;
        RECT 10.280000 57.480000 10.600000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 57.890000 10.600000 58.210000 ;
      LAYER met4 ;
        RECT 10.280000 57.890000 10.600000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 58.300000 10.600000 58.620000 ;
      LAYER met4 ;
        RECT 10.280000 58.300000 10.600000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 58.710000 10.600000 59.030000 ;
      LAYER met4 ;
        RECT 10.280000 58.710000 10.600000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 59.120000 10.600000 59.440000 ;
      LAYER met4 ;
        RECT 10.280000 59.120000 10.600000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 59.530000 10.600000 59.850000 ;
      LAYER met4 ;
        RECT 10.280000 59.530000 10.600000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 59.940000 10.600000 60.260000 ;
      LAYER met4 ;
        RECT 10.280000 59.940000 10.600000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 60.350000 10.600000 60.670000 ;
      LAYER met4 ;
        RECT 10.280000 60.350000 10.600000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 56.250000 11.005000 56.570000 ;
      LAYER met4 ;
        RECT 10.685000 56.250000 11.005000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 56.660000 11.005000 56.980000 ;
      LAYER met4 ;
        RECT 10.685000 56.660000 11.005000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 57.070000 11.005000 57.390000 ;
      LAYER met4 ;
        RECT 10.685000 57.070000 11.005000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 57.480000 11.005000 57.800000 ;
      LAYER met4 ;
        RECT 10.685000 57.480000 11.005000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 57.890000 11.005000 58.210000 ;
      LAYER met4 ;
        RECT 10.685000 57.890000 11.005000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 58.300000 11.005000 58.620000 ;
      LAYER met4 ;
        RECT 10.685000 58.300000 11.005000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 58.710000 11.005000 59.030000 ;
      LAYER met4 ;
        RECT 10.685000 58.710000 11.005000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 59.120000 11.005000 59.440000 ;
      LAYER met4 ;
        RECT 10.685000 59.120000 11.005000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 59.530000 11.005000 59.850000 ;
      LAYER met4 ;
        RECT 10.685000 59.530000 11.005000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 59.940000 11.005000 60.260000 ;
      LAYER met4 ;
        RECT 10.685000 59.940000 11.005000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 60.350000 11.005000 60.670000 ;
      LAYER met4 ;
        RECT 10.685000 60.350000 11.005000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 56.250000 11.410000 56.570000 ;
      LAYER met4 ;
        RECT 11.090000 56.250000 11.410000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 56.660000 11.410000 56.980000 ;
      LAYER met4 ;
        RECT 11.090000 56.660000 11.410000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 57.070000 11.410000 57.390000 ;
      LAYER met4 ;
        RECT 11.090000 57.070000 11.410000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 57.480000 11.410000 57.800000 ;
      LAYER met4 ;
        RECT 11.090000 57.480000 11.410000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 57.890000 11.410000 58.210000 ;
      LAYER met4 ;
        RECT 11.090000 57.890000 11.410000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 58.300000 11.410000 58.620000 ;
      LAYER met4 ;
        RECT 11.090000 58.300000 11.410000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 58.710000 11.410000 59.030000 ;
      LAYER met4 ;
        RECT 11.090000 58.710000 11.410000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 59.120000 11.410000 59.440000 ;
      LAYER met4 ;
        RECT 11.090000 59.120000 11.410000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 59.530000 11.410000 59.850000 ;
      LAYER met4 ;
        RECT 11.090000 59.530000 11.410000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 59.940000 11.410000 60.260000 ;
      LAYER met4 ;
        RECT 11.090000 59.940000 11.410000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 60.350000 11.410000 60.670000 ;
      LAYER met4 ;
        RECT 11.090000 60.350000 11.410000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 56.250000 11.815000 56.570000 ;
      LAYER met4 ;
        RECT 11.495000 56.250000 11.815000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 56.660000 11.815000 56.980000 ;
      LAYER met4 ;
        RECT 11.495000 56.660000 11.815000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 57.070000 11.815000 57.390000 ;
      LAYER met4 ;
        RECT 11.495000 57.070000 11.815000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 57.480000 11.815000 57.800000 ;
      LAYER met4 ;
        RECT 11.495000 57.480000 11.815000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 57.890000 11.815000 58.210000 ;
      LAYER met4 ;
        RECT 11.495000 57.890000 11.815000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 58.300000 11.815000 58.620000 ;
      LAYER met4 ;
        RECT 11.495000 58.300000 11.815000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 58.710000 11.815000 59.030000 ;
      LAYER met4 ;
        RECT 11.495000 58.710000 11.815000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 59.120000 11.815000 59.440000 ;
      LAYER met4 ;
        RECT 11.495000 59.120000 11.815000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 59.530000 11.815000 59.850000 ;
      LAYER met4 ;
        RECT 11.495000 59.530000 11.815000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 59.940000 11.815000 60.260000 ;
      LAYER met4 ;
        RECT 11.495000 59.940000 11.815000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 60.350000 11.815000 60.670000 ;
      LAYER met4 ;
        RECT 11.495000 60.350000 11.815000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 56.250000 12.220000 56.570000 ;
      LAYER met4 ;
        RECT 11.900000 56.250000 12.220000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 56.660000 12.220000 56.980000 ;
      LAYER met4 ;
        RECT 11.900000 56.660000 12.220000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 57.070000 12.220000 57.390000 ;
      LAYER met4 ;
        RECT 11.900000 57.070000 12.220000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 57.480000 12.220000 57.800000 ;
      LAYER met4 ;
        RECT 11.900000 57.480000 12.220000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 57.890000 12.220000 58.210000 ;
      LAYER met4 ;
        RECT 11.900000 57.890000 12.220000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 58.300000 12.220000 58.620000 ;
      LAYER met4 ;
        RECT 11.900000 58.300000 12.220000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 58.710000 12.220000 59.030000 ;
      LAYER met4 ;
        RECT 11.900000 58.710000 12.220000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 59.120000 12.220000 59.440000 ;
      LAYER met4 ;
        RECT 11.900000 59.120000 12.220000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 59.530000 12.220000 59.850000 ;
      LAYER met4 ;
        RECT 11.900000 59.530000 12.220000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 59.940000 12.220000 60.260000 ;
      LAYER met4 ;
        RECT 11.900000 59.940000 12.220000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 60.350000 12.220000 60.670000 ;
      LAYER met4 ;
        RECT 11.900000 60.350000 12.220000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 56.250000 12.625000 56.570000 ;
      LAYER met4 ;
        RECT 12.305000 56.250000 12.625000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 56.660000 12.625000 56.980000 ;
      LAYER met4 ;
        RECT 12.305000 56.660000 12.625000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 57.070000 12.625000 57.390000 ;
      LAYER met4 ;
        RECT 12.305000 57.070000 12.625000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 57.480000 12.625000 57.800000 ;
      LAYER met4 ;
        RECT 12.305000 57.480000 12.625000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 57.890000 12.625000 58.210000 ;
      LAYER met4 ;
        RECT 12.305000 57.890000 12.625000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 58.300000 12.625000 58.620000 ;
      LAYER met4 ;
        RECT 12.305000 58.300000 12.625000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 58.710000 12.625000 59.030000 ;
      LAYER met4 ;
        RECT 12.305000 58.710000 12.625000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 59.120000 12.625000 59.440000 ;
      LAYER met4 ;
        RECT 12.305000 59.120000 12.625000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 59.530000 12.625000 59.850000 ;
      LAYER met4 ;
        RECT 12.305000 59.530000 12.625000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 59.940000 12.625000 60.260000 ;
      LAYER met4 ;
        RECT 12.305000 59.940000 12.625000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 60.350000 12.625000 60.670000 ;
      LAYER met4 ;
        RECT 12.305000 60.350000 12.625000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 56.250000 13.030000 56.570000 ;
      LAYER met4 ;
        RECT 12.710000 56.250000 13.030000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 56.660000 13.030000 56.980000 ;
      LAYER met4 ;
        RECT 12.710000 56.660000 13.030000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 57.070000 13.030000 57.390000 ;
      LAYER met4 ;
        RECT 12.710000 57.070000 13.030000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 57.480000 13.030000 57.800000 ;
      LAYER met4 ;
        RECT 12.710000 57.480000 13.030000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 57.890000 13.030000 58.210000 ;
      LAYER met4 ;
        RECT 12.710000 57.890000 13.030000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 58.300000 13.030000 58.620000 ;
      LAYER met4 ;
        RECT 12.710000 58.300000 13.030000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 58.710000 13.030000 59.030000 ;
      LAYER met4 ;
        RECT 12.710000 58.710000 13.030000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 59.120000 13.030000 59.440000 ;
      LAYER met4 ;
        RECT 12.710000 59.120000 13.030000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 59.530000 13.030000 59.850000 ;
      LAYER met4 ;
        RECT 12.710000 59.530000 13.030000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 59.940000 13.030000 60.260000 ;
      LAYER met4 ;
        RECT 12.710000 59.940000 13.030000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 60.350000 13.030000 60.670000 ;
      LAYER met4 ;
        RECT 12.710000 60.350000 13.030000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 56.250000 13.435000 56.570000 ;
      LAYER met4 ;
        RECT 13.115000 56.250000 13.435000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 56.660000 13.435000 56.980000 ;
      LAYER met4 ;
        RECT 13.115000 56.660000 13.435000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 57.070000 13.435000 57.390000 ;
      LAYER met4 ;
        RECT 13.115000 57.070000 13.435000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 57.480000 13.435000 57.800000 ;
      LAYER met4 ;
        RECT 13.115000 57.480000 13.435000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 57.890000 13.435000 58.210000 ;
      LAYER met4 ;
        RECT 13.115000 57.890000 13.435000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 58.300000 13.435000 58.620000 ;
      LAYER met4 ;
        RECT 13.115000 58.300000 13.435000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 58.710000 13.435000 59.030000 ;
      LAYER met4 ;
        RECT 13.115000 58.710000 13.435000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 59.120000 13.435000 59.440000 ;
      LAYER met4 ;
        RECT 13.115000 59.120000 13.435000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 59.530000 13.435000 59.850000 ;
      LAYER met4 ;
        RECT 13.115000 59.530000 13.435000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 59.940000 13.435000 60.260000 ;
      LAYER met4 ;
        RECT 13.115000 59.940000 13.435000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 60.350000 13.435000 60.670000 ;
      LAYER met4 ;
        RECT 13.115000 60.350000 13.435000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 56.250000 13.840000 56.570000 ;
      LAYER met4 ;
        RECT 13.520000 56.250000 13.840000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 56.660000 13.840000 56.980000 ;
      LAYER met4 ;
        RECT 13.520000 56.660000 13.840000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 57.070000 13.840000 57.390000 ;
      LAYER met4 ;
        RECT 13.520000 57.070000 13.840000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 57.480000 13.840000 57.800000 ;
      LAYER met4 ;
        RECT 13.520000 57.480000 13.840000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 57.890000 13.840000 58.210000 ;
      LAYER met4 ;
        RECT 13.520000 57.890000 13.840000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 58.300000 13.840000 58.620000 ;
      LAYER met4 ;
        RECT 13.520000 58.300000 13.840000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 58.710000 13.840000 59.030000 ;
      LAYER met4 ;
        RECT 13.520000 58.710000 13.840000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 59.120000 13.840000 59.440000 ;
      LAYER met4 ;
        RECT 13.520000 59.120000 13.840000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 59.530000 13.840000 59.850000 ;
      LAYER met4 ;
        RECT 13.520000 59.530000 13.840000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 59.940000 13.840000 60.260000 ;
      LAYER met4 ;
        RECT 13.520000 59.940000 13.840000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 60.350000 13.840000 60.670000 ;
      LAYER met4 ;
        RECT 13.520000 60.350000 13.840000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 56.250000 14.245000 56.570000 ;
      LAYER met4 ;
        RECT 13.925000 56.250000 14.245000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 56.660000 14.245000 56.980000 ;
      LAYER met4 ;
        RECT 13.925000 56.660000 14.245000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 57.070000 14.245000 57.390000 ;
      LAYER met4 ;
        RECT 13.925000 57.070000 14.245000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 57.480000 14.245000 57.800000 ;
      LAYER met4 ;
        RECT 13.925000 57.480000 14.245000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 57.890000 14.245000 58.210000 ;
      LAYER met4 ;
        RECT 13.925000 57.890000 14.245000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 58.300000 14.245000 58.620000 ;
      LAYER met4 ;
        RECT 13.925000 58.300000 14.245000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 58.710000 14.245000 59.030000 ;
      LAYER met4 ;
        RECT 13.925000 58.710000 14.245000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 59.120000 14.245000 59.440000 ;
      LAYER met4 ;
        RECT 13.925000 59.120000 14.245000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 59.530000 14.245000 59.850000 ;
      LAYER met4 ;
        RECT 13.925000 59.530000 14.245000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 59.940000 14.245000 60.260000 ;
      LAYER met4 ;
        RECT 13.925000 59.940000 14.245000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 60.350000 14.245000 60.670000 ;
      LAYER met4 ;
        RECT 13.925000 60.350000 14.245000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 56.250000 14.650000 56.570000 ;
      LAYER met4 ;
        RECT 14.330000 56.250000 14.650000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 56.660000 14.650000 56.980000 ;
      LAYER met4 ;
        RECT 14.330000 56.660000 14.650000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 57.070000 14.650000 57.390000 ;
      LAYER met4 ;
        RECT 14.330000 57.070000 14.650000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 57.480000 14.650000 57.800000 ;
      LAYER met4 ;
        RECT 14.330000 57.480000 14.650000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 57.890000 14.650000 58.210000 ;
      LAYER met4 ;
        RECT 14.330000 57.890000 14.650000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 58.300000 14.650000 58.620000 ;
      LAYER met4 ;
        RECT 14.330000 58.300000 14.650000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 58.710000 14.650000 59.030000 ;
      LAYER met4 ;
        RECT 14.330000 58.710000 14.650000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 59.120000 14.650000 59.440000 ;
      LAYER met4 ;
        RECT 14.330000 59.120000 14.650000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 59.530000 14.650000 59.850000 ;
      LAYER met4 ;
        RECT 14.330000 59.530000 14.650000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 59.940000 14.650000 60.260000 ;
      LAYER met4 ;
        RECT 14.330000 59.940000 14.650000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 60.350000 14.650000 60.670000 ;
      LAYER met4 ;
        RECT 14.330000 60.350000 14.650000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 56.250000 15.055000 56.570000 ;
      LAYER met4 ;
        RECT 14.735000 56.250000 15.055000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 56.660000 15.055000 56.980000 ;
      LAYER met4 ;
        RECT 14.735000 56.660000 15.055000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 57.070000 15.055000 57.390000 ;
      LAYER met4 ;
        RECT 14.735000 57.070000 15.055000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 57.480000 15.055000 57.800000 ;
      LAYER met4 ;
        RECT 14.735000 57.480000 15.055000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 57.890000 15.055000 58.210000 ;
      LAYER met4 ;
        RECT 14.735000 57.890000 15.055000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 58.300000 15.055000 58.620000 ;
      LAYER met4 ;
        RECT 14.735000 58.300000 15.055000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 58.710000 15.055000 59.030000 ;
      LAYER met4 ;
        RECT 14.735000 58.710000 15.055000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 59.120000 15.055000 59.440000 ;
      LAYER met4 ;
        RECT 14.735000 59.120000 15.055000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 59.530000 15.055000 59.850000 ;
      LAYER met4 ;
        RECT 14.735000 59.530000 15.055000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 59.940000 15.055000 60.260000 ;
      LAYER met4 ;
        RECT 14.735000 59.940000 15.055000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 60.350000 15.055000 60.670000 ;
      LAYER met4 ;
        RECT 14.735000 60.350000 15.055000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 56.250000 15.460000 56.570000 ;
      LAYER met4 ;
        RECT 15.140000 56.250000 15.460000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 56.660000 15.460000 56.980000 ;
      LAYER met4 ;
        RECT 15.140000 56.660000 15.460000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 57.070000 15.460000 57.390000 ;
      LAYER met4 ;
        RECT 15.140000 57.070000 15.460000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 57.480000 15.460000 57.800000 ;
      LAYER met4 ;
        RECT 15.140000 57.480000 15.460000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 57.890000 15.460000 58.210000 ;
      LAYER met4 ;
        RECT 15.140000 57.890000 15.460000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 58.300000 15.460000 58.620000 ;
      LAYER met4 ;
        RECT 15.140000 58.300000 15.460000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 58.710000 15.460000 59.030000 ;
      LAYER met4 ;
        RECT 15.140000 58.710000 15.460000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 59.120000 15.460000 59.440000 ;
      LAYER met4 ;
        RECT 15.140000 59.120000 15.460000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 59.530000 15.460000 59.850000 ;
      LAYER met4 ;
        RECT 15.140000 59.530000 15.460000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 59.940000 15.460000 60.260000 ;
      LAYER met4 ;
        RECT 15.140000 59.940000 15.460000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 60.350000 15.460000 60.670000 ;
      LAYER met4 ;
        RECT 15.140000 60.350000 15.460000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 56.250000 15.865000 56.570000 ;
      LAYER met4 ;
        RECT 15.545000 56.250000 15.865000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 56.660000 15.865000 56.980000 ;
      LAYER met4 ;
        RECT 15.545000 56.660000 15.865000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 57.070000 15.865000 57.390000 ;
      LAYER met4 ;
        RECT 15.545000 57.070000 15.865000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 57.480000 15.865000 57.800000 ;
      LAYER met4 ;
        RECT 15.545000 57.480000 15.865000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 57.890000 15.865000 58.210000 ;
      LAYER met4 ;
        RECT 15.545000 57.890000 15.865000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 58.300000 15.865000 58.620000 ;
      LAYER met4 ;
        RECT 15.545000 58.300000 15.865000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 58.710000 15.865000 59.030000 ;
      LAYER met4 ;
        RECT 15.545000 58.710000 15.865000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 59.120000 15.865000 59.440000 ;
      LAYER met4 ;
        RECT 15.545000 59.120000 15.865000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 59.530000 15.865000 59.850000 ;
      LAYER met4 ;
        RECT 15.545000 59.530000 15.865000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 59.940000 15.865000 60.260000 ;
      LAYER met4 ;
        RECT 15.545000 59.940000 15.865000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 60.350000 15.865000 60.670000 ;
      LAYER met4 ;
        RECT 15.545000 60.350000 15.865000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 56.250000 16.270000 56.570000 ;
      LAYER met4 ;
        RECT 15.950000 56.250000 16.270000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 56.660000 16.270000 56.980000 ;
      LAYER met4 ;
        RECT 15.950000 56.660000 16.270000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 57.070000 16.270000 57.390000 ;
      LAYER met4 ;
        RECT 15.950000 57.070000 16.270000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 57.480000 16.270000 57.800000 ;
      LAYER met4 ;
        RECT 15.950000 57.480000 16.270000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 57.890000 16.270000 58.210000 ;
      LAYER met4 ;
        RECT 15.950000 57.890000 16.270000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 58.300000 16.270000 58.620000 ;
      LAYER met4 ;
        RECT 15.950000 58.300000 16.270000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 58.710000 16.270000 59.030000 ;
      LAYER met4 ;
        RECT 15.950000 58.710000 16.270000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 59.120000 16.270000 59.440000 ;
      LAYER met4 ;
        RECT 15.950000 59.120000 16.270000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 59.530000 16.270000 59.850000 ;
      LAYER met4 ;
        RECT 15.950000 59.530000 16.270000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 59.940000 16.270000 60.260000 ;
      LAYER met4 ;
        RECT 15.950000 59.940000 16.270000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 60.350000 16.270000 60.670000 ;
      LAYER met4 ;
        RECT 15.950000 60.350000 16.270000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 56.250000 16.675000 56.570000 ;
      LAYER met4 ;
        RECT 16.355000 56.250000 16.675000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 56.660000 16.675000 56.980000 ;
      LAYER met4 ;
        RECT 16.355000 56.660000 16.675000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 57.070000 16.675000 57.390000 ;
      LAYER met4 ;
        RECT 16.355000 57.070000 16.675000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 57.480000 16.675000 57.800000 ;
      LAYER met4 ;
        RECT 16.355000 57.480000 16.675000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 57.890000 16.675000 58.210000 ;
      LAYER met4 ;
        RECT 16.355000 57.890000 16.675000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 58.300000 16.675000 58.620000 ;
      LAYER met4 ;
        RECT 16.355000 58.300000 16.675000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 58.710000 16.675000 59.030000 ;
      LAYER met4 ;
        RECT 16.355000 58.710000 16.675000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 59.120000 16.675000 59.440000 ;
      LAYER met4 ;
        RECT 16.355000 59.120000 16.675000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 59.530000 16.675000 59.850000 ;
      LAYER met4 ;
        RECT 16.355000 59.530000 16.675000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 59.940000 16.675000 60.260000 ;
      LAYER met4 ;
        RECT 16.355000 59.940000 16.675000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 60.350000 16.675000 60.670000 ;
      LAYER met4 ;
        RECT 16.355000 60.350000 16.675000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 56.250000 17.080000 56.570000 ;
      LAYER met4 ;
        RECT 16.760000 56.250000 17.080000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 56.660000 17.080000 56.980000 ;
      LAYER met4 ;
        RECT 16.760000 56.660000 17.080000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 57.070000 17.080000 57.390000 ;
      LAYER met4 ;
        RECT 16.760000 57.070000 17.080000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 57.480000 17.080000 57.800000 ;
      LAYER met4 ;
        RECT 16.760000 57.480000 17.080000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 57.890000 17.080000 58.210000 ;
      LAYER met4 ;
        RECT 16.760000 57.890000 17.080000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 58.300000 17.080000 58.620000 ;
      LAYER met4 ;
        RECT 16.760000 58.300000 17.080000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 58.710000 17.080000 59.030000 ;
      LAYER met4 ;
        RECT 16.760000 58.710000 17.080000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 59.120000 17.080000 59.440000 ;
      LAYER met4 ;
        RECT 16.760000 59.120000 17.080000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 59.530000 17.080000 59.850000 ;
      LAYER met4 ;
        RECT 16.760000 59.530000 17.080000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 59.940000 17.080000 60.260000 ;
      LAYER met4 ;
        RECT 16.760000 59.940000 17.080000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 60.350000 17.080000 60.670000 ;
      LAYER met4 ;
        RECT 16.760000 60.350000 17.080000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 56.250000 17.485000 56.570000 ;
      LAYER met4 ;
        RECT 17.165000 56.250000 17.485000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 56.660000 17.485000 56.980000 ;
      LAYER met4 ;
        RECT 17.165000 56.660000 17.485000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 57.070000 17.485000 57.390000 ;
      LAYER met4 ;
        RECT 17.165000 57.070000 17.485000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 57.480000 17.485000 57.800000 ;
      LAYER met4 ;
        RECT 17.165000 57.480000 17.485000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 57.890000 17.485000 58.210000 ;
      LAYER met4 ;
        RECT 17.165000 57.890000 17.485000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 58.300000 17.485000 58.620000 ;
      LAYER met4 ;
        RECT 17.165000 58.300000 17.485000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 58.710000 17.485000 59.030000 ;
      LAYER met4 ;
        RECT 17.165000 58.710000 17.485000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 59.120000 17.485000 59.440000 ;
      LAYER met4 ;
        RECT 17.165000 59.120000 17.485000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 59.530000 17.485000 59.850000 ;
      LAYER met4 ;
        RECT 17.165000 59.530000 17.485000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 59.940000 17.485000 60.260000 ;
      LAYER met4 ;
        RECT 17.165000 59.940000 17.485000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 60.350000 17.485000 60.670000 ;
      LAYER met4 ;
        RECT 17.165000 60.350000 17.485000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 56.250000 17.890000 56.570000 ;
      LAYER met4 ;
        RECT 17.570000 56.250000 17.890000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 56.660000 17.890000 56.980000 ;
      LAYER met4 ;
        RECT 17.570000 56.660000 17.890000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 57.070000 17.890000 57.390000 ;
      LAYER met4 ;
        RECT 17.570000 57.070000 17.890000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 57.480000 17.890000 57.800000 ;
      LAYER met4 ;
        RECT 17.570000 57.480000 17.890000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 57.890000 17.890000 58.210000 ;
      LAYER met4 ;
        RECT 17.570000 57.890000 17.890000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 58.300000 17.890000 58.620000 ;
      LAYER met4 ;
        RECT 17.570000 58.300000 17.890000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 58.710000 17.890000 59.030000 ;
      LAYER met4 ;
        RECT 17.570000 58.710000 17.890000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 59.120000 17.890000 59.440000 ;
      LAYER met4 ;
        RECT 17.570000 59.120000 17.890000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 59.530000 17.890000 59.850000 ;
      LAYER met4 ;
        RECT 17.570000 59.530000 17.890000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 59.940000 17.890000 60.260000 ;
      LAYER met4 ;
        RECT 17.570000 59.940000 17.890000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 60.350000 17.890000 60.670000 ;
      LAYER met4 ;
        RECT 17.570000 60.350000 17.890000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 56.250000 18.295000 56.570000 ;
      LAYER met4 ;
        RECT 17.975000 56.250000 18.295000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 56.660000 18.295000 56.980000 ;
      LAYER met4 ;
        RECT 17.975000 56.660000 18.295000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 57.070000 18.295000 57.390000 ;
      LAYER met4 ;
        RECT 17.975000 57.070000 18.295000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 57.480000 18.295000 57.800000 ;
      LAYER met4 ;
        RECT 17.975000 57.480000 18.295000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 57.890000 18.295000 58.210000 ;
      LAYER met4 ;
        RECT 17.975000 57.890000 18.295000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 58.300000 18.295000 58.620000 ;
      LAYER met4 ;
        RECT 17.975000 58.300000 18.295000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 58.710000 18.295000 59.030000 ;
      LAYER met4 ;
        RECT 17.975000 58.710000 18.295000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 59.120000 18.295000 59.440000 ;
      LAYER met4 ;
        RECT 17.975000 59.120000 18.295000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 59.530000 18.295000 59.850000 ;
      LAYER met4 ;
        RECT 17.975000 59.530000 18.295000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 59.940000 18.295000 60.260000 ;
      LAYER met4 ;
        RECT 17.975000 59.940000 18.295000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 60.350000 18.295000 60.670000 ;
      LAYER met4 ;
        RECT 17.975000 60.350000 18.295000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 56.250000 18.700000 56.570000 ;
      LAYER met4 ;
        RECT 18.380000 56.250000 18.700000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 56.660000 18.700000 56.980000 ;
      LAYER met4 ;
        RECT 18.380000 56.660000 18.700000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 57.070000 18.700000 57.390000 ;
      LAYER met4 ;
        RECT 18.380000 57.070000 18.700000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 57.480000 18.700000 57.800000 ;
      LAYER met4 ;
        RECT 18.380000 57.480000 18.700000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 57.890000 18.700000 58.210000 ;
      LAYER met4 ;
        RECT 18.380000 57.890000 18.700000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 58.300000 18.700000 58.620000 ;
      LAYER met4 ;
        RECT 18.380000 58.300000 18.700000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 58.710000 18.700000 59.030000 ;
      LAYER met4 ;
        RECT 18.380000 58.710000 18.700000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 59.120000 18.700000 59.440000 ;
      LAYER met4 ;
        RECT 18.380000 59.120000 18.700000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 59.530000 18.700000 59.850000 ;
      LAYER met4 ;
        RECT 18.380000 59.530000 18.700000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 59.940000 18.700000 60.260000 ;
      LAYER met4 ;
        RECT 18.380000 59.940000 18.700000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 60.350000 18.700000 60.670000 ;
      LAYER met4 ;
        RECT 18.380000 60.350000 18.700000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 56.250000 19.105000 56.570000 ;
      LAYER met4 ;
        RECT 18.785000 56.250000 19.105000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 56.660000 19.105000 56.980000 ;
      LAYER met4 ;
        RECT 18.785000 56.660000 19.105000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 57.070000 19.105000 57.390000 ;
      LAYER met4 ;
        RECT 18.785000 57.070000 19.105000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 57.480000 19.105000 57.800000 ;
      LAYER met4 ;
        RECT 18.785000 57.480000 19.105000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 57.890000 19.105000 58.210000 ;
      LAYER met4 ;
        RECT 18.785000 57.890000 19.105000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 58.300000 19.105000 58.620000 ;
      LAYER met4 ;
        RECT 18.785000 58.300000 19.105000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 58.710000 19.105000 59.030000 ;
      LAYER met4 ;
        RECT 18.785000 58.710000 19.105000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 59.120000 19.105000 59.440000 ;
      LAYER met4 ;
        RECT 18.785000 59.120000 19.105000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 59.530000 19.105000 59.850000 ;
      LAYER met4 ;
        RECT 18.785000 59.530000 19.105000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 59.940000 19.105000 60.260000 ;
      LAYER met4 ;
        RECT 18.785000 59.940000 19.105000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 60.350000 19.105000 60.670000 ;
      LAYER met4 ;
        RECT 18.785000 60.350000 19.105000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 56.250000 19.510000 56.570000 ;
      LAYER met4 ;
        RECT 19.190000 56.250000 19.510000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 56.660000 19.510000 56.980000 ;
      LAYER met4 ;
        RECT 19.190000 56.660000 19.510000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 57.070000 19.510000 57.390000 ;
      LAYER met4 ;
        RECT 19.190000 57.070000 19.510000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 57.480000 19.510000 57.800000 ;
      LAYER met4 ;
        RECT 19.190000 57.480000 19.510000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 57.890000 19.510000 58.210000 ;
      LAYER met4 ;
        RECT 19.190000 57.890000 19.510000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 58.300000 19.510000 58.620000 ;
      LAYER met4 ;
        RECT 19.190000 58.300000 19.510000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 58.710000 19.510000 59.030000 ;
      LAYER met4 ;
        RECT 19.190000 58.710000 19.510000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 59.120000 19.510000 59.440000 ;
      LAYER met4 ;
        RECT 19.190000 59.120000 19.510000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 59.530000 19.510000 59.850000 ;
      LAYER met4 ;
        RECT 19.190000 59.530000 19.510000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 59.940000 19.510000 60.260000 ;
      LAYER met4 ;
        RECT 19.190000 59.940000 19.510000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 60.350000 19.510000 60.670000 ;
      LAYER met4 ;
        RECT 19.190000 60.350000 19.510000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 56.250000 19.915000 56.570000 ;
      LAYER met4 ;
        RECT 19.595000 56.250000 19.915000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 56.660000 19.915000 56.980000 ;
      LAYER met4 ;
        RECT 19.595000 56.660000 19.915000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 57.070000 19.915000 57.390000 ;
      LAYER met4 ;
        RECT 19.595000 57.070000 19.915000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 57.480000 19.915000 57.800000 ;
      LAYER met4 ;
        RECT 19.595000 57.480000 19.915000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 57.890000 19.915000 58.210000 ;
      LAYER met4 ;
        RECT 19.595000 57.890000 19.915000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 58.300000 19.915000 58.620000 ;
      LAYER met4 ;
        RECT 19.595000 58.300000 19.915000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 58.710000 19.915000 59.030000 ;
      LAYER met4 ;
        RECT 19.595000 58.710000 19.915000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 59.120000 19.915000 59.440000 ;
      LAYER met4 ;
        RECT 19.595000 59.120000 19.915000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 59.530000 19.915000 59.850000 ;
      LAYER met4 ;
        RECT 19.595000 59.530000 19.915000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 59.940000 19.915000 60.260000 ;
      LAYER met4 ;
        RECT 19.595000 59.940000 19.915000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 60.350000 19.915000 60.670000 ;
      LAYER met4 ;
        RECT 19.595000 60.350000 19.915000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 56.250000 2.490000 56.570000 ;
      LAYER met4 ;
        RECT 2.170000 56.250000 2.490000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 56.660000 2.490000 56.980000 ;
      LAYER met4 ;
        RECT 2.170000 56.660000 2.490000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 57.070000 2.490000 57.390000 ;
      LAYER met4 ;
        RECT 2.170000 57.070000 2.490000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 57.480000 2.490000 57.800000 ;
      LAYER met4 ;
        RECT 2.170000 57.480000 2.490000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 57.890000 2.490000 58.210000 ;
      LAYER met4 ;
        RECT 2.170000 57.890000 2.490000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 58.300000 2.490000 58.620000 ;
      LAYER met4 ;
        RECT 2.170000 58.300000 2.490000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 58.710000 2.490000 59.030000 ;
      LAYER met4 ;
        RECT 2.170000 58.710000 2.490000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 59.120000 2.490000 59.440000 ;
      LAYER met4 ;
        RECT 2.170000 59.120000 2.490000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 59.530000 2.490000 59.850000 ;
      LAYER met4 ;
        RECT 2.170000 59.530000 2.490000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 59.940000 2.490000 60.260000 ;
      LAYER met4 ;
        RECT 2.170000 59.940000 2.490000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 60.350000 2.490000 60.670000 ;
      LAYER met4 ;
        RECT 2.170000 60.350000 2.490000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 56.250000 2.900000 56.570000 ;
      LAYER met4 ;
        RECT 2.580000 56.250000 2.900000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 56.660000 2.900000 56.980000 ;
      LAYER met4 ;
        RECT 2.580000 56.660000 2.900000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 57.070000 2.900000 57.390000 ;
      LAYER met4 ;
        RECT 2.580000 57.070000 2.900000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 57.480000 2.900000 57.800000 ;
      LAYER met4 ;
        RECT 2.580000 57.480000 2.900000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 57.890000 2.900000 58.210000 ;
      LAYER met4 ;
        RECT 2.580000 57.890000 2.900000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 58.300000 2.900000 58.620000 ;
      LAYER met4 ;
        RECT 2.580000 58.300000 2.900000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 58.710000 2.900000 59.030000 ;
      LAYER met4 ;
        RECT 2.580000 58.710000 2.900000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 59.120000 2.900000 59.440000 ;
      LAYER met4 ;
        RECT 2.580000 59.120000 2.900000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 59.530000 2.900000 59.850000 ;
      LAYER met4 ;
        RECT 2.580000 59.530000 2.900000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 59.940000 2.900000 60.260000 ;
      LAYER met4 ;
        RECT 2.580000 59.940000 2.900000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 60.350000 2.900000 60.670000 ;
      LAYER met4 ;
        RECT 2.580000 60.350000 2.900000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 56.250000 3.310000 56.570000 ;
      LAYER met4 ;
        RECT 2.990000 56.250000 3.310000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 56.660000 3.310000 56.980000 ;
      LAYER met4 ;
        RECT 2.990000 56.660000 3.310000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 57.070000 3.310000 57.390000 ;
      LAYER met4 ;
        RECT 2.990000 57.070000 3.310000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 57.480000 3.310000 57.800000 ;
      LAYER met4 ;
        RECT 2.990000 57.480000 3.310000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 57.890000 3.310000 58.210000 ;
      LAYER met4 ;
        RECT 2.990000 57.890000 3.310000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 58.300000 3.310000 58.620000 ;
      LAYER met4 ;
        RECT 2.990000 58.300000 3.310000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 58.710000 3.310000 59.030000 ;
      LAYER met4 ;
        RECT 2.990000 58.710000 3.310000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 59.120000 3.310000 59.440000 ;
      LAYER met4 ;
        RECT 2.990000 59.120000 3.310000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 59.530000 3.310000 59.850000 ;
      LAYER met4 ;
        RECT 2.990000 59.530000 3.310000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 59.940000 3.310000 60.260000 ;
      LAYER met4 ;
        RECT 2.990000 59.940000 3.310000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 60.350000 3.310000 60.670000 ;
      LAYER met4 ;
        RECT 2.990000 60.350000 3.310000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 56.250000 20.320000 56.570000 ;
      LAYER met4 ;
        RECT 20.000000 56.250000 20.320000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 56.660000 20.320000 56.980000 ;
      LAYER met4 ;
        RECT 20.000000 56.660000 20.320000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 57.070000 20.320000 57.390000 ;
      LAYER met4 ;
        RECT 20.000000 57.070000 20.320000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 57.480000 20.320000 57.800000 ;
      LAYER met4 ;
        RECT 20.000000 57.480000 20.320000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 57.890000 20.320000 58.210000 ;
      LAYER met4 ;
        RECT 20.000000 57.890000 20.320000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 58.300000 20.320000 58.620000 ;
      LAYER met4 ;
        RECT 20.000000 58.300000 20.320000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 58.710000 20.320000 59.030000 ;
      LAYER met4 ;
        RECT 20.000000 58.710000 20.320000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 59.120000 20.320000 59.440000 ;
      LAYER met4 ;
        RECT 20.000000 59.120000 20.320000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 59.530000 20.320000 59.850000 ;
      LAYER met4 ;
        RECT 20.000000 59.530000 20.320000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 59.940000 20.320000 60.260000 ;
      LAYER met4 ;
        RECT 20.000000 59.940000 20.320000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 60.350000 20.320000 60.670000 ;
      LAYER met4 ;
        RECT 20.000000 60.350000 20.320000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 56.250000 20.725000 56.570000 ;
      LAYER met4 ;
        RECT 20.405000 56.250000 20.725000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 56.660000 20.725000 56.980000 ;
      LAYER met4 ;
        RECT 20.405000 56.660000 20.725000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 57.070000 20.725000 57.390000 ;
      LAYER met4 ;
        RECT 20.405000 57.070000 20.725000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 57.480000 20.725000 57.800000 ;
      LAYER met4 ;
        RECT 20.405000 57.480000 20.725000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 57.890000 20.725000 58.210000 ;
      LAYER met4 ;
        RECT 20.405000 57.890000 20.725000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 58.300000 20.725000 58.620000 ;
      LAYER met4 ;
        RECT 20.405000 58.300000 20.725000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 58.710000 20.725000 59.030000 ;
      LAYER met4 ;
        RECT 20.405000 58.710000 20.725000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 59.120000 20.725000 59.440000 ;
      LAYER met4 ;
        RECT 20.405000 59.120000 20.725000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 59.530000 20.725000 59.850000 ;
      LAYER met4 ;
        RECT 20.405000 59.530000 20.725000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 59.940000 20.725000 60.260000 ;
      LAYER met4 ;
        RECT 20.405000 59.940000 20.725000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 60.350000 20.725000 60.670000 ;
      LAYER met4 ;
        RECT 20.405000 60.350000 20.725000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 56.250000 21.130000 56.570000 ;
      LAYER met4 ;
        RECT 20.810000 56.250000 21.130000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 56.660000 21.130000 56.980000 ;
      LAYER met4 ;
        RECT 20.810000 56.660000 21.130000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 57.070000 21.130000 57.390000 ;
      LAYER met4 ;
        RECT 20.810000 57.070000 21.130000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 57.480000 21.130000 57.800000 ;
      LAYER met4 ;
        RECT 20.810000 57.480000 21.130000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 57.890000 21.130000 58.210000 ;
      LAYER met4 ;
        RECT 20.810000 57.890000 21.130000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 58.300000 21.130000 58.620000 ;
      LAYER met4 ;
        RECT 20.810000 58.300000 21.130000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 58.710000 21.130000 59.030000 ;
      LAYER met4 ;
        RECT 20.810000 58.710000 21.130000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 59.120000 21.130000 59.440000 ;
      LAYER met4 ;
        RECT 20.810000 59.120000 21.130000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 59.530000 21.130000 59.850000 ;
      LAYER met4 ;
        RECT 20.810000 59.530000 21.130000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 59.940000 21.130000 60.260000 ;
      LAYER met4 ;
        RECT 20.810000 59.940000 21.130000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 60.350000 21.130000 60.670000 ;
      LAYER met4 ;
        RECT 20.810000 60.350000 21.130000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 56.250000 21.535000 56.570000 ;
      LAYER met4 ;
        RECT 21.215000 56.250000 21.535000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 56.660000 21.535000 56.980000 ;
      LAYER met4 ;
        RECT 21.215000 56.660000 21.535000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 57.070000 21.535000 57.390000 ;
      LAYER met4 ;
        RECT 21.215000 57.070000 21.535000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 57.480000 21.535000 57.800000 ;
      LAYER met4 ;
        RECT 21.215000 57.480000 21.535000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 57.890000 21.535000 58.210000 ;
      LAYER met4 ;
        RECT 21.215000 57.890000 21.535000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 58.300000 21.535000 58.620000 ;
      LAYER met4 ;
        RECT 21.215000 58.300000 21.535000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 58.710000 21.535000 59.030000 ;
      LAYER met4 ;
        RECT 21.215000 58.710000 21.535000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 59.120000 21.535000 59.440000 ;
      LAYER met4 ;
        RECT 21.215000 59.120000 21.535000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 59.530000 21.535000 59.850000 ;
      LAYER met4 ;
        RECT 21.215000 59.530000 21.535000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 59.940000 21.535000 60.260000 ;
      LAYER met4 ;
        RECT 21.215000 59.940000 21.535000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 60.350000 21.535000 60.670000 ;
      LAYER met4 ;
        RECT 21.215000 60.350000 21.535000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 56.250000 21.940000 56.570000 ;
      LAYER met4 ;
        RECT 21.620000 56.250000 21.940000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 56.660000 21.940000 56.980000 ;
      LAYER met4 ;
        RECT 21.620000 56.660000 21.940000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 57.070000 21.940000 57.390000 ;
      LAYER met4 ;
        RECT 21.620000 57.070000 21.940000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 57.480000 21.940000 57.800000 ;
      LAYER met4 ;
        RECT 21.620000 57.480000 21.940000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 57.890000 21.940000 58.210000 ;
      LAYER met4 ;
        RECT 21.620000 57.890000 21.940000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 58.300000 21.940000 58.620000 ;
      LAYER met4 ;
        RECT 21.620000 58.300000 21.940000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 58.710000 21.940000 59.030000 ;
      LAYER met4 ;
        RECT 21.620000 58.710000 21.940000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 59.120000 21.940000 59.440000 ;
      LAYER met4 ;
        RECT 21.620000 59.120000 21.940000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 59.530000 21.940000 59.850000 ;
      LAYER met4 ;
        RECT 21.620000 59.530000 21.940000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 59.940000 21.940000 60.260000 ;
      LAYER met4 ;
        RECT 21.620000 59.940000 21.940000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 60.350000 21.940000 60.670000 ;
      LAYER met4 ;
        RECT 21.620000 60.350000 21.940000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 56.250000 22.345000 56.570000 ;
      LAYER met4 ;
        RECT 22.025000 56.250000 22.345000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 56.660000 22.345000 56.980000 ;
      LAYER met4 ;
        RECT 22.025000 56.660000 22.345000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 57.070000 22.345000 57.390000 ;
      LAYER met4 ;
        RECT 22.025000 57.070000 22.345000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 57.480000 22.345000 57.800000 ;
      LAYER met4 ;
        RECT 22.025000 57.480000 22.345000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 57.890000 22.345000 58.210000 ;
      LAYER met4 ;
        RECT 22.025000 57.890000 22.345000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 58.300000 22.345000 58.620000 ;
      LAYER met4 ;
        RECT 22.025000 58.300000 22.345000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 58.710000 22.345000 59.030000 ;
      LAYER met4 ;
        RECT 22.025000 58.710000 22.345000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 59.120000 22.345000 59.440000 ;
      LAYER met4 ;
        RECT 22.025000 59.120000 22.345000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 59.530000 22.345000 59.850000 ;
      LAYER met4 ;
        RECT 22.025000 59.530000 22.345000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 59.940000 22.345000 60.260000 ;
      LAYER met4 ;
        RECT 22.025000 59.940000 22.345000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 60.350000 22.345000 60.670000 ;
      LAYER met4 ;
        RECT 22.025000 60.350000 22.345000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 56.250000 22.750000 56.570000 ;
      LAYER met4 ;
        RECT 22.430000 56.250000 22.750000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 56.660000 22.750000 56.980000 ;
      LAYER met4 ;
        RECT 22.430000 56.660000 22.750000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 57.070000 22.750000 57.390000 ;
      LAYER met4 ;
        RECT 22.430000 57.070000 22.750000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 57.480000 22.750000 57.800000 ;
      LAYER met4 ;
        RECT 22.430000 57.480000 22.750000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 57.890000 22.750000 58.210000 ;
      LAYER met4 ;
        RECT 22.430000 57.890000 22.750000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 58.300000 22.750000 58.620000 ;
      LAYER met4 ;
        RECT 22.430000 58.300000 22.750000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 58.710000 22.750000 59.030000 ;
      LAYER met4 ;
        RECT 22.430000 58.710000 22.750000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 59.120000 22.750000 59.440000 ;
      LAYER met4 ;
        RECT 22.430000 59.120000 22.750000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 59.530000 22.750000 59.850000 ;
      LAYER met4 ;
        RECT 22.430000 59.530000 22.750000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 59.940000 22.750000 60.260000 ;
      LAYER met4 ;
        RECT 22.430000 59.940000 22.750000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 60.350000 22.750000 60.670000 ;
      LAYER met4 ;
        RECT 22.430000 60.350000 22.750000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 56.250000 23.155000 56.570000 ;
      LAYER met4 ;
        RECT 22.835000 56.250000 23.155000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 56.660000 23.155000 56.980000 ;
      LAYER met4 ;
        RECT 22.835000 56.660000 23.155000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 57.070000 23.155000 57.390000 ;
      LAYER met4 ;
        RECT 22.835000 57.070000 23.155000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 57.480000 23.155000 57.800000 ;
      LAYER met4 ;
        RECT 22.835000 57.480000 23.155000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 57.890000 23.155000 58.210000 ;
      LAYER met4 ;
        RECT 22.835000 57.890000 23.155000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 58.300000 23.155000 58.620000 ;
      LAYER met4 ;
        RECT 22.835000 58.300000 23.155000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 58.710000 23.155000 59.030000 ;
      LAYER met4 ;
        RECT 22.835000 58.710000 23.155000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 59.120000 23.155000 59.440000 ;
      LAYER met4 ;
        RECT 22.835000 59.120000 23.155000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 59.530000 23.155000 59.850000 ;
      LAYER met4 ;
        RECT 22.835000 59.530000 23.155000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 59.940000 23.155000 60.260000 ;
      LAYER met4 ;
        RECT 22.835000 59.940000 23.155000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 60.350000 23.155000 60.670000 ;
      LAYER met4 ;
        RECT 22.835000 60.350000 23.155000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 56.250000 23.560000 56.570000 ;
      LAYER met4 ;
        RECT 23.240000 56.250000 23.560000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 56.660000 23.560000 56.980000 ;
      LAYER met4 ;
        RECT 23.240000 56.660000 23.560000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 57.070000 23.560000 57.390000 ;
      LAYER met4 ;
        RECT 23.240000 57.070000 23.560000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 57.480000 23.560000 57.800000 ;
      LAYER met4 ;
        RECT 23.240000 57.480000 23.560000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 57.890000 23.560000 58.210000 ;
      LAYER met4 ;
        RECT 23.240000 57.890000 23.560000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 58.300000 23.560000 58.620000 ;
      LAYER met4 ;
        RECT 23.240000 58.300000 23.560000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 58.710000 23.560000 59.030000 ;
      LAYER met4 ;
        RECT 23.240000 58.710000 23.560000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 59.120000 23.560000 59.440000 ;
      LAYER met4 ;
        RECT 23.240000 59.120000 23.560000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 59.530000 23.560000 59.850000 ;
      LAYER met4 ;
        RECT 23.240000 59.530000 23.560000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 59.940000 23.560000 60.260000 ;
      LAYER met4 ;
        RECT 23.240000 59.940000 23.560000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 60.350000 23.560000 60.670000 ;
      LAYER met4 ;
        RECT 23.240000 60.350000 23.560000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 56.250000 23.965000 56.570000 ;
      LAYER met4 ;
        RECT 23.645000 56.250000 23.965000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 56.660000 23.965000 56.980000 ;
      LAYER met4 ;
        RECT 23.645000 56.660000 23.965000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 57.070000 23.965000 57.390000 ;
      LAYER met4 ;
        RECT 23.645000 57.070000 23.965000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 57.480000 23.965000 57.800000 ;
      LAYER met4 ;
        RECT 23.645000 57.480000 23.965000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 57.890000 23.965000 58.210000 ;
      LAYER met4 ;
        RECT 23.645000 57.890000 23.965000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 58.300000 23.965000 58.620000 ;
      LAYER met4 ;
        RECT 23.645000 58.300000 23.965000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 58.710000 23.965000 59.030000 ;
      LAYER met4 ;
        RECT 23.645000 58.710000 23.965000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 59.120000 23.965000 59.440000 ;
      LAYER met4 ;
        RECT 23.645000 59.120000 23.965000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 59.530000 23.965000 59.850000 ;
      LAYER met4 ;
        RECT 23.645000 59.530000 23.965000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 59.940000 23.965000 60.260000 ;
      LAYER met4 ;
        RECT 23.645000 59.940000 23.965000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 60.350000 23.965000 60.670000 ;
      LAYER met4 ;
        RECT 23.645000 60.350000 23.965000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 56.250000 24.370000 56.570000 ;
      LAYER met4 ;
        RECT 24.050000 56.250000 24.370000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 56.660000 24.370000 56.980000 ;
      LAYER met4 ;
        RECT 24.050000 56.660000 24.370000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 57.070000 24.370000 57.390000 ;
      LAYER met4 ;
        RECT 24.050000 57.070000 24.370000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 57.480000 24.370000 57.800000 ;
      LAYER met4 ;
        RECT 24.050000 57.480000 24.370000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 57.890000 24.370000 58.210000 ;
      LAYER met4 ;
        RECT 24.050000 57.890000 24.370000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 58.300000 24.370000 58.620000 ;
      LAYER met4 ;
        RECT 24.050000 58.300000 24.370000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 58.710000 24.370000 59.030000 ;
      LAYER met4 ;
        RECT 24.050000 58.710000 24.370000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 59.120000 24.370000 59.440000 ;
      LAYER met4 ;
        RECT 24.050000 59.120000 24.370000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 59.530000 24.370000 59.850000 ;
      LAYER met4 ;
        RECT 24.050000 59.530000 24.370000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 59.940000 24.370000 60.260000 ;
      LAYER met4 ;
        RECT 24.050000 59.940000 24.370000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 60.350000 24.370000 60.670000 ;
      LAYER met4 ;
        RECT 24.050000 60.350000 24.370000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 56.250000 3.715000 56.570000 ;
      LAYER met4 ;
        RECT 3.395000 56.250000 3.715000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 56.660000 3.715000 56.980000 ;
      LAYER met4 ;
        RECT 3.395000 56.660000 3.715000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 57.070000 3.715000 57.390000 ;
      LAYER met4 ;
        RECT 3.395000 57.070000 3.715000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 57.480000 3.715000 57.800000 ;
      LAYER met4 ;
        RECT 3.395000 57.480000 3.715000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 57.890000 3.715000 58.210000 ;
      LAYER met4 ;
        RECT 3.395000 57.890000 3.715000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 58.300000 3.715000 58.620000 ;
      LAYER met4 ;
        RECT 3.395000 58.300000 3.715000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 58.710000 3.715000 59.030000 ;
      LAYER met4 ;
        RECT 3.395000 58.710000 3.715000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 59.120000 3.715000 59.440000 ;
      LAYER met4 ;
        RECT 3.395000 59.120000 3.715000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 59.530000 3.715000 59.850000 ;
      LAYER met4 ;
        RECT 3.395000 59.530000 3.715000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 59.940000 3.715000 60.260000 ;
      LAYER met4 ;
        RECT 3.395000 59.940000 3.715000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 60.350000 3.715000 60.670000 ;
      LAYER met4 ;
        RECT 3.395000 60.350000 3.715000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 56.250000 4.120000 56.570000 ;
      LAYER met4 ;
        RECT 3.800000 56.250000 4.120000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 56.660000 4.120000 56.980000 ;
      LAYER met4 ;
        RECT 3.800000 56.660000 4.120000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 57.070000 4.120000 57.390000 ;
      LAYER met4 ;
        RECT 3.800000 57.070000 4.120000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 57.480000 4.120000 57.800000 ;
      LAYER met4 ;
        RECT 3.800000 57.480000 4.120000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 57.890000 4.120000 58.210000 ;
      LAYER met4 ;
        RECT 3.800000 57.890000 4.120000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 58.300000 4.120000 58.620000 ;
      LAYER met4 ;
        RECT 3.800000 58.300000 4.120000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 58.710000 4.120000 59.030000 ;
      LAYER met4 ;
        RECT 3.800000 58.710000 4.120000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 59.120000 4.120000 59.440000 ;
      LAYER met4 ;
        RECT 3.800000 59.120000 4.120000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 59.530000 4.120000 59.850000 ;
      LAYER met4 ;
        RECT 3.800000 59.530000 4.120000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 59.940000 4.120000 60.260000 ;
      LAYER met4 ;
        RECT 3.800000 59.940000 4.120000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 60.350000 4.120000 60.670000 ;
      LAYER met4 ;
        RECT 3.800000 60.350000 4.120000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 56.250000 4.525000 56.570000 ;
      LAYER met4 ;
        RECT 4.205000 56.250000 4.525000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 56.660000 4.525000 56.980000 ;
      LAYER met4 ;
        RECT 4.205000 56.660000 4.525000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 57.070000 4.525000 57.390000 ;
      LAYER met4 ;
        RECT 4.205000 57.070000 4.525000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 57.480000 4.525000 57.800000 ;
      LAYER met4 ;
        RECT 4.205000 57.480000 4.525000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 57.890000 4.525000 58.210000 ;
      LAYER met4 ;
        RECT 4.205000 57.890000 4.525000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 58.300000 4.525000 58.620000 ;
      LAYER met4 ;
        RECT 4.205000 58.300000 4.525000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 58.710000 4.525000 59.030000 ;
      LAYER met4 ;
        RECT 4.205000 58.710000 4.525000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 59.120000 4.525000 59.440000 ;
      LAYER met4 ;
        RECT 4.205000 59.120000 4.525000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 59.530000 4.525000 59.850000 ;
      LAYER met4 ;
        RECT 4.205000 59.530000 4.525000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 59.940000 4.525000 60.260000 ;
      LAYER met4 ;
        RECT 4.205000 59.940000 4.525000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 60.350000 4.525000 60.670000 ;
      LAYER met4 ;
        RECT 4.205000 60.350000 4.525000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 56.250000 4.930000 56.570000 ;
      LAYER met4 ;
        RECT 4.610000 56.250000 4.930000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 56.660000 4.930000 56.980000 ;
      LAYER met4 ;
        RECT 4.610000 56.660000 4.930000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 57.070000 4.930000 57.390000 ;
      LAYER met4 ;
        RECT 4.610000 57.070000 4.930000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 57.480000 4.930000 57.800000 ;
      LAYER met4 ;
        RECT 4.610000 57.480000 4.930000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 57.890000 4.930000 58.210000 ;
      LAYER met4 ;
        RECT 4.610000 57.890000 4.930000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 58.300000 4.930000 58.620000 ;
      LAYER met4 ;
        RECT 4.610000 58.300000 4.930000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 58.710000 4.930000 59.030000 ;
      LAYER met4 ;
        RECT 4.610000 58.710000 4.930000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 59.120000 4.930000 59.440000 ;
      LAYER met4 ;
        RECT 4.610000 59.120000 4.930000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 59.530000 4.930000 59.850000 ;
      LAYER met4 ;
        RECT 4.610000 59.530000 4.930000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 59.940000 4.930000 60.260000 ;
      LAYER met4 ;
        RECT 4.610000 59.940000 4.930000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 60.350000 4.930000 60.670000 ;
      LAYER met4 ;
        RECT 4.610000 60.350000 4.930000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 56.250000 5.335000 56.570000 ;
      LAYER met4 ;
        RECT 5.015000 56.250000 5.335000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 56.660000 5.335000 56.980000 ;
      LAYER met4 ;
        RECT 5.015000 56.660000 5.335000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 57.070000 5.335000 57.390000 ;
      LAYER met4 ;
        RECT 5.015000 57.070000 5.335000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 57.480000 5.335000 57.800000 ;
      LAYER met4 ;
        RECT 5.015000 57.480000 5.335000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 57.890000 5.335000 58.210000 ;
      LAYER met4 ;
        RECT 5.015000 57.890000 5.335000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 58.300000 5.335000 58.620000 ;
      LAYER met4 ;
        RECT 5.015000 58.300000 5.335000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 58.710000 5.335000 59.030000 ;
      LAYER met4 ;
        RECT 5.015000 58.710000 5.335000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 59.120000 5.335000 59.440000 ;
      LAYER met4 ;
        RECT 5.015000 59.120000 5.335000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 59.530000 5.335000 59.850000 ;
      LAYER met4 ;
        RECT 5.015000 59.530000 5.335000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 59.940000 5.335000 60.260000 ;
      LAYER met4 ;
        RECT 5.015000 59.940000 5.335000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 60.350000 5.335000 60.670000 ;
      LAYER met4 ;
        RECT 5.015000 60.350000 5.335000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 56.250000 5.740000 56.570000 ;
      LAYER met4 ;
        RECT 5.420000 56.250000 5.740000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 56.660000 5.740000 56.980000 ;
      LAYER met4 ;
        RECT 5.420000 56.660000 5.740000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 57.070000 5.740000 57.390000 ;
      LAYER met4 ;
        RECT 5.420000 57.070000 5.740000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 57.480000 5.740000 57.800000 ;
      LAYER met4 ;
        RECT 5.420000 57.480000 5.740000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 57.890000 5.740000 58.210000 ;
      LAYER met4 ;
        RECT 5.420000 57.890000 5.740000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 58.300000 5.740000 58.620000 ;
      LAYER met4 ;
        RECT 5.420000 58.300000 5.740000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 58.710000 5.740000 59.030000 ;
      LAYER met4 ;
        RECT 5.420000 58.710000 5.740000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 59.120000 5.740000 59.440000 ;
      LAYER met4 ;
        RECT 5.420000 59.120000 5.740000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 59.530000 5.740000 59.850000 ;
      LAYER met4 ;
        RECT 5.420000 59.530000 5.740000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 59.940000 5.740000 60.260000 ;
      LAYER met4 ;
        RECT 5.420000 59.940000 5.740000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 60.350000 5.740000 60.670000 ;
      LAYER met4 ;
        RECT 5.420000 60.350000 5.740000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 56.250000 6.145000 56.570000 ;
      LAYER met4 ;
        RECT 5.825000 56.250000 6.145000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 56.660000 6.145000 56.980000 ;
      LAYER met4 ;
        RECT 5.825000 56.660000 6.145000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 57.070000 6.145000 57.390000 ;
      LAYER met4 ;
        RECT 5.825000 57.070000 6.145000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 57.480000 6.145000 57.800000 ;
      LAYER met4 ;
        RECT 5.825000 57.480000 6.145000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 57.890000 6.145000 58.210000 ;
      LAYER met4 ;
        RECT 5.825000 57.890000 6.145000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 58.300000 6.145000 58.620000 ;
      LAYER met4 ;
        RECT 5.825000 58.300000 6.145000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 58.710000 6.145000 59.030000 ;
      LAYER met4 ;
        RECT 5.825000 58.710000 6.145000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 59.120000 6.145000 59.440000 ;
      LAYER met4 ;
        RECT 5.825000 59.120000 6.145000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 59.530000 6.145000 59.850000 ;
      LAYER met4 ;
        RECT 5.825000 59.530000 6.145000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 59.940000 6.145000 60.260000 ;
      LAYER met4 ;
        RECT 5.825000 59.940000 6.145000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 60.350000 6.145000 60.670000 ;
      LAYER met4 ;
        RECT 5.825000 60.350000 6.145000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 56.250000 51.105000 56.570000 ;
      LAYER met4 ;
        RECT 50.785000 56.250000 51.105000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 56.660000 51.105000 56.980000 ;
      LAYER met4 ;
        RECT 50.785000 56.660000 51.105000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 57.070000 51.105000 57.390000 ;
      LAYER met4 ;
        RECT 50.785000 57.070000 51.105000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 57.480000 51.105000 57.800000 ;
      LAYER met4 ;
        RECT 50.785000 57.480000 51.105000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 57.890000 51.105000 58.210000 ;
      LAYER met4 ;
        RECT 50.785000 57.890000 51.105000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 58.300000 51.105000 58.620000 ;
      LAYER met4 ;
        RECT 50.785000 58.300000 51.105000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 58.710000 51.105000 59.030000 ;
      LAYER met4 ;
        RECT 50.785000 58.710000 51.105000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 59.120000 51.105000 59.440000 ;
      LAYER met4 ;
        RECT 50.785000 59.120000 51.105000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 59.530000 51.105000 59.850000 ;
      LAYER met4 ;
        RECT 50.785000 59.530000 51.105000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 59.940000 51.105000 60.260000 ;
      LAYER met4 ;
        RECT 50.785000 59.940000 51.105000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 60.350000 51.105000 60.670000 ;
      LAYER met4 ;
        RECT 50.785000 60.350000 51.105000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 56.250000 51.515000 56.570000 ;
      LAYER met4 ;
        RECT 51.195000 56.250000 51.515000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 56.660000 51.515000 56.980000 ;
      LAYER met4 ;
        RECT 51.195000 56.660000 51.515000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 57.070000 51.515000 57.390000 ;
      LAYER met4 ;
        RECT 51.195000 57.070000 51.515000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 57.480000 51.515000 57.800000 ;
      LAYER met4 ;
        RECT 51.195000 57.480000 51.515000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 57.890000 51.515000 58.210000 ;
      LAYER met4 ;
        RECT 51.195000 57.890000 51.515000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 58.300000 51.515000 58.620000 ;
      LAYER met4 ;
        RECT 51.195000 58.300000 51.515000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 58.710000 51.515000 59.030000 ;
      LAYER met4 ;
        RECT 51.195000 58.710000 51.515000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 59.120000 51.515000 59.440000 ;
      LAYER met4 ;
        RECT 51.195000 59.120000 51.515000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 59.530000 51.515000 59.850000 ;
      LAYER met4 ;
        RECT 51.195000 59.530000 51.515000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 59.940000 51.515000 60.260000 ;
      LAYER met4 ;
        RECT 51.195000 59.940000 51.515000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 60.350000 51.515000 60.670000 ;
      LAYER met4 ;
        RECT 51.195000 60.350000 51.515000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 56.250000 51.925000 56.570000 ;
      LAYER met4 ;
        RECT 51.605000 56.250000 51.925000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 56.660000 51.925000 56.980000 ;
      LAYER met4 ;
        RECT 51.605000 56.660000 51.925000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 57.070000 51.925000 57.390000 ;
      LAYER met4 ;
        RECT 51.605000 57.070000 51.925000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 57.480000 51.925000 57.800000 ;
      LAYER met4 ;
        RECT 51.605000 57.480000 51.925000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 57.890000 51.925000 58.210000 ;
      LAYER met4 ;
        RECT 51.605000 57.890000 51.925000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 58.300000 51.925000 58.620000 ;
      LAYER met4 ;
        RECT 51.605000 58.300000 51.925000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 58.710000 51.925000 59.030000 ;
      LAYER met4 ;
        RECT 51.605000 58.710000 51.925000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 59.120000 51.925000 59.440000 ;
      LAYER met4 ;
        RECT 51.605000 59.120000 51.925000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 59.530000 51.925000 59.850000 ;
      LAYER met4 ;
        RECT 51.605000 59.530000 51.925000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 59.940000 51.925000 60.260000 ;
      LAYER met4 ;
        RECT 51.605000 59.940000 51.925000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 60.350000 51.925000 60.670000 ;
      LAYER met4 ;
        RECT 51.605000 60.350000 51.925000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 56.250000 52.335000 56.570000 ;
      LAYER met4 ;
        RECT 52.015000 56.250000 52.335000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 56.660000 52.335000 56.980000 ;
      LAYER met4 ;
        RECT 52.015000 56.660000 52.335000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 57.070000 52.335000 57.390000 ;
      LAYER met4 ;
        RECT 52.015000 57.070000 52.335000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 57.480000 52.335000 57.800000 ;
      LAYER met4 ;
        RECT 52.015000 57.480000 52.335000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 57.890000 52.335000 58.210000 ;
      LAYER met4 ;
        RECT 52.015000 57.890000 52.335000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 58.300000 52.335000 58.620000 ;
      LAYER met4 ;
        RECT 52.015000 58.300000 52.335000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 58.710000 52.335000 59.030000 ;
      LAYER met4 ;
        RECT 52.015000 58.710000 52.335000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 59.120000 52.335000 59.440000 ;
      LAYER met4 ;
        RECT 52.015000 59.120000 52.335000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 59.530000 52.335000 59.850000 ;
      LAYER met4 ;
        RECT 52.015000 59.530000 52.335000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 59.940000 52.335000 60.260000 ;
      LAYER met4 ;
        RECT 52.015000 59.940000 52.335000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 60.350000 52.335000 60.670000 ;
      LAYER met4 ;
        RECT 52.015000 60.350000 52.335000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 56.250000 52.745000 56.570000 ;
      LAYER met4 ;
        RECT 52.425000 56.250000 52.745000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 56.660000 52.745000 56.980000 ;
      LAYER met4 ;
        RECT 52.425000 56.660000 52.745000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 57.070000 52.745000 57.390000 ;
      LAYER met4 ;
        RECT 52.425000 57.070000 52.745000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 57.480000 52.745000 57.800000 ;
      LAYER met4 ;
        RECT 52.425000 57.480000 52.745000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 57.890000 52.745000 58.210000 ;
      LAYER met4 ;
        RECT 52.425000 57.890000 52.745000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 58.300000 52.745000 58.620000 ;
      LAYER met4 ;
        RECT 52.425000 58.300000 52.745000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 58.710000 52.745000 59.030000 ;
      LAYER met4 ;
        RECT 52.425000 58.710000 52.745000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 59.120000 52.745000 59.440000 ;
      LAYER met4 ;
        RECT 52.425000 59.120000 52.745000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 59.530000 52.745000 59.850000 ;
      LAYER met4 ;
        RECT 52.425000 59.530000 52.745000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 59.940000 52.745000 60.260000 ;
      LAYER met4 ;
        RECT 52.425000 59.940000 52.745000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 60.350000 52.745000 60.670000 ;
      LAYER met4 ;
        RECT 52.425000 60.350000 52.745000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 56.250000 53.155000 56.570000 ;
      LAYER met4 ;
        RECT 52.835000 56.250000 53.155000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 56.660000 53.155000 56.980000 ;
      LAYER met4 ;
        RECT 52.835000 56.660000 53.155000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 57.070000 53.155000 57.390000 ;
      LAYER met4 ;
        RECT 52.835000 57.070000 53.155000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 57.480000 53.155000 57.800000 ;
      LAYER met4 ;
        RECT 52.835000 57.480000 53.155000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 57.890000 53.155000 58.210000 ;
      LAYER met4 ;
        RECT 52.835000 57.890000 53.155000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 58.300000 53.155000 58.620000 ;
      LAYER met4 ;
        RECT 52.835000 58.300000 53.155000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 58.710000 53.155000 59.030000 ;
      LAYER met4 ;
        RECT 52.835000 58.710000 53.155000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 59.120000 53.155000 59.440000 ;
      LAYER met4 ;
        RECT 52.835000 59.120000 53.155000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 59.530000 53.155000 59.850000 ;
      LAYER met4 ;
        RECT 52.835000 59.530000 53.155000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 59.940000 53.155000 60.260000 ;
      LAYER met4 ;
        RECT 52.835000 59.940000 53.155000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 60.350000 53.155000 60.670000 ;
      LAYER met4 ;
        RECT 52.835000 60.350000 53.155000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 56.250000 53.565000 56.570000 ;
      LAYER met4 ;
        RECT 53.245000 56.250000 53.565000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 56.660000 53.565000 56.980000 ;
      LAYER met4 ;
        RECT 53.245000 56.660000 53.565000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 57.070000 53.565000 57.390000 ;
      LAYER met4 ;
        RECT 53.245000 57.070000 53.565000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 57.480000 53.565000 57.800000 ;
      LAYER met4 ;
        RECT 53.245000 57.480000 53.565000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 57.890000 53.565000 58.210000 ;
      LAYER met4 ;
        RECT 53.245000 57.890000 53.565000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 58.300000 53.565000 58.620000 ;
      LAYER met4 ;
        RECT 53.245000 58.300000 53.565000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 58.710000 53.565000 59.030000 ;
      LAYER met4 ;
        RECT 53.245000 58.710000 53.565000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 59.120000 53.565000 59.440000 ;
      LAYER met4 ;
        RECT 53.245000 59.120000 53.565000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 59.530000 53.565000 59.850000 ;
      LAYER met4 ;
        RECT 53.245000 59.530000 53.565000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 59.940000 53.565000 60.260000 ;
      LAYER met4 ;
        RECT 53.245000 59.940000 53.565000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 60.350000 53.565000 60.670000 ;
      LAYER met4 ;
        RECT 53.245000 60.350000 53.565000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 56.250000 53.975000 56.570000 ;
      LAYER met4 ;
        RECT 53.655000 56.250000 53.975000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 56.660000 53.975000 56.980000 ;
      LAYER met4 ;
        RECT 53.655000 56.660000 53.975000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 57.070000 53.975000 57.390000 ;
      LAYER met4 ;
        RECT 53.655000 57.070000 53.975000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 57.480000 53.975000 57.800000 ;
      LAYER met4 ;
        RECT 53.655000 57.480000 53.975000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 57.890000 53.975000 58.210000 ;
      LAYER met4 ;
        RECT 53.655000 57.890000 53.975000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 58.300000 53.975000 58.620000 ;
      LAYER met4 ;
        RECT 53.655000 58.300000 53.975000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 58.710000 53.975000 59.030000 ;
      LAYER met4 ;
        RECT 53.655000 58.710000 53.975000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 59.120000 53.975000 59.440000 ;
      LAYER met4 ;
        RECT 53.655000 59.120000 53.975000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 59.530000 53.975000 59.850000 ;
      LAYER met4 ;
        RECT 53.655000 59.530000 53.975000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 59.940000 53.975000 60.260000 ;
      LAYER met4 ;
        RECT 53.655000 59.940000 53.975000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.655000 60.350000 53.975000 60.670000 ;
      LAYER met4 ;
        RECT 53.655000 60.350000 53.975000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 56.250000 54.385000 56.570000 ;
      LAYER met4 ;
        RECT 54.065000 56.250000 54.385000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 56.660000 54.385000 56.980000 ;
      LAYER met4 ;
        RECT 54.065000 56.660000 54.385000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 57.070000 54.385000 57.390000 ;
      LAYER met4 ;
        RECT 54.065000 57.070000 54.385000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 57.480000 54.385000 57.800000 ;
      LAYER met4 ;
        RECT 54.065000 57.480000 54.385000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 57.890000 54.385000 58.210000 ;
      LAYER met4 ;
        RECT 54.065000 57.890000 54.385000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 58.300000 54.385000 58.620000 ;
      LAYER met4 ;
        RECT 54.065000 58.300000 54.385000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 58.710000 54.385000 59.030000 ;
      LAYER met4 ;
        RECT 54.065000 58.710000 54.385000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 59.120000 54.385000 59.440000 ;
      LAYER met4 ;
        RECT 54.065000 59.120000 54.385000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 59.530000 54.385000 59.850000 ;
      LAYER met4 ;
        RECT 54.065000 59.530000 54.385000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 59.940000 54.385000 60.260000 ;
      LAYER met4 ;
        RECT 54.065000 59.940000 54.385000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 60.350000 54.385000 60.670000 ;
      LAYER met4 ;
        RECT 54.065000 60.350000 54.385000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 56.250000 54.795000 56.570000 ;
      LAYER met4 ;
        RECT 54.475000 56.250000 54.795000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 56.660000 54.795000 56.980000 ;
      LAYER met4 ;
        RECT 54.475000 56.660000 54.795000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 57.070000 54.795000 57.390000 ;
      LAYER met4 ;
        RECT 54.475000 57.070000 54.795000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 57.480000 54.795000 57.800000 ;
      LAYER met4 ;
        RECT 54.475000 57.480000 54.795000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 57.890000 54.795000 58.210000 ;
      LAYER met4 ;
        RECT 54.475000 57.890000 54.795000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 58.300000 54.795000 58.620000 ;
      LAYER met4 ;
        RECT 54.475000 58.300000 54.795000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 58.710000 54.795000 59.030000 ;
      LAYER met4 ;
        RECT 54.475000 58.710000 54.795000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 59.120000 54.795000 59.440000 ;
      LAYER met4 ;
        RECT 54.475000 59.120000 54.795000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 59.530000 54.795000 59.850000 ;
      LAYER met4 ;
        RECT 54.475000 59.530000 54.795000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 59.940000 54.795000 60.260000 ;
      LAYER met4 ;
        RECT 54.475000 59.940000 54.795000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.475000 60.350000 54.795000 60.670000 ;
      LAYER met4 ;
        RECT 54.475000 60.350000 54.795000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 56.250000 55.205000 56.570000 ;
      LAYER met4 ;
        RECT 54.885000 56.250000 55.205000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 56.660000 55.205000 56.980000 ;
      LAYER met4 ;
        RECT 54.885000 56.660000 55.205000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 57.070000 55.205000 57.390000 ;
      LAYER met4 ;
        RECT 54.885000 57.070000 55.205000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 57.480000 55.205000 57.800000 ;
      LAYER met4 ;
        RECT 54.885000 57.480000 55.205000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 57.890000 55.205000 58.210000 ;
      LAYER met4 ;
        RECT 54.885000 57.890000 55.205000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 58.300000 55.205000 58.620000 ;
      LAYER met4 ;
        RECT 54.885000 58.300000 55.205000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 58.710000 55.205000 59.030000 ;
      LAYER met4 ;
        RECT 54.885000 58.710000 55.205000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 59.120000 55.205000 59.440000 ;
      LAYER met4 ;
        RECT 54.885000 59.120000 55.205000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 59.530000 55.205000 59.850000 ;
      LAYER met4 ;
        RECT 54.885000 59.530000 55.205000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 59.940000 55.205000 60.260000 ;
      LAYER met4 ;
        RECT 54.885000 59.940000 55.205000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.885000 60.350000 55.205000 60.670000 ;
      LAYER met4 ;
        RECT 54.885000 60.350000 55.205000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 56.250000 55.615000 56.570000 ;
      LAYER met4 ;
        RECT 55.295000 56.250000 55.615000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 56.660000 55.615000 56.980000 ;
      LAYER met4 ;
        RECT 55.295000 56.660000 55.615000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 57.070000 55.615000 57.390000 ;
      LAYER met4 ;
        RECT 55.295000 57.070000 55.615000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 57.480000 55.615000 57.800000 ;
      LAYER met4 ;
        RECT 55.295000 57.480000 55.615000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 57.890000 55.615000 58.210000 ;
      LAYER met4 ;
        RECT 55.295000 57.890000 55.615000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 58.300000 55.615000 58.620000 ;
      LAYER met4 ;
        RECT 55.295000 58.300000 55.615000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 58.710000 55.615000 59.030000 ;
      LAYER met4 ;
        RECT 55.295000 58.710000 55.615000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 59.120000 55.615000 59.440000 ;
      LAYER met4 ;
        RECT 55.295000 59.120000 55.615000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 59.530000 55.615000 59.850000 ;
      LAYER met4 ;
        RECT 55.295000 59.530000 55.615000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 59.940000 55.615000 60.260000 ;
      LAYER met4 ;
        RECT 55.295000 59.940000 55.615000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.295000 60.350000 55.615000 60.670000 ;
      LAYER met4 ;
        RECT 55.295000 60.350000 55.615000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 56.250000 56.025000 56.570000 ;
      LAYER met4 ;
        RECT 55.705000 56.250000 56.025000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 56.660000 56.025000 56.980000 ;
      LAYER met4 ;
        RECT 55.705000 56.660000 56.025000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 57.070000 56.025000 57.390000 ;
      LAYER met4 ;
        RECT 55.705000 57.070000 56.025000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 57.480000 56.025000 57.800000 ;
      LAYER met4 ;
        RECT 55.705000 57.480000 56.025000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 57.890000 56.025000 58.210000 ;
      LAYER met4 ;
        RECT 55.705000 57.890000 56.025000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 58.300000 56.025000 58.620000 ;
      LAYER met4 ;
        RECT 55.705000 58.300000 56.025000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 58.710000 56.025000 59.030000 ;
      LAYER met4 ;
        RECT 55.705000 58.710000 56.025000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 59.120000 56.025000 59.440000 ;
      LAYER met4 ;
        RECT 55.705000 59.120000 56.025000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 59.530000 56.025000 59.850000 ;
      LAYER met4 ;
        RECT 55.705000 59.530000 56.025000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 59.940000 56.025000 60.260000 ;
      LAYER met4 ;
        RECT 55.705000 59.940000 56.025000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705000 60.350000 56.025000 60.670000 ;
      LAYER met4 ;
        RECT 55.705000 60.350000 56.025000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 56.250000 56.435000 56.570000 ;
      LAYER met4 ;
        RECT 56.115000 56.250000 56.435000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 56.660000 56.435000 56.980000 ;
      LAYER met4 ;
        RECT 56.115000 56.660000 56.435000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 57.070000 56.435000 57.390000 ;
      LAYER met4 ;
        RECT 56.115000 57.070000 56.435000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 57.480000 56.435000 57.800000 ;
      LAYER met4 ;
        RECT 56.115000 57.480000 56.435000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 57.890000 56.435000 58.210000 ;
      LAYER met4 ;
        RECT 56.115000 57.890000 56.435000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 58.300000 56.435000 58.620000 ;
      LAYER met4 ;
        RECT 56.115000 58.300000 56.435000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 58.710000 56.435000 59.030000 ;
      LAYER met4 ;
        RECT 56.115000 58.710000 56.435000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 59.120000 56.435000 59.440000 ;
      LAYER met4 ;
        RECT 56.115000 59.120000 56.435000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 59.530000 56.435000 59.850000 ;
      LAYER met4 ;
        RECT 56.115000 59.530000 56.435000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 59.940000 56.435000 60.260000 ;
      LAYER met4 ;
        RECT 56.115000 59.940000 56.435000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.115000 60.350000 56.435000 60.670000 ;
      LAYER met4 ;
        RECT 56.115000 60.350000 56.435000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 56.250000 56.845000 56.570000 ;
      LAYER met4 ;
        RECT 56.525000 56.250000 56.845000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 56.660000 56.845000 56.980000 ;
      LAYER met4 ;
        RECT 56.525000 56.660000 56.845000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 57.070000 56.845000 57.390000 ;
      LAYER met4 ;
        RECT 56.525000 57.070000 56.845000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 57.480000 56.845000 57.800000 ;
      LAYER met4 ;
        RECT 56.525000 57.480000 56.845000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 57.890000 56.845000 58.210000 ;
      LAYER met4 ;
        RECT 56.525000 57.890000 56.845000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 58.300000 56.845000 58.620000 ;
      LAYER met4 ;
        RECT 56.525000 58.300000 56.845000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 58.710000 56.845000 59.030000 ;
      LAYER met4 ;
        RECT 56.525000 58.710000 56.845000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 59.120000 56.845000 59.440000 ;
      LAYER met4 ;
        RECT 56.525000 59.120000 56.845000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 59.530000 56.845000 59.850000 ;
      LAYER met4 ;
        RECT 56.525000 59.530000 56.845000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 59.940000 56.845000 60.260000 ;
      LAYER met4 ;
        RECT 56.525000 59.940000 56.845000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 60.350000 56.845000 60.670000 ;
      LAYER met4 ;
        RECT 56.525000 60.350000 56.845000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 56.250000 57.250000 56.570000 ;
      LAYER met4 ;
        RECT 56.930000 56.250000 57.250000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 56.660000 57.250000 56.980000 ;
      LAYER met4 ;
        RECT 56.930000 56.660000 57.250000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 57.070000 57.250000 57.390000 ;
      LAYER met4 ;
        RECT 56.930000 57.070000 57.250000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 57.480000 57.250000 57.800000 ;
      LAYER met4 ;
        RECT 56.930000 57.480000 57.250000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 57.890000 57.250000 58.210000 ;
      LAYER met4 ;
        RECT 56.930000 57.890000 57.250000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 58.300000 57.250000 58.620000 ;
      LAYER met4 ;
        RECT 56.930000 58.300000 57.250000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 58.710000 57.250000 59.030000 ;
      LAYER met4 ;
        RECT 56.930000 58.710000 57.250000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 59.120000 57.250000 59.440000 ;
      LAYER met4 ;
        RECT 56.930000 59.120000 57.250000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 59.530000 57.250000 59.850000 ;
      LAYER met4 ;
        RECT 56.930000 59.530000 57.250000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 59.940000 57.250000 60.260000 ;
      LAYER met4 ;
        RECT 56.930000 59.940000 57.250000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 60.350000 57.250000 60.670000 ;
      LAYER met4 ;
        RECT 56.930000 60.350000 57.250000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 56.250000 57.655000 56.570000 ;
      LAYER met4 ;
        RECT 57.335000 56.250000 57.655000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 56.660000 57.655000 56.980000 ;
      LAYER met4 ;
        RECT 57.335000 56.660000 57.655000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 57.070000 57.655000 57.390000 ;
      LAYER met4 ;
        RECT 57.335000 57.070000 57.655000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 57.480000 57.655000 57.800000 ;
      LAYER met4 ;
        RECT 57.335000 57.480000 57.655000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 57.890000 57.655000 58.210000 ;
      LAYER met4 ;
        RECT 57.335000 57.890000 57.655000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 58.300000 57.655000 58.620000 ;
      LAYER met4 ;
        RECT 57.335000 58.300000 57.655000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 58.710000 57.655000 59.030000 ;
      LAYER met4 ;
        RECT 57.335000 58.710000 57.655000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 59.120000 57.655000 59.440000 ;
      LAYER met4 ;
        RECT 57.335000 59.120000 57.655000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 59.530000 57.655000 59.850000 ;
      LAYER met4 ;
        RECT 57.335000 59.530000 57.655000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 59.940000 57.655000 60.260000 ;
      LAYER met4 ;
        RECT 57.335000 59.940000 57.655000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 60.350000 57.655000 60.670000 ;
      LAYER met4 ;
        RECT 57.335000 60.350000 57.655000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 56.250000 58.060000 56.570000 ;
      LAYER met4 ;
        RECT 57.740000 56.250000 58.060000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 56.660000 58.060000 56.980000 ;
      LAYER met4 ;
        RECT 57.740000 56.660000 58.060000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 57.070000 58.060000 57.390000 ;
      LAYER met4 ;
        RECT 57.740000 57.070000 58.060000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 57.480000 58.060000 57.800000 ;
      LAYER met4 ;
        RECT 57.740000 57.480000 58.060000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 57.890000 58.060000 58.210000 ;
      LAYER met4 ;
        RECT 57.740000 57.890000 58.060000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 58.300000 58.060000 58.620000 ;
      LAYER met4 ;
        RECT 57.740000 58.300000 58.060000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 58.710000 58.060000 59.030000 ;
      LAYER met4 ;
        RECT 57.740000 58.710000 58.060000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 59.120000 58.060000 59.440000 ;
      LAYER met4 ;
        RECT 57.740000 59.120000 58.060000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 59.530000 58.060000 59.850000 ;
      LAYER met4 ;
        RECT 57.740000 59.530000 58.060000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 59.940000 58.060000 60.260000 ;
      LAYER met4 ;
        RECT 57.740000 59.940000 58.060000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 60.350000 58.060000 60.670000 ;
      LAYER met4 ;
        RECT 57.740000 60.350000 58.060000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 56.250000 58.465000 56.570000 ;
      LAYER met4 ;
        RECT 58.145000 56.250000 58.465000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 56.660000 58.465000 56.980000 ;
      LAYER met4 ;
        RECT 58.145000 56.660000 58.465000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 57.070000 58.465000 57.390000 ;
      LAYER met4 ;
        RECT 58.145000 57.070000 58.465000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 57.480000 58.465000 57.800000 ;
      LAYER met4 ;
        RECT 58.145000 57.480000 58.465000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 57.890000 58.465000 58.210000 ;
      LAYER met4 ;
        RECT 58.145000 57.890000 58.465000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 58.300000 58.465000 58.620000 ;
      LAYER met4 ;
        RECT 58.145000 58.300000 58.465000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 58.710000 58.465000 59.030000 ;
      LAYER met4 ;
        RECT 58.145000 58.710000 58.465000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 59.120000 58.465000 59.440000 ;
      LAYER met4 ;
        RECT 58.145000 59.120000 58.465000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 59.530000 58.465000 59.850000 ;
      LAYER met4 ;
        RECT 58.145000 59.530000 58.465000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 59.940000 58.465000 60.260000 ;
      LAYER met4 ;
        RECT 58.145000 59.940000 58.465000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 60.350000 58.465000 60.670000 ;
      LAYER met4 ;
        RECT 58.145000 60.350000 58.465000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 56.250000 58.870000 56.570000 ;
      LAYER met4 ;
        RECT 58.550000 56.250000 58.870000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 56.660000 58.870000 56.980000 ;
      LAYER met4 ;
        RECT 58.550000 56.660000 58.870000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 57.070000 58.870000 57.390000 ;
      LAYER met4 ;
        RECT 58.550000 57.070000 58.870000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 57.480000 58.870000 57.800000 ;
      LAYER met4 ;
        RECT 58.550000 57.480000 58.870000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 57.890000 58.870000 58.210000 ;
      LAYER met4 ;
        RECT 58.550000 57.890000 58.870000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 58.300000 58.870000 58.620000 ;
      LAYER met4 ;
        RECT 58.550000 58.300000 58.870000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 58.710000 58.870000 59.030000 ;
      LAYER met4 ;
        RECT 58.550000 58.710000 58.870000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 59.120000 58.870000 59.440000 ;
      LAYER met4 ;
        RECT 58.550000 59.120000 58.870000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 59.530000 58.870000 59.850000 ;
      LAYER met4 ;
        RECT 58.550000 59.530000 58.870000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 59.940000 58.870000 60.260000 ;
      LAYER met4 ;
        RECT 58.550000 59.940000 58.870000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 60.350000 58.870000 60.670000 ;
      LAYER met4 ;
        RECT 58.550000 60.350000 58.870000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 56.250000 59.275000 56.570000 ;
      LAYER met4 ;
        RECT 58.955000 56.250000 59.275000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 56.660000 59.275000 56.980000 ;
      LAYER met4 ;
        RECT 58.955000 56.660000 59.275000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 57.070000 59.275000 57.390000 ;
      LAYER met4 ;
        RECT 58.955000 57.070000 59.275000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 57.480000 59.275000 57.800000 ;
      LAYER met4 ;
        RECT 58.955000 57.480000 59.275000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 57.890000 59.275000 58.210000 ;
      LAYER met4 ;
        RECT 58.955000 57.890000 59.275000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 58.300000 59.275000 58.620000 ;
      LAYER met4 ;
        RECT 58.955000 58.300000 59.275000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 58.710000 59.275000 59.030000 ;
      LAYER met4 ;
        RECT 58.955000 58.710000 59.275000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 59.120000 59.275000 59.440000 ;
      LAYER met4 ;
        RECT 58.955000 59.120000 59.275000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 59.530000 59.275000 59.850000 ;
      LAYER met4 ;
        RECT 58.955000 59.530000 59.275000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 59.940000 59.275000 60.260000 ;
      LAYER met4 ;
        RECT 58.955000 59.940000 59.275000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 60.350000 59.275000 60.670000 ;
      LAYER met4 ;
        RECT 58.955000 60.350000 59.275000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 56.250000 59.680000 56.570000 ;
      LAYER met4 ;
        RECT 59.360000 56.250000 59.680000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 56.660000 59.680000 56.980000 ;
      LAYER met4 ;
        RECT 59.360000 56.660000 59.680000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 57.070000 59.680000 57.390000 ;
      LAYER met4 ;
        RECT 59.360000 57.070000 59.680000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 57.480000 59.680000 57.800000 ;
      LAYER met4 ;
        RECT 59.360000 57.480000 59.680000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 57.890000 59.680000 58.210000 ;
      LAYER met4 ;
        RECT 59.360000 57.890000 59.680000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 58.300000 59.680000 58.620000 ;
      LAYER met4 ;
        RECT 59.360000 58.300000 59.680000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 58.710000 59.680000 59.030000 ;
      LAYER met4 ;
        RECT 59.360000 58.710000 59.680000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 59.120000 59.680000 59.440000 ;
      LAYER met4 ;
        RECT 59.360000 59.120000 59.680000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 59.530000 59.680000 59.850000 ;
      LAYER met4 ;
        RECT 59.360000 59.530000 59.680000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 59.940000 59.680000 60.260000 ;
      LAYER met4 ;
        RECT 59.360000 59.940000 59.680000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 60.350000 59.680000 60.670000 ;
      LAYER met4 ;
        RECT 59.360000 60.350000 59.680000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 56.250000 60.085000 56.570000 ;
      LAYER met4 ;
        RECT 59.765000 56.250000 60.085000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 56.660000 60.085000 56.980000 ;
      LAYER met4 ;
        RECT 59.765000 56.660000 60.085000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 57.070000 60.085000 57.390000 ;
      LAYER met4 ;
        RECT 59.765000 57.070000 60.085000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 57.480000 60.085000 57.800000 ;
      LAYER met4 ;
        RECT 59.765000 57.480000 60.085000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 57.890000 60.085000 58.210000 ;
      LAYER met4 ;
        RECT 59.765000 57.890000 60.085000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 58.300000 60.085000 58.620000 ;
      LAYER met4 ;
        RECT 59.765000 58.300000 60.085000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 58.710000 60.085000 59.030000 ;
      LAYER met4 ;
        RECT 59.765000 58.710000 60.085000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 59.120000 60.085000 59.440000 ;
      LAYER met4 ;
        RECT 59.765000 59.120000 60.085000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 59.530000 60.085000 59.850000 ;
      LAYER met4 ;
        RECT 59.765000 59.530000 60.085000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 59.940000 60.085000 60.260000 ;
      LAYER met4 ;
        RECT 59.765000 59.940000 60.085000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 60.350000 60.085000 60.670000 ;
      LAYER met4 ;
        RECT 59.765000 60.350000 60.085000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 56.250000 6.550000 56.570000 ;
      LAYER met4 ;
        RECT 6.230000 56.250000 6.550000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 56.660000 6.550000 56.980000 ;
      LAYER met4 ;
        RECT 6.230000 56.660000 6.550000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 57.070000 6.550000 57.390000 ;
      LAYER met4 ;
        RECT 6.230000 57.070000 6.550000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 57.480000 6.550000 57.800000 ;
      LAYER met4 ;
        RECT 6.230000 57.480000 6.550000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 57.890000 6.550000 58.210000 ;
      LAYER met4 ;
        RECT 6.230000 57.890000 6.550000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 58.300000 6.550000 58.620000 ;
      LAYER met4 ;
        RECT 6.230000 58.300000 6.550000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 58.710000 6.550000 59.030000 ;
      LAYER met4 ;
        RECT 6.230000 58.710000 6.550000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 59.120000 6.550000 59.440000 ;
      LAYER met4 ;
        RECT 6.230000 59.120000 6.550000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 59.530000 6.550000 59.850000 ;
      LAYER met4 ;
        RECT 6.230000 59.530000 6.550000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 59.940000 6.550000 60.260000 ;
      LAYER met4 ;
        RECT 6.230000 59.940000 6.550000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 60.350000 6.550000 60.670000 ;
      LAYER met4 ;
        RECT 6.230000 60.350000 6.550000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 56.250000 6.955000 56.570000 ;
      LAYER met4 ;
        RECT 6.635000 56.250000 6.955000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 56.660000 6.955000 56.980000 ;
      LAYER met4 ;
        RECT 6.635000 56.660000 6.955000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 57.070000 6.955000 57.390000 ;
      LAYER met4 ;
        RECT 6.635000 57.070000 6.955000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 57.480000 6.955000 57.800000 ;
      LAYER met4 ;
        RECT 6.635000 57.480000 6.955000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 57.890000 6.955000 58.210000 ;
      LAYER met4 ;
        RECT 6.635000 57.890000 6.955000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 58.300000 6.955000 58.620000 ;
      LAYER met4 ;
        RECT 6.635000 58.300000 6.955000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 58.710000 6.955000 59.030000 ;
      LAYER met4 ;
        RECT 6.635000 58.710000 6.955000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 59.120000 6.955000 59.440000 ;
      LAYER met4 ;
        RECT 6.635000 59.120000 6.955000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 59.530000 6.955000 59.850000 ;
      LAYER met4 ;
        RECT 6.635000 59.530000 6.955000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 59.940000 6.955000 60.260000 ;
      LAYER met4 ;
        RECT 6.635000 59.940000 6.955000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 60.350000 6.955000 60.670000 ;
      LAYER met4 ;
        RECT 6.635000 60.350000 6.955000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 56.250000 60.490000 56.570000 ;
      LAYER met4 ;
        RECT 60.170000 56.250000 60.490000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 56.660000 60.490000 56.980000 ;
      LAYER met4 ;
        RECT 60.170000 56.660000 60.490000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 57.070000 60.490000 57.390000 ;
      LAYER met4 ;
        RECT 60.170000 57.070000 60.490000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 57.480000 60.490000 57.800000 ;
      LAYER met4 ;
        RECT 60.170000 57.480000 60.490000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 57.890000 60.490000 58.210000 ;
      LAYER met4 ;
        RECT 60.170000 57.890000 60.490000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 58.300000 60.490000 58.620000 ;
      LAYER met4 ;
        RECT 60.170000 58.300000 60.490000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 58.710000 60.490000 59.030000 ;
      LAYER met4 ;
        RECT 60.170000 58.710000 60.490000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 59.120000 60.490000 59.440000 ;
      LAYER met4 ;
        RECT 60.170000 59.120000 60.490000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 59.530000 60.490000 59.850000 ;
      LAYER met4 ;
        RECT 60.170000 59.530000 60.490000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 59.940000 60.490000 60.260000 ;
      LAYER met4 ;
        RECT 60.170000 59.940000 60.490000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 60.350000 60.490000 60.670000 ;
      LAYER met4 ;
        RECT 60.170000 60.350000 60.490000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 56.250000 60.895000 56.570000 ;
      LAYER met4 ;
        RECT 60.575000 56.250000 60.895000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 56.660000 60.895000 56.980000 ;
      LAYER met4 ;
        RECT 60.575000 56.660000 60.895000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 57.070000 60.895000 57.390000 ;
      LAYER met4 ;
        RECT 60.575000 57.070000 60.895000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 57.480000 60.895000 57.800000 ;
      LAYER met4 ;
        RECT 60.575000 57.480000 60.895000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 57.890000 60.895000 58.210000 ;
      LAYER met4 ;
        RECT 60.575000 57.890000 60.895000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 58.300000 60.895000 58.620000 ;
      LAYER met4 ;
        RECT 60.575000 58.300000 60.895000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 58.710000 60.895000 59.030000 ;
      LAYER met4 ;
        RECT 60.575000 58.710000 60.895000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 59.120000 60.895000 59.440000 ;
      LAYER met4 ;
        RECT 60.575000 59.120000 60.895000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 59.530000 60.895000 59.850000 ;
      LAYER met4 ;
        RECT 60.575000 59.530000 60.895000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 59.940000 60.895000 60.260000 ;
      LAYER met4 ;
        RECT 60.575000 59.940000 60.895000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 60.350000 60.895000 60.670000 ;
      LAYER met4 ;
        RECT 60.575000 60.350000 60.895000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 56.250000 61.300000 56.570000 ;
      LAYER met4 ;
        RECT 60.980000 56.250000 61.300000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 56.660000 61.300000 56.980000 ;
      LAYER met4 ;
        RECT 60.980000 56.660000 61.300000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 57.070000 61.300000 57.390000 ;
      LAYER met4 ;
        RECT 60.980000 57.070000 61.300000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 57.480000 61.300000 57.800000 ;
      LAYER met4 ;
        RECT 60.980000 57.480000 61.300000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 57.890000 61.300000 58.210000 ;
      LAYER met4 ;
        RECT 60.980000 57.890000 61.300000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 58.300000 61.300000 58.620000 ;
      LAYER met4 ;
        RECT 60.980000 58.300000 61.300000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 58.710000 61.300000 59.030000 ;
      LAYER met4 ;
        RECT 60.980000 58.710000 61.300000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 59.120000 61.300000 59.440000 ;
      LAYER met4 ;
        RECT 60.980000 59.120000 61.300000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 59.530000 61.300000 59.850000 ;
      LAYER met4 ;
        RECT 60.980000 59.530000 61.300000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 59.940000 61.300000 60.260000 ;
      LAYER met4 ;
        RECT 60.980000 59.940000 61.300000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 60.350000 61.300000 60.670000 ;
      LAYER met4 ;
        RECT 60.980000 60.350000 61.300000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 56.250000 61.705000 56.570000 ;
      LAYER met4 ;
        RECT 61.385000 56.250000 61.705000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 56.660000 61.705000 56.980000 ;
      LAYER met4 ;
        RECT 61.385000 56.660000 61.705000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 57.070000 61.705000 57.390000 ;
      LAYER met4 ;
        RECT 61.385000 57.070000 61.705000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 57.480000 61.705000 57.800000 ;
      LAYER met4 ;
        RECT 61.385000 57.480000 61.705000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 57.890000 61.705000 58.210000 ;
      LAYER met4 ;
        RECT 61.385000 57.890000 61.705000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 58.300000 61.705000 58.620000 ;
      LAYER met4 ;
        RECT 61.385000 58.300000 61.705000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 58.710000 61.705000 59.030000 ;
      LAYER met4 ;
        RECT 61.385000 58.710000 61.705000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 59.120000 61.705000 59.440000 ;
      LAYER met4 ;
        RECT 61.385000 59.120000 61.705000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 59.530000 61.705000 59.850000 ;
      LAYER met4 ;
        RECT 61.385000 59.530000 61.705000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 59.940000 61.705000 60.260000 ;
      LAYER met4 ;
        RECT 61.385000 59.940000 61.705000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 60.350000 61.705000 60.670000 ;
      LAYER met4 ;
        RECT 61.385000 60.350000 61.705000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 56.250000 62.110000 56.570000 ;
      LAYER met4 ;
        RECT 61.790000 56.250000 62.110000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 56.660000 62.110000 56.980000 ;
      LAYER met4 ;
        RECT 61.790000 56.660000 62.110000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 57.070000 62.110000 57.390000 ;
      LAYER met4 ;
        RECT 61.790000 57.070000 62.110000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 57.480000 62.110000 57.800000 ;
      LAYER met4 ;
        RECT 61.790000 57.480000 62.110000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 57.890000 62.110000 58.210000 ;
      LAYER met4 ;
        RECT 61.790000 57.890000 62.110000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 58.300000 62.110000 58.620000 ;
      LAYER met4 ;
        RECT 61.790000 58.300000 62.110000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 58.710000 62.110000 59.030000 ;
      LAYER met4 ;
        RECT 61.790000 58.710000 62.110000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 59.120000 62.110000 59.440000 ;
      LAYER met4 ;
        RECT 61.790000 59.120000 62.110000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 59.530000 62.110000 59.850000 ;
      LAYER met4 ;
        RECT 61.790000 59.530000 62.110000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 59.940000 62.110000 60.260000 ;
      LAYER met4 ;
        RECT 61.790000 59.940000 62.110000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 60.350000 62.110000 60.670000 ;
      LAYER met4 ;
        RECT 61.790000 60.350000 62.110000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 56.250000 62.515000 56.570000 ;
      LAYER met4 ;
        RECT 62.195000 56.250000 62.515000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 56.660000 62.515000 56.980000 ;
      LAYER met4 ;
        RECT 62.195000 56.660000 62.515000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 57.070000 62.515000 57.390000 ;
      LAYER met4 ;
        RECT 62.195000 57.070000 62.515000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 57.480000 62.515000 57.800000 ;
      LAYER met4 ;
        RECT 62.195000 57.480000 62.515000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 57.890000 62.515000 58.210000 ;
      LAYER met4 ;
        RECT 62.195000 57.890000 62.515000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 58.300000 62.515000 58.620000 ;
      LAYER met4 ;
        RECT 62.195000 58.300000 62.515000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 58.710000 62.515000 59.030000 ;
      LAYER met4 ;
        RECT 62.195000 58.710000 62.515000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 59.120000 62.515000 59.440000 ;
      LAYER met4 ;
        RECT 62.195000 59.120000 62.515000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 59.530000 62.515000 59.850000 ;
      LAYER met4 ;
        RECT 62.195000 59.530000 62.515000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 59.940000 62.515000 60.260000 ;
      LAYER met4 ;
        RECT 62.195000 59.940000 62.515000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 60.350000 62.515000 60.670000 ;
      LAYER met4 ;
        RECT 62.195000 60.350000 62.515000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 56.250000 62.920000 56.570000 ;
      LAYER met4 ;
        RECT 62.600000 56.250000 62.920000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 56.660000 62.920000 56.980000 ;
      LAYER met4 ;
        RECT 62.600000 56.660000 62.920000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 57.070000 62.920000 57.390000 ;
      LAYER met4 ;
        RECT 62.600000 57.070000 62.920000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 57.480000 62.920000 57.800000 ;
      LAYER met4 ;
        RECT 62.600000 57.480000 62.920000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 57.890000 62.920000 58.210000 ;
      LAYER met4 ;
        RECT 62.600000 57.890000 62.920000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 58.300000 62.920000 58.620000 ;
      LAYER met4 ;
        RECT 62.600000 58.300000 62.920000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 58.710000 62.920000 59.030000 ;
      LAYER met4 ;
        RECT 62.600000 58.710000 62.920000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 59.120000 62.920000 59.440000 ;
      LAYER met4 ;
        RECT 62.600000 59.120000 62.920000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 59.530000 62.920000 59.850000 ;
      LAYER met4 ;
        RECT 62.600000 59.530000 62.920000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 59.940000 62.920000 60.260000 ;
      LAYER met4 ;
        RECT 62.600000 59.940000 62.920000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 60.350000 62.920000 60.670000 ;
      LAYER met4 ;
        RECT 62.600000 60.350000 62.920000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 56.250000 63.325000 56.570000 ;
      LAYER met4 ;
        RECT 63.005000 56.250000 63.325000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 56.660000 63.325000 56.980000 ;
      LAYER met4 ;
        RECT 63.005000 56.660000 63.325000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 57.070000 63.325000 57.390000 ;
      LAYER met4 ;
        RECT 63.005000 57.070000 63.325000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 57.480000 63.325000 57.800000 ;
      LAYER met4 ;
        RECT 63.005000 57.480000 63.325000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 57.890000 63.325000 58.210000 ;
      LAYER met4 ;
        RECT 63.005000 57.890000 63.325000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 58.300000 63.325000 58.620000 ;
      LAYER met4 ;
        RECT 63.005000 58.300000 63.325000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 58.710000 63.325000 59.030000 ;
      LAYER met4 ;
        RECT 63.005000 58.710000 63.325000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 59.120000 63.325000 59.440000 ;
      LAYER met4 ;
        RECT 63.005000 59.120000 63.325000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 59.530000 63.325000 59.850000 ;
      LAYER met4 ;
        RECT 63.005000 59.530000 63.325000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 59.940000 63.325000 60.260000 ;
      LAYER met4 ;
        RECT 63.005000 59.940000 63.325000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 60.350000 63.325000 60.670000 ;
      LAYER met4 ;
        RECT 63.005000 60.350000 63.325000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 56.250000 63.730000 56.570000 ;
      LAYER met4 ;
        RECT 63.410000 56.250000 63.730000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 56.660000 63.730000 56.980000 ;
      LAYER met4 ;
        RECT 63.410000 56.660000 63.730000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 57.070000 63.730000 57.390000 ;
      LAYER met4 ;
        RECT 63.410000 57.070000 63.730000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 57.480000 63.730000 57.800000 ;
      LAYER met4 ;
        RECT 63.410000 57.480000 63.730000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 57.890000 63.730000 58.210000 ;
      LAYER met4 ;
        RECT 63.410000 57.890000 63.730000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 58.300000 63.730000 58.620000 ;
      LAYER met4 ;
        RECT 63.410000 58.300000 63.730000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 58.710000 63.730000 59.030000 ;
      LAYER met4 ;
        RECT 63.410000 58.710000 63.730000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 59.120000 63.730000 59.440000 ;
      LAYER met4 ;
        RECT 63.410000 59.120000 63.730000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 59.530000 63.730000 59.850000 ;
      LAYER met4 ;
        RECT 63.410000 59.530000 63.730000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 59.940000 63.730000 60.260000 ;
      LAYER met4 ;
        RECT 63.410000 59.940000 63.730000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 60.350000 63.730000 60.670000 ;
      LAYER met4 ;
        RECT 63.410000 60.350000 63.730000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 56.250000 64.135000 56.570000 ;
      LAYER met4 ;
        RECT 63.815000 56.250000 64.135000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 56.660000 64.135000 56.980000 ;
      LAYER met4 ;
        RECT 63.815000 56.660000 64.135000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 57.070000 64.135000 57.390000 ;
      LAYER met4 ;
        RECT 63.815000 57.070000 64.135000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 57.480000 64.135000 57.800000 ;
      LAYER met4 ;
        RECT 63.815000 57.480000 64.135000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 57.890000 64.135000 58.210000 ;
      LAYER met4 ;
        RECT 63.815000 57.890000 64.135000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 58.300000 64.135000 58.620000 ;
      LAYER met4 ;
        RECT 63.815000 58.300000 64.135000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 58.710000 64.135000 59.030000 ;
      LAYER met4 ;
        RECT 63.815000 58.710000 64.135000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 59.120000 64.135000 59.440000 ;
      LAYER met4 ;
        RECT 63.815000 59.120000 64.135000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 59.530000 64.135000 59.850000 ;
      LAYER met4 ;
        RECT 63.815000 59.530000 64.135000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 59.940000 64.135000 60.260000 ;
      LAYER met4 ;
        RECT 63.815000 59.940000 64.135000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 60.350000 64.135000 60.670000 ;
      LAYER met4 ;
        RECT 63.815000 60.350000 64.135000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 56.250000 64.540000 56.570000 ;
      LAYER met4 ;
        RECT 64.220000 56.250000 64.540000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 56.660000 64.540000 56.980000 ;
      LAYER met4 ;
        RECT 64.220000 56.660000 64.540000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 57.070000 64.540000 57.390000 ;
      LAYER met4 ;
        RECT 64.220000 57.070000 64.540000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 57.480000 64.540000 57.800000 ;
      LAYER met4 ;
        RECT 64.220000 57.480000 64.540000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 57.890000 64.540000 58.210000 ;
      LAYER met4 ;
        RECT 64.220000 57.890000 64.540000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 58.300000 64.540000 58.620000 ;
      LAYER met4 ;
        RECT 64.220000 58.300000 64.540000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 58.710000 64.540000 59.030000 ;
      LAYER met4 ;
        RECT 64.220000 58.710000 64.540000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 59.120000 64.540000 59.440000 ;
      LAYER met4 ;
        RECT 64.220000 59.120000 64.540000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 59.530000 64.540000 59.850000 ;
      LAYER met4 ;
        RECT 64.220000 59.530000 64.540000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 59.940000 64.540000 60.260000 ;
      LAYER met4 ;
        RECT 64.220000 59.940000 64.540000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 60.350000 64.540000 60.670000 ;
      LAYER met4 ;
        RECT 64.220000 60.350000 64.540000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 56.250000 64.945000 56.570000 ;
      LAYER met4 ;
        RECT 64.625000 56.250000 64.945000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 56.660000 64.945000 56.980000 ;
      LAYER met4 ;
        RECT 64.625000 56.660000 64.945000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 57.070000 64.945000 57.390000 ;
      LAYER met4 ;
        RECT 64.625000 57.070000 64.945000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 57.480000 64.945000 57.800000 ;
      LAYER met4 ;
        RECT 64.625000 57.480000 64.945000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 57.890000 64.945000 58.210000 ;
      LAYER met4 ;
        RECT 64.625000 57.890000 64.945000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 58.300000 64.945000 58.620000 ;
      LAYER met4 ;
        RECT 64.625000 58.300000 64.945000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 58.710000 64.945000 59.030000 ;
      LAYER met4 ;
        RECT 64.625000 58.710000 64.945000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 59.120000 64.945000 59.440000 ;
      LAYER met4 ;
        RECT 64.625000 59.120000 64.945000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 59.530000 64.945000 59.850000 ;
      LAYER met4 ;
        RECT 64.625000 59.530000 64.945000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 59.940000 64.945000 60.260000 ;
      LAYER met4 ;
        RECT 64.625000 59.940000 64.945000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 60.350000 64.945000 60.670000 ;
      LAYER met4 ;
        RECT 64.625000 60.350000 64.945000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 56.250000 65.350000 56.570000 ;
      LAYER met4 ;
        RECT 65.030000 56.250000 65.350000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 56.660000 65.350000 56.980000 ;
      LAYER met4 ;
        RECT 65.030000 56.660000 65.350000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 57.070000 65.350000 57.390000 ;
      LAYER met4 ;
        RECT 65.030000 57.070000 65.350000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 57.480000 65.350000 57.800000 ;
      LAYER met4 ;
        RECT 65.030000 57.480000 65.350000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 57.890000 65.350000 58.210000 ;
      LAYER met4 ;
        RECT 65.030000 57.890000 65.350000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 58.300000 65.350000 58.620000 ;
      LAYER met4 ;
        RECT 65.030000 58.300000 65.350000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 58.710000 65.350000 59.030000 ;
      LAYER met4 ;
        RECT 65.030000 58.710000 65.350000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 59.120000 65.350000 59.440000 ;
      LAYER met4 ;
        RECT 65.030000 59.120000 65.350000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 59.530000 65.350000 59.850000 ;
      LAYER met4 ;
        RECT 65.030000 59.530000 65.350000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 59.940000 65.350000 60.260000 ;
      LAYER met4 ;
        RECT 65.030000 59.940000 65.350000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 60.350000 65.350000 60.670000 ;
      LAYER met4 ;
        RECT 65.030000 60.350000 65.350000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 56.250000 65.755000 56.570000 ;
      LAYER met4 ;
        RECT 65.435000 56.250000 65.755000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 56.660000 65.755000 56.980000 ;
      LAYER met4 ;
        RECT 65.435000 56.660000 65.755000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 57.070000 65.755000 57.390000 ;
      LAYER met4 ;
        RECT 65.435000 57.070000 65.755000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 57.480000 65.755000 57.800000 ;
      LAYER met4 ;
        RECT 65.435000 57.480000 65.755000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 57.890000 65.755000 58.210000 ;
      LAYER met4 ;
        RECT 65.435000 57.890000 65.755000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 58.300000 65.755000 58.620000 ;
      LAYER met4 ;
        RECT 65.435000 58.300000 65.755000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 58.710000 65.755000 59.030000 ;
      LAYER met4 ;
        RECT 65.435000 58.710000 65.755000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 59.120000 65.755000 59.440000 ;
      LAYER met4 ;
        RECT 65.435000 59.120000 65.755000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 59.530000 65.755000 59.850000 ;
      LAYER met4 ;
        RECT 65.435000 59.530000 65.755000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 59.940000 65.755000 60.260000 ;
      LAYER met4 ;
        RECT 65.435000 59.940000 65.755000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 60.350000 65.755000 60.670000 ;
      LAYER met4 ;
        RECT 65.435000 60.350000 65.755000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 56.250000 66.160000 56.570000 ;
      LAYER met4 ;
        RECT 65.840000 56.250000 66.160000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 56.660000 66.160000 56.980000 ;
      LAYER met4 ;
        RECT 65.840000 56.660000 66.160000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 57.070000 66.160000 57.390000 ;
      LAYER met4 ;
        RECT 65.840000 57.070000 66.160000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 57.480000 66.160000 57.800000 ;
      LAYER met4 ;
        RECT 65.840000 57.480000 66.160000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 57.890000 66.160000 58.210000 ;
      LAYER met4 ;
        RECT 65.840000 57.890000 66.160000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 58.300000 66.160000 58.620000 ;
      LAYER met4 ;
        RECT 65.840000 58.300000 66.160000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 58.710000 66.160000 59.030000 ;
      LAYER met4 ;
        RECT 65.840000 58.710000 66.160000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 59.120000 66.160000 59.440000 ;
      LAYER met4 ;
        RECT 65.840000 59.120000 66.160000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 59.530000 66.160000 59.850000 ;
      LAYER met4 ;
        RECT 65.840000 59.530000 66.160000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 59.940000 66.160000 60.260000 ;
      LAYER met4 ;
        RECT 65.840000 59.940000 66.160000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 60.350000 66.160000 60.670000 ;
      LAYER met4 ;
        RECT 65.840000 60.350000 66.160000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 56.250000 66.565000 56.570000 ;
      LAYER met4 ;
        RECT 66.245000 56.250000 66.565000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 56.660000 66.565000 56.980000 ;
      LAYER met4 ;
        RECT 66.245000 56.660000 66.565000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 57.070000 66.565000 57.390000 ;
      LAYER met4 ;
        RECT 66.245000 57.070000 66.565000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 57.480000 66.565000 57.800000 ;
      LAYER met4 ;
        RECT 66.245000 57.480000 66.565000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 57.890000 66.565000 58.210000 ;
      LAYER met4 ;
        RECT 66.245000 57.890000 66.565000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 58.300000 66.565000 58.620000 ;
      LAYER met4 ;
        RECT 66.245000 58.300000 66.565000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 58.710000 66.565000 59.030000 ;
      LAYER met4 ;
        RECT 66.245000 58.710000 66.565000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 59.120000 66.565000 59.440000 ;
      LAYER met4 ;
        RECT 66.245000 59.120000 66.565000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 59.530000 66.565000 59.850000 ;
      LAYER met4 ;
        RECT 66.245000 59.530000 66.565000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 59.940000 66.565000 60.260000 ;
      LAYER met4 ;
        RECT 66.245000 59.940000 66.565000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 60.350000 66.565000 60.670000 ;
      LAYER met4 ;
        RECT 66.245000 60.350000 66.565000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 56.250000 66.970000 56.570000 ;
      LAYER met4 ;
        RECT 66.650000 56.250000 66.970000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 56.660000 66.970000 56.980000 ;
      LAYER met4 ;
        RECT 66.650000 56.660000 66.970000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 57.070000 66.970000 57.390000 ;
      LAYER met4 ;
        RECT 66.650000 57.070000 66.970000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 57.480000 66.970000 57.800000 ;
      LAYER met4 ;
        RECT 66.650000 57.480000 66.970000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 57.890000 66.970000 58.210000 ;
      LAYER met4 ;
        RECT 66.650000 57.890000 66.970000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 58.300000 66.970000 58.620000 ;
      LAYER met4 ;
        RECT 66.650000 58.300000 66.970000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 58.710000 66.970000 59.030000 ;
      LAYER met4 ;
        RECT 66.650000 58.710000 66.970000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 59.120000 66.970000 59.440000 ;
      LAYER met4 ;
        RECT 66.650000 59.120000 66.970000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 59.530000 66.970000 59.850000 ;
      LAYER met4 ;
        RECT 66.650000 59.530000 66.970000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 59.940000 66.970000 60.260000 ;
      LAYER met4 ;
        RECT 66.650000 59.940000 66.970000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 60.350000 66.970000 60.670000 ;
      LAYER met4 ;
        RECT 66.650000 60.350000 66.970000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 56.250000 67.375000 56.570000 ;
      LAYER met4 ;
        RECT 67.055000 56.250000 67.375000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 56.660000 67.375000 56.980000 ;
      LAYER met4 ;
        RECT 67.055000 56.660000 67.375000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 57.070000 67.375000 57.390000 ;
      LAYER met4 ;
        RECT 67.055000 57.070000 67.375000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 57.480000 67.375000 57.800000 ;
      LAYER met4 ;
        RECT 67.055000 57.480000 67.375000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 57.890000 67.375000 58.210000 ;
      LAYER met4 ;
        RECT 67.055000 57.890000 67.375000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 58.300000 67.375000 58.620000 ;
      LAYER met4 ;
        RECT 67.055000 58.300000 67.375000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 58.710000 67.375000 59.030000 ;
      LAYER met4 ;
        RECT 67.055000 58.710000 67.375000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 59.120000 67.375000 59.440000 ;
      LAYER met4 ;
        RECT 67.055000 59.120000 67.375000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 59.530000 67.375000 59.850000 ;
      LAYER met4 ;
        RECT 67.055000 59.530000 67.375000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 59.940000 67.375000 60.260000 ;
      LAYER met4 ;
        RECT 67.055000 59.940000 67.375000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 60.350000 67.375000 60.670000 ;
      LAYER met4 ;
        RECT 67.055000 60.350000 67.375000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 56.250000 67.780000 56.570000 ;
      LAYER met4 ;
        RECT 67.460000 56.250000 67.780000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 56.660000 67.780000 56.980000 ;
      LAYER met4 ;
        RECT 67.460000 56.660000 67.780000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 57.070000 67.780000 57.390000 ;
      LAYER met4 ;
        RECT 67.460000 57.070000 67.780000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 57.480000 67.780000 57.800000 ;
      LAYER met4 ;
        RECT 67.460000 57.480000 67.780000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 57.890000 67.780000 58.210000 ;
      LAYER met4 ;
        RECT 67.460000 57.890000 67.780000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 58.300000 67.780000 58.620000 ;
      LAYER met4 ;
        RECT 67.460000 58.300000 67.780000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 58.710000 67.780000 59.030000 ;
      LAYER met4 ;
        RECT 67.460000 58.710000 67.780000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 59.120000 67.780000 59.440000 ;
      LAYER met4 ;
        RECT 67.460000 59.120000 67.780000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 59.530000 67.780000 59.850000 ;
      LAYER met4 ;
        RECT 67.460000 59.530000 67.780000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 59.940000 67.780000 60.260000 ;
      LAYER met4 ;
        RECT 67.460000 59.940000 67.780000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 60.350000 67.780000 60.670000 ;
      LAYER met4 ;
        RECT 67.460000 60.350000 67.780000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 56.250000 68.185000 56.570000 ;
      LAYER met4 ;
        RECT 67.865000 56.250000 68.185000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 56.660000 68.185000 56.980000 ;
      LAYER met4 ;
        RECT 67.865000 56.660000 68.185000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 57.070000 68.185000 57.390000 ;
      LAYER met4 ;
        RECT 67.865000 57.070000 68.185000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 57.480000 68.185000 57.800000 ;
      LAYER met4 ;
        RECT 67.865000 57.480000 68.185000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 57.890000 68.185000 58.210000 ;
      LAYER met4 ;
        RECT 67.865000 57.890000 68.185000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 58.300000 68.185000 58.620000 ;
      LAYER met4 ;
        RECT 67.865000 58.300000 68.185000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 58.710000 68.185000 59.030000 ;
      LAYER met4 ;
        RECT 67.865000 58.710000 68.185000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 59.120000 68.185000 59.440000 ;
      LAYER met4 ;
        RECT 67.865000 59.120000 68.185000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 59.530000 68.185000 59.850000 ;
      LAYER met4 ;
        RECT 67.865000 59.530000 68.185000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 59.940000 68.185000 60.260000 ;
      LAYER met4 ;
        RECT 67.865000 59.940000 68.185000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 60.350000 68.185000 60.670000 ;
      LAYER met4 ;
        RECT 67.865000 60.350000 68.185000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 56.250000 68.590000 56.570000 ;
      LAYER met4 ;
        RECT 68.270000 56.250000 68.590000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 56.660000 68.590000 56.980000 ;
      LAYER met4 ;
        RECT 68.270000 56.660000 68.590000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 57.070000 68.590000 57.390000 ;
      LAYER met4 ;
        RECT 68.270000 57.070000 68.590000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 57.480000 68.590000 57.800000 ;
      LAYER met4 ;
        RECT 68.270000 57.480000 68.590000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 57.890000 68.590000 58.210000 ;
      LAYER met4 ;
        RECT 68.270000 57.890000 68.590000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 58.300000 68.590000 58.620000 ;
      LAYER met4 ;
        RECT 68.270000 58.300000 68.590000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 58.710000 68.590000 59.030000 ;
      LAYER met4 ;
        RECT 68.270000 58.710000 68.590000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 59.120000 68.590000 59.440000 ;
      LAYER met4 ;
        RECT 68.270000 59.120000 68.590000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 59.530000 68.590000 59.850000 ;
      LAYER met4 ;
        RECT 68.270000 59.530000 68.590000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 59.940000 68.590000 60.260000 ;
      LAYER met4 ;
        RECT 68.270000 59.940000 68.590000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 60.350000 68.590000 60.670000 ;
      LAYER met4 ;
        RECT 68.270000 60.350000 68.590000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 56.250000 68.995000 56.570000 ;
      LAYER met4 ;
        RECT 68.675000 56.250000 68.995000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 56.660000 68.995000 56.980000 ;
      LAYER met4 ;
        RECT 68.675000 56.660000 68.995000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 57.070000 68.995000 57.390000 ;
      LAYER met4 ;
        RECT 68.675000 57.070000 68.995000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 57.480000 68.995000 57.800000 ;
      LAYER met4 ;
        RECT 68.675000 57.480000 68.995000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 57.890000 68.995000 58.210000 ;
      LAYER met4 ;
        RECT 68.675000 57.890000 68.995000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 58.300000 68.995000 58.620000 ;
      LAYER met4 ;
        RECT 68.675000 58.300000 68.995000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 58.710000 68.995000 59.030000 ;
      LAYER met4 ;
        RECT 68.675000 58.710000 68.995000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 59.120000 68.995000 59.440000 ;
      LAYER met4 ;
        RECT 68.675000 59.120000 68.995000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 59.530000 68.995000 59.850000 ;
      LAYER met4 ;
        RECT 68.675000 59.530000 68.995000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 59.940000 68.995000 60.260000 ;
      LAYER met4 ;
        RECT 68.675000 59.940000 68.995000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 60.350000 68.995000 60.670000 ;
      LAYER met4 ;
        RECT 68.675000 60.350000 68.995000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 56.250000 69.400000 56.570000 ;
      LAYER met4 ;
        RECT 69.080000 56.250000 69.400000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 56.660000 69.400000 56.980000 ;
      LAYER met4 ;
        RECT 69.080000 56.660000 69.400000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 57.070000 69.400000 57.390000 ;
      LAYER met4 ;
        RECT 69.080000 57.070000 69.400000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 57.480000 69.400000 57.800000 ;
      LAYER met4 ;
        RECT 69.080000 57.480000 69.400000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 57.890000 69.400000 58.210000 ;
      LAYER met4 ;
        RECT 69.080000 57.890000 69.400000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 58.300000 69.400000 58.620000 ;
      LAYER met4 ;
        RECT 69.080000 58.300000 69.400000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 58.710000 69.400000 59.030000 ;
      LAYER met4 ;
        RECT 69.080000 58.710000 69.400000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 59.120000 69.400000 59.440000 ;
      LAYER met4 ;
        RECT 69.080000 59.120000 69.400000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 59.530000 69.400000 59.850000 ;
      LAYER met4 ;
        RECT 69.080000 59.530000 69.400000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 59.940000 69.400000 60.260000 ;
      LAYER met4 ;
        RECT 69.080000 59.940000 69.400000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 60.350000 69.400000 60.670000 ;
      LAYER met4 ;
        RECT 69.080000 60.350000 69.400000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 56.250000 69.805000 56.570000 ;
      LAYER met4 ;
        RECT 69.485000 56.250000 69.805000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 56.660000 69.805000 56.980000 ;
      LAYER met4 ;
        RECT 69.485000 56.660000 69.805000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 57.070000 69.805000 57.390000 ;
      LAYER met4 ;
        RECT 69.485000 57.070000 69.805000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 57.480000 69.805000 57.800000 ;
      LAYER met4 ;
        RECT 69.485000 57.480000 69.805000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 57.890000 69.805000 58.210000 ;
      LAYER met4 ;
        RECT 69.485000 57.890000 69.805000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 58.300000 69.805000 58.620000 ;
      LAYER met4 ;
        RECT 69.485000 58.300000 69.805000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 58.710000 69.805000 59.030000 ;
      LAYER met4 ;
        RECT 69.485000 58.710000 69.805000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 59.120000 69.805000 59.440000 ;
      LAYER met4 ;
        RECT 69.485000 59.120000 69.805000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 59.530000 69.805000 59.850000 ;
      LAYER met4 ;
        RECT 69.485000 59.530000 69.805000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 59.940000 69.805000 60.260000 ;
      LAYER met4 ;
        RECT 69.485000 59.940000 69.805000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 60.350000 69.805000 60.670000 ;
      LAYER met4 ;
        RECT 69.485000 60.350000 69.805000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 56.250000 70.210000 56.570000 ;
      LAYER met4 ;
        RECT 69.890000 56.250000 70.210000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 56.660000 70.210000 56.980000 ;
      LAYER met4 ;
        RECT 69.890000 56.660000 70.210000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 57.070000 70.210000 57.390000 ;
      LAYER met4 ;
        RECT 69.890000 57.070000 70.210000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 57.480000 70.210000 57.800000 ;
      LAYER met4 ;
        RECT 69.890000 57.480000 70.210000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 57.890000 70.210000 58.210000 ;
      LAYER met4 ;
        RECT 69.890000 57.890000 70.210000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 58.300000 70.210000 58.620000 ;
      LAYER met4 ;
        RECT 69.890000 58.300000 70.210000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 58.710000 70.210000 59.030000 ;
      LAYER met4 ;
        RECT 69.890000 58.710000 70.210000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 59.120000 70.210000 59.440000 ;
      LAYER met4 ;
        RECT 69.890000 59.120000 70.210000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 59.530000 70.210000 59.850000 ;
      LAYER met4 ;
        RECT 69.890000 59.530000 70.210000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 59.940000 70.210000 60.260000 ;
      LAYER met4 ;
        RECT 69.890000 59.940000 70.210000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 60.350000 70.210000 60.670000 ;
      LAYER met4 ;
        RECT 69.890000 60.350000 70.210000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 56.250000 7.360000 56.570000 ;
      LAYER met4 ;
        RECT 7.040000 56.250000 7.360000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 56.660000 7.360000 56.980000 ;
      LAYER met4 ;
        RECT 7.040000 56.660000 7.360000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 57.070000 7.360000 57.390000 ;
      LAYER met4 ;
        RECT 7.040000 57.070000 7.360000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 57.480000 7.360000 57.800000 ;
      LAYER met4 ;
        RECT 7.040000 57.480000 7.360000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 57.890000 7.360000 58.210000 ;
      LAYER met4 ;
        RECT 7.040000 57.890000 7.360000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 58.300000 7.360000 58.620000 ;
      LAYER met4 ;
        RECT 7.040000 58.300000 7.360000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 58.710000 7.360000 59.030000 ;
      LAYER met4 ;
        RECT 7.040000 58.710000 7.360000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 59.120000 7.360000 59.440000 ;
      LAYER met4 ;
        RECT 7.040000 59.120000 7.360000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 59.530000 7.360000 59.850000 ;
      LAYER met4 ;
        RECT 7.040000 59.530000 7.360000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 59.940000 7.360000 60.260000 ;
      LAYER met4 ;
        RECT 7.040000 59.940000 7.360000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 60.350000 7.360000 60.670000 ;
      LAYER met4 ;
        RECT 7.040000 60.350000 7.360000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 56.250000 7.765000 56.570000 ;
      LAYER met4 ;
        RECT 7.445000 56.250000 7.765000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 56.660000 7.765000 56.980000 ;
      LAYER met4 ;
        RECT 7.445000 56.660000 7.765000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 57.070000 7.765000 57.390000 ;
      LAYER met4 ;
        RECT 7.445000 57.070000 7.765000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 57.480000 7.765000 57.800000 ;
      LAYER met4 ;
        RECT 7.445000 57.480000 7.765000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 57.890000 7.765000 58.210000 ;
      LAYER met4 ;
        RECT 7.445000 57.890000 7.765000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 58.300000 7.765000 58.620000 ;
      LAYER met4 ;
        RECT 7.445000 58.300000 7.765000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 58.710000 7.765000 59.030000 ;
      LAYER met4 ;
        RECT 7.445000 58.710000 7.765000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 59.120000 7.765000 59.440000 ;
      LAYER met4 ;
        RECT 7.445000 59.120000 7.765000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 59.530000 7.765000 59.850000 ;
      LAYER met4 ;
        RECT 7.445000 59.530000 7.765000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 59.940000 7.765000 60.260000 ;
      LAYER met4 ;
        RECT 7.445000 59.940000 7.765000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 60.350000 7.765000 60.670000 ;
      LAYER met4 ;
        RECT 7.445000 60.350000 7.765000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 56.250000 8.170000 56.570000 ;
      LAYER met4 ;
        RECT 7.850000 56.250000 8.170000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 56.660000 8.170000 56.980000 ;
      LAYER met4 ;
        RECT 7.850000 56.660000 8.170000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 57.070000 8.170000 57.390000 ;
      LAYER met4 ;
        RECT 7.850000 57.070000 8.170000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 57.480000 8.170000 57.800000 ;
      LAYER met4 ;
        RECT 7.850000 57.480000 8.170000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 57.890000 8.170000 58.210000 ;
      LAYER met4 ;
        RECT 7.850000 57.890000 8.170000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 58.300000 8.170000 58.620000 ;
      LAYER met4 ;
        RECT 7.850000 58.300000 8.170000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 58.710000 8.170000 59.030000 ;
      LAYER met4 ;
        RECT 7.850000 58.710000 8.170000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 59.120000 8.170000 59.440000 ;
      LAYER met4 ;
        RECT 7.850000 59.120000 8.170000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 59.530000 8.170000 59.850000 ;
      LAYER met4 ;
        RECT 7.850000 59.530000 8.170000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 59.940000 8.170000 60.260000 ;
      LAYER met4 ;
        RECT 7.850000 59.940000 8.170000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 60.350000 8.170000 60.670000 ;
      LAYER met4 ;
        RECT 7.850000 60.350000 8.170000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 56.250000 70.615000 56.570000 ;
      LAYER met4 ;
        RECT 70.295000 56.250000 70.615000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 56.660000 70.615000 56.980000 ;
      LAYER met4 ;
        RECT 70.295000 56.660000 70.615000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 57.070000 70.615000 57.390000 ;
      LAYER met4 ;
        RECT 70.295000 57.070000 70.615000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 57.480000 70.615000 57.800000 ;
      LAYER met4 ;
        RECT 70.295000 57.480000 70.615000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 57.890000 70.615000 58.210000 ;
      LAYER met4 ;
        RECT 70.295000 57.890000 70.615000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 58.300000 70.615000 58.620000 ;
      LAYER met4 ;
        RECT 70.295000 58.300000 70.615000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 58.710000 70.615000 59.030000 ;
      LAYER met4 ;
        RECT 70.295000 58.710000 70.615000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 59.120000 70.615000 59.440000 ;
      LAYER met4 ;
        RECT 70.295000 59.120000 70.615000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 59.530000 70.615000 59.850000 ;
      LAYER met4 ;
        RECT 70.295000 59.530000 70.615000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 59.940000 70.615000 60.260000 ;
      LAYER met4 ;
        RECT 70.295000 59.940000 70.615000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 60.350000 70.615000 60.670000 ;
      LAYER met4 ;
        RECT 70.295000 60.350000 70.615000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 56.250000 71.020000 56.570000 ;
      LAYER met4 ;
        RECT 70.700000 56.250000 71.020000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 56.660000 71.020000 56.980000 ;
      LAYER met4 ;
        RECT 70.700000 56.660000 71.020000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 57.070000 71.020000 57.390000 ;
      LAYER met4 ;
        RECT 70.700000 57.070000 71.020000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 57.480000 71.020000 57.800000 ;
      LAYER met4 ;
        RECT 70.700000 57.480000 71.020000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 57.890000 71.020000 58.210000 ;
      LAYER met4 ;
        RECT 70.700000 57.890000 71.020000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 58.300000 71.020000 58.620000 ;
      LAYER met4 ;
        RECT 70.700000 58.300000 71.020000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 58.710000 71.020000 59.030000 ;
      LAYER met4 ;
        RECT 70.700000 58.710000 71.020000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 59.120000 71.020000 59.440000 ;
      LAYER met4 ;
        RECT 70.700000 59.120000 71.020000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 59.530000 71.020000 59.850000 ;
      LAYER met4 ;
        RECT 70.700000 59.530000 71.020000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 59.940000 71.020000 60.260000 ;
      LAYER met4 ;
        RECT 70.700000 59.940000 71.020000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 60.350000 71.020000 60.670000 ;
      LAYER met4 ;
        RECT 70.700000 60.350000 71.020000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 56.250000 71.425000 56.570000 ;
      LAYER met4 ;
        RECT 71.105000 56.250000 71.425000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 56.660000 71.425000 56.980000 ;
      LAYER met4 ;
        RECT 71.105000 56.660000 71.425000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 57.070000 71.425000 57.390000 ;
      LAYER met4 ;
        RECT 71.105000 57.070000 71.425000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 57.480000 71.425000 57.800000 ;
      LAYER met4 ;
        RECT 71.105000 57.480000 71.425000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 57.890000 71.425000 58.210000 ;
      LAYER met4 ;
        RECT 71.105000 57.890000 71.425000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 58.300000 71.425000 58.620000 ;
      LAYER met4 ;
        RECT 71.105000 58.300000 71.425000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 58.710000 71.425000 59.030000 ;
      LAYER met4 ;
        RECT 71.105000 58.710000 71.425000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 59.120000 71.425000 59.440000 ;
      LAYER met4 ;
        RECT 71.105000 59.120000 71.425000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 59.530000 71.425000 59.850000 ;
      LAYER met4 ;
        RECT 71.105000 59.530000 71.425000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 59.940000 71.425000 60.260000 ;
      LAYER met4 ;
        RECT 71.105000 59.940000 71.425000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 60.350000 71.425000 60.670000 ;
      LAYER met4 ;
        RECT 71.105000 60.350000 71.425000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 56.250000 71.830000 56.570000 ;
      LAYER met4 ;
        RECT 71.510000 56.250000 71.830000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 56.660000 71.830000 56.980000 ;
      LAYER met4 ;
        RECT 71.510000 56.660000 71.830000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 57.070000 71.830000 57.390000 ;
      LAYER met4 ;
        RECT 71.510000 57.070000 71.830000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 57.480000 71.830000 57.800000 ;
      LAYER met4 ;
        RECT 71.510000 57.480000 71.830000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 57.890000 71.830000 58.210000 ;
      LAYER met4 ;
        RECT 71.510000 57.890000 71.830000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 58.300000 71.830000 58.620000 ;
      LAYER met4 ;
        RECT 71.510000 58.300000 71.830000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 58.710000 71.830000 59.030000 ;
      LAYER met4 ;
        RECT 71.510000 58.710000 71.830000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 59.120000 71.830000 59.440000 ;
      LAYER met4 ;
        RECT 71.510000 59.120000 71.830000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 59.530000 71.830000 59.850000 ;
      LAYER met4 ;
        RECT 71.510000 59.530000 71.830000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 59.940000 71.830000 60.260000 ;
      LAYER met4 ;
        RECT 71.510000 59.940000 71.830000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 60.350000 71.830000 60.670000 ;
      LAYER met4 ;
        RECT 71.510000 60.350000 71.830000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 56.250000 72.235000 56.570000 ;
      LAYER met4 ;
        RECT 71.915000 56.250000 72.235000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 56.660000 72.235000 56.980000 ;
      LAYER met4 ;
        RECT 71.915000 56.660000 72.235000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 57.070000 72.235000 57.390000 ;
      LAYER met4 ;
        RECT 71.915000 57.070000 72.235000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 57.480000 72.235000 57.800000 ;
      LAYER met4 ;
        RECT 71.915000 57.480000 72.235000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 57.890000 72.235000 58.210000 ;
      LAYER met4 ;
        RECT 71.915000 57.890000 72.235000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 58.300000 72.235000 58.620000 ;
      LAYER met4 ;
        RECT 71.915000 58.300000 72.235000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 58.710000 72.235000 59.030000 ;
      LAYER met4 ;
        RECT 71.915000 58.710000 72.235000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 59.120000 72.235000 59.440000 ;
      LAYER met4 ;
        RECT 71.915000 59.120000 72.235000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 59.530000 72.235000 59.850000 ;
      LAYER met4 ;
        RECT 71.915000 59.530000 72.235000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 59.940000 72.235000 60.260000 ;
      LAYER met4 ;
        RECT 71.915000 59.940000 72.235000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 60.350000 72.235000 60.670000 ;
      LAYER met4 ;
        RECT 71.915000 60.350000 72.235000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 56.250000 72.640000 56.570000 ;
      LAYER met4 ;
        RECT 72.320000 56.250000 72.640000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 56.660000 72.640000 56.980000 ;
      LAYER met4 ;
        RECT 72.320000 56.660000 72.640000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 57.070000 72.640000 57.390000 ;
      LAYER met4 ;
        RECT 72.320000 57.070000 72.640000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 57.480000 72.640000 57.800000 ;
      LAYER met4 ;
        RECT 72.320000 57.480000 72.640000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 57.890000 72.640000 58.210000 ;
      LAYER met4 ;
        RECT 72.320000 57.890000 72.640000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 58.300000 72.640000 58.620000 ;
      LAYER met4 ;
        RECT 72.320000 58.300000 72.640000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 58.710000 72.640000 59.030000 ;
      LAYER met4 ;
        RECT 72.320000 58.710000 72.640000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 59.120000 72.640000 59.440000 ;
      LAYER met4 ;
        RECT 72.320000 59.120000 72.640000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 59.530000 72.640000 59.850000 ;
      LAYER met4 ;
        RECT 72.320000 59.530000 72.640000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 59.940000 72.640000 60.260000 ;
      LAYER met4 ;
        RECT 72.320000 59.940000 72.640000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 60.350000 72.640000 60.670000 ;
      LAYER met4 ;
        RECT 72.320000 60.350000 72.640000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 56.250000 73.045000 56.570000 ;
      LAYER met4 ;
        RECT 72.725000 56.250000 73.045000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 56.660000 73.045000 56.980000 ;
      LAYER met4 ;
        RECT 72.725000 56.660000 73.045000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 57.070000 73.045000 57.390000 ;
      LAYER met4 ;
        RECT 72.725000 57.070000 73.045000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 57.480000 73.045000 57.800000 ;
      LAYER met4 ;
        RECT 72.725000 57.480000 73.045000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 57.890000 73.045000 58.210000 ;
      LAYER met4 ;
        RECT 72.725000 57.890000 73.045000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 58.300000 73.045000 58.620000 ;
      LAYER met4 ;
        RECT 72.725000 58.300000 73.045000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 58.710000 73.045000 59.030000 ;
      LAYER met4 ;
        RECT 72.725000 58.710000 73.045000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 59.120000 73.045000 59.440000 ;
      LAYER met4 ;
        RECT 72.725000 59.120000 73.045000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 59.530000 73.045000 59.850000 ;
      LAYER met4 ;
        RECT 72.725000 59.530000 73.045000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 59.940000 73.045000 60.260000 ;
      LAYER met4 ;
        RECT 72.725000 59.940000 73.045000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 60.350000 73.045000 60.670000 ;
      LAYER met4 ;
        RECT 72.725000 60.350000 73.045000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 56.250000 73.450000 56.570000 ;
      LAYER met4 ;
        RECT 73.130000 56.250000 73.450000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 56.660000 73.450000 56.980000 ;
      LAYER met4 ;
        RECT 73.130000 56.660000 73.450000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 57.070000 73.450000 57.390000 ;
      LAYER met4 ;
        RECT 73.130000 57.070000 73.450000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 57.480000 73.450000 57.800000 ;
      LAYER met4 ;
        RECT 73.130000 57.480000 73.450000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 57.890000 73.450000 58.210000 ;
      LAYER met4 ;
        RECT 73.130000 57.890000 73.450000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 58.300000 73.450000 58.620000 ;
      LAYER met4 ;
        RECT 73.130000 58.300000 73.450000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 58.710000 73.450000 59.030000 ;
      LAYER met4 ;
        RECT 73.130000 58.710000 73.450000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 59.120000 73.450000 59.440000 ;
      LAYER met4 ;
        RECT 73.130000 59.120000 73.450000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 59.530000 73.450000 59.850000 ;
      LAYER met4 ;
        RECT 73.130000 59.530000 73.450000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 59.940000 73.450000 60.260000 ;
      LAYER met4 ;
        RECT 73.130000 59.940000 73.450000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 60.350000 73.450000 60.670000 ;
      LAYER met4 ;
        RECT 73.130000 60.350000 73.450000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 56.250000 73.855000 56.570000 ;
      LAYER met4 ;
        RECT 73.535000 56.250000 73.855000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 56.660000 73.855000 56.980000 ;
      LAYER met4 ;
        RECT 73.535000 56.660000 73.855000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 57.070000 73.855000 57.390000 ;
      LAYER met4 ;
        RECT 73.535000 57.070000 73.855000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 57.480000 73.855000 57.800000 ;
      LAYER met4 ;
        RECT 73.535000 57.480000 73.855000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 57.890000 73.855000 58.210000 ;
      LAYER met4 ;
        RECT 73.535000 57.890000 73.855000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 58.300000 73.855000 58.620000 ;
      LAYER met4 ;
        RECT 73.535000 58.300000 73.855000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 58.710000 73.855000 59.030000 ;
      LAYER met4 ;
        RECT 73.535000 58.710000 73.855000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 59.120000 73.855000 59.440000 ;
      LAYER met4 ;
        RECT 73.535000 59.120000 73.855000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 59.530000 73.855000 59.850000 ;
      LAYER met4 ;
        RECT 73.535000 59.530000 73.855000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 59.940000 73.855000 60.260000 ;
      LAYER met4 ;
        RECT 73.535000 59.940000 73.855000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 60.350000 73.855000 60.670000 ;
      LAYER met4 ;
        RECT 73.535000 60.350000 73.855000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 56.250000 74.260000 56.570000 ;
      LAYER met4 ;
        RECT 73.940000 56.250000 74.260000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 56.660000 74.260000 56.980000 ;
      LAYER met4 ;
        RECT 73.940000 56.660000 74.260000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 57.070000 74.260000 57.390000 ;
      LAYER met4 ;
        RECT 73.940000 57.070000 74.260000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 57.480000 74.260000 57.800000 ;
      LAYER met4 ;
        RECT 73.940000 57.480000 74.260000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 57.890000 74.260000 58.210000 ;
      LAYER met4 ;
        RECT 73.940000 57.890000 74.260000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 58.300000 74.260000 58.620000 ;
      LAYER met4 ;
        RECT 73.940000 58.300000 74.260000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 58.710000 74.260000 59.030000 ;
      LAYER met4 ;
        RECT 73.940000 58.710000 74.260000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 59.120000 74.260000 59.440000 ;
      LAYER met4 ;
        RECT 73.940000 59.120000 74.260000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 59.530000 74.260000 59.850000 ;
      LAYER met4 ;
        RECT 73.940000 59.530000 74.260000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 59.940000 74.260000 60.260000 ;
      LAYER met4 ;
        RECT 73.940000 59.940000 74.260000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 60.350000 74.260000 60.670000 ;
      LAYER met4 ;
        RECT 73.940000 60.350000 74.260000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 56.250000 8.575000 56.570000 ;
      LAYER met4 ;
        RECT 8.255000 56.250000 8.575000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 56.660000 8.575000 56.980000 ;
      LAYER met4 ;
        RECT 8.255000 56.660000 8.575000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 57.070000 8.575000 57.390000 ;
      LAYER met4 ;
        RECT 8.255000 57.070000 8.575000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 57.480000 8.575000 57.800000 ;
      LAYER met4 ;
        RECT 8.255000 57.480000 8.575000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 57.890000 8.575000 58.210000 ;
      LAYER met4 ;
        RECT 8.255000 57.890000 8.575000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 58.300000 8.575000 58.620000 ;
      LAYER met4 ;
        RECT 8.255000 58.300000 8.575000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 58.710000 8.575000 59.030000 ;
      LAYER met4 ;
        RECT 8.255000 58.710000 8.575000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 59.120000 8.575000 59.440000 ;
      LAYER met4 ;
        RECT 8.255000 59.120000 8.575000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 59.530000 8.575000 59.850000 ;
      LAYER met4 ;
        RECT 8.255000 59.530000 8.575000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 59.940000 8.575000 60.260000 ;
      LAYER met4 ;
        RECT 8.255000 59.940000 8.575000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 60.350000 8.575000 60.670000 ;
      LAYER met4 ;
        RECT 8.255000 60.350000 8.575000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 56.250000 8.980000 56.570000 ;
      LAYER met4 ;
        RECT 8.660000 56.250000 8.980000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 56.660000 8.980000 56.980000 ;
      LAYER met4 ;
        RECT 8.660000 56.660000 8.980000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 57.070000 8.980000 57.390000 ;
      LAYER met4 ;
        RECT 8.660000 57.070000 8.980000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 57.480000 8.980000 57.800000 ;
      LAYER met4 ;
        RECT 8.660000 57.480000 8.980000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 57.890000 8.980000 58.210000 ;
      LAYER met4 ;
        RECT 8.660000 57.890000 8.980000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 58.300000 8.980000 58.620000 ;
      LAYER met4 ;
        RECT 8.660000 58.300000 8.980000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 58.710000 8.980000 59.030000 ;
      LAYER met4 ;
        RECT 8.660000 58.710000 8.980000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 59.120000 8.980000 59.440000 ;
      LAYER met4 ;
        RECT 8.660000 59.120000 8.980000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 59.530000 8.980000 59.850000 ;
      LAYER met4 ;
        RECT 8.660000 59.530000 8.980000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 59.940000 8.980000 60.260000 ;
      LAYER met4 ;
        RECT 8.660000 59.940000 8.980000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 60.350000 8.980000 60.670000 ;
      LAYER met4 ;
        RECT 8.660000 60.350000 8.980000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 56.250000 9.385000 56.570000 ;
      LAYER met4 ;
        RECT 9.065000 56.250000 9.385000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 56.660000 9.385000 56.980000 ;
      LAYER met4 ;
        RECT 9.065000 56.660000 9.385000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 57.070000 9.385000 57.390000 ;
      LAYER met4 ;
        RECT 9.065000 57.070000 9.385000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 57.480000 9.385000 57.800000 ;
      LAYER met4 ;
        RECT 9.065000 57.480000 9.385000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 57.890000 9.385000 58.210000 ;
      LAYER met4 ;
        RECT 9.065000 57.890000 9.385000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 58.300000 9.385000 58.620000 ;
      LAYER met4 ;
        RECT 9.065000 58.300000 9.385000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 58.710000 9.385000 59.030000 ;
      LAYER met4 ;
        RECT 9.065000 58.710000 9.385000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 59.120000 9.385000 59.440000 ;
      LAYER met4 ;
        RECT 9.065000 59.120000 9.385000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 59.530000 9.385000 59.850000 ;
      LAYER met4 ;
        RECT 9.065000 59.530000 9.385000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 59.940000 9.385000 60.260000 ;
      LAYER met4 ;
        RECT 9.065000 59.940000 9.385000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 60.350000 9.385000 60.670000 ;
      LAYER met4 ;
        RECT 9.065000 60.350000 9.385000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 56.250000 9.790000 56.570000 ;
      LAYER met4 ;
        RECT 9.470000 56.250000 9.790000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 56.660000 9.790000 56.980000 ;
      LAYER met4 ;
        RECT 9.470000 56.660000 9.790000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 57.070000 9.790000 57.390000 ;
      LAYER met4 ;
        RECT 9.470000 57.070000 9.790000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 57.480000 9.790000 57.800000 ;
      LAYER met4 ;
        RECT 9.470000 57.480000 9.790000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 57.890000 9.790000 58.210000 ;
      LAYER met4 ;
        RECT 9.470000 57.890000 9.790000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 58.300000 9.790000 58.620000 ;
      LAYER met4 ;
        RECT 9.470000 58.300000 9.790000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 58.710000 9.790000 59.030000 ;
      LAYER met4 ;
        RECT 9.470000 58.710000 9.790000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 59.120000 9.790000 59.440000 ;
      LAYER met4 ;
        RECT 9.470000 59.120000 9.790000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 59.530000 9.790000 59.850000 ;
      LAYER met4 ;
        RECT 9.470000 59.530000 9.790000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 59.940000 9.790000 60.260000 ;
      LAYER met4 ;
        RECT 9.470000 59.940000 9.790000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 60.350000 9.790000 60.670000 ;
      LAYER met4 ;
        RECT 9.470000 60.350000 9.790000 60.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 56.250000 10.195000 56.570000 ;
      LAYER met4 ;
        RECT 9.875000 56.250000 10.195000 56.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 56.660000 10.195000 56.980000 ;
      LAYER met4 ;
        RECT 9.875000 56.660000 10.195000 56.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 57.070000 10.195000 57.390000 ;
      LAYER met4 ;
        RECT 9.875000 57.070000 10.195000 57.390000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 57.480000 10.195000 57.800000 ;
      LAYER met4 ;
        RECT 9.875000 57.480000 10.195000 57.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 57.890000 10.195000 58.210000 ;
      LAYER met4 ;
        RECT 9.875000 57.890000 10.195000 58.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 58.300000 10.195000 58.620000 ;
      LAYER met4 ;
        RECT 9.875000 58.300000 10.195000 58.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 58.710000 10.195000 59.030000 ;
      LAYER met4 ;
        RECT 9.875000 58.710000 10.195000 59.030000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 59.120000 10.195000 59.440000 ;
      LAYER met4 ;
        RECT 9.875000 59.120000 10.195000 59.440000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 59.530000 10.195000 59.850000 ;
      LAYER met4 ;
        RECT 9.875000 59.530000 10.195000 59.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 59.940000 10.195000 60.260000 ;
      LAYER met4 ;
        RECT 9.875000 59.940000 10.195000 60.260000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 60.350000 10.195000 60.670000 ;
      LAYER met4 ;
        RECT 9.875000 60.350000 10.195000 60.670000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met3 ;
      RECT 0.500000 23.840000 74.700000 198.000000 ;
    LAYER met4 ;
      RECT 0.000000  0.035000 75.000000  45.965000 ;
      RECT 0.000000 49.745000 75.000000  50.725000 ;
      RECT 0.000000 54.505000 75.000000 198.000000 ;
    LAYER met5 ;
      RECT 0.000000  0.135000 72.130000  13.035000 ;
      RECT 0.000000 13.035000 72.435000  17.885000 ;
      RECT 0.000000 17.885000 75.000000  28.385000 ;
      RECT 0.000000 28.385000 72.130000  34.835000 ;
      RECT 0.000000 34.835000 75.000000  38.085000 ;
      RECT 0.000000 38.085000 72.130000  56.335000 ;
      RECT 0.000000 56.335000 75.000000  60.585000 ;
      RECT 0.000000 60.585000 72.130000  94.585000 ;
      RECT 0.000000 94.585000 75.000000 198.000000 ;
  END
END sky130_fd_io__overlay_vssio_lvc
END LIBRARY
