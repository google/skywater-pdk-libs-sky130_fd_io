# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__overlay_vssa_lvc
  CLASS BLOCK ;
  FOREIGN sky130_fd_io__overlay_vssa_lvc ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  75.00000 BY  198.0000 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.530000 34.760000 0.850000 35.080000 ;
      LAYER met4 ;
        RECT 0.530000 34.760000 0.850000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 35.200000 0.850000 35.520000 ;
      LAYER met4 ;
        RECT 0.530000 35.200000 0.850000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 35.640000 0.850000 35.960000 ;
      LAYER met4 ;
        RECT 0.530000 35.640000 0.850000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 36.080000 0.850000 36.400000 ;
      LAYER met4 ;
        RECT 0.530000 36.080000 0.850000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 36.520000 0.850000 36.840000 ;
      LAYER met4 ;
        RECT 0.530000 36.520000 0.850000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 36.960000 0.850000 37.280000 ;
      LAYER met4 ;
        RECT 0.530000 36.960000 0.850000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 37.400000 0.850000 37.720000 ;
      LAYER met4 ;
        RECT 0.530000 37.400000 0.850000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 37.840000 0.850000 38.160000 ;
      LAYER met4 ;
        RECT 0.530000 37.840000 0.850000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 49.655000 0.850000 49.975000 ;
      LAYER met4 ;
        RECT 0.530000 49.655000 0.850000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 50.075000 0.850000 50.395000 ;
      LAYER met4 ;
        RECT 0.530000 50.075000 0.850000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530000 50.495000 0.850000 50.815000 ;
      LAYER met4 ;
        RECT 0.530000 50.495000 0.850000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 34.760000 1.260000 35.080000 ;
      LAYER met4 ;
        RECT 0.940000 34.760000 1.260000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 35.200000 1.260000 35.520000 ;
      LAYER met4 ;
        RECT 0.940000 35.200000 1.260000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 35.640000 1.260000 35.960000 ;
      LAYER met4 ;
        RECT 0.940000 35.640000 1.260000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 36.080000 1.260000 36.400000 ;
      LAYER met4 ;
        RECT 0.940000 36.080000 1.260000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 36.520000 1.260000 36.840000 ;
      LAYER met4 ;
        RECT 0.940000 36.520000 1.260000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 36.960000 1.260000 37.280000 ;
      LAYER met4 ;
        RECT 0.940000 36.960000 1.260000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 37.400000 1.260000 37.720000 ;
      LAYER met4 ;
        RECT 0.940000 37.400000 1.260000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 37.840000 1.260000 38.160000 ;
      LAYER met4 ;
        RECT 0.940000 37.840000 1.260000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 49.655000 1.260000 49.975000 ;
      LAYER met4 ;
        RECT 0.940000 49.655000 1.260000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 50.075000 1.260000 50.395000 ;
      LAYER met4 ;
        RECT 0.940000 50.075000 1.260000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940000 50.495000 1.260000 50.815000 ;
      LAYER met4 ;
        RECT 0.940000 50.495000 1.260000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 34.760000 1.670000 35.080000 ;
      LAYER met4 ;
        RECT 1.350000 34.760000 1.670000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 35.200000 1.670000 35.520000 ;
      LAYER met4 ;
        RECT 1.350000 35.200000 1.670000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 35.640000 1.670000 35.960000 ;
      LAYER met4 ;
        RECT 1.350000 35.640000 1.670000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 36.080000 1.670000 36.400000 ;
      LAYER met4 ;
        RECT 1.350000 36.080000 1.670000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 36.520000 1.670000 36.840000 ;
      LAYER met4 ;
        RECT 1.350000 36.520000 1.670000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 36.960000 1.670000 37.280000 ;
      LAYER met4 ;
        RECT 1.350000 36.960000 1.670000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 37.400000 1.670000 37.720000 ;
      LAYER met4 ;
        RECT 1.350000 37.400000 1.670000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 37.840000 1.670000 38.160000 ;
      LAYER met4 ;
        RECT 1.350000 37.840000 1.670000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 49.655000 1.670000 49.975000 ;
      LAYER met4 ;
        RECT 1.350000 49.655000 1.670000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 50.075000 1.670000 50.395000 ;
      LAYER met4 ;
        RECT 1.350000 50.075000 1.670000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350000 50.495000 1.670000 50.815000 ;
      LAYER met4 ;
        RECT 1.350000 50.495000 1.670000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 34.760000 2.080000 35.080000 ;
      LAYER met4 ;
        RECT 1.760000 34.760000 2.080000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 35.200000 2.080000 35.520000 ;
      LAYER met4 ;
        RECT 1.760000 35.200000 2.080000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 35.640000 2.080000 35.960000 ;
      LAYER met4 ;
        RECT 1.760000 35.640000 2.080000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 36.080000 2.080000 36.400000 ;
      LAYER met4 ;
        RECT 1.760000 36.080000 2.080000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 36.520000 2.080000 36.840000 ;
      LAYER met4 ;
        RECT 1.760000 36.520000 2.080000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 36.960000 2.080000 37.280000 ;
      LAYER met4 ;
        RECT 1.760000 36.960000 2.080000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 37.400000 2.080000 37.720000 ;
      LAYER met4 ;
        RECT 1.760000 37.400000 2.080000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 37.840000 2.080000 38.160000 ;
      LAYER met4 ;
        RECT 1.760000 37.840000 2.080000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 49.655000 2.080000 49.975000 ;
      LAYER met4 ;
        RECT 1.760000 49.655000 2.080000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 50.075000 2.080000 50.395000 ;
      LAYER met4 ;
        RECT 1.760000 50.075000 2.080000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760000 50.495000 2.080000 50.815000 ;
      LAYER met4 ;
        RECT 1.760000 50.495000 2.080000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 34.760000 10.600000 35.080000 ;
      LAYER met4 ;
        RECT 10.280000 34.760000 10.600000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 35.200000 10.600000 35.520000 ;
      LAYER met4 ;
        RECT 10.280000 35.200000 10.600000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 35.640000 10.600000 35.960000 ;
      LAYER met4 ;
        RECT 10.280000 35.640000 10.600000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 36.080000 10.600000 36.400000 ;
      LAYER met4 ;
        RECT 10.280000 36.080000 10.600000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 36.520000 10.600000 36.840000 ;
      LAYER met4 ;
        RECT 10.280000 36.520000 10.600000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 36.960000 10.600000 37.280000 ;
      LAYER met4 ;
        RECT 10.280000 36.960000 10.600000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 37.400000 10.600000 37.720000 ;
      LAYER met4 ;
        RECT 10.280000 37.400000 10.600000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 37.840000 10.600000 38.160000 ;
      LAYER met4 ;
        RECT 10.280000 37.840000 10.600000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 49.655000 10.600000 49.975000 ;
      LAYER met4 ;
        RECT 10.280000 49.655000 10.600000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 50.075000 10.600000 50.395000 ;
      LAYER met4 ;
        RECT 10.280000 50.075000 10.600000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 50.495000 10.600000 50.815000 ;
      LAYER met4 ;
        RECT 10.280000 50.495000 10.600000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 34.760000 11.005000 35.080000 ;
      LAYER met4 ;
        RECT 10.685000 34.760000 11.005000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 35.200000 11.005000 35.520000 ;
      LAYER met4 ;
        RECT 10.685000 35.200000 11.005000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 35.640000 11.005000 35.960000 ;
      LAYER met4 ;
        RECT 10.685000 35.640000 11.005000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 36.080000 11.005000 36.400000 ;
      LAYER met4 ;
        RECT 10.685000 36.080000 11.005000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 36.520000 11.005000 36.840000 ;
      LAYER met4 ;
        RECT 10.685000 36.520000 11.005000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 36.960000 11.005000 37.280000 ;
      LAYER met4 ;
        RECT 10.685000 36.960000 11.005000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 37.400000 11.005000 37.720000 ;
      LAYER met4 ;
        RECT 10.685000 37.400000 11.005000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 37.840000 11.005000 38.160000 ;
      LAYER met4 ;
        RECT 10.685000 37.840000 11.005000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 49.655000 11.005000 49.975000 ;
      LAYER met4 ;
        RECT 10.685000 49.655000 11.005000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 50.075000 11.005000 50.395000 ;
      LAYER met4 ;
        RECT 10.685000 50.075000 11.005000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 50.495000 11.005000 50.815000 ;
      LAYER met4 ;
        RECT 10.685000 50.495000 11.005000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 34.760000 11.410000 35.080000 ;
      LAYER met4 ;
        RECT 11.090000 34.760000 11.410000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 35.200000 11.410000 35.520000 ;
      LAYER met4 ;
        RECT 11.090000 35.200000 11.410000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 35.640000 11.410000 35.960000 ;
      LAYER met4 ;
        RECT 11.090000 35.640000 11.410000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 36.080000 11.410000 36.400000 ;
      LAYER met4 ;
        RECT 11.090000 36.080000 11.410000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 36.520000 11.410000 36.840000 ;
      LAYER met4 ;
        RECT 11.090000 36.520000 11.410000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 36.960000 11.410000 37.280000 ;
      LAYER met4 ;
        RECT 11.090000 36.960000 11.410000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 37.400000 11.410000 37.720000 ;
      LAYER met4 ;
        RECT 11.090000 37.400000 11.410000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 37.840000 11.410000 38.160000 ;
      LAYER met4 ;
        RECT 11.090000 37.840000 11.410000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 49.655000 11.410000 49.975000 ;
      LAYER met4 ;
        RECT 11.090000 49.655000 11.410000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 50.075000 11.410000 50.395000 ;
      LAYER met4 ;
        RECT 11.090000 50.075000 11.410000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 50.495000 11.410000 50.815000 ;
      LAYER met4 ;
        RECT 11.090000 50.495000 11.410000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 34.760000 11.815000 35.080000 ;
      LAYER met4 ;
        RECT 11.495000 34.760000 11.815000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 35.200000 11.815000 35.520000 ;
      LAYER met4 ;
        RECT 11.495000 35.200000 11.815000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 35.640000 11.815000 35.960000 ;
      LAYER met4 ;
        RECT 11.495000 35.640000 11.815000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 36.080000 11.815000 36.400000 ;
      LAYER met4 ;
        RECT 11.495000 36.080000 11.815000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 36.520000 11.815000 36.840000 ;
      LAYER met4 ;
        RECT 11.495000 36.520000 11.815000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 36.960000 11.815000 37.280000 ;
      LAYER met4 ;
        RECT 11.495000 36.960000 11.815000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 37.400000 11.815000 37.720000 ;
      LAYER met4 ;
        RECT 11.495000 37.400000 11.815000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 37.840000 11.815000 38.160000 ;
      LAYER met4 ;
        RECT 11.495000 37.840000 11.815000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 49.655000 11.815000 49.975000 ;
      LAYER met4 ;
        RECT 11.495000 49.655000 11.815000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 50.075000 11.815000 50.395000 ;
      LAYER met4 ;
        RECT 11.495000 50.075000 11.815000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 50.495000 11.815000 50.815000 ;
      LAYER met4 ;
        RECT 11.495000 50.495000 11.815000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 34.760000 12.220000 35.080000 ;
      LAYER met4 ;
        RECT 11.900000 34.760000 12.220000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 35.200000 12.220000 35.520000 ;
      LAYER met4 ;
        RECT 11.900000 35.200000 12.220000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 35.640000 12.220000 35.960000 ;
      LAYER met4 ;
        RECT 11.900000 35.640000 12.220000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 36.080000 12.220000 36.400000 ;
      LAYER met4 ;
        RECT 11.900000 36.080000 12.220000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 36.520000 12.220000 36.840000 ;
      LAYER met4 ;
        RECT 11.900000 36.520000 12.220000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 36.960000 12.220000 37.280000 ;
      LAYER met4 ;
        RECT 11.900000 36.960000 12.220000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 37.400000 12.220000 37.720000 ;
      LAYER met4 ;
        RECT 11.900000 37.400000 12.220000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 37.840000 12.220000 38.160000 ;
      LAYER met4 ;
        RECT 11.900000 37.840000 12.220000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 49.655000 12.220000 49.975000 ;
      LAYER met4 ;
        RECT 11.900000 49.655000 12.220000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 50.075000 12.220000 50.395000 ;
      LAYER met4 ;
        RECT 11.900000 50.075000 12.220000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 50.495000 12.220000 50.815000 ;
      LAYER met4 ;
        RECT 11.900000 50.495000 12.220000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 34.760000 12.625000 35.080000 ;
      LAYER met4 ;
        RECT 12.305000 34.760000 12.625000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 35.200000 12.625000 35.520000 ;
      LAYER met4 ;
        RECT 12.305000 35.200000 12.625000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 35.640000 12.625000 35.960000 ;
      LAYER met4 ;
        RECT 12.305000 35.640000 12.625000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 36.080000 12.625000 36.400000 ;
      LAYER met4 ;
        RECT 12.305000 36.080000 12.625000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 36.520000 12.625000 36.840000 ;
      LAYER met4 ;
        RECT 12.305000 36.520000 12.625000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 36.960000 12.625000 37.280000 ;
      LAYER met4 ;
        RECT 12.305000 36.960000 12.625000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 37.400000 12.625000 37.720000 ;
      LAYER met4 ;
        RECT 12.305000 37.400000 12.625000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 37.840000 12.625000 38.160000 ;
      LAYER met4 ;
        RECT 12.305000 37.840000 12.625000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 49.655000 12.625000 49.975000 ;
      LAYER met4 ;
        RECT 12.305000 49.655000 12.625000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 50.075000 12.625000 50.395000 ;
      LAYER met4 ;
        RECT 12.305000 50.075000 12.625000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 50.495000 12.625000 50.815000 ;
      LAYER met4 ;
        RECT 12.305000 50.495000 12.625000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 34.760000 13.030000 35.080000 ;
      LAYER met4 ;
        RECT 12.710000 34.760000 13.030000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 35.200000 13.030000 35.520000 ;
      LAYER met4 ;
        RECT 12.710000 35.200000 13.030000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 35.640000 13.030000 35.960000 ;
      LAYER met4 ;
        RECT 12.710000 35.640000 13.030000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 36.080000 13.030000 36.400000 ;
      LAYER met4 ;
        RECT 12.710000 36.080000 13.030000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 36.520000 13.030000 36.840000 ;
      LAYER met4 ;
        RECT 12.710000 36.520000 13.030000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 36.960000 13.030000 37.280000 ;
      LAYER met4 ;
        RECT 12.710000 36.960000 13.030000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 37.400000 13.030000 37.720000 ;
      LAYER met4 ;
        RECT 12.710000 37.400000 13.030000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 37.840000 13.030000 38.160000 ;
      LAYER met4 ;
        RECT 12.710000 37.840000 13.030000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 49.655000 13.030000 49.975000 ;
      LAYER met4 ;
        RECT 12.710000 49.655000 13.030000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 50.075000 13.030000 50.395000 ;
      LAYER met4 ;
        RECT 12.710000 50.075000 13.030000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 50.495000 13.030000 50.815000 ;
      LAYER met4 ;
        RECT 12.710000 50.495000 13.030000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 34.760000 13.435000 35.080000 ;
      LAYER met4 ;
        RECT 13.115000 34.760000 13.435000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 35.200000 13.435000 35.520000 ;
      LAYER met4 ;
        RECT 13.115000 35.200000 13.435000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 35.640000 13.435000 35.960000 ;
      LAYER met4 ;
        RECT 13.115000 35.640000 13.435000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 36.080000 13.435000 36.400000 ;
      LAYER met4 ;
        RECT 13.115000 36.080000 13.435000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 36.520000 13.435000 36.840000 ;
      LAYER met4 ;
        RECT 13.115000 36.520000 13.435000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 36.960000 13.435000 37.280000 ;
      LAYER met4 ;
        RECT 13.115000 36.960000 13.435000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 37.400000 13.435000 37.720000 ;
      LAYER met4 ;
        RECT 13.115000 37.400000 13.435000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 37.840000 13.435000 38.160000 ;
      LAYER met4 ;
        RECT 13.115000 37.840000 13.435000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 49.655000 13.435000 49.975000 ;
      LAYER met4 ;
        RECT 13.115000 49.655000 13.435000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 50.075000 13.435000 50.395000 ;
      LAYER met4 ;
        RECT 13.115000 50.075000 13.435000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 50.495000 13.435000 50.815000 ;
      LAYER met4 ;
        RECT 13.115000 50.495000 13.435000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 34.760000 13.840000 35.080000 ;
      LAYER met4 ;
        RECT 13.520000 34.760000 13.840000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 35.200000 13.840000 35.520000 ;
      LAYER met4 ;
        RECT 13.520000 35.200000 13.840000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 35.640000 13.840000 35.960000 ;
      LAYER met4 ;
        RECT 13.520000 35.640000 13.840000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 36.080000 13.840000 36.400000 ;
      LAYER met4 ;
        RECT 13.520000 36.080000 13.840000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 36.520000 13.840000 36.840000 ;
      LAYER met4 ;
        RECT 13.520000 36.520000 13.840000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 36.960000 13.840000 37.280000 ;
      LAYER met4 ;
        RECT 13.520000 36.960000 13.840000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 37.400000 13.840000 37.720000 ;
      LAYER met4 ;
        RECT 13.520000 37.400000 13.840000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 37.840000 13.840000 38.160000 ;
      LAYER met4 ;
        RECT 13.520000 37.840000 13.840000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 49.655000 13.840000 49.975000 ;
      LAYER met4 ;
        RECT 13.520000 49.655000 13.840000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 50.075000 13.840000 50.395000 ;
      LAYER met4 ;
        RECT 13.520000 50.075000 13.840000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 50.495000 13.840000 50.815000 ;
      LAYER met4 ;
        RECT 13.520000 50.495000 13.840000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 34.760000 14.245000 35.080000 ;
      LAYER met4 ;
        RECT 13.925000 34.760000 14.245000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 35.200000 14.245000 35.520000 ;
      LAYER met4 ;
        RECT 13.925000 35.200000 14.245000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 35.640000 14.245000 35.960000 ;
      LAYER met4 ;
        RECT 13.925000 35.640000 14.245000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 36.080000 14.245000 36.400000 ;
      LAYER met4 ;
        RECT 13.925000 36.080000 14.245000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 36.520000 14.245000 36.840000 ;
      LAYER met4 ;
        RECT 13.925000 36.520000 14.245000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 36.960000 14.245000 37.280000 ;
      LAYER met4 ;
        RECT 13.925000 36.960000 14.245000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 37.400000 14.245000 37.720000 ;
      LAYER met4 ;
        RECT 13.925000 37.400000 14.245000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 37.840000 14.245000 38.160000 ;
      LAYER met4 ;
        RECT 13.925000 37.840000 14.245000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 49.655000 14.245000 49.975000 ;
      LAYER met4 ;
        RECT 13.925000 49.655000 14.245000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 50.075000 14.245000 50.395000 ;
      LAYER met4 ;
        RECT 13.925000 50.075000 14.245000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 50.495000 14.245000 50.815000 ;
      LAYER met4 ;
        RECT 13.925000 50.495000 14.245000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 34.760000 14.650000 35.080000 ;
      LAYER met4 ;
        RECT 14.330000 34.760000 14.650000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 35.200000 14.650000 35.520000 ;
      LAYER met4 ;
        RECT 14.330000 35.200000 14.650000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 35.640000 14.650000 35.960000 ;
      LAYER met4 ;
        RECT 14.330000 35.640000 14.650000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 36.080000 14.650000 36.400000 ;
      LAYER met4 ;
        RECT 14.330000 36.080000 14.650000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 36.520000 14.650000 36.840000 ;
      LAYER met4 ;
        RECT 14.330000 36.520000 14.650000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 36.960000 14.650000 37.280000 ;
      LAYER met4 ;
        RECT 14.330000 36.960000 14.650000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 37.400000 14.650000 37.720000 ;
      LAYER met4 ;
        RECT 14.330000 37.400000 14.650000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 37.840000 14.650000 38.160000 ;
      LAYER met4 ;
        RECT 14.330000 37.840000 14.650000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 49.655000 14.650000 49.975000 ;
      LAYER met4 ;
        RECT 14.330000 49.655000 14.650000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 50.075000 14.650000 50.395000 ;
      LAYER met4 ;
        RECT 14.330000 50.075000 14.650000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 50.495000 14.650000 50.815000 ;
      LAYER met4 ;
        RECT 14.330000 50.495000 14.650000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 34.760000 15.055000 35.080000 ;
      LAYER met4 ;
        RECT 14.735000 34.760000 15.055000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 35.200000 15.055000 35.520000 ;
      LAYER met4 ;
        RECT 14.735000 35.200000 15.055000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 35.640000 15.055000 35.960000 ;
      LAYER met4 ;
        RECT 14.735000 35.640000 15.055000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 36.080000 15.055000 36.400000 ;
      LAYER met4 ;
        RECT 14.735000 36.080000 15.055000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 36.520000 15.055000 36.840000 ;
      LAYER met4 ;
        RECT 14.735000 36.520000 15.055000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 36.960000 15.055000 37.280000 ;
      LAYER met4 ;
        RECT 14.735000 36.960000 15.055000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 37.400000 15.055000 37.720000 ;
      LAYER met4 ;
        RECT 14.735000 37.400000 15.055000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 37.840000 15.055000 38.160000 ;
      LAYER met4 ;
        RECT 14.735000 37.840000 15.055000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 49.655000 15.055000 49.975000 ;
      LAYER met4 ;
        RECT 14.735000 49.655000 15.055000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 50.075000 15.055000 50.395000 ;
      LAYER met4 ;
        RECT 14.735000 50.075000 15.055000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 50.495000 15.055000 50.815000 ;
      LAYER met4 ;
        RECT 14.735000 50.495000 15.055000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 34.760000 15.460000 35.080000 ;
      LAYER met4 ;
        RECT 15.140000 34.760000 15.460000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 35.200000 15.460000 35.520000 ;
      LAYER met4 ;
        RECT 15.140000 35.200000 15.460000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 35.640000 15.460000 35.960000 ;
      LAYER met4 ;
        RECT 15.140000 35.640000 15.460000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 36.080000 15.460000 36.400000 ;
      LAYER met4 ;
        RECT 15.140000 36.080000 15.460000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 36.520000 15.460000 36.840000 ;
      LAYER met4 ;
        RECT 15.140000 36.520000 15.460000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 36.960000 15.460000 37.280000 ;
      LAYER met4 ;
        RECT 15.140000 36.960000 15.460000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 37.400000 15.460000 37.720000 ;
      LAYER met4 ;
        RECT 15.140000 37.400000 15.460000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 37.840000 15.460000 38.160000 ;
      LAYER met4 ;
        RECT 15.140000 37.840000 15.460000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 49.655000 15.460000 49.975000 ;
      LAYER met4 ;
        RECT 15.140000 49.655000 15.460000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 50.075000 15.460000 50.395000 ;
      LAYER met4 ;
        RECT 15.140000 50.075000 15.460000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 50.495000 15.460000 50.815000 ;
      LAYER met4 ;
        RECT 15.140000 50.495000 15.460000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 34.760000 15.865000 35.080000 ;
      LAYER met4 ;
        RECT 15.545000 34.760000 15.865000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 35.200000 15.865000 35.520000 ;
      LAYER met4 ;
        RECT 15.545000 35.200000 15.865000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 35.640000 15.865000 35.960000 ;
      LAYER met4 ;
        RECT 15.545000 35.640000 15.865000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 36.080000 15.865000 36.400000 ;
      LAYER met4 ;
        RECT 15.545000 36.080000 15.865000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 36.520000 15.865000 36.840000 ;
      LAYER met4 ;
        RECT 15.545000 36.520000 15.865000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 36.960000 15.865000 37.280000 ;
      LAYER met4 ;
        RECT 15.545000 36.960000 15.865000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 37.400000 15.865000 37.720000 ;
      LAYER met4 ;
        RECT 15.545000 37.400000 15.865000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 37.840000 15.865000 38.160000 ;
      LAYER met4 ;
        RECT 15.545000 37.840000 15.865000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 49.655000 15.865000 49.975000 ;
      LAYER met4 ;
        RECT 15.545000 49.655000 15.865000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 50.075000 15.865000 50.395000 ;
      LAYER met4 ;
        RECT 15.545000 50.075000 15.865000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 50.495000 15.865000 50.815000 ;
      LAYER met4 ;
        RECT 15.545000 50.495000 15.865000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 34.760000 16.270000 35.080000 ;
      LAYER met4 ;
        RECT 15.950000 34.760000 16.270000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 35.200000 16.270000 35.520000 ;
      LAYER met4 ;
        RECT 15.950000 35.200000 16.270000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 35.640000 16.270000 35.960000 ;
      LAYER met4 ;
        RECT 15.950000 35.640000 16.270000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 36.080000 16.270000 36.400000 ;
      LAYER met4 ;
        RECT 15.950000 36.080000 16.270000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 36.520000 16.270000 36.840000 ;
      LAYER met4 ;
        RECT 15.950000 36.520000 16.270000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 36.960000 16.270000 37.280000 ;
      LAYER met4 ;
        RECT 15.950000 36.960000 16.270000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 37.400000 16.270000 37.720000 ;
      LAYER met4 ;
        RECT 15.950000 37.400000 16.270000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 37.840000 16.270000 38.160000 ;
      LAYER met4 ;
        RECT 15.950000 37.840000 16.270000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 49.655000 16.270000 49.975000 ;
      LAYER met4 ;
        RECT 15.950000 49.655000 16.270000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 50.075000 16.270000 50.395000 ;
      LAYER met4 ;
        RECT 15.950000 50.075000 16.270000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 50.495000 16.270000 50.815000 ;
      LAYER met4 ;
        RECT 15.950000 50.495000 16.270000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 34.760000 16.675000 35.080000 ;
      LAYER met4 ;
        RECT 16.355000 34.760000 16.675000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 35.200000 16.675000 35.520000 ;
      LAYER met4 ;
        RECT 16.355000 35.200000 16.675000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 35.640000 16.675000 35.960000 ;
      LAYER met4 ;
        RECT 16.355000 35.640000 16.675000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 36.080000 16.675000 36.400000 ;
      LAYER met4 ;
        RECT 16.355000 36.080000 16.675000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 36.520000 16.675000 36.840000 ;
      LAYER met4 ;
        RECT 16.355000 36.520000 16.675000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 36.960000 16.675000 37.280000 ;
      LAYER met4 ;
        RECT 16.355000 36.960000 16.675000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 37.400000 16.675000 37.720000 ;
      LAYER met4 ;
        RECT 16.355000 37.400000 16.675000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 37.840000 16.675000 38.160000 ;
      LAYER met4 ;
        RECT 16.355000 37.840000 16.675000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 49.655000 16.675000 49.975000 ;
      LAYER met4 ;
        RECT 16.355000 49.655000 16.675000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 50.075000 16.675000 50.395000 ;
      LAYER met4 ;
        RECT 16.355000 50.075000 16.675000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 50.495000 16.675000 50.815000 ;
      LAYER met4 ;
        RECT 16.355000 50.495000 16.675000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 34.760000 17.080000 35.080000 ;
      LAYER met4 ;
        RECT 16.760000 34.760000 17.080000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 35.200000 17.080000 35.520000 ;
      LAYER met4 ;
        RECT 16.760000 35.200000 17.080000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 35.640000 17.080000 35.960000 ;
      LAYER met4 ;
        RECT 16.760000 35.640000 17.080000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 36.080000 17.080000 36.400000 ;
      LAYER met4 ;
        RECT 16.760000 36.080000 17.080000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 36.520000 17.080000 36.840000 ;
      LAYER met4 ;
        RECT 16.760000 36.520000 17.080000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 36.960000 17.080000 37.280000 ;
      LAYER met4 ;
        RECT 16.760000 36.960000 17.080000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 37.400000 17.080000 37.720000 ;
      LAYER met4 ;
        RECT 16.760000 37.400000 17.080000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 37.840000 17.080000 38.160000 ;
      LAYER met4 ;
        RECT 16.760000 37.840000 17.080000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 49.655000 17.080000 49.975000 ;
      LAYER met4 ;
        RECT 16.760000 49.655000 17.080000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 50.075000 17.080000 50.395000 ;
      LAYER met4 ;
        RECT 16.760000 50.075000 17.080000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 50.495000 17.080000 50.815000 ;
      LAYER met4 ;
        RECT 16.760000 50.495000 17.080000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 34.760000 17.485000 35.080000 ;
      LAYER met4 ;
        RECT 17.165000 34.760000 17.485000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 35.200000 17.485000 35.520000 ;
      LAYER met4 ;
        RECT 17.165000 35.200000 17.485000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 35.640000 17.485000 35.960000 ;
      LAYER met4 ;
        RECT 17.165000 35.640000 17.485000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 36.080000 17.485000 36.400000 ;
      LAYER met4 ;
        RECT 17.165000 36.080000 17.485000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 36.520000 17.485000 36.840000 ;
      LAYER met4 ;
        RECT 17.165000 36.520000 17.485000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 36.960000 17.485000 37.280000 ;
      LAYER met4 ;
        RECT 17.165000 36.960000 17.485000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 37.400000 17.485000 37.720000 ;
      LAYER met4 ;
        RECT 17.165000 37.400000 17.485000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 37.840000 17.485000 38.160000 ;
      LAYER met4 ;
        RECT 17.165000 37.840000 17.485000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 49.655000 17.485000 49.975000 ;
      LAYER met4 ;
        RECT 17.165000 49.655000 17.485000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 50.075000 17.485000 50.395000 ;
      LAYER met4 ;
        RECT 17.165000 50.075000 17.485000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 50.495000 17.485000 50.815000 ;
      LAYER met4 ;
        RECT 17.165000 50.495000 17.485000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 34.760000 17.890000 35.080000 ;
      LAYER met4 ;
        RECT 17.570000 34.760000 17.890000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 35.200000 17.890000 35.520000 ;
      LAYER met4 ;
        RECT 17.570000 35.200000 17.890000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 35.640000 17.890000 35.960000 ;
      LAYER met4 ;
        RECT 17.570000 35.640000 17.890000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 36.080000 17.890000 36.400000 ;
      LAYER met4 ;
        RECT 17.570000 36.080000 17.890000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 36.520000 17.890000 36.840000 ;
      LAYER met4 ;
        RECT 17.570000 36.520000 17.890000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 36.960000 17.890000 37.280000 ;
      LAYER met4 ;
        RECT 17.570000 36.960000 17.890000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 37.400000 17.890000 37.720000 ;
      LAYER met4 ;
        RECT 17.570000 37.400000 17.890000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 37.840000 17.890000 38.160000 ;
      LAYER met4 ;
        RECT 17.570000 37.840000 17.890000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 49.655000 17.890000 49.975000 ;
      LAYER met4 ;
        RECT 17.570000 49.655000 17.890000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 50.075000 17.890000 50.395000 ;
      LAYER met4 ;
        RECT 17.570000 50.075000 17.890000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 50.495000 17.890000 50.815000 ;
      LAYER met4 ;
        RECT 17.570000 50.495000 17.890000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 34.760000 18.295000 35.080000 ;
      LAYER met4 ;
        RECT 17.975000 34.760000 18.295000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 35.200000 18.295000 35.520000 ;
      LAYER met4 ;
        RECT 17.975000 35.200000 18.295000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 35.640000 18.295000 35.960000 ;
      LAYER met4 ;
        RECT 17.975000 35.640000 18.295000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 36.080000 18.295000 36.400000 ;
      LAYER met4 ;
        RECT 17.975000 36.080000 18.295000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 36.520000 18.295000 36.840000 ;
      LAYER met4 ;
        RECT 17.975000 36.520000 18.295000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 36.960000 18.295000 37.280000 ;
      LAYER met4 ;
        RECT 17.975000 36.960000 18.295000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 37.400000 18.295000 37.720000 ;
      LAYER met4 ;
        RECT 17.975000 37.400000 18.295000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 37.840000 18.295000 38.160000 ;
      LAYER met4 ;
        RECT 17.975000 37.840000 18.295000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 49.655000 18.295000 49.975000 ;
      LAYER met4 ;
        RECT 17.975000 49.655000 18.295000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 50.075000 18.295000 50.395000 ;
      LAYER met4 ;
        RECT 17.975000 50.075000 18.295000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 50.495000 18.295000 50.815000 ;
      LAYER met4 ;
        RECT 17.975000 50.495000 18.295000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 34.760000 18.700000 35.080000 ;
      LAYER met4 ;
        RECT 18.380000 34.760000 18.700000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 35.200000 18.700000 35.520000 ;
      LAYER met4 ;
        RECT 18.380000 35.200000 18.700000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 35.640000 18.700000 35.960000 ;
      LAYER met4 ;
        RECT 18.380000 35.640000 18.700000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 36.080000 18.700000 36.400000 ;
      LAYER met4 ;
        RECT 18.380000 36.080000 18.700000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 36.520000 18.700000 36.840000 ;
      LAYER met4 ;
        RECT 18.380000 36.520000 18.700000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 36.960000 18.700000 37.280000 ;
      LAYER met4 ;
        RECT 18.380000 36.960000 18.700000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 37.400000 18.700000 37.720000 ;
      LAYER met4 ;
        RECT 18.380000 37.400000 18.700000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 37.840000 18.700000 38.160000 ;
      LAYER met4 ;
        RECT 18.380000 37.840000 18.700000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 49.655000 18.700000 49.975000 ;
      LAYER met4 ;
        RECT 18.380000 49.655000 18.700000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 50.075000 18.700000 50.395000 ;
      LAYER met4 ;
        RECT 18.380000 50.075000 18.700000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 50.495000 18.700000 50.815000 ;
      LAYER met4 ;
        RECT 18.380000 50.495000 18.700000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 34.760000 19.105000 35.080000 ;
      LAYER met4 ;
        RECT 18.785000 34.760000 19.105000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 35.200000 19.105000 35.520000 ;
      LAYER met4 ;
        RECT 18.785000 35.200000 19.105000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 35.640000 19.105000 35.960000 ;
      LAYER met4 ;
        RECT 18.785000 35.640000 19.105000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 36.080000 19.105000 36.400000 ;
      LAYER met4 ;
        RECT 18.785000 36.080000 19.105000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 36.520000 19.105000 36.840000 ;
      LAYER met4 ;
        RECT 18.785000 36.520000 19.105000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 36.960000 19.105000 37.280000 ;
      LAYER met4 ;
        RECT 18.785000 36.960000 19.105000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 37.400000 19.105000 37.720000 ;
      LAYER met4 ;
        RECT 18.785000 37.400000 19.105000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 37.840000 19.105000 38.160000 ;
      LAYER met4 ;
        RECT 18.785000 37.840000 19.105000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 49.655000 19.105000 49.975000 ;
      LAYER met4 ;
        RECT 18.785000 49.655000 19.105000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 50.075000 19.105000 50.395000 ;
      LAYER met4 ;
        RECT 18.785000 50.075000 19.105000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 50.495000 19.105000 50.815000 ;
      LAYER met4 ;
        RECT 18.785000 50.495000 19.105000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 34.760000 19.510000 35.080000 ;
      LAYER met4 ;
        RECT 19.190000 34.760000 19.510000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 35.200000 19.510000 35.520000 ;
      LAYER met4 ;
        RECT 19.190000 35.200000 19.510000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 35.640000 19.510000 35.960000 ;
      LAYER met4 ;
        RECT 19.190000 35.640000 19.510000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 36.080000 19.510000 36.400000 ;
      LAYER met4 ;
        RECT 19.190000 36.080000 19.510000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 36.520000 19.510000 36.840000 ;
      LAYER met4 ;
        RECT 19.190000 36.520000 19.510000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 36.960000 19.510000 37.280000 ;
      LAYER met4 ;
        RECT 19.190000 36.960000 19.510000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 37.400000 19.510000 37.720000 ;
      LAYER met4 ;
        RECT 19.190000 37.400000 19.510000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 37.840000 19.510000 38.160000 ;
      LAYER met4 ;
        RECT 19.190000 37.840000 19.510000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 49.655000 19.510000 49.975000 ;
      LAYER met4 ;
        RECT 19.190000 49.655000 19.510000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 50.075000 19.510000 50.395000 ;
      LAYER met4 ;
        RECT 19.190000 50.075000 19.510000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 50.495000 19.510000 50.815000 ;
      LAYER met4 ;
        RECT 19.190000 50.495000 19.510000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 34.760000 19.915000 35.080000 ;
      LAYER met4 ;
        RECT 19.595000 34.760000 19.915000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 35.200000 19.915000 35.520000 ;
      LAYER met4 ;
        RECT 19.595000 35.200000 19.915000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 35.640000 19.915000 35.960000 ;
      LAYER met4 ;
        RECT 19.595000 35.640000 19.915000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 36.080000 19.915000 36.400000 ;
      LAYER met4 ;
        RECT 19.595000 36.080000 19.915000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 36.520000 19.915000 36.840000 ;
      LAYER met4 ;
        RECT 19.595000 36.520000 19.915000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 36.960000 19.915000 37.280000 ;
      LAYER met4 ;
        RECT 19.595000 36.960000 19.915000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 37.400000 19.915000 37.720000 ;
      LAYER met4 ;
        RECT 19.595000 37.400000 19.915000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 37.840000 19.915000 38.160000 ;
      LAYER met4 ;
        RECT 19.595000 37.840000 19.915000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 49.655000 19.915000 49.975000 ;
      LAYER met4 ;
        RECT 19.595000 49.655000 19.915000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 50.075000 19.915000 50.395000 ;
      LAYER met4 ;
        RECT 19.595000 50.075000 19.915000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 50.495000 19.915000 50.815000 ;
      LAYER met4 ;
        RECT 19.595000 50.495000 19.915000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 34.760000 2.490000 35.080000 ;
      LAYER met4 ;
        RECT 2.170000 34.760000 2.490000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 35.200000 2.490000 35.520000 ;
      LAYER met4 ;
        RECT 2.170000 35.200000 2.490000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 35.640000 2.490000 35.960000 ;
      LAYER met4 ;
        RECT 2.170000 35.640000 2.490000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 36.080000 2.490000 36.400000 ;
      LAYER met4 ;
        RECT 2.170000 36.080000 2.490000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 36.520000 2.490000 36.840000 ;
      LAYER met4 ;
        RECT 2.170000 36.520000 2.490000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 36.960000 2.490000 37.280000 ;
      LAYER met4 ;
        RECT 2.170000 36.960000 2.490000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 37.400000 2.490000 37.720000 ;
      LAYER met4 ;
        RECT 2.170000 37.400000 2.490000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 37.840000 2.490000 38.160000 ;
      LAYER met4 ;
        RECT 2.170000 37.840000 2.490000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 49.655000 2.490000 49.975000 ;
      LAYER met4 ;
        RECT 2.170000 49.655000 2.490000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 50.075000 2.490000 50.395000 ;
      LAYER met4 ;
        RECT 2.170000 50.075000 2.490000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170000 50.495000 2.490000 50.815000 ;
      LAYER met4 ;
        RECT 2.170000 50.495000 2.490000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 34.760000 2.900000 35.080000 ;
      LAYER met4 ;
        RECT 2.580000 34.760000 2.900000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 35.200000 2.900000 35.520000 ;
      LAYER met4 ;
        RECT 2.580000 35.200000 2.900000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 35.640000 2.900000 35.960000 ;
      LAYER met4 ;
        RECT 2.580000 35.640000 2.900000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 36.080000 2.900000 36.400000 ;
      LAYER met4 ;
        RECT 2.580000 36.080000 2.900000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 36.520000 2.900000 36.840000 ;
      LAYER met4 ;
        RECT 2.580000 36.520000 2.900000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 36.960000 2.900000 37.280000 ;
      LAYER met4 ;
        RECT 2.580000 36.960000 2.900000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 37.400000 2.900000 37.720000 ;
      LAYER met4 ;
        RECT 2.580000 37.400000 2.900000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 37.840000 2.900000 38.160000 ;
      LAYER met4 ;
        RECT 2.580000 37.840000 2.900000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 49.655000 2.900000 49.975000 ;
      LAYER met4 ;
        RECT 2.580000 49.655000 2.900000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 50.075000 2.900000 50.395000 ;
      LAYER met4 ;
        RECT 2.580000 50.075000 2.900000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580000 50.495000 2.900000 50.815000 ;
      LAYER met4 ;
        RECT 2.580000 50.495000 2.900000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 34.760000 3.310000 35.080000 ;
      LAYER met4 ;
        RECT 2.990000 34.760000 3.310000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 35.200000 3.310000 35.520000 ;
      LAYER met4 ;
        RECT 2.990000 35.200000 3.310000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 35.640000 3.310000 35.960000 ;
      LAYER met4 ;
        RECT 2.990000 35.640000 3.310000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 36.080000 3.310000 36.400000 ;
      LAYER met4 ;
        RECT 2.990000 36.080000 3.310000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 36.520000 3.310000 36.840000 ;
      LAYER met4 ;
        RECT 2.990000 36.520000 3.310000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 36.960000 3.310000 37.280000 ;
      LAYER met4 ;
        RECT 2.990000 36.960000 3.310000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 37.400000 3.310000 37.720000 ;
      LAYER met4 ;
        RECT 2.990000 37.400000 3.310000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 37.840000 3.310000 38.160000 ;
      LAYER met4 ;
        RECT 2.990000 37.840000 3.310000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 49.655000 3.310000 49.975000 ;
      LAYER met4 ;
        RECT 2.990000 49.655000 3.310000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 50.075000 3.310000 50.395000 ;
      LAYER met4 ;
        RECT 2.990000 50.075000 3.310000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 50.495000 3.310000 50.815000 ;
      LAYER met4 ;
        RECT 2.990000 50.495000 3.310000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 34.760000 20.320000 35.080000 ;
      LAYER met4 ;
        RECT 20.000000 34.760000 20.320000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 35.200000 20.320000 35.520000 ;
      LAYER met4 ;
        RECT 20.000000 35.200000 20.320000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 35.640000 20.320000 35.960000 ;
      LAYER met4 ;
        RECT 20.000000 35.640000 20.320000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 36.080000 20.320000 36.400000 ;
      LAYER met4 ;
        RECT 20.000000 36.080000 20.320000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 36.520000 20.320000 36.840000 ;
      LAYER met4 ;
        RECT 20.000000 36.520000 20.320000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 36.960000 20.320000 37.280000 ;
      LAYER met4 ;
        RECT 20.000000 36.960000 20.320000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 37.400000 20.320000 37.720000 ;
      LAYER met4 ;
        RECT 20.000000 37.400000 20.320000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 37.840000 20.320000 38.160000 ;
      LAYER met4 ;
        RECT 20.000000 37.840000 20.320000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 49.655000 20.320000 49.975000 ;
      LAYER met4 ;
        RECT 20.000000 49.655000 20.320000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 50.075000 20.320000 50.395000 ;
      LAYER met4 ;
        RECT 20.000000 50.075000 20.320000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 50.495000 20.320000 50.815000 ;
      LAYER met4 ;
        RECT 20.000000 50.495000 20.320000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 34.760000 20.725000 35.080000 ;
      LAYER met4 ;
        RECT 20.405000 34.760000 20.725000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 35.200000 20.725000 35.520000 ;
      LAYER met4 ;
        RECT 20.405000 35.200000 20.725000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 35.640000 20.725000 35.960000 ;
      LAYER met4 ;
        RECT 20.405000 35.640000 20.725000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 36.080000 20.725000 36.400000 ;
      LAYER met4 ;
        RECT 20.405000 36.080000 20.725000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 36.520000 20.725000 36.840000 ;
      LAYER met4 ;
        RECT 20.405000 36.520000 20.725000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 36.960000 20.725000 37.280000 ;
      LAYER met4 ;
        RECT 20.405000 36.960000 20.725000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 37.400000 20.725000 37.720000 ;
      LAYER met4 ;
        RECT 20.405000 37.400000 20.725000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 37.840000 20.725000 38.160000 ;
      LAYER met4 ;
        RECT 20.405000 37.840000 20.725000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 49.655000 20.725000 49.975000 ;
      LAYER met4 ;
        RECT 20.405000 49.655000 20.725000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 50.075000 20.725000 50.395000 ;
      LAYER met4 ;
        RECT 20.405000 50.075000 20.725000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 50.495000 20.725000 50.815000 ;
      LAYER met4 ;
        RECT 20.405000 50.495000 20.725000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 34.760000 21.130000 35.080000 ;
      LAYER met4 ;
        RECT 20.810000 34.760000 21.130000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 35.200000 21.130000 35.520000 ;
      LAYER met4 ;
        RECT 20.810000 35.200000 21.130000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 35.640000 21.130000 35.960000 ;
      LAYER met4 ;
        RECT 20.810000 35.640000 21.130000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 36.080000 21.130000 36.400000 ;
      LAYER met4 ;
        RECT 20.810000 36.080000 21.130000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 36.520000 21.130000 36.840000 ;
      LAYER met4 ;
        RECT 20.810000 36.520000 21.130000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 36.960000 21.130000 37.280000 ;
      LAYER met4 ;
        RECT 20.810000 36.960000 21.130000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 37.400000 21.130000 37.720000 ;
      LAYER met4 ;
        RECT 20.810000 37.400000 21.130000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 37.840000 21.130000 38.160000 ;
      LAYER met4 ;
        RECT 20.810000 37.840000 21.130000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 49.655000 21.130000 49.975000 ;
      LAYER met4 ;
        RECT 20.810000 49.655000 21.130000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 50.075000 21.130000 50.395000 ;
      LAYER met4 ;
        RECT 20.810000 50.075000 21.130000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 50.495000 21.130000 50.815000 ;
      LAYER met4 ;
        RECT 20.810000 50.495000 21.130000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 34.760000 21.535000 35.080000 ;
      LAYER met4 ;
        RECT 21.215000 34.760000 21.535000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 35.200000 21.535000 35.520000 ;
      LAYER met4 ;
        RECT 21.215000 35.200000 21.535000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 35.640000 21.535000 35.960000 ;
      LAYER met4 ;
        RECT 21.215000 35.640000 21.535000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 36.080000 21.535000 36.400000 ;
      LAYER met4 ;
        RECT 21.215000 36.080000 21.535000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 36.520000 21.535000 36.840000 ;
      LAYER met4 ;
        RECT 21.215000 36.520000 21.535000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 36.960000 21.535000 37.280000 ;
      LAYER met4 ;
        RECT 21.215000 36.960000 21.535000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 37.400000 21.535000 37.720000 ;
      LAYER met4 ;
        RECT 21.215000 37.400000 21.535000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 37.840000 21.535000 38.160000 ;
      LAYER met4 ;
        RECT 21.215000 37.840000 21.535000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 49.655000 21.535000 49.975000 ;
      LAYER met4 ;
        RECT 21.215000 49.655000 21.535000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 50.075000 21.535000 50.395000 ;
      LAYER met4 ;
        RECT 21.215000 50.075000 21.535000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 50.495000 21.535000 50.815000 ;
      LAYER met4 ;
        RECT 21.215000 50.495000 21.535000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 34.760000 21.940000 35.080000 ;
      LAYER met4 ;
        RECT 21.620000 34.760000 21.940000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 35.200000 21.940000 35.520000 ;
      LAYER met4 ;
        RECT 21.620000 35.200000 21.940000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 35.640000 21.940000 35.960000 ;
      LAYER met4 ;
        RECT 21.620000 35.640000 21.940000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 36.080000 21.940000 36.400000 ;
      LAYER met4 ;
        RECT 21.620000 36.080000 21.940000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 36.520000 21.940000 36.840000 ;
      LAYER met4 ;
        RECT 21.620000 36.520000 21.940000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 36.960000 21.940000 37.280000 ;
      LAYER met4 ;
        RECT 21.620000 36.960000 21.940000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 37.400000 21.940000 37.720000 ;
      LAYER met4 ;
        RECT 21.620000 37.400000 21.940000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 37.840000 21.940000 38.160000 ;
      LAYER met4 ;
        RECT 21.620000 37.840000 21.940000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 49.655000 21.940000 49.975000 ;
      LAYER met4 ;
        RECT 21.620000 49.655000 21.940000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 50.075000 21.940000 50.395000 ;
      LAYER met4 ;
        RECT 21.620000 50.075000 21.940000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 50.495000 21.940000 50.815000 ;
      LAYER met4 ;
        RECT 21.620000 50.495000 21.940000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 34.760000 22.345000 35.080000 ;
      LAYER met4 ;
        RECT 22.025000 34.760000 22.345000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 35.200000 22.345000 35.520000 ;
      LAYER met4 ;
        RECT 22.025000 35.200000 22.345000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 35.640000 22.345000 35.960000 ;
      LAYER met4 ;
        RECT 22.025000 35.640000 22.345000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 36.080000 22.345000 36.400000 ;
      LAYER met4 ;
        RECT 22.025000 36.080000 22.345000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 36.520000 22.345000 36.840000 ;
      LAYER met4 ;
        RECT 22.025000 36.520000 22.345000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 36.960000 22.345000 37.280000 ;
      LAYER met4 ;
        RECT 22.025000 36.960000 22.345000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 37.400000 22.345000 37.720000 ;
      LAYER met4 ;
        RECT 22.025000 37.400000 22.345000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 37.840000 22.345000 38.160000 ;
      LAYER met4 ;
        RECT 22.025000 37.840000 22.345000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 49.655000 22.345000 49.975000 ;
      LAYER met4 ;
        RECT 22.025000 49.655000 22.345000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 50.075000 22.345000 50.395000 ;
      LAYER met4 ;
        RECT 22.025000 50.075000 22.345000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 50.495000 22.345000 50.815000 ;
      LAYER met4 ;
        RECT 22.025000 50.495000 22.345000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 34.760000 22.750000 35.080000 ;
      LAYER met4 ;
        RECT 22.430000 34.760000 22.750000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 35.200000 22.750000 35.520000 ;
      LAYER met4 ;
        RECT 22.430000 35.200000 22.750000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 35.640000 22.750000 35.960000 ;
      LAYER met4 ;
        RECT 22.430000 35.640000 22.750000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 36.080000 22.750000 36.400000 ;
      LAYER met4 ;
        RECT 22.430000 36.080000 22.750000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 36.520000 22.750000 36.840000 ;
      LAYER met4 ;
        RECT 22.430000 36.520000 22.750000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 36.960000 22.750000 37.280000 ;
      LAYER met4 ;
        RECT 22.430000 36.960000 22.750000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 37.400000 22.750000 37.720000 ;
      LAYER met4 ;
        RECT 22.430000 37.400000 22.750000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 37.840000 22.750000 38.160000 ;
      LAYER met4 ;
        RECT 22.430000 37.840000 22.750000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 49.655000 22.750000 49.975000 ;
      LAYER met4 ;
        RECT 22.430000 49.655000 22.750000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 50.075000 22.750000 50.395000 ;
      LAYER met4 ;
        RECT 22.430000 50.075000 22.750000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 50.495000 22.750000 50.815000 ;
      LAYER met4 ;
        RECT 22.430000 50.495000 22.750000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 34.760000 23.155000 35.080000 ;
      LAYER met4 ;
        RECT 22.835000 34.760000 23.155000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 35.200000 23.155000 35.520000 ;
      LAYER met4 ;
        RECT 22.835000 35.200000 23.155000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 35.640000 23.155000 35.960000 ;
      LAYER met4 ;
        RECT 22.835000 35.640000 23.155000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 36.080000 23.155000 36.400000 ;
      LAYER met4 ;
        RECT 22.835000 36.080000 23.155000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 36.520000 23.155000 36.840000 ;
      LAYER met4 ;
        RECT 22.835000 36.520000 23.155000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 36.960000 23.155000 37.280000 ;
      LAYER met4 ;
        RECT 22.835000 36.960000 23.155000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 37.400000 23.155000 37.720000 ;
      LAYER met4 ;
        RECT 22.835000 37.400000 23.155000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 37.840000 23.155000 38.160000 ;
      LAYER met4 ;
        RECT 22.835000 37.840000 23.155000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 49.655000 23.155000 49.975000 ;
      LAYER met4 ;
        RECT 22.835000 49.655000 23.155000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 50.075000 23.155000 50.395000 ;
      LAYER met4 ;
        RECT 22.835000 50.075000 23.155000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 50.495000 23.155000 50.815000 ;
      LAYER met4 ;
        RECT 22.835000 50.495000 23.155000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 34.760000 23.560000 35.080000 ;
      LAYER met4 ;
        RECT 23.240000 34.760000 23.560000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 35.200000 23.560000 35.520000 ;
      LAYER met4 ;
        RECT 23.240000 35.200000 23.560000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 35.640000 23.560000 35.960000 ;
      LAYER met4 ;
        RECT 23.240000 35.640000 23.560000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 36.080000 23.560000 36.400000 ;
      LAYER met4 ;
        RECT 23.240000 36.080000 23.560000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 36.520000 23.560000 36.840000 ;
      LAYER met4 ;
        RECT 23.240000 36.520000 23.560000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 36.960000 23.560000 37.280000 ;
      LAYER met4 ;
        RECT 23.240000 36.960000 23.560000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 37.400000 23.560000 37.720000 ;
      LAYER met4 ;
        RECT 23.240000 37.400000 23.560000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 37.840000 23.560000 38.160000 ;
      LAYER met4 ;
        RECT 23.240000 37.840000 23.560000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 49.655000 23.560000 49.975000 ;
      LAYER met4 ;
        RECT 23.240000 49.655000 23.560000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 50.075000 23.560000 50.395000 ;
      LAYER met4 ;
        RECT 23.240000 50.075000 23.560000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 50.495000 23.560000 50.815000 ;
      LAYER met4 ;
        RECT 23.240000 50.495000 23.560000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 34.760000 23.965000 35.080000 ;
      LAYER met4 ;
        RECT 23.645000 34.760000 23.965000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 35.200000 23.965000 35.520000 ;
      LAYER met4 ;
        RECT 23.645000 35.200000 23.965000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 35.640000 23.965000 35.960000 ;
      LAYER met4 ;
        RECT 23.645000 35.640000 23.965000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 36.080000 23.965000 36.400000 ;
      LAYER met4 ;
        RECT 23.645000 36.080000 23.965000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 36.520000 23.965000 36.840000 ;
      LAYER met4 ;
        RECT 23.645000 36.520000 23.965000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 36.960000 23.965000 37.280000 ;
      LAYER met4 ;
        RECT 23.645000 36.960000 23.965000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 37.400000 23.965000 37.720000 ;
      LAYER met4 ;
        RECT 23.645000 37.400000 23.965000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 37.840000 23.965000 38.160000 ;
      LAYER met4 ;
        RECT 23.645000 37.840000 23.965000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 49.655000 23.965000 49.975000 ;
      LAYER met4 ;
        RECT 23.645000 49.655000 23.965000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 50.075000 23.965000 50.395000 ;
      LAYER met4 ;
        RECT 23.645000 50.075000 23.965000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 50.495000 23.965000 50.815000 ;
      LAYER met4 ;
        RECT 23.645000 50.495000 23.965000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 34.760000 24.370000 35.080000 ;
      LAYER met4 ;
        RECT 24.050000 34.760000 24.370000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 35.200000 24.370000 35.520000 ;
      LAYER met4 ;
        RECT 24.050000 35.200000 24.370000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 35.640000 24.370000 35.960000 ;
      LAYER met4 ;
        RECT 24.050000 35.640000 24.370000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 36.080000 24.370000 36.400000 ;
      LAYER met4 ;
        RECT 24.050000 36.080000 24.370000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 36.520000 24.370000 36.840000 ;
      LAYER met4 ;
        RECT 24.050000 36.520000 24.370000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 36.960000 24.370000 37.280000 ;
      LAYER met4 ;
        RECT 24.050000 36.960000 24.370000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 37.400000 24.370000 37.720000 ;
      LAYER met4 ;
        RECT 24.050000 37.400000 24.370000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 37.840000 24.370000 38.160000 ;
      LAYER met4 ;
        RECT 24.050000 37.840000 24.370000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 49.655000 24.370000 49.975000 ;
      LAYER met4 ;
        RECT 24.050000 49.655000 24.370000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 50.075000 24.370000 50.395000 ;
      LAYER met4 ;
        RECT 24.050000 50.075000 24.370000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050000 50.495000 24.370000 50.815000 ;
      LAYER met4 ;
        RECT 24.050000 50.495000 24.370000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 34.760000 3.715000 35.080000 ;
      LAYER met4 ;
        RECT 3.395000 34.760000 3.715000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 35.200000 3.715000 35.520000 ;
      LAYER met4 ;
        RECT 3.395000 35.200000 3.715000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 35.640000 3.715000 35.960000 ;
      LAYER met4 ;
        RECT 3.395000 35.640000 3.715000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 36.080000 3.715000 36.400000 ;
      LAYER met4 ;
        RECT 3.395000 36.080000 3.715000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 36.520000 3.715000 36.840000 ;
      LAYER met4 ;
        RECT 3.395000 36.520000 3.715000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 36.960000 3.715000 37.280000 ;
      LAYER met4 ;
        RECT 3.395000 36.960000 3.715000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 37.400000 3.715000 37.720000 ;
      LAYER met4 ;
        RECT 3.395000 37.400000 3.715000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 37.840000 3.715000 38.160000 ;
      LAYER met4 ;
        RECT 3.395000 37.840000 3.715000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 49.655000 3.715000 49.975000 ;
      LAYER met4 ;
        RECT 3.395000 49.655000 3.715000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 50.075000 3.715000 50.395000 ;
      LAYER met4 ;
        RECT 3.395000 50.075000 3.715000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 50.495000 3.715000 50.815000 ;
      LAYER met4 ;
        RECT 3.395000 50.495000 3.715000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 34.760000 4.120000 35.080000 ;
      LAYER met4 ;
        RECT 3.800000 34.760000 4.120000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 35.200000 4.120000 35.520000 ;
      LAYER met4 ;
        RECT 3.800000 35.200000 4.120000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 35.640000 4.120000 35.960000 ;
      LAYER met4 ;
        RECT 3.800000 35.640000 4.120000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 36.080000 4.120000 36.400000 ;
      LAYER met4 ;
        RECT 3.800000 36.080000 4.120000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 36.520000 4.120000 36.840000 ;
      LAYER met4 ;
        RECT 3.800000 36.520000 4.120000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 36.960000 4.120000 37.280000 ;
      LAYER met4 ;
        RECT 3.800000 36.960000 4.120000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 37.400000 4.120000 37.720000 ;
      LAYER met4 ;
        RECT 3.800000 37.400000 4.120000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 37.840000 4.120000 38.160000 ;
      LAYER met4 ;
        RECT 3.800000 37.840000 4.120000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 49.655000 4.120000 49.975000 ;
      LAYER met4 ;
        RECT 3.800000 49.655000 4.120000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 50.075000 4.120000 50.395000 ;
      LAYER met4 ;
        RECT 3.800000 50.075000 4.120000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 50.495000 4.120000 50.815000 ;
      LAYER met4 ;
        RECT 3.800000 50.495000 4.120000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 34.760000 4.525000 35.080000 ;
      LAYER met4 ;
        RECT 4.205000 34.760000 4.525000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 35.200000 4.525000 35.520000 ;
      LAYER met4 ;
        RECT 4.205000 35.200000 4.525000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 35.640000 4.525000 35.960000 ;
      LAYER met4 ;
        RECT 4.205000 35.640000 4.525000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 36.080000 4.525000 36.400000 ;
      LAYER met4 ;
        RECT 4.205000 36.080000 4.525000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 36.520000 4.525000 36.840000 ;
      LAYER met4 ;
        RECT 4.205000 36.520000 4.525000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 36.960000 4.525000 37.280000 ;
      LAYER met4 ;
        RECT 4.205000 36.960000 4.525000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 37.400000 4.525000 37.720000 ;
      LAYER met4 ;
        RECT 4.205000 37.400000 4.525000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 37.840000 4.525000 38.160000 ;
      LAYER met4 ;
        RECT 4.205000 37.840000 4.525000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 49.655000 4.525000 49.975000 ;
      LAYER met4 ;
        RECT 4.205000 49.655000 4.525000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 50.075000 4.525000 50.395000 ;
      LAYER met4 ;
        RECT 4.205000 50.075000 4.525000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 50.495000 4.525000 50.815000 ;
      LAYER met4 ;
        RECT 4.205000 50.495000 4.525000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 34.760000 4.930000 35.080000 ;
      LAYER met4 ;
        RECT 4.610000 34.760000 4.930000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 35.200000 4.930000 35.520000 ;
      LAYER met4 ;
        RECT 4.610000 35.200000 4.930000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 35.640000 4.930000 35.960000 ;
      LAYER met4 ;
        RECT 4.610000 35.640000 4.930000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 36.080000 4.930000 36.400000 ;
      LAYER met4 ;
        RECT 4.610000 36.080000 4.930000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 36.520000 4.930000 36.840000 ;
      LAYER met4 ;
        RECT 4.610000 36.520000 4.930000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 36.960000 4.930000 37.280000 ;
      LAYER met4 ;
        RECT 4.610000 36.960000 4.930000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 37.400000 4.930000 37.720000 ;
      LAYER met4 ;
        RECT 4.610000 37.400000 4.930000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 37.840000 4.930000 38.160000 ;
      LAYER met4 ;
        RECT 4.610000 37.840000 4.930000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 49.655000 4.930000 49.975000 ;
      LAYER met4 ;
        RECT 4.610000 49.655000 4.930000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 50.075000 4.930000 50.395000 ;
      LAYER met4 ;
        RECT 4.610000 50.075000 4.930000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 50.495000 4.930000 50.815000 ;
      LAYER met4 ;
        RECT 4.610000 50.495000 4.930000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 34.760000 5.335000 35.080000 ;
      LAYER met4 ;
        RECT 5.015000 34.760000 5.335000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 35.200000 5.335000 35.520000 ;
      LAYER met4 ;
        RECT 5.015000 35.200000 5.335000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 35.640000 5.335000 35.960000 ;
      LAYER met4 ;
        RECT 5.015000 35.640000 5.335000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 36.080000 5.335000 36.400000 ;
      LAYER met4 ;
        RECT 5.015000 36.080000 5.335000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 36.520000 5.335000 36.840000 ;
      LAYER met4 ;
        RECT 5.015000 36.520000 5.335000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 36.960000 5.335000 37.280000 ;
      LAYER met4 ;
        RECT 5.015000 36.960000 5.335000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 37.400000 5.335000 37.720000 ;
      LAYER met4 ;
        RECT 5.015000 37.400000 5.335000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 37.840000 5.335000 38.160000 ;
      LAYER met4 ;
        RECT 5.015000 37.840000 5.335000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 49.655000 5.335000 49.975000 ;
      LAYER met4 ;
        RECT 5.015000 49.655000 5.335000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 50.075000 5.335000 50.395000 ;
      LAYER met4 ;
        RECT 5.015000 50.075000 5.335000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 50.495000 5.335000 50.815000 ;
      LAYER met4 ;
        RECT 5.015000 50.495000 5.335000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 34.760000 5.740000 35.080000 ;
      LAYER met4 ;
        RECT 5.420000 34.760000 5.740000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 35.200000 5.740000 35.520000 ;
      LAYER met4 ;
        RECT 5.420000 35.200000 5.740000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 35.640000 5.740000 35.960000 ;
      LAYER met4 ;
        RECT 5.420000 35.640000 5.740000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 36.080000 5.740000 36.400000 ;
      LAYER met4 ;
        RECT 5.420000 36.080000 5.740000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 36.520000 5.740000 36.840000 ;
      LAYER met4 ;
        RECT 5.420000 36.520000 5.740000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 36.960000 5.740000 37.280000 ;
      LAYER met4 ;
        RECT 5.420000 36.960000 5.740000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 37.400000 5.740000 37.720000 ;
      LAYER met4 ;
        RECT 5.420000 37.400000 5.740000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 37.840000 5.740000 38.160000 ;
      LAYER met4 ;
        RECT 5.420000 37.840000 5.740000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 49.655000 5.740000 49.975000 ;
      LAYER met4 ;
        RECT 5.420000 49.655000 5.740000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 50.075000 5.740000 50.395000 ;
      LAYER met4 ;
        RECT 5.420000 50.075000 5.740000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 50.495000 5.740000 50.815000 ;
      LAYER met4 ;
        RECT 5.420000 50.495000 5.740000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 34.760000 6.145000 35.080000 ;
      LAYER met4 ;
        RECT 5.825000 34.760000 6.145000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 35.200000 6.145000 35.520000 ;
      LAYER met4 ;
        RECT 5.825000 35.200000 6.145000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 35.640000 6.145000 35.960000 ;
      LAYER met4 ;
        RECT 5.825000 35.640000 6.145000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 36.080000 6.145000 36.400000 ;
      LAYER met4 ;
        RECT 5.825000 36.080000 6.145000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 36.520000 6.145000 36.840000 ;
      LAYER met4 ;
        RECT 5.825000 36.520000 6.145000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 36.960000 6.145000 37.280000 ;
      LAYER met4 ;
        RECT 5.825000 36.960000 6.145000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 37.400000 6.145000 37.720000 ;
      LAYER met4 ;
        RECT 5.825000 37.400000 6.145000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 37.840000 6.145000 38.160000 ;
      LAYER met4 ;
        RECT 5.825000 37.840000 6.145000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 49.655000 6.145000 49.975000 ;
      LAYER met4 ;
        RECT 5.825000 49.655000 6.145000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 50.075000 6.145000 50.395000 ;
      LAYER met4 ;
        RECT 5.825000 50.075000 6.145000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 50.495000 6.145000 50.815000 ;
      LAYER met4 ;
        RECT 5.825000 50.495000 6.145000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 34.760000 51.105000 35.080000 ;
      LAYER met4 ;
        RECT 50.785000 34.760000 51.105000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 35.200000 51.105000 35.520000 ;
      LAYER met4 ;
        RECT 50.785000 35.200000 51.105000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 35.640000 51.105000 35.960000 ;
      LAYER met4 ;
        RECT 50.785000 35.640000 51.105000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 36.080000 51.105000 36.400000 ;
      LAYER met4 ;
        RECT 50.785000 36.080000 51.105000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 36.520000 51.105000 36.840000 ;
      LAYER met4 ;
        RECT 50.785000 36.520000 51.105000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 36.960000 51.105000 37.280000 ;
      LAYER met4 ;
        RECT 50.785000 36.960000 51.105000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 37.400000 51.105000 37.720000 ;
      LAYER met4 ;
        RECT 50.785000 37.400000 51.105000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 37.840000 51.105000 38.160000 ;
      LAYER met4 ;
        RECT 50.785000 37.840000 51.105000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 49.655000 51.105000 49.975000 ;
      LAYER met4 ;
        RECT 50.785000 49.655000 51.105000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 50.075000 51.105000 50.395000 ;
      LAYER met4 ;
        RECT 50.785000 50.075000 51.105000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 50.495000 51.105000 50.815000 ;
      LAYER met4 ;
        RECT 50.785000 50.495000 51.105000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 34.760000 51.515000 35.080000 ;
      LAYER met4 ;
        RECT 51.195000 34.760000 51.515000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 35.200000 51.515000 35.520000 ;
      LAYER met4 ;
        RECT 51.195000 35.200000 51.515000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 35.640000 51.515000 35.960000 ;
      LAYER met4 ;
        RECT 51.195000 35.640000 51.515000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 36.080000 51.515000 36.400000 ;
      LAYER met4 ;
        RECT 51.195000 36.080000 51.515000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 36.520000 51.515000 36.840000 ;
      LAYER met4 ;
        RECT 51.195000 36.520000 51.515000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 36.960000 51.515000 37.280000 ;
      LAYER met4 ;
        RECT 51.195000 36.960000 51.515000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 37.400000 51.515000 37.720000 ;
      LAYER met4 ;
        RECT 51.195000 37.400000 51.515000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 37.840000 51.515000 38.160000 ;
      LAYER met4 ;
        RECT 51.195000 37.840000 51.515000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 49.655000 51.515000 49.975000 ;
      LAYER met4 ;
        RECT 51.195000 49.655000 51.515000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 50.075000 51.515000 50.395000 ;
      LAYER met4 ;
        RECT 51.195000 50.075000 51.515000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 50.495000 51.515000 50.815000 ;
      LAYER met4 ;
        RECT 51.195000 50.495000 51.515000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 34.760000 51.925000 35.080000 ;
      LAYER met4 ;
        RECT 51.605000 34.760000 51.925000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 35.200000 51.925000 35.520000 ;
      LAYER met4 ;
        RECT 51.605000 35.200000 51.925000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 35.640000 51.925000 35.960000 ;
      LAYER met4 ;
        RECT 51.605000 35.640000 51.925000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 36.080000 51.925000 36.400000 ;
      LAYER met4 ;
        RECT 51.605000 36.080000 51.925000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 36.520000 51.925000 36.840000 ;
      LAYER met4 ;
        RECT 51.605000 36.520000 51.925000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 36.960000 51.925000 37.280000 ;
      LAYER met4 ;
        RECT 51.605000 36.960000 51.925000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 37.400000 51.925000 37.720000 ;
      LAYER met4 ;
        RECT 51.605000 37.400000 51.925000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 37.840000 51.925000 38.160000 ;
      LAYER met4 ;
        RECT 51.605000 37.840000 51.925000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 49.655000 51.925000 49.975000 ;
      LAYER met4 ;
        RECT 51.605000 49.655000 51.925000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 50.075000 51.925000 50.395000 ;
      LAYER met4 ;
        RECT 51.605000 50.075000 51.925000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 50.495000 51.925000 50.815000 ;
      LAYER met4 ;
        RECT 51.605000 50.495000 51.925000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 34.760000 52.335000 35.080000 ;
      LAYER met4 ;
        RECT 52.015000 34.760000 52.335000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 35.200000 52.335000 35.520000 ;
      LAYER met4 ;
        RECT 52.015000 35.200000 52.335000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 35.640000 52.335000 35.960000 ;
      LAYER met4 ;
        RECT 52.015000 35.640000 52.335000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 36.080000 52.335000 36.400000 ;
      LAYER met4 ;
        RECT 52.015000 36.080000 52.335000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 36.520000 52.335000 36.840000 ;
      LAYER met4 ;
        RECT 52.015000 36.520000 52.335000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 36.960000 52.335000 37.280000 ;
      LAYER met4 ;
        RECT 52.015000 36.960000 52.335000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 37.400000 52.335000 37.720000 ;
      LAYER met4 ;
        RECT 52.015000 37.400000 52.335000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 37.840000 52.335000 38.160000 ;
      LAYER met4 ;
        RECT 52.015000 37.840000 52.335000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 49.655000 52.335000 49.975000 ;
      LAYER met4 ;
        RECT 52.015000 49.655000 52.335000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 50.075000 52.335000 50.395000 ;
      LAYER met4 ;
        RECT 52.015000 50.075000 52.335000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 50.495000 52.335000 50.815000 ;
      LAYER met4 ;
        RECT 52.015000 50.495000 52.335000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 34.760000 52.745000 35.080000 ;
      LAYER met4 ;
        RECT 52.425000 34.760000 52.745000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 35.200000 52.745000 35.520000 ;
      LAYER met4 ;
        RECT 52.425000 35.200000 52.745000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 35.640000 52.745000 35.960000 ;
      LAYER met4 ;
        RECT 52.425000 35.640000 52.745000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 36.080000 52.745000 36.400000 ;
      LAYER met4 ;
        RECT 52.425000 36.080000 52.745000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 36.520000 52.745000 36.840000 ;
      LAYER met4 ;
        RECT 52.425000 36.520000 52.745000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 36.960000 52.745000 37.280000 ;
      LAYER met4 ;
        RECT 52.425000 36.960000 52.745000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 37.400000 52.745000 37.720000 ;
      LAYER met4 ;
        RECT 52.425000 37.400000 52.745000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 37.840000 52.745000 38.160000 ;
      LAYER met4 ;
        RECT 52.425000 37.840000 52.745000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 49.655000 52.745000 49.975000 ;
      LAYER met4 ;
        RECT 52.425000 49.655000 52.745000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 50.075000 52.745000 50.395000 ;
      LAYER met4 ;
        RECT 52.425000 50.075000 52.745000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 50.495000 52.745000 50.815000 ;
      LAYER met4 ;
        RECT 52.425000 50.495000 52.745000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 34.760000 53.155000 35.080000 ;
      LAYER met4 ;
        RECT 52.835000 34.760000 53.155000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 35.200000 53.155000 35.520000 ;
      LAYER met4 ;
        RECT 52.835000 35.200000 53.155000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 35.640000 53.155000 35.960000 ;
      LAYER met4 ;
        RECT 52.835000 35.640000 53.155000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 36.080000 53.155000 36.400000 ;
      LAYER met4 ;
        RECT 52.835000 36.080000 53.155000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 36.520000 53.155000 36.840000 ;
      LAYER met4 ;
        RECT 52.835000 36.520000 53.155000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 36.960000 53.155000 37.280000 ;
      LAYER met4 ;
        RECT 52.835000 36.960000 53.155000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 37.400000 53.155000 37.720000 ;
      LAYER met4 ;
        RECT 52.835000 37.400000 53.155000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 37.840000 53.155000 38.160000 ;
      LAYER met4 ;
        RECT 52.835000 37.840000 53.155000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 49.655000 53.155000 49.975000 ;
      LAYER met4 ;
        RECT 52.835000 49.655000 53.155000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 50.075000 53.155000 50.395000 ;
      LAYER met4 ;
        RECT 52.835000 50.075000 53.155000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 50.495000 53.155000 50.815000 ;
      LAYER met4 ;
        RECT 52.835000 50.495000 53.155000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 34.760000 53.565000 35.080000 ;
      LAYER met4 ;
        RECT 53.245000 34.760000 53.565000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 35.200000 53.565000 35.520000 ;
      LAYER met4 ;
        RECT 53.245000 35.200000 53.565000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 35.640000 53.565000 35.960000 ;
      LAYER met4 ;
        RECT 53.245000 35.640000 53.565000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 36.080000 53.565000 36.400000 ;
      LAYER met4 ;
        RECT 53.245000 36.080000 53.565000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 36.520000 53.565000 36.840000 ;
      LAYER met4 ;
        RECT 53.245000 36.520000 53.565000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 36.960000 53.565000 37.280000 ;
      LAYER met4 ;
        RECT 53.245000 36.960000 53.565000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 37.400000 53.565000 37.720000 ;
      LAYER met4 ;
        RECT 53.245000 37.400000 53.565000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 37.840000 53.565000 38.160000 ;
      LAYER met4 ;
        RECT 53.245000 37.840000 53.565000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 49.655000 53.565000 49.975000 ;
      LAYER met4 ;
        RECT 53.245000 49.655000 53.565000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 50.075000 53.565000 50.395000 ;
      LAYER met4 ;
        RECT 53.245000 50.075000 53.565000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 50.495000 53.565000 50.815000 ;
      LAYER met4 ;
        RECT 53.245000 50.495000 53.565000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 34.760000 53.970000 35.080000 ;
      LAYER met4 ;
        RECT 53.650000 34.760000 53.970000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 35.200000 53.970000 35.520000 ;
      LAYER met4 ;
        RECT 53.650000 35.200000 53.970000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 35.640000 53.970000 35.960000 ;
      LAYER met4 ;
        RECT 53.650000 35.640000 53.970000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 36.080000 53.970000 36.400000 ;
      LAYER met4 ;
        RECT 53.650000 36.080000 53.970000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 36.520000 53.970000 36.840000 ;
      LAYER met4 ;
        RECT 53.650000 36.520000 53.970000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 36.960000 53.970000 37.280000 ;
      LAYER met4 ;
        RECT 53.650000 36.960000 53.970000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 37.400000 53.970000 37.720000 ;
      LAYER met4 ;
        RECT 53.650000 37.400000 53.970000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 37.840000 53.970000 38.160000 ;
      LAYER met4 ;
        RECT 53.650000 37.840000 53.970000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 49.655000 53.970000 49.975000 ;
      LAYER met4 ;
        RECT 53.650000 49.655000 53.970000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 50.075000 53.970000 50.395000 ;
      LAYER met4 ;
        RECT 53.650000 50.075000 53.970000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 50.495000 53.970000 50.815000 ;
      LAYER met4 ;
        RECT 53.650000 50.495000 53.970000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 34.760000 54.375000 35.080000 ;
      LAYER met4 ;
        RECT 54.055000 34.760000 54.375000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 35.200000 54.375000 35.520000 ;
      LAYER met4 ;
        RECT 54.055000 35.200000 54.375000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 35.640000 54.375000 35.960000 ;
      LAYER met4 ;
        RECT 54.055000 35.640000 54.375000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 36.080000 54.375000 36.400000 ;
      LAYER met4 ;
        RECT 54.055000 36.080000 54.375000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 36.520000 54.375000 36.840000 ;
      LAYER met4 ;
        RECT 54.055000 36.520000 54.375000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 36.960000 54.375000 37.280000 ;
      LAYER met4 ;
        RECT 54.055000 36.960000 54.375000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 37.400000 54.375000 37.720000 ;
      LAYER met4 ;
        RECT 54.055000 37.400000 54.375000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 37.840000 54.375000 38.160000 ;
      LAYER met4 ;
        RECT 54.055000 37.840000 54.375000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 49.655000 54.375000 49.975000 ;
      LAYER met4 ;
        RECT 54.055000 49.655000 54.375000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 50.075000 54.375000 50.395000 ;
      LAYER met4 ;
        RECT 54.055000 50.075000 54.375000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 50.495000 54.375000 50.815000 ;
      LAYER met4 ;
        RECT 54.055000 50.495000 54.375000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 34.760000 54.780000 35.080000 ;
      LAYER met4 ;
        RECT 54.460000 34.760000 54.780000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 35.200000 54.780000 35.520000 ;
      LAYER met4 ;
        RECT 54.460000 35.200000 54.780000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 35.640000 54.780000 35.960000 ;
      LAYER met4 ;
        RECT 54.460000 35.640000 54.780000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 36.080000 54.780000 36.400000 ;
      LAYER met4 ;
        RECT 54.460000 36.080000 54.780000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 36.520000 54.780000 36.840000 ;
      LAYER met4 ;
        RECT 54.460000 36.520000 54.780000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 36.960000 54.780000 37.280000 ;
      LAYER met4 ;
        RECT 54.460000 36.960000 54.780000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 37.400000 54.780000 37.720000 ;
      LAYER met4 ;
        RECT 54.460000 37.400000 54.780000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 37.840000 54.780000 38.160000 ;
      LAYER met4 ;
        RECT 54.460000 37.840000 54.780000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 49.655000 54.780000 49.975000 ;
      LAYER met4 ;
        RECT 54.460000 49.655000 54.780000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 50.075000 54.780000 50.395000 ;
      LAYER met4 ;
        RECT 54.460000 50.075000 54.780000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 50.495000 54.780000 50.815000 ;
      LAYER met4 ;
        RECT 54.460000 50.495000 54.780000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 34.760000 55.185000 35.080000 ;
      LAYER met4 ;
        RECT 54.865000 34.760000 55.185000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 35.200000 55.185000 35.520000 ;
      LAYER met4 ;
        RECT 54.865000 35.200000 55.185000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 35.640000 55.185000 35.960000 ;
      LAYER met4 ;
        RECT 54.865000 35.640000 55.185000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 36.080000 55.185000 36.400000 ;
      LAYER met4 ;
        RECT 54.865000 36.080000 55.185000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 36.520000 55.185000 36.840000 ;
      LAYER met4 ;
        RECT 54.865000 36.520000 55.185000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 36.960000 55.185000 37.280000 ;
      LAYER met4 ;
        RECT 54.865000 36.960000 55.185000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 37.400000 55.185000 37.720000 ;
      LAYER met4 ;
        RECT 54.865000 37.400000 55.185000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 37.840000 55.185000 38.160000 ;
      LAYER met4 ;
        RECT 54.865000 37.840000 55.185000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 49.655000 55.185000 49.975000 ;
      LAYER met4 ;
        RECT 54.865000 49.655000 55.185000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 50.075000 55.185000 50.395000 ;
      LAYER met4 ;
        RECT 54.865000 50.075000 55.185000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 50.495000 55.185000 50.815000 ;
      LAYER met4 ;
        RECT 54.865000 50.495000 55.185000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 34.760000 55.590000 35.080000 ;
      LAYER met4 ;
        RECT 55.270000 34.760000 55.590000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 35.200000 55.590000 35.520000 ;
      LAYER met4 ;
        RECT 55.270000 35.200000 55.590000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 35.640000 55.590000 35.960000 ;
      LAYER met4 ;
        RECT 55.270000 35.640000 55.590000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 36.080000 55.590000 36.400000 ;
      LAYER met4 ;
        RECT 55.270000 36.080000 55.590000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 36.520000 55.590000 36.840000 ;
      LAYER met4 ;
        RECT 55.270000 36.520000 55.590000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 36.960000 55.590000 37.280000 ;
      LAYER met4 ;
        RECT 55.270000 36.960000 55.590000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 37.400000 55.590000 37.720000 ;
      LAYER met4 ;
        RECT 55.270000 37.400000 55.590000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 37.840000 55.590000 38.160000 ;
      LAYER met4 ;
        RECT 55.270000 37.840000 55.590000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 49.655000 55.590000 49.975000 ;
      LAYER met4 ;
        RECT 55.270000 49.655000 55.590000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 50.075000 55.590000 50.395000 ;
      LAYER met4 ;
        RECT 55.270000 50.075000 55.590000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 50.495000 55.590000 50.815000 ;
      LAYER met4 ;
        RECT 55.270000 50.495000 55.590000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 34.760000 55.995000 35.080000 ;
      LAYER met4 ;
        RECT 55.675000 34.760000 55.995000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 35.200000 55.995000 35.520000 ;
      LAYER met4 ;
        RECT 55.675000 35.200000 55.995000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 35.640000 55.995000 35.960000 ;
      LAYER met4 ;
        RECT 55.675000 35.640000 55.995000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 36.080000 55.995000 36.400000 ;
      LAYER met4 ;
        RECT 55.675000 36.080000 55.995000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 36.520000 55.995000 36.840000 ;
      LAYER met4 ;
        RECT 55.675000 36.520000 55.995000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 36.960000 55.995000 37.280000 ;
      LAYER met4 ;
        RECT 55.675000 36.960000 55.995000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 37.400000 55.995000 37.720000 ;
      LAYER met4 ;
        RECT 55.675000 37.400000 55.995000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 37.840000 55.995000 38.160000 ;
      LAYER met4 ;
        RECT 55.675000 37.840000 55.995000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 49.655000 55.995000 49.975000 ;
      LAYER met4 ;
        RECT 55.675000 49.655000 55.995000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 50.075000 55.995000 50.395000 ;
      LAYER met4 ;
        RECT 55.675000 50.075000 55.995000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 50.495000 55.995000 50.815000 ;
      LAYER met4 ;
        RECT 55.675000 50.495000 55.995000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 34.760000 56.400000 35.080000 ;
      LAYER met4 ;
        RECT 56.080000 34.760000 56.400000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 35.200000 56.400000 35.520000 ;
      LAYER met4 ;
        RECT 56.080000 35.200000 56.400000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 35.640000 56.400000 35.960000 ;
      LAYER met4 ;
        RECT 56.080000 35.640000 56.400000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 36.080000 56.400000 36.400000 ;
      LAYER met4 ;
        RECT 56.080000 36.080000 56.400000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 36.520000 56.400000 36.840000 ;
      LAYER met4 ;
        RECT 56.080000 36.520000 56.400000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 36.960000 56.400000 37.280000 ;
      LAYER met4 ;
        RECT 56.080000 36.960000 56.400000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 37.400000 56.400000 37.720000 ;
      LAYER met4 ;
        RECT 56.080000 37.400000 56.400000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 37.840000 56.400000 38.160000 ;
      LAYER met4 ;
        RECT 56.080000 37.840000 56.400000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 49.655000 56.400000 49.975000 ;
      LAYER met4 ;
        RECT 56.080000 49.655000 56.400000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 50.075000 56.400000 50.395000 ;
      LAYER met4 ;
        RECT 56.080000 50.075000 56.400000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 50.495000 56.400000 50.815000 ;
      LAYER met4 ;
        RECT 56.080000 50.495000 56.400000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 34.760000 56.805000 35.080000 ;
      LAYER met4 ;
        RECT 56.485000 34.760000 56.805000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 35.200000 56.805000 35.520000 ;
      LAYER met4 ;
        RECT 56.485000 35.200000 56.805000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 35.640000 56.805000 35.960000 ;
      LAYER met4 ;
        RECT 56.485000 35.640000 56.805000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 36.080000 56.805000 36.400000 ;
      LAYER met4 ;
        RECT 56.485000 36.080000 56.805000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 36.520000 56.805000 36.840000 ;
      LAYER met4 ;
        RECT 56.485000 36.520000 56.805000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 36.960000 56.805000 37.280000 ;
      LAYER met4 ;
        RECT 56.485000 36.960000 56.805000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 37.400000 56.805000 37.720000 ;
      LAYER met4 ;
        RECT 56.485000 37.400000 56.805000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 37.840000 56.805000 38.160000 ;
      LAYER met4 ;
        RECT 56.485000 37.840000 56.805000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 49.655000 56.805000 49.975000 ;
      LAYER met4 ;
        RECT 56.485000 49.655000 56.805000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 50.075000 56.805000 50.395000 ;
      LAYER met4 ;
        RECT 56.485000 50.075000 56.805000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 50.495000 56.805000 50.815000 ;
      LAYER met4 ;
        RECT 56.485000 50.495000 56.805000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 34.760000 57.210000 35.080000 ;
      LAYER met4 ;
        RECT 56.890000 34.760000 57.210000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 35.200000 57.210000 35.520000 ;
      LAYER met4 ;
        RECT 56.890000 35.200000 57.210000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 35.640000 57.210000 35.960000 ;
      LAYER met4 ;
        RECT 56.890000 35.640000 57.210000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 36.080000 57.210000 36.400000 ;
      LAYER met4 ;
        RECT 56.890000 36.080000 57.210000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 36.520000 57.210000 36.840000 ;
      LAYER met4 ;
        RECT 56.890000 36.520000 57.210000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 36.960000 57.210000 37.280000 ;
      LAYER met4 ;
        RECT 56.890000 36.960000 57.210000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 37.400000 57.210000 37.720000 ;
      LAYER met4 ;
        RECT 56.890000 37.400000 57.210000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 37.840000 57.210000 38.160000 ;
      LAYER met4 ;
        RECT 56.890000 37.840000 57.210000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 49.655000 57.210000 49.975000 ;
      LAYER met4 ;
        RECT 56.890000 49.655000 57.210000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 50.075000 57.210000 50.395000 ;
      LAYER met4 ;
        RECT 56.890000 50.075000 57.210000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 50.495000 57.210000 50.815000 ;
      LAYER met4 ;
        RECT 56.890000 50.495000 57.210000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 34.760000 57.615000 35.080000 ;
      LAYER met4 ;
        RECT 57.295000 34.760000 57.615000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 35.200000 57.615000 35.520000 ;
      LAYER met4 ;
        RECT 57.295000 35.200000 57.615000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 35.640000 57.615000 35.960000 ;
      LAYER met4 ;
        RECT 57.295000 35.640000 57.615000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 36.080000 57.615000 36.400000 ;
      LAYER met4 ;
        RECT 57.295000 36.080000 57.615000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 36.520000 57.615000 36.840000 ;
      LAYER met4 ;
        RECT 57.295000 36.520000 57.615000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 36.960000 57.615000 37.280000 ;
      LAYER met4 ;
        RECT 57.295000 36.960000 57.615000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 37.400000 57.615000 37.720000 ;
      LAYER met4 ;
        RECT 57.295000 37.400000 57.615000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 37.840000 57.615000 38.160000 ;
      LAYER met4 ;
        RECT 57.295000 37.840000 57.615000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 49.655000 57.615000 49.975000 ;
      LAYER met4 ;
        RECT 57.295000 49.655000 57.615000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 50.075000 57.615000 50.395000 ;
      LAYER met4 ;
        RECT 57.295000 50.075000 57.615000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 50.495000 57.615000 50.815000 ;
      LAYER met4 ;
        RECT 57.295000 50.495000 57.615000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 34.760000 58.020000 35.080000 ;
      LAYER met4 ;
        RECT 57.700000 34.760000 58.020000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 35.200000 58.020000 35.520000 ;
      LAYER met4 ;
        RECT 57.700000 35.200000 58.020000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 35.640000 58.020000 35.960000 ;
      LAYER met4 ;
        RECT 57.700000 35.640000 58.020000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 36.080000 58.020000 36.400000 ;
      LAYER met4 ;
        RECT 57.700000 36.080000 58.020000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 36.520000 58.020000 36.840000 ;
      LAYER met4 ;
        RECT 57.700000 36.520000 58.020000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 36.960000 58.020000 37.280000 ;
      LAYER met4 ;
        RECT 57.700000 36.960000 58.020000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 37.400000 58.020000 37.720000 ;
      LAYER met4 ;
        RECT 57.700000 37.400000 58.020000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 37.840000 58.020000 38.160000 ;
      LAYER met4 ;
        RECT 57.700000 37.840000 58.020000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 49.655000 58.020000 49.975000 ;
      LAYER met4 ;
        RECT 57.700000 49.655000 58.020000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 50.075000 58.020000 50.395000 ;
      LAYER met4 ;
        RECT 57.700000 50.075000 58.020000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 50.495000 58.020000 50.815000 ;
      LAYER met4 ;
        RECT 57.700000 50.495000 58.020000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 34.760000 58.425000 35.080000 ;
      LAYER met4 ;
        RECT 58.105000 34.760000 58.425000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 35.200000 58.425000 35.520000 ;
      LAYER met4 ;
        RECT 58.105000 35.200000 58.425000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 35.640000 58.425000 35.960000 ;
      LAYER met4 ;
        RECT 58.105000 35.640000 58.425000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 36.080000 58.425000 36.400000 ;
      LAYER met4 ;
        RECT 58.105000 36.080000 58.425000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 36.520000 58.425000 36.840000 ;
      LAYER met4 ;
        RECT 58.105000 36.520000 58.425000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 36.960000 58.425000 37.280000 ;
      LAYER met4 ;
        RECT 58.105000 36.960000 58.425000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 37.400000 58.425000 37.720000 ;
      LAYER met4 ;
        RECT 58.105000 37.400000 58.425000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 37.840000 58.425000 38.160000 ;
      LAYER met4 ;
        RECT 58.105000 37.840000 58.425000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 49.655000 58.425000 49.975000 ;
      LAYER met4 ;
        RECT 58.105000 49.655000 58.425000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 50.075000 58.425000 50.395000 ;
      LAYER met4 ;
        RECT 58.105000 50.075000 58.425000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 50.495000 58.425000 50.815000 ;
      LAYER met4 ;
        RECT 58.105000 50.495000 58.425000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 34.760000 58.830000 35.080000 ;
      LAYER met4 ;
        RECT 58.510000 34.760000 58.830000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 35.200000 58.830000 35.520000 ;
      LAYER met4 ;
        RECT 58.510000 35.200000 58.830000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 35.640000 58.830000 35.960000 ;
      LAYER met4 ;
        RECT 58.510000 35.640000 58.830000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 36.080000 58.830000 36.400000 ;
      LAYER met4 ;
        RECT 58.510000 36.080000 58.830000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 36.520000 58.830000 36.840000 ;
      LAYER met4 ;
        RECT 58.510000 36.520000 58.830000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 36.960000 58.830000 37.280000 ;
      LAYER met4 ;
        RECT 58.510000 36.960000 58.830000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 37.400000 58.830000 37.720000 ;
      LAYER met4 ;
        RECT 58.510000 37.400000 58.830000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 37.840000 58.830000 38.160000 ;
      LAYER met4 ;
        RECT 58.510000 37.840000 58.830000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 49.655000 58.830000 49.975000 ;
      LAYER met4 ;
        RECT 58.510000 49.655000 58.830000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 50.075000 58.830000 50.395000 ;
      LAYER met4 ;
        RECT 58.510000 50.075000 58.830000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 50.495000 58.830000 50.815000 ;
      LAYER met4 ;
        RECT 58.510000 50.495000 58.830000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 34.760000 59.235000 35.080000 ;
      LAYER met4 ;
        RECT 58.915000 34.760000 59.235000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 35.200000 59.235000 35.520000 ;
      LAYER met4 ;
        RECT 58.915000 35.200000 59.235000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 35.640000 59.235000 35.960000 ;
      LAYER met4 ;
        RECT 58.915000 35.640000 59.235000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 36.080000 59.235000 36.400000 ;
      LAYER met4 ;
        RECT 58.915000 36.080000 59.235000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 36.520000 59.235000 36.840000 ;
      LAYER met4 ;
        RECT 58.915000 36.520000 59.235000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 36.960000 59.235000 37.280000 ;
      LAYER met4 ;
        RECT 58.915000 36.960000 59.235000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 37.400000 59.235000 37.720000 ;
      LAYER met4 ;
        RECT 58.915000 37.400000 59.235000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 37.840000 59.235000 38.160000 ;
      LAYER met4 ;
        RECT 58.915000 37.840000 59.235000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 49.655000 59.235000 49.975000 ;
      LAYER met4 ;
        RECT 58.915000 49.655000 59.235000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 50.075000 59.235000 50.395000 ;
      LAYER met4 ;
        RECT 58.915000 50.075000 59.235000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 50.495000 59.235000 50.815000 ;
      LAYER met4 ;
        RECT 58.915000 50.495000 59.235000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 34.760000 59.640000 35.080000 ;
      LAYER met4 ;
        RECT 59.320000 34.760000 59.640000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 35.200000 59.640000 35.520000 ;
      LAYER met4 ;
        RECT 59.320000 35.200000 59.640000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 35.640000 59.640000 35.960000 ;
      LAYER met4 ;
        RECT 59.320000 35.640000 59.640000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 36.080000 59.640000 36.400000 ;
      LAYER met4 ;
        RECT 59.320000 36.080000 59.640000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 36.520000 59.640000 36.840000 ;
      LAYER met4 ;
        RECT 59.320000 36.520000 59.640000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 36.960000 59.640000 37.280000 ;
      LAYER met4 ;
        RECT 59.320000 36.960000 59.640000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 37.400000 59.640000 37.720000 ;
      LAYER met4 ;
        RECT 59.320000 37.400000 59.640000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 37.840000 59.640000 38.160000 ;
      LAYER met4 ;
        RECT 59.320000 37.840000 59.640000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 49.655000 59.640000 49.975000 ;
      LAYER met4 ;
        RECT 59.320000 49.655000 59.640000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 50.075000 59.640000 50.395000 ;
      LAYER met4 ;
        RECT 59.320000 50.075000 59.640000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 50.495000 59.640000 50.815000 ;
      LAYER met4 ;
        RECT 59.320000 50.495000 59.640000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 34.760000 60.045000 35.080000 ;
      LAYER met4 ;
        RECT 59.725000 34.760000 60.045000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 35.200000 60.045000 35.520000 ;
      LAYER met4 ;
        RECT 59.725000 35.200000 60.045000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 35.640000 60.045000 35.960000 ;
      LAYER met4 ;
        RECT 59.725000 35.640000 60.045000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 36.080000 60.045000 36.400000 ;
      LAYER met4 ;
        RECT 59.725000 36.080000 60.045000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 36.520000 60.045000 36.840000 ;
      LAYER met4 ;
        RECT 59.725000 36.520000 60.045000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 36.960000 60.045000 37.280000 ;
      LAYER met4 ;
        RECT 59.725000 36.960000 60.045000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 37.400000 60.045000 37.720000 ;
      LAYER met4 ;
        RECT 59.725000 37.400000 60.045000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 37.840000 60.045000 38.160000 ;
      LAYER met4 ;
        RECT 59.725000 37.840000 60.045000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 49.655000 60.045000 49.975000 ;
      LAYER met4 ;
        RECT 59.725000 49.655000 60.045000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 50.075000 60.045000 50.395000 ;
      LAYER met4 ;
        RECT 59.725000 50.075000 60.045000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 50.495000 60.045000 50.815000 ;
      LAYER met4 ;
        RECT 59.725000 50.495000 60.045000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 34.760000 6.550000 35.080000 ;
      LAYER met4 ;
        RECT 6.230000 34.760000 6.550000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 35.200000 6.550000 35.520000 ;
      LAYER met4 ;
        RECT 6.230000 35.200000 6.550000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 35.640000 6.550000 35.960000 ;
      LAYER met4 ;
        RECT 6.230000 35.640000 6.550000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 36.080000 6.550000 36.400000 ;
      LAYER met4 ;
        RECT 6.230000 36.080000 6.550000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 36.520000 6.550000 36.840000 ;
      LAYER met4 ;
        RECT 6.230000 36.520000 6.550000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 36.960000 6.550000 37.280000 ;
      LAYER met4 ;
        RECT 6.230000 36.960000 6.550000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 37.400000 6.550000 37.720000 ;
      LAYER met4 ;
        RECT 6.230000 37.400000 6.550000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 37.840000 6.550000 38.160000 ;
      LAYER met4 ;
        RECT 6.230000 37.840000 6.550000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 49.655000 6.550000 49.975000 ;
      LAYER met4 ;
        RECT 6.230000 49.655000 6.550000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 50.075000 6.550000 50.395000 ;
      LAYER met4 ;
        RECT 6.230000 50.075000 6.550000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 50.495000 6.550000 50.815000 ;
      LAYER met4 ;
        RECT 6.230000 50.495000 6.550000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 34.760000 6.955000 35.080000 ;
      LAYER met4 ;
        RECT 6.635000 34.760000 6.955000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 35.200000 6.955000 35.520000 ;
      LAYER met4 ;
        RECT 6.635000 35.200000 6.955000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 35.640000 6.955000 35.960000 ;
      LAYER met4 ;
        RECT 6.635000 35.640000 6.955000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 36.080000 6.955000 36.400000 ;
      LAYER met4 ;
        RECT 6.635000 36.080000 6.955000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 36.520000 6.955000 36.840000 ;
      LAYER met4 ;
        RECT 6.635000 36.520000 6.955000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 36.960000 6.955000 37.280000 ;
      LAYER met4 ;
        RECT 6.635000 36.960000 6.955000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 37.400000 6.955000 37.720000 ;
      LAYER met4 ;
        RECT 6.635000 37.400000 6.955000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 37.840000 6.955000 38.160000 ;
      LAYER met4 ;
        RECT 6.635000 37.840000 6.955000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 49.655000 6.955000 49.975000 ;
      LAYER met4 ;
        RECT 6.635000 49.655000 6.955000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 50.075000 6.955000 50.395000 ;
      LAYER met4 ;
        RECT 6.635000 50.075000 6.955000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 50.495000 6.955000 50.815000 ;
      LAYER met4 ;
        RECT 6.635000 50.495000 6.955000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 34.760000 60.450000 35.080000 ;
      LAYER met4 ;
        RECT 60.130000 34.760000 60.450000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 35.200000 60.450000 35.520000 ;
      LAYER met4 ;
        RECT 60.130000 35.200000 60.450000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 35.640000 60.450000 35.960000 ;
      LAYER met4 ;
        RECT 60.130000 35.640000 60.450000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 36.080000 60.450000 36.400000 ;
      LAYER met4 ;
        RECT 60.130000 36.080000 60.450000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 36.520000 60.450000 36.840000 ;
      LAYER met4 ;
        RECT 60.130000 36.520000 60.450000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 36.960000 60.450000 37.280000 ;
      LAYER met4 ;
        RECT 60.130000 36.960000 60.450000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 37.400000 60.450000 37.720000 ;
      LAYER met4 ;
        RECT 60.130000 37.400000 60.450000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 37.840000 60.450000 38.160000 ;
      LAYER met4 ;
        RECT 60.130000 37.840000 60.450000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 49.655000 60.450000 49.975000 ;
      LAYER met4 ;
        RECT 60.130000 49.655000 60.450000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 50.075000 60.450000 50.395000 ;
      LAYER met4 ;
        RECT 60.130000 50.075000 60.450000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 50.495000 60.450000 50.815000 ;
      LAYER met4 ;
        RECT 60.130000 50.495000 60.450000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 34.760000 60.855000 35.080000 ;
      LAYER met4 ;
        RECT 60.535000 34.760000 60.855000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 35.200000 60.855000 35.520000 ;
      LAYER met4 ;
        RECT 60.535000 35.200000 60.855000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 35.640000 60.855000 35.960000 ;
      LAYER met4 ;
        RECT 60.535000 35.640000 60.855000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 36.080000 60.855000 36.400000 ;
      LAYER met4 ;
        RECT 60.535000 36.080000 60.855000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 36.520000 60.855000 36.840000 ;
      LAYER met4 ;
        RECT 60.535000 36.520000 60.855000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 36.960000 60.855000 37.280000 ;
      LAYER met4 ;
        RECT 60.535000 36.960000 60.855000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 37.400000 60.855000 37.720000 ;
      LAYER met4 ;
        RECT 60.535000 37.400000 60.855000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 37.840000 60.855000 38.160000 ;
      LAYER met4 ;
        RECT 60.535000 37.840000 60.855000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 49.655000 60.855000 49.975000 ;
      LAYER met4 ;
        RECT 60.535000 49.655000 60.855000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 50.075000 60.855000 50.395000 ;
      LAYER met4 ;
        RECT 60.535000 50.075000 60.855000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 50.495000 60.855000 50.815000 ;
      LAYER met4 ;
        RECT 60.535000 50.495000 60.855000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 34.760000 61.260000 35.080000 ;
      LAYER met4 ;
        RECT 60.940000 34.760000 61.260000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 35.200000 61.260000 35.520000 ;
      LAYER met4 ;
        RECT 60.940000 35.200000 61.260000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 35.640000 61.260000 35.960000 ;
      LAYER met4 ;
        RECT 60.940000 35.640000 61.260000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 36.080000 61.260000 36.400000 ;
      LAYER met4 ;
        RECT 60.940000 36.080000 61.260000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 36.520000 61.260000 36.840000 ;
      LAYER met4 ;
        RECT 60.940000 36.520000 61.260000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 36.960000 61.260000 37.280000 ;
      LAYER met4 ;
        RECT 60.940000 36.960000 61.260000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 37.400000 61.260000 37.720000 ;
      LAYER met4 ;
        RECT 60.940000 37.400000 61.260000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 37.840000 61.260000 38.160000 ;
      LAYER met4 ;
        RECT 60.940000 37.840000 61.260000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 49.655000 61.260000 49.975000 ;
      LAYER met4 ;
        RECT 60.940000 49.655000 61.260000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 50.075000 61.260000 50.395000 ;
      LAYER met4 ;
        RECT 60.940000 50.075000 61.260000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 50.495000 61.260000 50.815000 ;
      LAYER met4 ;
        RECT 60.940000 50.495000 61.260000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 34.760000 61.665000 35.080000 ;
      LAYER met4 ;
        RECT 61.345000 34.760000 61.665000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 35.200000 61.665000 35.520000 ;
      LAYER met4 ;
        RECT 61.345000 35.200000 61.665000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 35.640000 61.665000 35.960000 ;
      LAYER met4 ;
        RECT 61.345000 35.640000 61.665000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 36.080000 61.665000 36.400000 ;
      LAYER met4 ;
        RECT 61.345000 36.080000 61.665000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 36.520000 61.665000 36.840000 ;
      LAYER met4 ;
        RECT 61.345000 36.520000 61.665000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 36.960000 61.665000 37.280000 ;
      LAYER met4 ;
        RECT 61.345000 36.960000 61.665000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 37.400000 61.665000 37.720000 ;
      LAYER met4 ;
        RECT 61.345000 37.400000 61.665000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 37.840000 61.665000 38.160000 ;
      LAYER met4 ;
        RECT 61.345000 37.840000 61.665000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 49.655000 61.665000 49.975000 ;
      LAYER met4 ;
        RECT 61.345000 49.655000 61.665000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 50.075000 61.665000 50.395000 ;
      LAYER met4 ;
        RECT 61.345000 50.075000 61.665000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 50.495000 61.665000 50.815000 ;
      LAYER met4 ;
        RECT 61.345000 50.495000 61.665000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 34.760000 62.070000 35.080000 ;
      LAYER met4 ;
        RECT 61.750000 34.760000 62.070000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 35.200000 62.070000 35.520000 ;
      LAYER met4 ;
        RECT 61.750000 35.200000 62.070000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 35.640000 62.070000 35.960000 ;
      LAYER met4 ;
        RECT 61.750000 35.640000 62.070000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 36.080000 62.070000 36.400000 ;
      LAYER met4 ;
        RECT 61.750000 36.080000 62.070000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 36.520000 62.070000 36.840000 ;
      LAYER met4 ;
        RECT 61.750000 36.520000 62.070000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 36.960000 62.070000 37.280000 ;
      LAYER met4 ;
        RECT 61.750000 36.960000 62.070000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 37.400000 62.070000 37.720000 ;
      LAYER met4 ;
        RECT 61.750000 37.400000 62.070000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 37.840000 62.070000 38.160000 ;
      LAYER met4 ;
        RECT 61.750000 37.840000 62.070000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 49.655000 62.070000 49.975000 ;
      LAYER met4 ;
        RECT 61.750000 49.655000 62.070000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 50.075000 62.070000 50.395000 ;
      LAYER met4 ;
        RECT 61.750000 50.075000 62.070000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 50.495000 62.070000 50.815000 ;
      LAYER met4 ;
        RECT 61.750000 50.495000 62.070000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 34.760000 62.475000 35.080000 ;
      LAYER met4 ;
        RECT 62.155000 34.760000 62.475000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 35.200000 62.475000 35.520000 ;
      LAYER met4 ;
        RECT 62.155000 35.200000 62.475000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 35.640000 62.475000 35.960000 ;
      LAYER met4 ;
        RECT 62.155000 35.640000 62.475000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 36.080000 62.475000 36.400000 ;
      LAYER met4 ;
        RECT 62.155000 36.080000 62.475000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 36.520000 62.475000 36.840000 ;
      LAYER met4 ;
        RECT 62.155000 36.520000 62.475000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 36.960000 62.475000 37.280000 ;
      LAYER met4 ;
        RECT 62.155000 36.960000 62.475000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 37.400000 62.475000 37.720000 ;
      LAYER met4 ;
        RECT 62.155000 37.400000 62.475000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 37.840000 62.475000 38.160000 ;
      LAYER met4 ;
        RECT 62.155000 37.840000 62.475000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 49.655000 62.475000 49.975000 ;
      LAYER met4 ;
        RECT 62.155000 49.655000 62.475000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 50.075000 62.475000 50.395000 ;
      LAYER met4 ;
        RECT 62.155000 50.075000 62.475000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 50.495000 62.475000 50.815000 ;
      LAYER met4 ;
        RECT 62.155000 50.495000 62.475000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 34.760000 62.880000 35.080000 ;
      LAYER met4 ;
        RECT 62.560000 34.760000 62.880000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 35.200000 62.880000 35.520000 ;
      LAYER met4 ;
        RECT 62.560000 35.200000 62.880000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 35.640000 62.880000 35.960000 ;
      LAYER met4 ;
        RECT 62.560000 35.640000 62.880000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 36.080000 62.880000 36.400000 ;
      LAYER met4 ;
        RECT 62.560000 36.080000 62.880000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 36.520000 62.880000 36.840000 ;
      LAYER met4 ;
        RECT 62.560000 36.520000 62.880000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 36.960000 62.880000 37.280000 ;
      LAYER met4 ;
        RECT 62.560000 36.960000 62.880000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 37.400000 62.880000 37.720000 ;
      LAYER met4 ;
        RECT 62.560000 37.400000 62.880000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 37.840000 62.880000 38.160000 ;
      LAYER met4 ;
        RECT 62.560000 37.840000 62.880000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 49.655000 62.880000 49.975000 ;
      LAYER met4 ;
        RECT 62.560000 49.655000 62.880000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 50.075000 62.880000 50.395000 ;
      LAYER met4 ;
        RECT 62.560000 50.075000 62.880000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 50.495000 62.880000 50.815000 ;
      LAYER met4 ;
        RECT 62.560000 50.495000 62.880000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 34.760000 63.285000 35.080000 ;
      LAYER met4 ;
        RECT 62.965000 34.760000 63.285000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 35.200000 63.285000 35.520000 ;
      LAYER met4 ;
        RECT 62.965000 35.200000 63.285000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 35.640000 63.285000 35.960000 ;
      LAYER met4 ;
        RECT 62.965000 35.640000 63.285000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 36.080000 63.285000 36.400000 ;
      LAYER met4 ;
        RECT 62.965000 36.080000 63.285000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 36.520000 63.285000 36.840000 ;
      LAYER met4 ;
        RECT 62.965000 36.520000 63.285000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 36.960000 63.285000 37.280000 ;
      LAYER met4 ;
        RECT 62.965000 36.960000 63.285000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 37.400000 63.285000 37.720000 ;
      LAYER met4 ;
        RECT 62.965000 37.400000 63.285000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 37.840000 63.285000 38.160000 ;
      LAYER met4 ;
        RECT 62.965000 37.840000 63.285000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 49.655000 63.285000 49.975000 ;
      LAYER met4 ;
        RECT 62.965000 49.655000 63.285000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 50.075000 63.285000 50.395000 ;
      LAYER met4 ;
        RECT 62.965000 50.075000 63.285000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 50.495000 63.285000 50.815000 ;
      LAYER met4 ;
        RECT 62.965000 50.495000 63.285000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 34.760000 63.690000 35.080000 ;
      LAYER met4 ;
        RECT 63.370000 34.760000 63.690000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 35.200000 63.690000 35.520000 ;
      LAYER met4 ;
        RECT 63.370000 35.200000 63.690000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 35.640000 63.690000 35.960000 ;
      LAYER met4 ;
        RECT 63.370000 35.640000 63.690000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 36.080000 63.690000 36.400000 ;
      LAYER met4 ;
        RECT 63.370000 36.080000 63.690000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 36.520000 63.690000 36.840000 ;
      LAYER met4 ;
        RECT 63.370000 36.520000 63.690000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 36.960000 63.690000 37.280000 ;
      LAYER met4 ;
        RECT 63.370000 36.960000 63.690000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 37.400000 63.690000 37.720000 ;
      LAYER met4 ;
        RECT 63.370000 37.400000 63.690000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 37.840000 63.690000 38.160000 ;
      LAYER met4 ;
        RECT 63.370000 37.840000 63.690000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 49.655000 63.690000 49.975000 ;
      LAYER met4 ;
        RECT 63.370000 49.655000 63.690000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 50.075000 63.690000 50.395000 ;
      LAYER met4 ;
        RECT 63.370000 50.075000 63.690000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 50.495000 63.690000 50.815000 ;
      LAYER met4 ;
        RECT 63.370000 50.495000 63.690000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 34.760000 64.095000 35.080000 ;
      LAYER met4 ;
        RECT 63.775000 34.760000 64.095000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 35.200000 64.095000 35.520000 ;
      LAYER met4 ;
        RECT 63.775000 35.200000 64.095000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 35.640000 64.095000 35.960000 ;
      LAYER met4 ;
        RECT 63.775000 35.640000 64.095000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 36.080000 64.095000 36.400000 ;
      LAYER met4 ;
        RECT 63.775000 36.080000 64.095000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 36.520000 64.095000 36.840000 ;
      LAYER met4 ;
        RECT 63.775000 36.520000 64.095000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 36.960000 64.095000 37.280000 ;
      LAYER met4 ;
        RECT 63.775000 36.960000 64.095000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 37.400000 64.095000 37.720000 ;
      LAYER met4 ;
        RECT 63.775000 37.400000 64.095000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 37.840000 64.095000 38.160000 ;
      LAYER met4 ;
        RECT 63.775000 37.840000 64.095000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 49.655000 64.095000 49.975000 ;
      LAYER met4 ;
        RECT 63.775000 49.655000 64.095000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 50.075000 64.095000 50.395000 ;
      LAYER met4 ;
        RECT 63.775000 50.075000 64.095000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 50.495000 64.095000 50.815000 ;
      LAYER met4 ;
        RECT 63.775000 50.495000 64.095000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 34.760000 64.500000 35.080000 ;
      LAYER met4 ;
        RECT 64.180000 34.760000 64.500000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 35.200000 64.500000 35.520000 ;
      LAYER met4 ;
        RECT 64.180000 35.200000 64.500000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 35.640000 64.500000 35.960000 ;
      LAYER met4 ;
        RECT 64.180000 35.640000 64.500000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 36.080000 64.500000 36.400000 ;
      LAYER met4 ;
        RECT 64.180000 36.080000 64.500000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 36.520000 64.500000 36.840000 ;
      LAYER met4 ;
        RECT 64.180000 36.520000 64.500000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 36.960000 64.500000 37.280000 ;
      LAYER met4 ;
        RECT 64.180000 36.960000 64.500000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 37.400000 64.500000 37.720000 ;
      LAYER met4 ;
        RECT 64.180000 37.400000 64.500000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 37.840000 64.500000 38.160000 ;
      LAYER met4 ;
        RECT 64.180000 37.840000 64.500000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 49.655000 64.500000 49.975000 ;
      LAYER met4 ;
        RECT 64.180000 49.655000 64.500000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 50.075000 64.500000 50.395000 ;
      LAYER met4 ;
        RECT 64.180000 50.075000 64.500000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 50.495000 64.500000 50.815000 ;
      LAYER met4 ;
        RECT 64.180000 50.495000 64.500000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 34.760000 64.905000 35.080000 ;
      LAYER met4 ;
        RECT 64.585000 34.760000 64.905000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 35.200000 64.905000 35.520000 ;
      LAYER met4 ;
        RECT 64.585000 35.200000 64.905000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 35.640000 64.905000 35.960000 ;
      LAYER met4 ;
        RECT 64.585000 35.640000 64.905000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 36.080000 64.905000 36.400000 ;
      LAYER met4 ;
        RECT 64.585000 36.080000 64.905000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 36.520000 64.905000 36.840000 ;
      LAYER met4 ;
        RECT 64.585000 36.520000 64.905000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 36.960000 64.905000 37.280000 ;
      LAYER met4 ;
        RECT 64.585000 36.960000 64.905000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 37.400000 64.905000 37.720000 ;
      LAYER met4 ;
        RECT 64.585000 37.400000 64.905000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 37.840000 64.905000 38.160000 ;
      LAYER met4 ;
        RECT 64.585000 37.840000 64.905000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 49.655000 64.905000 49.975000 ;
      LAYER met4 ;
        RECT 64.585000 49.655000 64.905000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 50.075000 64.905000 50.395000 ;
      LAYER met4 ;
        RECT 64.585000 50.075000 64.905000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 50.495000 64.905000 50.815000 ;
      LAYER met4 ;
        RECT 64.585000 50.495000 64.905000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 34.760000 65.310000 35.080000 ;
      LAYER met4 ;
        RECT 64.990000 34.760000 65.310000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 35.200000 65.310000 35.520000 ;
      LAYER met4 ;
        RECT 64.990000 35.200000 65.310000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 35.640000 65.310000 35.960000 ;
      LAYER met4 ;
        RECT 64.990000 35.640000 65.310000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 36.080000 65.310000 36.400000 ;
      LAYER met4 ;
        RECT 64.990000 36.080000 65.310000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 36.520000 65.310000 36.840000 ;
      LAYER met4 ;
        RECT 64.990000 36.520000 65.310000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 36.960000 65.310000 37.280000 ;
      LAYER met4 ;
        RECT 64.990000 36.960000 65.310000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 37.400000 65.310000 37.720000 ;
      LAYER met4 ;
        RECT 64.990000 37.400000 65.310000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 37.840000 65.310000 38.160000 ;
      LAYER met4 ;
        RECT 64.990000 37.840000 65.310000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 49.655000 65.310000 49.975000 ;
      LAYER met4 ;
        RECT 64.990000 49.655000 65.310000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 50.075000 65.310000 50.395000 ;
      LAYER met4 ;
        RECT 64.990000 50.075000 65.310000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 50.495000 65.310000 50.815000 ;
      LAYER met4 ;
        RECT 64.990000 50.495000 65.310000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 34.760000 65.715000 35.080000 ;
      LAYER met4 ;
        RECT 65.395000 34.760000 65.715000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 35.200000 65.715000 35.520000 ;
      LAYER met4 ;
        RECT 65.395000 35.200000 65.715000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 35.640000 65.715000 35.960000 ;
      LAYER met4 ;
        RECT 65.395000 35.640000 65.715000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 36.080000 65.715000 36.400000 ;
      LAYER met4 ;
        RECT 65.395000 36.080000 65.715000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 36.520000 65.715000 36.840000 ;
      LAYER met4 ;
        RECT 65.395000 36.520000 65.715000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 36.960000 65.715000 37.280000 ;
      LAYER met4 ;
        RECT 65.395000 36.960000 65.715000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 37.400000 65.715000 37.720000 ;
      LAYER met4 ;
        RECT 65.395000 37.400000 65.715000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 37.840000 65.715000 38.160000 ;
      LAYER met4 ;
        RECT 65.395000 37.840000 65.715000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 49.655000 65.715000 49.975000 ;
      LAYER met4 ;
        RECT 65.395000 49.655000 65.715000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 50.075000 65.715000 50.395000 ;
      LAYER met4 ;
        RECT 65.395000 50.075000 65.715000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 50.495000 65.715000 50.815000 ;
      LAYER met4 ;
        RECT 65.395000 50.495000 65.715000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 34.760000 66.120000 35.080000 ;
      LAYER met4 ;
        RECT 65.800000 34.760000 66.120000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 35.200000 66.120000 35.520000 ;
      LAYER met4 ;
        RECT 65.800000 35.200000 66.120000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 35.640000 66.120000 35.960000 ;
      LAYER met4 ;
        RECT 65.800000 35.640000 66.120000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 36.080000 66.120000 36.400000 ;
      LAYER met4 ;
        RECT 65.800000 36.080000 66.120000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 36.520000 66.120000 36.840000 ;
      LAYER met4 ;
        RECT 65.800000 36.520000 66.120000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 36.960000 66.120000 37.280000 ;
      LAYER met4 ;
        RECT 65.800000 36.960000 66.120000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 37.400000 66.120000 37.720000 ;
      LAYER met4 ;
        RECT 65.800000 37.400000 66.120000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 37.840000 66.120000 38.160000 ;
      LAYER met4 ;
        RECT 65.800000 37.840000 66.120000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 49.655000 66.120000 49.975000 ;
      LAYER met4 ;
        RECT 65.800000 49.655000 66.120000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 50.075000 66.120000 50.395000 ;
      LAYER met4 ;
        RECT 65.800000 50.075000 66.120000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 50.495000 66.120000 50.815000 ;
      LAYER met4 ;
        RECT 65.800000 50.495000 66.120000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 34.760000 66.525000 35.080000 ;
      LAYER met4 ;
        RECT 66.205000 34.760000 66.525000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 35.200000 66.525000 35.520000 ;
      LAYER met4 ;
        RECT 66.205000 35.200000 66.525000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 35.640000 66.525000 35.960000 ;
      LAYER met4 ;
        RECT 66.205000 35.640000 66.525000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 36.080000 66.525000 36.400000 ;
      LAYER met4 ;
        RECT 66.205000 36.080000 66.525000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 36.520000 66.525000 36.840000 ;
      LAYER met4 ;
        RECT 66.205000 36.520000 66.525000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 36.960000 66.525000 37.280000 ;
      LAYER met4 ;
        RECT 66.205000 36.960000 66.525000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 37.400000 66.525000 37.720000 ;
      LAYER met4 ;
        RECT 66.205000 37.400000 66.525000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 37.840000 66.525000 38.160000 ;
      LAYER met4 ;
        RECT 66.205000 37.840000 66.525000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 49.655000 66.525000 49.975000 ;
      LAYER met4 ;
        RECT 66.205000 49.655000 66.525000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 50.075000 66.525000 50.395000 ;
      LAYER met4 ;
        RECT 66.205000 50.075000 66.525000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 50.495000 66.525000 50.815000 ;
      LAYER met4 ;
        RECT 66.205000 50.495000 66.525000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 34.760000 66.930000 35.080000 ;
      LAYER met4 ;
        RECT 66.610000 34.760000 66.930000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 35.200000 66.930000 35.520000 ;
      LAYER met4 ;
        RECT 66.610000 35.200000 66.930000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 35.640000 66.930000 35.960000 ;
      LAYER met4 ;
        RECT 66.610000 35.640000 66.930000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 36.080000 66.930000 36.400000 ;
      LAYER met4 ;
        RECT 66.610000 36.080000 66.930000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 36.520000 66.930000 36.840000 ;
      LAYER met4 ;
        RECT 66.610000 36.520000 66.930000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 36.960000 66.930000 37.280000 ;
      LAYER met4 ;
        RECT 66.610000 36.960000 66.930000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 37.400000 66.930000 37.720000 ;
      LAYER met4 ;
        RECT 66.610000 37.400000 66.930000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 37.840000 66.930000 38.160000 ;
      LAYER met4 ;
        RECT 66.610000 37.840000 66.930000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 49.655000 66.930000 49.975000 ;
      LAYER met4 ;
        RECT 66.610000 49.655000 66.930000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 50.075000 66.930000 50.395000 ;
      LAYER met4 ;
        RECT 66.610000 50.075000 66.930000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 50.495000 66.930000 50.815000 ;
      LAYER met4 ;
        RECT 66.610000 50.495000 66.930000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 34.760000 67.335000 35.080000 ;
      LAYER met4 ;
        RECT 67.015000 34.760000 67.335000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 35.200000 67.335000 35.520000 ;
      LAYER met4 ;
        RECT 67.015000 35.200000 67.335000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 35.640000 67.335000 35.960000 ;
      LAYER met4 ;
        RECT 67.015000 35.640000 67.335000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 36.080000 67.335000 36.400000 ;
      LAYER met4 ;
        RECT 67.015000 36.080000 67.335000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 36.520000 67.335000 36.840000 ;
      LAYER met4 ;
        RECT 67.015000 36.520000 67.335000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 36.960000 67.335000 37.280000 ;
      LAYER met4 ;
        RECT 67.015000 36.960000 67.335000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 37.400000 67.335000 37.720000 ;
      LAYER met4 ;
        RECT 67.015000 37.400000 67.335000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 37.840000 67.335000 38.160000 ;
      LAYER met4 ;
        RECT 67.015000 37.840000 67.335000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 49.655000 67.335000 49.975000 ;
      LAYER met4 ;
        RECT 67.015000 49.655000 67.335000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 50.075000 67.335000 50.395000 ;
      LAYER met4 ;
        RECT 67.015000 50.075000 67.335000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 50.495000 67.335000 50.815000 ;
      LAYER met4 ;
        RECT 67.015000 50.495000 67.335000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 34.760000 67.740000 35.080000 ;
      LAYER met4 ;
        RECT 67.420000 34.760000 67.740000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 35.200000 67.740000 35.520000 ;
      LAYER met4 ;
        RECT 67.420000 35.200000 67.740000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 35.640000 67.740000 35.960000 ;
      LAYER met4 ;
        RECT 67.420000 35.640000 67.740000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 36.080000 67.740000 36.400000 ;
      LAYER met4 ;
        RECT 67.420000 36.080000 67.740000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 36.520000 67.740000 36.840000 ;
      LAYER met4 ;
        RECT 67.420000 36.520000 67.740000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 36.960000 67.740000 37.280000 ;
      LAYER met4 ;
        RECT 67.420000 36.960000 67.740000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 37.400000 67.740000 37.720000 ;
      LAYER met4 ;
        RECT 67.420000 37.400000 67.740000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 37.840000 67.740000 38.160000 ;
      LAYER met4 ;
        RECT 67.420000 37.840000 67.740000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 49.655000 67.740000 49.975000 ;
      LAYER met4 ;
        RECT 67.420000 49.655000 67.740000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 50.075000 67.740000 50.395000 ;
      LAYER met4 ;
        RECT 67.420000 50.075000 67.740000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 50.495000 67.740000 50.815000 ;
      LAYER met4 ;
        RECT 67.420000 50.495000 67.740000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 34.760000 68.145000 35.080000 ;
      LAYER met4 ;
        RECT 67.825000 34.760000 68.145000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 35.200000 68.145000 35.520000 ;
      LAYER met4 ;
        RECT 67.825000 35.200000 68.145000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 35.640000 68.145000 35.960000 ;
      LAYER met4 ;
        RECT 67.825000 35.640000 68.145000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 36.080000 68.145000 36.400000 ;
      LAYER met4 ;
        RECT 67.825000 36.080000 68.145000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 36.520000 68.145000 36.840000 ;
      LAYER met4 ;
        RECT 67.825000 36.520000 68.145000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 36.960000 68.145000 37.280000 ;
      LAYER met4 ;
        RECT 67.825000 36.960000 68.145000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 37.400000 68.145000 37.720000 ;
      LAYER met4 ;
        RECT 67.825000 37.400000 68.145000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 37.840000 68.145000 38.160000 ;
      LAYER met4 ;
        RECT 67.825000 37.840000 68.145000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 49.655000 68.145000 49.975000 ;
      LAYER met4 ;
        RECT 67.825000 49.655000 68.145000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 50.075000 68.145000 50.395000 ;
      LAYER met4 ;
        RECT 67.825000 50.075000 68.145000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 50.495000 68.145000 50.815000 ;
      LAYER met4 ;
        RECT 67.825000 50.495000 68.145000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 34.760000 68.550000 35.080000 ;
      LAYER met4 ;
        RECT 68.230000 34.760000 68.550000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 35.200000 68.550000 35.520000 ;
      LAYER met4 ;
        RECT 68.230000 35.200000 68.550000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 35.640000 68.550000 35.960000 ;
      LAYER met4 ;
        RECT 68.230000 35.640000 68.550000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 36.080000 68.550000 36.400000 ;
      LAYER met4 ;
        RECT 68.230000 36.080000 68.550000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 36.520000 68.550000 36.840000 ;
      LAYER met4 ;
        RECT 68.230000 36.520000 68.550000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 36.960000 68.550000 37.280000 ;
      LAYER met4 ;
        RECT 68.230000 36.960000 68.550000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 37.400000 68.550000 37.720000 ;
      LAYER met4 ;
        RECT 68.230000 37.400000 68.550000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 37.840000 68.550000 38.160000 ;
      LAYER met4 ;
        RECT 68.230000 37.840000 68.550000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 49.655000 68.550000 49.975000 ;
      LAYER met4 ;
        RECT 68.230000 49.655000 68.550000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 50.075000 68.550000 50.395000 ;
      LAYER met4 ;
        RECT 68.230000 50.075000 68.550000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 50.495000 68.550000 50.815000 ;
      LAYER met4 ;
        RECT 68.230000 50.495000 68.550000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 34.760000 68.955000 35.080000 ;
      LAYER met4 ;
        RECT 68.635000 34.760000 68.955000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 35.200000 68.955000 35.520000 ;
      LAYER met4 ;
        RECT 68.635000 35.200000 68.955000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 35.640000 68.955000 35.960000 ;
      LAYER met4 ;
        RECT 68.635000 35.640000 68.955000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 36.080000 68.955000 36.400000 ;
      LAYER met4 ;
        RECT 68.635000 36.080000 68.955000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 36.520000 68.955000 36.840000 ;
      LAYER met4 ;
        RECT 68.635000 36.520000 68.955000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 36.960000 68.955000 37.280000 ;
      LAYER met4 ;
        RECT 68.635000 36.960000 68.955000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 37.400000 68.955000 37.720000 ;
      LAYER met4 ;
        RECT 68.635000 37.400000 68.955000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 37.840000 68.955000 38.160000 ;
      LAYER met4 ;
        RECT 68.635000 37.840000 68.955000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 49.655000 68.955000 49.975000 ;
      LAYER met4 ;
        RECT 68.635000 49.655000 68.955000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 50.075000 68.955000 50.395000 ;
      LAYER met4 ;
        RECT 68.635000 50.075000 68.955000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 50.495000 68.955000 50.815000 ;
      LAYER met4 ;
        RECT 68.635000 50.495000 68.955000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 34.760000 69.360000 35.080000 ;
      LAYER met4 ;
        RECT 69.040000 34.760000 69.360000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 35.200000 69.360000 35.520000 ;
      LAYER met4 ;
        RECT 69.040000 35.200000 69.360000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 35.640000 69.360000 35.960000 ;
      LAYER met4 ;
        RECT 69.040000 35.640000 69.360000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 36.080000 69.360000 36.400000 ;
      LAYER met4 ;
        RECT 69.040000 36.080000 69.360000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 36.520000 69.360000 36.840000 ;
      LAYER met4 ;
        RECT 69.040000 36.520000 69.360000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 36.960000 69.360000 37.280000 ;
      LAYER met4 ;
        RECT 69.040000 36.960000 69.360000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 37.400000 69.360000 37.720000 ;
      LAYER met4 ;
        RECT 69.040000 37.400000 69.360000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 37.840000 69.360000 38.160000 ;
      LAYER met4 ;
        RECT 69.040000 37.840000 69.360000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 49.655000 69.360000 49.975000 ;
      LAYER met4 ;
        RECT 69.040000 49.655000 69.360000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 50.075000 69.360000 50.395000 ;
      LAYER met4 ;
        RECT 69.040000 50.075000 69.360000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 50.495000 69.360000 50.815000 ;
      LAYER met4 ;
        RECT 69.040000 50.495000 69.360000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 34.760000 69.765000 35.080000 ;
      LAYER met4 ;
        RECT 69.445000 34.760000 69.765000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 35.200000 69.765000 35.520000 ;
      LAYER met4 ;
        RECT 69.445000 35.200000 69.765000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 35.640000 69.765000 35.960000 ;
      LAYER met4 ;
        RECT 69.445000 35.640000 69.765000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 36.080000 69.765000 36.400000 ;
      LAYER met4 ;
        RECT 69.445000 36.080000 69.765000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 36.520000 69.765000 36.840000 ;
      LAYER met4 ;
        RECT 69.445000 36.520000 69.765000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 36.960000 69.765000 37.280000 ;
      LAYER met4 ;
        RECT 69.445000 36.960000 69.765000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 37.400000 69.765000 37.720000 ;
      LAYER met4 ;
        RECT 69.445000 37.400000 69.765000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 37.840000 69.765000 38.160000 ;
      LAYER met4 ;
        RECT 69.445000 37.840000 69.765000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 49.655000 69.765000 49.975000 ;
      LAYER met4 ;
        RECT 69.445000 49.655000 69.765000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 50.075000 69.765000 50.395000 ;
      LAYER met4 ;
        RECT 69.445000 50.075000 69.765000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 50.495000 69.765000 50.815000 ;
      LAYER met4 ;
        RECT 69.445000 50.495000 69.765000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 34.760000 70.170000 35.080000 ;
      LAYER met4 ;
        RECT 69.850000 34.760000 70.170000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 35.200000 70.170000 35.520000 ;
      LAYER met4 ;
        RECT 69.850000 35.200000 70.170000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 35.640000 70.170000 35.960000 ;
      LAYER met4 ;
        RECT 69.850000 35.640000 70.170000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 36.080000 70.170000 36.400000 ;
      LAYER met4 ;
        RECT 69.850000 36.080000 70.170000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 36.520000 70.170000 36.840000 ;
      LAYER met4 ;
        RECT 69.850000 36.520000 70.170000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 36.960000 70.170000 37.280000 ;
      LAYER met4 ;
        RECT 69.850000 36.960000 70.170000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 37.400000 70.170000 37.720000 ;
      LAYER met4 ;
        RECT 69.850000 37.400000 70.170000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 37.840000 70.170000 38.160000 ;
      LAYER met4 ;
        RECT 69.850000 37.840000 70.170000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 49.655000 70.170000 49.975000 ;
      LAYER met4 ;
        RECT 69.850000 49.655000 70.170000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 50.075000 70.170000 50.395000 ;
      LAYER met4 ;
        RECT 69.850000 50.075000 70.170000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 50.495000 70.170000 50.815000 ;
      LAYER met4 ;
        RECT 69.850000 50.495000 70.170000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 34.760000 7.360000 35.080000 ;
      LAYER met4 ;
        RECT 7.040000 34.760000 7.360000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 35.200000 7.360000 35.520000 ;
      LAYER met4 ;
        RECT 7.040000 35.200000 7.360000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 35.640000 7.360000 35.960000 ;
      LAYER met4 ;
        RECT 7.040000 35.640000 7.360000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 36.080000 7.360000 36.400000 ;
      LAYER met4 ;
        RECT 7.040000 36.080000 7.360000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 36.520000 7.360000 36.840000 ;
      LAYER met4 ;
        RECT 7.040000 36.520000 7.360000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 36.960000 7.360000 37.280000 ;
      LAYER met4 ;
        RECT 7.040000 36.960000 7.360000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 37.400000 7.360000 37.720000 ;
      LAYER met4 ;
        RECT 7.040000 37.400000 7.360000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 37.840000 7.360000 38.160000 ;
      LAYER met4 ;
        RECT 7.040000 37.840000 7.360000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 49.655000 7.360000 49.975000 ;
      LAYER met4 ;
        RECT 7.040000 49.655000 7.360000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 50.075000 7.360000 50.395000 ;
      LAYER met4 ;
        RECT 7.040000 50.075000 7.360000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 50.495000 7.360000 50.815000 ;
      LAYER met4 ;
        RECT 7.040000 50.495000 7.360000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 34.760000 7.765000 35.080000 ;
      LAYER met4 ;
        RECT 7.445000 34.760000 7.765000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 35.200000 7.765000 35.520000 ;
      LAYER met4 ;
        RECT 7.445000 35.200000 7.765000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 35.640000 7.765000 35.960000 ;
      LAYER met4 ;
        RECT 7.445000 35.640000 7.765000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 36.080000 7.765000 36.400000 ;
      LAYER met4 ;
        RECT 7.445000 36.080000 7.765000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 36.520000 7.765000 36.840000 ;
      LAYER met4 ;
        RECT 7.445000 36.520000 7.765000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 36.960000 7.765000 37.280000 ;
      LAYER met4 ;
        RECT 7.445000 36.960000 7.765000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 37.400000 7.765000 37.720000 ;
      LAYER met4 ;
        RECT 7.445000 37.400000 7.765000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 37.840000 7.765000 38.160000 ;
      LAYER met4 ;
        RECT 7.445000 37.840000 7.765000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 49.655000 7.765000 49.975000 ;
      LAYER met4 ;
        RECT 7.445000 49.655000 7.765000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 50.075000 7.765000 50.395000 ;
      LAYER met4 ;
        RECT 7.445000 50.075000 7.765000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 50.495000 7.765000 50.815000 ;
      LAYER met4 ;
        RECT 7.445000 50.495000 7.765000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 34.760000 8.170000 35.080000 ;
      LAYER met4 ;
        RECT 7.850000 34.760000 8.170000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 35.200000 8.170000 35.520000 ;
      LAYER met4 ;
        RECT 7.850000 35.200000 8.170000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 35.640000 8.170000 35.960000 ;
      LAYER met4 ;
        RECT 7.850000 35.640000 8.170000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 36.080000 8.170000 36.400000 ;
      LAYER met4 ;
        RECT 7.850000 36.080000 8.170000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 36.520000 8.170000 36.840000 ;
      LAYER met4 ;
        RECT 7.850000 36.520000 8.170000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 36.960000 8.170000 37.280000 ;
      LAYER met4 ;
        RECT 7.850000 36.960000 8.170000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 37.400000 8.170000 37.720000 ;
      LAYER met4 ;
        RECT 7.850000 37.400000 8.170000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 37.840000 8.170000 38.160000 ;
      LAYER met4 ;
        RECT 7.850000 37.840000 8.170000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 49.655000 8.170000 49.975000 ;
      LAYER met4 ;
        RECT 7.850000 49.655000 8.170000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 50.075000 8.170000 50.395000 ;
      LAYER met4 ;
        RECT 7.850000 50.075000 8.170000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 50.495000 8.170000 50.815000 ;
      LAYER met4 ;
        RECT 7.850000 50.495000 8.170000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 34.760000 70.575000 35.080000 ;
      LAYER met4 ;
        RECT 70.255000 34.760000 70.575000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 35.200000 70.575000 35.520000 ;
      LAYER met4 ;
        RECT 70.255000 35.200000 70.575000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 35.640000 70.575000 35.960000 ;
      LAYER met4 ;
        RECT 70.255000 35.640000 70.575000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 36.080000 70.575000 36.400000 ;
      LAYER met4 ;
        RECT 70.255000 36.080000 70.575000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 36.520000 70.575000 36.840000 ;
      LAYER met4 ;
        RECT 70.255000 36.520000 70.575000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 36.960000 70.575000 37.280000 ;
      LAYER met4 ;
        RECT 70.255000 36.960000 70.575000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 37.400000 70.575000 37.720000 ;
      LAYER met4 ;
        RECT 70.255000 37.400000 70.575000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 37.840000 70.575000 38.160000 ;
      LAYER met4 ;
        RECT 70.255000 37.840000 70.575000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 49.655000 70.575000 49.975000 ;
      LAYER met4 ;
        RECT 70.255000 49.655000 70.575000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 50.075000 70.575000 50.395000 ;
      LAYER met4 ;
        RECT 70.255000 50.075000 70.575000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 50.495000 70.575000 50.815000 ;
      LAYER met4 ;
        RECT 70.255000 50.495000 70.575000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 34.760000 70.980000 35.080000 ;
      LAYER met4 ;
        RECT 70.660000 34.760000 70.980000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 35.200000 70.980000 35.520000 ;
      LAYER met4 ;
        RECT 70.660000 35.200000 70.980000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 35.640000 70.980000 35.960000 ;
      LAYER met4 ;
        RECT 70.660000 35.640000 70.980000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 36.080000 70.980000 36.400000 ;
      LAYER met4 ;
        RECT 70.660000 36.080000 70.980000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 36.520000 70.980000 36.840000 ;
      LAYER met4 ;
        RECT 70.660000 36.520000 70.980000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 36.960000 70.980000 37.280000 ;
      LAYER met4 ;
        RECT 70.660000 36.960000 70.980000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 37.400000 70.980000 37.720000 ;
      LAYER met4 ;
        RECT 70.660000 37.400000 70.980000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 37.840000 70.980000 38.160000 ;
      LAYER met4 ;
        RECT 70.660000 37.840000 70.980000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 49.655000 70.980000 49.975000 ;
      LAYER met4 ;
        RECT 70.660000 49.655000 70.980000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 50.075000 70.980000 50.395000 ;
      LAYER met4 ;
        RECT 70.660000 50.075000 70.980000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 50.495000 70.980000 50.815000 ;
      LAYER met4 ;
        RECT 70.660000 50.495000 70.980000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 34.760000 71.385000 35.080000 ;
      LAYER met4 ;
        RECT 71.065000 34.760000 71.385000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 35.200000 71.385000 35.520000 ;
      LAYER met4 ;
        RECT 71.065000 35.200000 71.385000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 35.640000 71.385000 35.960000 ;
      LAYER met4 ;
        RECT 71.065000 35.640000 71.385000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 36.080000 71.385000 36.400000 ;
      LAYER met4 ;
        RECT 71.065000 36.080000 71.385000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 36.520000 71.385000 36.840000 ;
      LAYER met4 ;
        RECT 71.065000 36.520000 71.385000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 36.960000 71.385000 37.280000 ;
      LAYER met4 ;
        RECT 71.065000 36.960000 71.385000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 37.400000 71.385000 37.720000 ;
      LAYER met4 ;
        RECT 71.065000 37.400000 71.385000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 37.840000 71.385000 38.160000 ;
      LAYER met4 ;
        RECT 71.065000 37.840000 71.385000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 49.655000 71.385000 49.975000 ;
      LAYER met4 ;
        RECT 71.065000 49.655000 71.385000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 50.075000 71.385000 50.395000 ;
      LAYER met4 ;
        RECT 71.065000 50.075000 71.385000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 50.495000 71.385000 50.815000 ;
      LAYER met4 ;
        RECT 71.065000 50.495000 71.385000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 34.760000 71.790000 35.080000 ;
      LAYER met4 ;
        RECT 71.470000 34.760000 71.790000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 35.200000 71.790000 35.520000 ;
      LAYER met4 ;
        RECT 71.470000 35.200000 71.790000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 35.640000 71.790000 35.960000 ;
      LAYER met4 ;
        RECT 71.470000 35.640000 71.790000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 36.080000 71.790000 36.400000 ;
      LAYER met4 ;
        RECT 71.470000 36.080000 71.790000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 36.520000 71.790000 36.840000 ;
      LAYER met4 ;
        RECT 71.470000 36.520000 71.790000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 36.960000 71.790000 37.280000 ;
      LAYER met4 ;
        RECT 71.470000 36.960000 71.790000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 37.400000 71.790000 37.720000 ;
      LAYER met4 ;
        RECT 71.470000 37.400000 71.790000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 37.840000 71.790000 38.160000 ;
      LAYER met4 ;
        RECT 71.470000 37.840000 71.790000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 49.655000 71.790000 49.975000 ;
      LAYER met4 ;
        RECT 71.470000 49.655000 71.790000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 50.075000 71.790000 50.395000 ;
      LAYER met4 ;
        RECT 71.470000 50.075000 71.790000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 50.495000 71.790000 50.815000 ;
      LAYER met4 ;
        RECT 71.470000 50.495000 71.790000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 34.760000 72.195000 35.080000 ;
      LAYER met4 ;
        RECT 71.875000 34.760000 72.195000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 35.200000 72.195000 35.520000 ;
      LAYER met4 ;
        RECT 71.875000 35.200000 72.195000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 35.640000 72.195000 35.960000 ;
      LAYER met4 ;
        RECT 71.875000 35.640000 72.195000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 36.080000 72.195000 36.400000 ;
      LAYER met4 ;
        RECT 71.875000 36.080000 72.195000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 36.520000 72.195000 36.840000 ;
      LAYER met4 ;
        RECT 71.875000 36.520000 72.195000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 36.960000 72.195000 37.280000 ;
      LAYER met4 ;
        RECT 71.875000 36.960000 72.195000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 37.400000 72.195000 37.720000 ;
      LAYER met4 ;
        RECT 71.875000 37.400000 72.195000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 37.840000 72.195000 38.160000 ;
      LAYER met4 ;
        RECT 71.875000 37.840000 72.195000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 49.655000 72.195000 49.975000 ;
      LAYER met4 ;
        RECT 71.875000 49.655000 72.195000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 50.075000 72.195000 50.395000 ;
      LAYER met4 ;
        RECT 71.875000 50.075000 72.195000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 50.495000 72.195000 50.815000 ;
      LAYER met4 ;
        RECT 71.875000 50.495000 72.195000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 34.760000 72.600000 35.080000 ;
      LAYER met4 ;
        RECT 72.280000 34.760000 72.600000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 35.200000 72.600000 35.520000 ;
      LAYER met4 ;
        RECT 72.280000 35.200000 72.600000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 35.640000 72.600000 35.960000 ;
      LAYER met4 ;
        RECT 72.280000 35.640000 72.600000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 36.080000 72.600000 36.400000 ;
      LAYER met4 ;
        RECT 72.280000 36.080000 72.600000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 36.520000 72.600000 36.840000 ;
      LAYER met4 ;
        RECT 72.280000 36.520000 72.600000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 36.960000 72.600000 37.280000 ;
      LAYER met4 ;
        RECT 72.280000 36.960000 72.600000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 37.400000 72.600000 37.720000 ;
      LAYER met4 ;
        RECT 72.280000 37.400000 72.600000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 37.840000 72.600000 38.160000 ;
      LAYER met4 ;
        RECT 72.280000 37.840000 72.600000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 49.655000 72.600000 49.975000 ;
      LAYER met4 ;
        RECT 72.280000 49.655000 72.600000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 50.075000 72.600000 50.395000 ;
      LAYER met4 ;
        RECT 72.280000 50.075000 72.600000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 50.495000 72.600000 50.815000 ;
      LAYER met4 ;
        RECT 72.280000 50.495000 72.600000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 34.760000 73.005000 35.080000 ;
      LAYER met4 ;
        RECT 72.685000 34.760000 73.005000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 35.200000 73.005000 35.520000 ;
      LAYER met4 ;
        RECT 72.685000 35.200000 73.005000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 35.640000 73.005000 35.960000 ;
      LAYER met4 ;
        RECT 72.685000 35.640000 73.005000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 36.080000 73.005000 36.400000 ;
      LAYER met4 ;
        RECT 72.685000 36.080000 73.005000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 36.520000 73.005000 36.840000 ;
      LAYER met4 ;
        RECT 72.685000 36.520000 73.005000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 36.960000 73.005000 37.280000 ;
      LAYER met4 ;
        RECT 72.685000 36.960000 73.005000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 37.400000 73.005000 37.720000 ;
      LAYER met4 ;
        RECT 72.685000 37.400000 73.005000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 37.840000 73.005000 38.160000 ;
      LAYER met4 ;
        RECT 72.685000 37.840000 73.005000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 49.655000 73.005000 49.975000 ;
      LAYER met4 ;
        RECT 72.685000 49.655000 73.005000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 50.075000 73.005000 50.395000 ;
      LAYER met4 ;
        RECT 72.685000 50.075000 73.005000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 50.495000 73.005000 50.815000 ;
      LAYER met4 ;
        RECT 72.685000 50.495000 73.005000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 34.760000 73.410000 35.080000 ;
      LAYER met4 ;
        RECT 73.090000 34.760000 73.410000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 35.200000 73.410000 35.520000 ;
      LAYER met4 ;
        RECT 73.090000 35.200000 73.410000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 35.640000 73.410000 35.960000 ;
      LAYER met4 ;
        RECT 73.090000 35.640000 73.410000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 36.080000 73.410000 36.400000 ;
      LAYER met4 ;
        RECT 73.090000 36.080000 73.410000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 36.520000 73.410000 36.840000 ;
      LAYER met4 ;
        RECT 73.090000 36.520000 73.410000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 36.960000 73.410000 37.280000 ;
      LAYER met4 ;
        RECT 73.090000 36.960000 73.410000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 37.400000 73.410000 37.720000 ;
      LAYER met4 ;
        RECT 73.090000 37.400000 73.410000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 37.840000 73.410000 38.160000 ;
      LAYER met4 ;
        RECT 73.090000 37.840000 73.410000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 49.655000 73.410000 49.975000 ;
      LAYER met4 ;
        RECT 73.090000 49.655000 73.410000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 50.075000 73.410000 50.395000 ;
      LAYER met4 ;
        RECT 73.090000 50.075000 73.410000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 50.495000 73.410000 50.815000 ;
      LAYER met4 ;
        RECT 73.090000 50.495000 73.410000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 34.760000 73.815000 35.080000 ;
      LAYER met4 ;
        RECT 73.495000 34.760000 73.815000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 35.200000 73.815000 35.520000 ;
      LAYER met4 ;
        RECT 73.495000 35.200000 73.815000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 35.640000 73.815000 35.960000 ;
      LAYER met4 ;
        RECT 73.495000 35.640000 73.815000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 36.080000 73.815000 36.400000 ;
      LAYER met4 ;
        RECT 73.495000 36.080000 73.815000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 36.520000 73.815000 36.840000 ;
      LAYER met4 ;
        RECT 73.495000 36.520000 73.815000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 36.960000 73.815000 37.280000 ;
      LAYER met4 ;
        RECT 73.495000 36.960000 73.815000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 37.400000 73.815000 37.720000 ;
      LAYER met4 ;
        RECT 73.495000 37.400000 73.815000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 37.840000 73.815000 38.160000 ;
      LAYER met4 ;
        RECT 73.495000 37.840000 73.815000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 49.655000 73.815000 49.975000 ;
      LAYER met4 ;
        RECT 73.495000 49.655000 73.815000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 50.075000 73.815000 50.395000 ;
      LAYER met4 ;
        RECT 73.495000 50.075000 73.815000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 50.495000 73.815000 50.815000 ;
      LAYER met4 ;
        RECT 73.495000 50.495000 73.815000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 34.760000 74.220000 35.080000 ;
      LAYER met4 ;
        RECT 73.900000 34.760000 74.220000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 35.200000 74.220000 35.520000 ;
      LAYER met4 ;
        RECT 73.900000 35.200000 74.220000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 35.640000 74.220000 35.960000 ;
      LAYER met4 ;
        RECT 73.900000 35.640000 74.220000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 36.080000 74.220000 36.400000 ;
      LAYER met4 ;
        RECT 73.900000 36.080000 74.220000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 36.520000 74.220000 36.840000 ;
      LAYER met4 ;
        RECT 73.900000 36.520000 74.220000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 36.960000 74.220000 37.280000 ;
      LAYER met4 ;
        RECT 73.900000 36.960000 74.220000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 37.400000 74.220000 37.720000 ;
      LAYER met4 ;
        RECT 73.900000 37.400000 74.220000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 37.840000 74.220000 38.160000 ;
      LAYER met4 ;
        RECT 73.900000 37.840000 74.220000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 49.655000 74.220000 49.975000 ;
      LAYER met4 ;
        RECT 73.900000 49.655000 74.220000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 50.075000 74.220000 50.395000 ;
      LAYER met4 ;
        RECT 73.900000 50.075000 74.220000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 50.495000 74.220000 50.815000 ;
      LAYER met4 ;
        RECT 73.900000 50.495000 74.220000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 34.760000 74.625000 35.080000 ;
      LAYER met4 ;
        RECT 74.305000 34.760000 74.625000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 35.200000 74.625000 35.520000 ;
      LAYER met4 ;
        RECT 74.305000 35.200000 74.625000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 35.640000 74.625000 35.960000 ;
      LAYER met4 ;
        RECT 74.305000 35.640000 74.625000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 36.080000 74.625000 36.400000 ;
      LAYER met4 ;
        RECT 74.305000 36.080000 74.625000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 36.520000 74.625000 36.840000 ;
      LAYER met4 ;
        RECT 74.305000 36.520000 74.625000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 36.960000 74.625000 37.280000 ;
      LAYER met4 ;
        RECT 74.305000 36.960000 74.625000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 37.400000 74.625000 37.720000 ;
      LAYER met4 ;
        RECT 74.305000 37.400000 74.625000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 37.840000 74.625000 38.160000 ;
      LAYER met4 ;
        RECT 74.305000 37.840000 74.625000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 49.655000 74.625000 49.975000 ;
      LAYER met4 ;
        RECT 74.305000 49.655000 74.625000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 50.075000 74.625000 50.395000 ;
      LAYER met4 ;
        RECT 74.305000 50.075000 74.625000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 50.495000 74.625000 50.815000 ;
      LAYER met4 ;
        RECT 74.305000 50.495000 74.625000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 34.760000 8.575000 35.080000 ;
      LAYER met4 ;
        RECT 8.255000 34.760000 8.575000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 35.200000 8.575000 35.520000 ;
      LAYER met4 ;
        RECT 8.255000 35.200000 8.575000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 35.640000 8.575000 35.960000 ;
      LAYER met4 ;
        RECT 8.255000 35.640000 8.575000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 36.080000 8.575000 36.400000 ;
      LAYER met4 ;
        RECT 8.255000 36.080000 8.575000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 36.520000 8.575000 36.840000 ;
      LAYER met4 ;
        RECT 8.255000 36.520000 8.575000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 36.960000 8.575000 37.280000 ;
      LAYER met4 ;
        RECT 8.255000 36.960000 8.575000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 37.400000 8.575000 37.720000 ;
      LAYER met4 ;
        RECT 8.255000 37.400000 8.575000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 37.840000 8.575000 38.160000 ;
      LAYER met4 ;
        RECT 8.255000 37.840000 8.575000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 49.655000 8.575000 49.975000 ;
      LAYER met4 ;
        RECT 8.255000 49.655000 8.575000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 50.075000 8.575000 50.395000 ;
      LAYER met4 ;
        RECT 8.255000 50.075000 8.575000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 50.495000 8.575000 50.815000 ;
      LAYER met4 ;
        RECT 8.255000 50.495000 8.575000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 34.760000 8.980000 35.080000 ;
      LAYER met4 ;
        RECT 8.660000 34.760000 8.980000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 35.200000 8.980000 35.520000 ;
      LAYER met4 ;
        RECT 8.660000 35.200000 8.980000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 35.640000 8.980000 35.960000 ;
      LAYER met4 ;
        RECT 8.660000 35.640000 8.980000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 36.080000 8.980000 36.400000 ;
      LAYER met4 ;
        RECT 8.660000 36.080000 8.980000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 36.520000 8.980000 36.840000 ;
      LAYER met4 ;
        RECT 8.660000 36.520000 8.980000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 36.960000 8.980000 37.280000 ;
      LAYER met4 ;
        RECT 8.660000 36.960000 8.980000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 37.400000 8.980000 37.720000 ;
      LAYER met4 ;
        RECT 8.660000 37.400000 8.980000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 37.840000 8.980000 38.160000 ;
      LAYER met4 ;
        RECT 8.660000 37.840000 8.980000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 49.655000 8.980000 49.975000 ;
      LAYER met4 ;
        RECT 8.660000 49.655000 8.980000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 50.075000 8.980000 50.395000 ;
      LAYER met4 ;
        RECT 8.660000 50.075000 8.980000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 50.495000 8.980000 50.815000 ;
      LAYER met4 ;
        RECT 8.660000 50.495000 8.980000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 34.760000 9.385000 35.080000 ;
      LAYER met4 ;
        RECT 9.065000 34.760000 9.385000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 35.200000 9.385000 35.520000 ;
      LAYER met4 ;
        RECT 9.065000 35.200000 9.385000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 35.640000 9.385000 35.960000 ;
      LAYER met4 ;
        RECT 9.065000 35.640000 9.385000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 36.080000 9.385000 36.400000 ;
      LAYER met4 ;
        RECT 9.065000 36.080000 9.385000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 36.520000 9.385000 36.840000 ;
      LAYER met4 ;
        RECT 9.065000 36.520000 9.385000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 36.960000 9.385000 37.280000 ;
      LAYER met4 ;
        RECT 9.065000 36.960000 9.385000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 37.400000 9.385000 37.720000 ;
      LAYER met4 ;
        RECT 9.065000 37.400000 9.385000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 37.840000 9.385000 38.160000 ;
      LAYER met4 ;
        RECT 9.065000 37.840000 9.385000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 49.655000 9.385000 49.975000 ;
      LAYER met4 ;
        RECT 9.065000 49.655000 9.385000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 50.075000 9.385000 50.395000 ;
      LAYER met4 ;
        RECT 9.065000 50.075000 9.385000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 50.495000 9.385000 50.815000 ;
      LAYER met4 ;
        RECT 9.065000 50.495000 9.385000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 34.760000 9.790000 35.080000 ;
      LAYER met4 ;
        RECT 9.470000 34.760000 9.790000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 35.200000 9.790000 35.520000 ;
      LAYER met4 ;
        RECT 9.470000 35.200000 9.790000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 35.640000 9.790000 35.960000 ;
      LAYER met4 ;
        RECT 9.470000 35.640000 9.790000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 36.080000 9.790000 36.400000 ;
      LAYER met4 ;
        RECT 9.470000 36.080000 9.790000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 36.520000 9.790000 36.840000 ;
      LAYER met4 ;
        RECT 9.470000 36.520000 9.790000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 36.960000 9.790000 37.280000 ;
      LAYER met4 ;
        RECT 9.470000 36.960000 9.790000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 37.400000 9.790000 37.720000 ;
      LAYER met4 ;
        RECT 9.470000 37.400000 9.790000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 37.840000 9.790000 38.160000 ;
      LAYER met4 ;
        RECT 9.470000 37.840000 9.790000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 49.655000 9.790000 49.975000 ;
      LAYER met4 ;
        RECT 9.470000 49.655000 9.790000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 50.075000 9.790000 50.395000 ;
      LAYER met4 ;
        RECT 9.470000 50.075000 9.790000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 50.495000 9.790000 50.815000 ;
      LAYER met4 ;
        RECT 9.470000 50.495000 9.790000 50.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 34.760000 10.195000 35.080000 ;
      LAYER met4 ;
        RECT 9.875000 34.760000 10.195000 35.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 35.200000 10.195000 35.520000 ;
      LAYER met4 ;
        RECT 9.875000 35.200000 10.195000 35.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 35.640000 10.195000 35.960000 ;
      LAYER met4 ;
        RECT 9.875000 35.640000 10.195000 35.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 36.080000 10.195000 36.400000 ;
      LAYER met4 ;
        RECT 9.875000 36.080000 10.195000 36.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 36.520000 10.195000 36.840000 ;
      LAYER met4 ;
        RECT 9.875000 36.520000 10.195000 36.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 36.960000 10.195000 37.280000 ;
      LAYER met4 ;
        RECT 9.875000 36.960000 10.195000 37.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 37.400000 10.195000 37.720000 ;
      LAYER met4 ;
        RECT 9.875000 37.400000 10.195000 37.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 37.840000 10.195000 38.160000 ;
      LAYER met4 ;
        RECT 9.875000 37.840000 10.195000 38.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 49.655000 10.195000 49.975000 ;
      LAYER met4 ;
        RECT 9.875000 49.655000 10.195000 49.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 50.075000 10.195000 50.395000 ;
      LAYER met4 ;
        RECT 9.875000 50.075000 10.195000 50.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 50.495000 10.195000 50.815000 ;
      LAYER met4 ;
        RECT 9.875000 50.495000 10.195000 50.815000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met3 ;
      RECT 0.500000 34.740000 74.655000 50.820000 ;
    LAYER met4 ;
      RECT 0.000000  0.035000 75.000000  45.965000 ;
      RECT 0.000000 49.745000 75.000000  50.725000 ;
      RECT 0.000000 54.505000 75.000000 198.000000 ;
    LAYER met5 ;
      RECT 0.000000  0.135000 72.130000  13.035000 ;
      RECT 0.000000 13.035000 72.435000  17.885000 ;
      RECT 0.000000 17.885000 75.000000  22.335000 ;
      RECT 0.000000 22.335000 72.130000  34.835000 ;
      RECT 0.000000 34.835000 75.000000  38.085000 ;
      RECT 0.000000 38.085000 72.130000  45.735000 ;
      RECT 0.000000 45.735000 75.000000  54.735000 ;
      RECT 0.000000 54.735000 72.130000  94.585000 ;
      RECT 0.000000 94.585000 75.000000 198.000000 ;
  END
END sky130_fd_io__overlay_vssa_lvc
END LIBRARY
