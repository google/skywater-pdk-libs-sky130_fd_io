# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sky130_fd_io__top_lvclamp
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 47.895 BY 198 ;
  SYMMETRY X Y R90 ;

  PIN ogc_lvc
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 41.84 48.76 42.865 48.83 ;
        RECT 41.91 48.83 42.865 48.9 ;
        RECT 41.98 48.9 42.865 48.97 ;
        RECT 42.05 48.97 42.865 49.04 ;
        RECT 42.115 49.04 42.865 49.105 ;
        RECT 38.54 17.295 39.385 17.365 ;
        RECT 38.61 17.365 39.385 17.435 ;
        RECT 38.635 17.435 39.385 17.46 ;
        RECT 38.635 16.575 39.385 16.64 ;
        RECT 38.57 16.64 39.385 16.705 ;
        RECT 9.69 48.76 10.475 48.83 ;
        RECT 9.69 48.83 10.405 48.9 ;
        RECT 9.69 48.9 10.335 48.97 ;
        RECT 9.69 48.97 10.28 49.025 ;
        RECT 9.69 47.435 10.28 47.505 ;
        RECT 9.69 47.505 10.35 47.575 ;
        RECT 9.69 47.575 10.42 47.645 ;
        RECT 9.69 47.645 10.49 47.7 ;
        RECT 9.69 17.295 10.345 17.355 ;
        RECT 9.69 17.355 10.285 17.415 ;
        RECT 9.69 17.415 10.28 17.42 ;
        RECT 42.115 196.58 42.865 196.65 ;
        RECT 42.045 196.65 42.865 196.72 ;
        RECT 41.975 196.72 42.865 196.79 ;
        RECT 41.905 196.79 42.865 196.82 ;
        RECT 42.115 49.105 42.865 196.58 ;
        RECT 9.69 196.65 10.28 196.72 ;
        RECT 9.69 196.72 10.35 196.79 ;
        RECT 9.69 196.79 10.42 196.82 ;
        RECT 38.635 17.46 39.385 47.53 ;
        RECT 38.635 0 39.385 16.575 ;
        RECT 38.635 47.535 39.39 47.605 ;
        RECT 38.565 47.605 39.46 47.675 ;
        RECT 38.495 47.675 39.53 47.7 ;
        RECT 38.635 47.53 39.385 47.535 ;
        RECT 9.69 196.82 42.865 197.41 ;
        RECT 9.69 17.42 10.28 47.435 ;
        RECT 9.69 49.025 10.28 196.65 ;
        RECT 9.69 16.705 39.385 17.295 ;
        RECT 9.69 47.7 42.865 48.76 ;
    END
  END ogc_lvc

  PIN src_bdy_lvc
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 28.04 0 41.09 193.675 ;
    END
  END src_bdy_lvc

  PIN drn_lvc
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 13.62 0 26.54 189.96 ;
    END
  END drn_lvc
  OBS
    LAYER li1 ;
      RECT 9.985 8.035 16.945 8.205 ;
      RECT 17.635 7.575 24.595 7.745 ;
      RECT 9.985 7.575 16.945 7.745 ;
      RECT 17.635 9.415 24.595 9.585 ;
      RECT 9.985 9.415 16.945 9.585 ;
      RECT 17.635 8.955 24.425 9.125 ;
      RECT 9.985 8.955 16.945 9.125 ;
      RECT 13.2 28.055 35.24 28.225 ;
      RECT 15.115 58.92 38.635 59.09 ;
      RECT 15.115 50.11 38.645 50.28 ;
      RECT 15.175 50.08 38.585 50.11 ;
      RECT 12.34 46.53 36.9 46.7 ;
      RECT 12.4 46.7 36.84 46.705 ;
      RECT 12.34 37.53 36.9 37.7 ;
      RECT 15.115 69.11 38.635 69.28 ;
      RECT 26.195 95.425 38.645 95.595 ;
      RECT 26.195 86.055 38.645 86.225 ;
      RECT 15.115 77.76 38.645 77.93 ;
      RECT 26.195 125.39 38.645 125.56 ;
      RECT 26.195 115.45 38.645 115.62 ;
      RECT 26.195 105.245 38.645 105.415 ;
      RECT 26.195 135.355 38.645 135.525 ;
      RECT 15.115 155.215 38.645 155.385 ;
      RECT 15.115 146.08 38.645 146.25 ;
      RECT 15.115 194.1 38.645 194.27 ;
      RECT 15.115 185.155 38.645 185.325 ;
      RECT 15.115 175.325 38.645 175.495 ;
      RECT 15.115 165.33 38.645 165.5 ;
      RECT 26.615 146.9 27.145 153.57 ;
      RECT 26.625 153.57 27.135 153.63 ;
      RECT 26.625 146.84 27.135 146.9 ;
      RECT 33.36 146.84 34.25 153.63 ;
      RECT 30.59 146.84 31.48 153.63 ;
      RECT 33.36 156.84 34.25 163.63 ;
      RECT 30.59 156.84 31.48 163.63 ;
      RECT 33.36 166.84 34.25 173.63 ;
      RECT 30.59 166.84 31.48 173.63 ;
      RECT 32.155 156.9 32.685 163.57 ;
      RECT 32.165 163.57 32.675 163.63 ;
      RECT 32.165 156.84 32.675 156.9 ;
      RECT 32.155 166.9 32.685 173.57 ;
      RECT 32.165 173.57 32.675 173.63 ;
      RECT 32.165 166.84 32.675 166.9 ;
      RECT 32.155 146.9 32.685 153.57 ;
      RECT 32.165 153.57 32.675 153.63 ;
      RECT 32.165 146.84 32.675 146.9 ;
      RECT 36.13 146.84 37.02 153.63 ;
      RECT 36.13 156.84 37.02 163.63 ;
      RECT 36.13 166.84 37.02 173.63 ;
      RECT 37.695 146.84 38.225 153.63 ;
      RECT 37.695 156.84 38.225 163.63 ;
      RECT 37.695 166.84 38.225 173.63 ;
      RECT 34.925 146.9 35.455 153.57 ;
      RECT 34.935 153.57 35.445 153.63 ;
      RECT 34.935 146.84 35.445 146.9 ;
      RECT 34.925 156.9 35.455 163.57 ;
      RECT 34.935 163.57 35.445 163.63 ;
      RECT 34.935 156.84 35.445 156.9 ;
      RECT 34.925 166.9 35.455 173.57 ;
      RECT 34.935 173.57 35.445 173.63 ;
      RECT 34.935 166.84 35.445 166.9 ;
      RECT 38.9 146.84 39.79 153.63 ;
      RECT 38.9 156.84 39.79 163.63 ;
      RECT 38.9 166.84 39.79 173.63 ;
      RECT 16.74 186.84 17.63 193.63 ;
      RECT 13.97 186.84 14.86 193.63 ;
      RECT 16.74 176.84 17.63 183.63 ;
      RECT 13.97 176.84 14.86 183.63 ;
      RECT 15.535 176.9 16.065 183.57 ;
      RECT 15.545 183.57 16.055 183.63 ;
      RECT 15.545 176.84 16.055 176.9 ;
      RECT 15.535 186.9 16.065 193.57 ;
      RECT 15.545 193.57 16.055 193.63 ;
      RECT 15.545 186.84 16.055 186.9 ;
      RECT 19.51 186.84 20.4 193.63 ;
      RECT 19.51 176.84 20.4 183.63 ;
      RECT 18.305 176.9 18.835 183.57 ;
      RECT 18.315 183.57 18.825 183.63 ;
      RECT 18.315 176.84 18.825 176.9 ;
      RECT 21.075 176.9 21.605 183.57 ;
      RECT 21.085 183.57 21.595 183.63 ;
      RECT 21.085 176.84 21.595 176.9 ;
      RECT 21.075 186.9 21.605 193.57 ;
      RECT 21.085 193.57 21.595 193.63 ;
      RECT 21.085 186.84 21.595 186.9 ;
      RECT 18.305 186.9 18.835 193.57 ;
      RECT 18.315 193.57 18.825 193.63 ;
      RECT 18.315 186.84 18.825 186.9 ;
      RECT 25.05 186.84 25.94 193.63 ;
      RECT 22.28 186.84 23.17 193.63 ;
      RECT 25.05 176.84 25.94 183.63 ;
      RECT 22.28 176.84 23.17 183.63 ;
      RECT 23.845 186.9 24.375 193.57 ;
      RECT 23.855 193.57 24.365 193.63 ;
      RECT 23.855 186.84 24.365 186.9 ;
      RECT 23.845 176.9 24.375 183.57 ;
      RECT 23.855 183.57 24.365 183.63 ;
      RECT 23.855 176.84 24.365 176.9 ;
      RECT 27.82 186.84 28.71 193.63 ;
      RECT 27.82 176.84 28.71 183.63 ;
      RECT 29.385 186.9 29.915 193.57 ;
      RECT 29.395 193.57 29.905 193.63 ;
      RECT 29.395 186.84 29.905 186.9 ;
      RECT 26.615 186.9 27.145 193.57 ;
      RECT 26.625 193.57 27.135 193.63 ;
      RECT 26.625 186.84 27.135 186.9 ;
      RECT 26.615 176.9 27.145 183.57 ;
      RECT 26.625 183.57 27.135 183.63 ;
      RECT 26.625 176.84 27.135 176.9 ;
      RECT 29.385 176.9 29.915 183.57 ;
      RECT 29.395 183.57 29.905 183.63 ;
      RECT 29.395 176.84 29.905 176.9 ;
      RECT 30.59 186.84 31.48 193.63 ;
      RECT 33.36 176.84 34.25 183.63 ;
      RECT 30.59 176.84 31.48 183.63 ;
      RECT 33.36 186.84 34.25 193.63 ;
      RECT 32.155 186.9 32.685 193.57 ;
      RECT 32.505 193.57 32.675 193.63 ;
      RECT 32.505 186.84 32.675 186.9 ;
      RECT 32.165 193.57 32.335 193.63 ;
      RECT 32.165 186.84 32.335 186.9 ;
      RECT 32.155 176.9 32.685 183.57 ;
      RECT 32.505 183.57 32.675 183.63 ;
      RECT 32.505 176.84 32.675 176.9 ;
      RECT 32.165 183.57 32.335 183.63 ;
      RECT 32.165 176.84 32.335 176.9 ;
      RECT 36.13 176.84 37.02 183.63 ;
      RECT 36.13 186.84 37.02 193.63 ;
      RECT 37.695 176.84 38.225 183.63 ;
      RECT 37.695 186.84 38.225 193.63 ;
      RECT 34.925 176.9 35.455 183.57 ;
      RECT 34.935 183.57 35.445 183.63 ;
      RECT 34.935 176.84 35.445 176.9 ;
      RECT 34.925 186.9 35.455 193.57 ;
      RECT 34.935 193.57 35.445 193.63 ;
      RECT 34.935 186.84 35.445 186.9 ;
      RECT 38.9 176.84 39.79 183.63 ;
      RECT 38.9 186.84 39.79 193.63 ;
      RECT 26.7 1.76 37.97 11.975 ;
      RECT 9.155 11.975 39.52 15.635 ;
      RECT 17.635 5.735 24.595 5.905 ;
      RECT 9.985 5.735 16.945 5.905 ;
      RECT 17.635 5.275 24.425 5.445 ;
      RECT 9.985 5.275 16.945 5.445 ;
      RECT 17.635 4.815 24.595 4.985 ;
      RECT 9.985 4.815 16.945 4.985 ;
      RECT 17.635 7.115 24.425 7.285 ;
      RECT 9.985 7.115 16.945 7.285 ;
      RECT 17.635 6.655 24.595 6.825 ;
      RECT 9.985 6.655 16.945 6.825 ;
      RECT 17.635 6.195 24.425 6.365 ;
      RECT 9.985 6.195 16.945 6.365 ;
      RECT 17.635 8.495 24.595 8.665 ;
      RECT 9.985 8.495 16.945 8.665 ;
      RECT 17.635 8.035 24.425 8.205 ;
      RECT 32.165 103.57 32.675 103.63 ;
      RECT 32.165 96.84 32.675 96.9 ;
      RECT 36.13 116.84 37.02 123.63 ;
      RECT 36.13 106.84 37.02 113.63 ;
      RECT 36.13 96.84 37.02 103.63 ;
      RECT 34.925 96.9 35.455 103.57 ;
      RECT 34.935 103.57 35.445 103.63 ;
      RECT 34.935 96.84 35.445 96.9 ;
      RECT 34.925 106.9 35.455 113.57 ;
      RECT 34.935 113.57 35.445 113.63 ;
      RECT 34.935 106.84 35.445 106.9 ;
      RECT 34.925 116.9 35.455 123.57 ;
      RECT 34.935 123.57 35.445 123.63 ;
      RECT 34.935 116.84 35.445 116.9 ;
      RECT 37.695 96.84 38.225 103.63 ;
      RECT 37.695 106.84 38.225 113.63 ;
      RECT 37.695 116.84 38.225 123.63 ;
      RECT 38.9 116.84 39.79 123.63 ;
      RECT 38.9 106.84 39.79 113.63 ;
      RECT 38.9 96.84 39.79 103.63 ;
      RECT 25.05 126.84 25.94 133.63 ;
      RECT 25.05 136.84 25.94 143.63 ;
      RECT 27.82 126.84 28.71 133.63 ;
      RECT 27.82 136.84 28.71 143.63 ;
      RECT 26.615 126.9 27.145 133.57 ;
      RECT 26.625 133.57 27.135 133.63 ;
      RECT 26.625 126.84 27.135 126.9 ;
      RECT 29.385 126.9 29.915 133.57 ;
      RECT 29.395 133.57 29.905 133.63 ;
      RECT 29.395 126.84 29.905 126.9 ;
      RECT 26.615 136.9 27.145 143.57 ;
      RECT 26.625 143.57 27.135 143.63 ;
      RECT 26.625 136.84 27.135 136.9 ;
      RECT 29.385 136.9 29.915 143.57 ;
      RECT 29.395 143.57 29.905 143.63 ;
      RECT 29.395 136.84 29.905 136.9 ;
      RECT 33.36 126.84 34.25 133.63 ;
      RECT 30.59 126.84 31.48 133.63 ;
      RECT 33.36 136.84 34.25 143.63 ;
      RECT 30.59 136.84 31.48 143.63 ;
      RECT 32.155 126.9 32.685 133.57 ;
      RECT 32.165 133.57 32.675 133.63 ;
      RECT 32.165 126.84 32.675 126.9 ;
      RECT 32.155 136.9 32.685 143.57 ;
      RECT 32.165 143.57 32.675 143.63 ;
      RECT 32.165 136.84 32.675 136.9 ;
      RECT 36.13 126.84 37.02 133.63 ;
      RECT 36.13 136.84 37.02 143.63 ;
      RECT 37.695 126.84 38.225 133.63 ;
      RECT 37.695 136.84 38.225 143.63 ;
      RECT 34.925 126.9 35.455 133.57 ;
      RECT 34.935 133.57 35.445 133.63 ;
      RECT 34.935 126.84 35.445 126.9 ;
      RECT 34.925 136.9 35.455 143.57 ;
      RECT 34.935 143.57 35.445 143.63 ;
      RECT 34.935 136.84 35.445 136.9 ;
      RECT 38.9 126.84 39.79 133.63 ;
      RECT 38.9 136.84 39.79 143.63 ;
      RECT 16.74 146.84 17.63 153.63 ;
      RECT 13.97 146.84 14.86 153.63 ;
      RECT 16.74 156.84 17.63 163.63 ;
      RECT 13.97 156.84 14.86 163.63 ;
      RECT 16.74 166.84 17.63 173.63 ;
      RECT 13.97 166.84 14.86 173.63 ;
      RECT 15.535 156.9 16.065 163.57 ;
      RECT 15.545 163.57 16.055 163.63 ;
      RECT 15.545 156.84 16.055 156.9 ;
      RECT 15.535 166.9 16.065 173.57 ;
      RECT 15.545 173.57 16.055 173.63 ;
      RECT 15.545 166.84 16.055 166.9 ;
      RECT 15.535 146.9 16.065 153.57 ;
      RECT 15.545 153.57 16.055 153.63 ;
      RECT 15.545 146.84 16.055 146.9 ;
      RECT 19.51 146.84 20.4 153.63 ;
      RECT 19.51 156.84 20.4 163.63 ;
      RECT 19.51 166.84 20.4 173.63 ;
      RECT 18.305 156.9 18.835 163.57 ;
      RECT 18.315 163.57 18.825 163.63 ;
      RECT 18.315 156.84 18.825 156.9 ;
      RECT 18.305 166.9 18.835 173.57 ;
      RECT 18.315 173.57 18.825 173.63 ;
      RECT 18.315 166.84 18.825 166.9 ;
      RECT 21.075 166.9 21.605 173.57 ;
      RECT 21.085 173.57 21.595 173.63 ;
      RECT 21.085 166.84 21.595 166.9 ;
      RECT 21.075 156.9 21.605 163.57 ;
      RECT 21.085 163.57 21.595 163.63 ;
      RECT 21.085 156.84 21.595 156.9 ;
      RECT 21.075 146.9 21.605 153.57 ;
      RECT 21.085 153.57 21.595 153.63 ;
      RECT 21.085 146.84 21.595 146.9 ;
      RECT 18.305 146.9 18.835 153.57 ;
      RECT 18.315 153.57 18.825 153.63 ;
      RECT 18.315 146.84 18.825 146.9 ;
      RECT 25.05 146.84 25.94 153.63 ;
      RECT 22.28 146.84 23.17 153.63 ;
      RECT 25.05 156.84 25.94 163.63 ;
      RECT 22.28 156.84 23.17 163.63 ;
      RECT 25.05 166.84 25.94 173.63 ;
      RECT 22.28 166.84 23.17 173.63 ;
      RECT 23.845 166.9 24.375 173.57 ;
      RECT 23.855 173.57 24.365 173.63 ;
      RECT 23.855 166.84 24.365 166.9 ;
      RECT 23.845 156.9 24.375 163.57 ;
      RECT 23.855 163.57 24.365 163.63 ;
      RECT 23.855 156.84 24.365 156.9 ;
      RECT 23.845 146.9 24.375 153.57 ;
      RECT 23.855 153.57 24.365 153.63 ;
      RECT 23.855 146.84 24.365 146.9 ;
      RECT 27.82 146.84 28.71 153.63 ;
      RECT 27.82 156.84 28.71 163.63 ;
      RECT 27.82 166.84 28.71 173.63 ;
      RECT 26.615 156.9 27.145 163.57 ;
      RECT 26.625 163.57 27.135 163.63 ;
      RECT 26.625 156.84 27.135 156.9 ;
      RECT 26.615 166.9 27.145 173.57 ;
      RECT 26.625 173.57 27.135 173.63 ;
      RECT 26.625 166.84 27.135 166.9 ;
      RECT 29.385 156.9 29.915 163.57 ;
      RECT 29.395 163.57 29.905 163.63 ;
      RECT 29.395 156.84 29.905 156.9 ;
      RECT 29.385 166.9 29.915 173.57 ;
      RECT 29.395 173.57 29.905 173.63 ;
      RECT 29.395 166.84 29.905 166.9 ;
      RECT 29.385 146.9 29.915 153.57 ;
      RECT 29.395 153.57 29.905 153.63 ;
      RECT 29.395 146.84 29.905 146.9 ;
      RECT 27.82 60.5 28.71 67.29 ;
      RECT 27.82 50.5 28.71 57.29 ;
      RECT 29.385 50.56 29.915 57.23 ;
      RECT 29.395 57.23 29.905 57.29 ;
      RECT 29.395 50.5 29.905 50.56 ;
      RECT 26.615 60.56 27.145 67.23 ;
      RECT 26.625 67.23 27.135 67.29 ;
      RECT 26.625 60.5 27.135 60.56 ;
      RECT 26.615 50.56 27.145 57.23 ;
      RECT 26.625 57.23 27.135 57.29 ;
      RECT 26.625 50.5 27.135 50.56 ;
      RECT 29.385 60.56 29.915 67.23 ;
      RECT 29.395 67.23 29.905 67.29 ;
      RECT 29.395 60.5 29.905 60.56 ;
      RECT 33.36 60.5 34.25 67.29 ;
      RECT 30.59 60.5 31.48 67.29 ;
      RECT 33.36 50.5 34.25 57.29 ;
      RECT 30.59 50.5 31.48 57.29 ;
      RECT 32.155 60.56 32.685 67.23 ;
      RECT 32.165 67.23 32.675 67.29 ;
      RECT 32.165 60.5 32.675 60.56 ;
      RECT 32.155 50.56 32.685 57.23 ;
      RECT 32.165 57.23 32.675 57.29 ;
      RECT 32.165 50.5 32.675 50.56 ;
      RECT 36.13 60.5 37.02 67.29 ;
      RECT 36.13 50.5 37.02 57.29 ;
      RECT 34.925 50.56 35.455 57.23 ;
      RECT 34.935 57.23 35.445 57.29 ;
      RECT 34.935 50.5 35.445 50.56 ;
      RECT 34.925 60.56 35.455 67.23 ;
      RECT 34.935 67.23 35.445 67.29 ;
      RECT 34.935 60.5 35.445 60.56 ;
      RECT 37.695 50.5 38.225 57.29 ;
      RECT 37.695 60.5 38.225 67.29 ;
      RECT 38.9 60.5 39.79 67.29 ;
      RECT 38.9 50.5 39.79 57.29 ;
      RECT 16.74 70.5 17.63 77.29 ;
      RECT 13.97 70.5 14.86 77.29 ;
      RECT 15.535 70.56 16.065 77.23 ;
      RECT 15.545 77.23 16.055 77.29 ;
      RECT 15.545 70.5 16.055 70.56 ;
      RECT 19.51 70.5 20.4 77.29 ;
      RECT 21.075 70.56 21.605 77.23 ;
      RECT 21.085 77.23 21.595 77.29 ;
      RECT 21.085 70.5 21.595 70.56 ;
      RECT 18.305 70.56 18.835 77.23 ;
      RECT 18.315 77.23 18.825 77.29 ;
      RECT 18.315 70.5 18.825 70.56 ;
      RECT 25.05 70.5 25.94 77.29 ;
      RECT 22.28 70.5 23.17 77.29 ;
      RECT 25.05 86.84 25.94 93.63 ;
      RECT 23.845 70.56 24.375 77.23 ;
      RECT 23.855 77.23 24.365 77.29 ;
      RECT 23.855 70.5 24.365 70.56 ;
      RECT 27.82 70.5 28.71 77.29 ;
      RECT 27.82 86.84 28.71 93.63 ;
      RECT 26.615 70.56 27.145 77.23 ;
      RECT 26.625 77.23 27.135 77.29 ;
      RECT 26.625 70.5 27.135 70.56 ;
      RECT 26.615 86.9 27.145 93.57 ;
      RECT 26.625 93.57 27.135 93.63 ;
      RECT 26.625 86.84 27.135 86.9 ;
      RECT 29.385 86.9 29.915 93.57 ;
      RECT 29.395 93.57 29.905 93.63 ;
      RECT 29.395 86.84 29.905 86.9 ;
      RECT 29.385 70.56 29.915 77.23 ;
      RECT 29.395 77.23 29.905 77.29 ;
      RECT 29.395 70.5 29.905 70.56 ;
      RECT 33.36 70.5 34.25 77.29 ;
      RECT 30.59 70.5 31.48 77.29 ;
      RECT 33.36 86.84 34.25 93.63 ;
      RECT 30.59 86.84 31.48 93.63 ;
      RECT 32.155 86.9 32.685 93.57 ;
      RECT 32.165 93.57 32.675 93.63 ;
      RECT 32.165 86.84 32.675 86.9 ;
      RECT 32.155 70.56 32.685 77.23 ;
      RECT 32.165 77.23 32.675 77.29 ;
      RECT 32.165 70.5 32.675 70.56 ;
      RECT 36.13 70.5 37.02 77.29 ;
      RECT 36.13 86.84 37.02 93.63 ;
      RECT 34.925 70.56 35.455 77.23 ;
      RECT 34.935 77.23 35.445 77.29 ;
      RECT 34.935 70.5 35.445 70.56 ;
      RECT 34.925 86.9 35.455 93.57 ;
      RECT 34.935 93.57 35.445 93.63 ;
      RECT 34.935 86.84 35.445 86.9 ;
      RECT 37.695 70.5 38.225 77.29 ;
      RECT 37.695 86.84 38.225 93.63 ;
      RECT 38.9 70.5 39.79 77.29 ;
      RECT 38.9 86.84 39.79 93.63 ;
      RECT 25.05 116.84 25.94 123.63 ;
      RECT 25.05 106.84 25.94 113.63 ;
      RECT 25.05 96.84 25.94 103.63 ;
      RECT 27.82 116.84 28.71 123.63 ;
      RECT 27.82 106.84 28.71 113.63 ;
      RECT 27.82 96.84 28.71 103.63 ;
      RECT 26.615 116.9 27.145 123.57 ;
      RECT 26.625 123.57 27.135 123.63 ;
      RECT 26.625 116.84 27.135 116.9 ;
      RECT 26.615 106.9 27.145 113.57 ;
      RECT 26.625 113.57 27.135 113.63 ;
      RECT 26.625 106.84 27.135 106.9 ;
      RECT 26.615 96.9 27.145 103.57 ;
      RECT 26.625 103.57 27.135 103.63 ;
      RECT 26.625 96.84 27.135 96.9 ;
      RECT 29.385 116.9 29.915 123.57 ;
      RECT 29.395 123.57 29.905 123.63 ;
      RECT 29.395 116.84 29.905 116.9 ;
      RECT 29.385 106.9 29.915 113.57 ;
      RECT 29.395 113.57 29.905 113.63 ;
      RECT 29.395 106.84 29.905 106.9 ;
      RECT 29.385 96.9 29.915 103.57 ;
      RECT 29.395 103.57 29.905 103.63 ;
      RECT 29.395 96.84 29.905 96.9 ;
      RECT 33.36 116.84 34.25 123.63 ;
      RECT 30.59 116.84 31.48 123.63 ;
      RECT 33.36 106.84 34.25 113.63 ;
      RECT 30.59 106.84 31.48 113.63 ;
      RECT 33.36 96.84 34.25 103.63 ;
      RECT 30.59 96.84 31.48 103.63 ;
      RECT 32.155 116.9 32.685 123.57 ;
      RECT 32.165 123.57 32.675 123.63 ;
      RECT 32.165 116.84 32.675 116.9 ;
      RECT 32.155 106.9 32.685 113.57 ;
      RECT 32.165 113.57 32.675 113.63 ;
      RECT 32.165 106.84 32.675 106.9 ;
      RECT 32.155 96.9 32.685 103.57 ;
      RECT 13.52 144.825 23.46 144.91 ;
      RECT 13.24 85.36 23.46 144.825 ;
      RECT 13.24 79.675 39.54 85.36 ;
      RECT 13.52 79.56 39.54 79.675 ;
      RECT 11.37 49.595 12.22 194.86 ;
      RECT 11.37 49.15 41.095 49.595 ;
      RECT 11.37 194.86 41.095 195.71 ;
      RECT 40.245 49.595 41.095 194.86 ;
      RECT 9.73 16.735 39.195 17.265 ;
      RECT 42.145 48.73 42.675 196.85 ;
      RECT 38.665 17.265 39.195 47.68 ;
      RECT 9.73 17.265 10.28 17.295 ;
      RECT 38.665 48.525 42.675 48.73 ;
      RECT 38.665 47.68 42.675 47.935 ;
      RECT 9.69 17.295 10.28 47.935 ;
      RECT 9.69 196.85 42.675 197.38 ;
      RECT 9.69 48.525 10.28 196.85 ;
      RECT 9.69 47.935 42.675 48.525 ;
      RECT 0.405 1.3 1.1 1.47 ;
      RECT 0.405 1.47 1.095 1.48 ;
      RECT 0.405 0.48 1.095 1.3 ;
      RECT 6.79 0.515 8.39 1.495 ;
      RECT 6.79 1.495 8.345 1.705 ;
      RECT 9.005 4.49 9.175 9.91 ;
      RECT 9.005 4.32 25.195 4.49 ;
      RECT 9.005 9.91 25.195 10.08 ;
      RECT 25.025 4.49 25.195 9.91 ;
      RECT 9.595 5.04 9.765 9.36 ;
      RECT 17.245 5.04 17.415 9.36 ;
      RECT 13.435 20.795 13.605 27.73 ;
      RECT 12.975 20.795 13.145 27.585 ;
      RECT 12.085 30.27 12.305 37.06 ;
      RECT 12.085 39.27 12.305 46.06 ;
      RECT 10.705 19.185 38.065 19.715 ;
      RECT 10.705 38.435 11.67 46.98 ;
      RECT 37.435 29.235 38.065 38.205 ;
      RECT 10.705 19.715 11.67 29.005 ;
      RECT 37.435 38.435 38.065 46.98 ;
      RECT 10.705 29.235 11.67 38.205 ;
      RECT 37.435 19.715 38.065 29.005 ;
      RECT 10.705 46.98 38.065 47.275 ;
      RECT 10.705 29.005 38.065 29.235 ;
      RECT 10.705 38.205 38.065 38.435 ;
      RECT 13.895 20.795 14.065 27.585 ;
      RECT 18.135 20.795 18.355 26.595 ;
      RECT 18.175 26.595 18.345 27.585 ;
      RECT 20.37 30.27 20.59 37.06 ;
      RECT 20.37 39.27 20.59 46.06 ;
      RECT 22.43 20.795 22.65 26.595 ;
      RECT 22.455 26.595 22.625 27.585 ;
      RECT 26.71 20.795 26.93 26.595 ;
      RECT 26.735 26.595 26.905 27.585 ;
      RECT 28.66 30.27 28.88 37.06 ;
      RECT 28.66 39.27 28.88 46.06 ;
      RECT 31.005 20.795 31.225 26.595 ;
      RECT 31.015 26.595 31.185 27.585 ;
      RECT 35.27 20.795 35.49 26.595 ;
      RECT 35.295 26.595 35.465 27.585 ;
      RECT 36.905 30.27 37.125 37.06 ;
      RECT 36.905 39.27 37.125 46.06 ;
      RECT 16.74 60.5 17.63 67.29 ;
      RECT 13.97 60.5 14.86 67.29 ;
      RECT 16.74 50.5 17.63 57.29 ;
      RECT 13.97 50.5 14.86 57.29 ;
      RECT 15.535 60.56 16.065 67.23 ;
      RECT 15.545 67.23 16.055 67.29 ;
      RECT 15.545 60.5 16.055 60.56 ;
      RECT 15.535 50.56 16.065 57.23 ;
      RECT 15.545 57.23 16.055 57.29 ;
      RECT 15.545 50.5 16.055 50.56 ;
      RECT 19.51 60.5 20.4 67.29 ;
      RECT 19.51 50.5 20.4 57.29 ;
      RECT 21.075 60.56 21.605 67.23 ;
      RECT 21.085 67.23 21.595 67.29 ;
      RECT 21.085 60.5 21.595 60.56 ;
      RECT 21.075 50.56 21.605 57.23 ;
      RECT 21.085 57.23 21.595 57.29 ;
      RECT 21.085 50.5 21.595 50.56 ;
      RECT 18.305 60.56 18.835 67.23 ;
      RECT 18.315 67.23 18.825 67.29 ;
      RECT 18.315 60.5 18.825 60.56 ;
      RECT 18.305 50.56 18.835 57.23 ;
      RECT 18.315 57.23 18.825 57.29 ;
      RECT 18.315 50.5 18.825 50.56 ;
      RECT 25.05 60.5 25.94 67.29 ;
      RECT 22.28 60.5 23.17 67.29 ;
      RECT 25.05 50.5 25.94 57.29 ;
      RECT 22.28 50.5 23.17 57.29 ;
      RECT 23.845 60.56 24.375 67.23 ;
      RECT 23.855 67.23 24.365 67.29 ;
      RECT 23.855 60.5 24.365 60.56 ;
      RECT 23.845 50.56 24.375 57.23 ;
      RECT 23.855 57.23 24.365 57.29 ;
      RECT 23.855 50.5 24.365 50.56 ;
    LAYER met1 ;
      RECT 0 16.515 38.445 16.565 ;
      RECT 0 0 38.495 16.515 ;
      RECT 0 197.55 47.895 198 ;
      RECT 0 16.565 9.55 197.55 ;
      RECT 10.605 48.9 41.895 49.085 ;
      RECT 10.42 17.52 38.495 47.375 ;
      RECT 10.42 196.59 41.815 196.68 ;
      RECT 10.42 47.375 38.495 47.475 ;
      RECT 10.42 196.52 41.905 196.59 ;
      RECT 10.42 49.165 41.975 196.52 ;
      RECT 10.465 17.435 38.455 17.48 ;
      RECT 10.42 17.48 38.495 17.52 ;
      RECT 10.42 49.085 41.975 49.165 ;
      RECT 10.52 47.475 38.41 47.56 ;
      RECT 39.525 0 47.895 47.47 ;
      RECT 39.525 47.47 47.895 47.56 ;
      RECT 43.005 47.56 47.895 197.55 ;
      RECT 9.41 197.69 43.145 198 ;
      RECT 39.665 0 47.895 47.42 ;
      RECT 43.145 47.42 47.895 198 ;
      RECT 0 16.425 9.41 198 ;
      RECT 0 0 38.355 16.425 ;
      RECT 10.56 52.225 13.565 193.46 ;
      RECT 10.56 49.22 41.835 52.225 ;
      RECT 10.56 193.46 41.835 196.465 ;
      RECT 38.83 52.225 41.835 193.46 ;
      RECT 13.56 52.04 38.835 193.54 ;
      RECT 10.66 49.04 41.655 49.09 ;
      RECT 10.61 49.09 41.705 49.14 ;
      RECT 10.56 49.14 41.755 49.18 ;
      RECT 10.56 49.18 41.795 49.22 ;
      RECT 10.56 196.465 41.8 196.5 ;
      RECT 10.56 196.5 41.76 196.54 ;
      RECT 10.56 20.58 13.565 44.315 ;
      RECT 10.56 17.575 38.355 20.58 ;
      RECT 10.56 44.315 38.355 47.32 ;
      RECT 35.35 20.58 38.355 44.315 ;
      RECT 13.56 20.575 35.355 44.42 ;
      RECT 10.61 47.32 38.355 47.37 ;
      RECT 10.66 47.37 38.355 47.42 ;
    LAYER met5 ;
      RECT 0 0 47.895 198 ;
    LAYER met4 ;
      RECT 0 0 47.895 198 ;
    LAYER met3 ;
      RECT 26.94 0 27.64 190.36 ;
      RECT 41.49 0 47.895 194.075 ;
      RECT 0 194.075 47.895 198 ;
      RECT 0 190.36 27.64 194.075 ;
      RECT 0 0 13.22 190.36 ;
    LAYER met2 ;
      RECT 0 0 47.895 198 ;
  END
END sky130_fd_io__top_lvclamp
  
END LIBRARY
