# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_io__overlay_vdda_lvc
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 198 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 1.270000 54.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 1.270000 49.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 6.885000 1.270000 11.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 6.885000 75.000000 11.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 6.985000 1.270000 11.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 0.035000 1.270000 5.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 0.035000 75.000000 5.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 0.135000 1.270000 5.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.600000 12.940000 24.500000 16.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000 12.940000 74.655000 16.380000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 12.935000 24.475000 16.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.780000 12.935000 75.000000 16.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 13.035000 0.965000 16.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.690000 13.020000  0.890000 13.220000 ;
        RECT  0.690000 13.460000  0.890000 13.660000 ;
        RECT  0.690000 13.900000  0.890000 14.100000 ;
        RECT  0.690000 14.340000  0.890000 14.540000 ;
        RECT  0.690000 14.780000  0.890000 14.980000 ;
        RECT  0.690000 15.220000  0.890000 15.420000 ;
        RECT  0.690000 15.660000  0.890000 15.860000 ;
        RECT  0.690000 16.100000  0.890000 16.300000 ;
        RECT  1.100000 13.020000  1.300000 13.220000 ;
        RECT  1.100000 13.460000  1.300000 13.660000 ;
        RECT  1.100000 13.900000  1.300000 14.100000 ;
        RECT  1.100000 14.340000  1.300000 14.540000 ;
        RECT  1.100000 14.780000  1.300000 14.980000 ;
        RECT  1.100000 15.220000  1.300000 15.420000 ;
        RECT  1.100000 15.660000  1.300000 15.860000 ;
        RECT  1.100000 16.100000  1.300000 16.300000 ;
        RECT  1.510000 13.020000  1.710000 13.220000 ;
        RECT  1.510000 13.460000  1.710000 13.660000 ;
        RECT  1.510000 13.900000  1.710000 14.100000 ;
        RECT  1.510000 14.340000  1.710000 14.540000 ;
        RECT  1.510000 14.780000  1.710000 14.980000 ;
        RECT  1.510000 15.220000  1.710000 15.420000 ;
        RECT  1.510000 15.660000  1.710000 15.860000 ;
        RECT  1.510000 16.100000  1.710000 16.300000 ;
        RECT  1.920000 13.020000  2.120000 13.220000 ;
        RECT  1.920000 13.460000  2.120000 13.660000 ;
        RECT  1.920000 13.900000  2.120000 14.100000 ;
        RECT  1.920000 14.340000  2.120000 14.540000 ;
        RECT  1.920000 14.780000  2.120000 14.980000 ;
        RECT  1.920000 15.220000  2.120000 15.420000 ;
        RECT  1.920000 15.660000  2.120000 15.860000 ;
        RECT  1.920000 16.100000  2.120000 16.300000 ;
        RECT  2.330000 13.020000  2.530000 13.220000 ;
        RECT  2.330000 13.460000  2.530000 13.660000 ;
        RECT  2.330000 13.900000  2.530000 14.100000 ;
        RECT  2.330000 14.340000  2.530000 14.540000 ;
        RECT  2.330000 14.780000  2.530000 14.980000 ;
        RECT  2.330000 15.220000  2.530000 15.420000 ;
        RECT  2.330000 15.660000  2.530000 15.860000 ;
        RECT  2.330000 16.100000  2.530000 16.300000 ;
        RECT  2.740000 13.020000  2.940000 13.220000 ;
        RECT  2.740000 13.460000  2.940000 13.660000 ;
        RECT  2.740000 13.900000  2.940000 14.100000 ;
        RECT  2.740000 14.340000  2.940000 14.540000 ;
        RECT  2.740000 14.780000  2.940000 14.980000 ;
        RECT  2.740000 15.220000  2.940000 15.420000 ;
        RECT  2.740000 15.660000  2.940000 15.860000 ;
        RECT  2.740000 16.100000  2.940000 16.300000 ;
        RECT  3.150000 13.020000  3.350000 13.220000 ;
        RECT  3.150000 13.460000  3.350000 13.660000 ;
        RECT  3.150000 13.900000  3.350000 14.100000 ;
        RECT  3.150000 14.340000  3.350000 14.540000 ;
        RECT  3.150000 14.780000  3.350000 14.980000 ;
        RECT  3.150000 15.220000  3.350000 15.420000 ;
        RECT  3.150000 15.660000  3.350000 15.860000 ;
        RECT  3.150000 16.100000  3.350000 16.300000 ;
        RECT  3.555000 13.020000  3.755000 13.220000 ;
        RECT  3.555000 13.460000  3.755000 13.660000 ;
        RECT  3.555000 13.900000  3.755000 14.100000 ;
        RECT  3.555000 14.340000  3.755000 14.540000 ;
        RECT  3.555000 14.780000  3.755000 14.980000 ;
        RECT  3.555000 15.220000  3.755000 15.420000 ;
        RECT  3.555000 15.660000  3.755000 15.860000 ;
        RECT  3.555000 16.100000  3.755000 16.300000 ;
        RECT  3.960000 13.020000  4.160000 13.220000 ;
        RECT  3.960000 13.460000  4.160000 13.660000 ;
        RECT  3.960000 13.900000  4.160000 14.100000 ;
        RECT  3.960000 14.340000  4.160000 14.540000 ;
        RECT  3.960000 14.780000  4.160000 14.980000 ;
        RECT  3.960000 15.220000  4.160000 15.420000 ;
        RECT  3.960000 15.660000  4.160000 15.860000 ;
        RECT  3.960000 16.100000  4.160000 16.300000 ;
        RECT  4.365000 13.020000  4.565000 13.220000 ;
        RECT  4.365000 13.460000  4.565000 13.660000 ;
        RECT  4.365000 13.900000  4.565000 14.100000 ;
        RECT  4.365000 14.340000  4.565000 14.540000 ;
        RECT  4.365000 14.780000  4.565000 14.980000 ;
        RECT  4.365000 15.220000  4.565000 15.420000 ;
        RECT  4.365000 15.660000  4.565000 15.860000 ;
        RECT  4.365000 16.100000  4.565000 16.300000 ;
        RECT  4.770000 13.020000  4.970000 13.220000 ;
        RECT  4.770000 13.460000  4.970000 13.660000 ;
        RECT  4.770000 13.900000  4.970000 14.100000 ;
        RECT  4.770000 14.340000  4.970000 14.540000 ;
        RECT  4.770000 14.780000  4.970000 14.980000 ;
        RECT  4.770000 15.220000  4.970000 15.420000 ;
        RECT  4.770000 15.660000  4.970000 15.860000 ;
        RECT  4.770000 16.100000  4.970000 16.300000 ;
        RECT  5.175000 13.020000  5.375000 13.220000 ;
        RECT  5.175000 13.460000  5.375000 13.660000 ;
        RECT  5.175000 13.900000  5.375000 14.100000 ;
        RECT  5.175000 14.340000  5.375000 14.540000 ;
        RECT  5.175000 14.780000  5.375000 14.980000 ;
        RECT  5.175000 15.220000  5.375000 15.420000 ;
        RECT  5.175000 15.660000  5.375000 15.860000 ;
        RECT  5.175000 16.100000  5.375000 16.300000 ;
        RECT  5.580000 13.020000  5.780000 13.220000 ;
        RECT  5.580000 13.460000  5.780000 13.660000 ;
        RECT  5.580000 13.900000  5.780000 14.100000 ;
        RECT  5.580000 14.340000  5.780000 14.540000 ;
        RECT  5.580000 14.780000  5.780000 14.980000 ;
        RECT  5.580000 15.220000  5.780000 15.420000 ;
        RECT  5.580000 15.660000  5.780000 15.860000 ;
        RECT  5.580000 16.100000  5.780000 16.300000 ;
        RECT  5.985000 13.020000  6.185000 13.220000 ;
        RECT  5.985000 13.460000  6.185000 13.660000 ;
        RECT  5.985000 13.900000  6.185000 14.100000 ;
        RECT  5.985000 14.340000  6.185000 14.540000 ;
        RECT  5.985000 14.780000  6.185000 14.980000 ;
        RECT  5.985000 15.220000  6.185000 15.420000 ;
        RECT  5.985000 15.660000  6.185000 15.860000 ;
        RECT  5.985000 16.100000  6.185000 16.300000 ;
        RECT  6.390000 13.020000  6.590000 13.220000 ;
        RECT  6.390000 13.460000  6.590000 13.660000 ;
        RECT  6.390000 13.900000  6.590000 14.100000 ;
        RECT  6.390000 14.340000  6.590000 14.540000 ;
        RECT  6.390000 14.780000  6.590000 14.980000 ;
        RECT  6.390000 15.220000  6.590000 15.420000 ;
        RECT  6.390000 15.660000  6.590000 15.860000 ;
        RECT  6.390000 16.100000  6.590000 16.300000 ;
        RECT  6.795000 13.020000  6.995000 13.220000 ;
        RECT  6.795000 13.460000  6.995000 13.660000 ;
        RECT  6.795000 13.900000  6.995000 14.100000 ;
        RECT  6.795000 14.340000  6.995000 14.540000 ;
        RECT  6.795000 14.780000  6.995000 14.980000 ;
        RECT  6.795000 15.220000  6.995000 15.420000 ;
        RECT  6.795000 15.660000  6.995000 15.860000 ;
        RECT  6.795000 16.100000  6.995000 16.300000 ;
        RECT  7.200000 13.020000  7.400000 13.220000 ;
        RECT  7.200000 13.460000  7.400000 13.660000 ;
        RECT  7.200000 13.900000  7.400000 14.100000 ;
        RECT  7.200000 14.340000  7.400000 14.540000 ;
        RECT  7.200000 14.780000  7.400000 14.980000 ;
        RECT  7.200000 15.220000  7.400000 15.420000 ;
        RECT  7.200000 15.660000  7.400000 15.860000 ;
        RECT  7.200000 16.100000  7.400000 16.300000 ;
        RECT  7.605000 13.020000  7.805000 13.220000 ;
        RECT  7.605000 13.460000  7.805000 13.660000 ;
        RECT  7.605000 13.900000  7.805000 14.100000 ;
        RECT  7.605000 14.340000  7.805000 14.540000 ;
        RECT  7.605000 14.780000  7.805000 14.980000 ;
        RECT  7.605000 15.220000  7.805000 15.420000 ;
        RECT  7.605000 15.660000  7.805000 15.860000 ;
        RECT  7.605000 16.100000  7.805000 16.300000 ;
        RECT  8.010000 13.020000  8.210000 13.220000 ;
        RECT  8.010000 13.460000  8.210000 13.660000 ;
        RECT  8.010000 13.900000  8.210000 14.100000 ;
        RECT  8.010000 14.340000  8.210000 14.540000 ;
        RECT  8.010000 14.780000  8.210000 14.980000 ;
        RECT  8.010000 15.220000  8.210000 15.420000 ;
        RECT  8.010000 15.660000  8.210000 15.860000 ;
        RECT  8.010000 16.100000  8.210000 16.300000 ;
        RECT  8.415000 13.020000  8.615000 13.220000 ;
        RECT  8.415000 13.460000  8.615000 13.660000 ;
        RECT  8.415000 13.900000  8.615000 14.100000 ;
        RECT  8.415000 14.340000  8.615000 14.540000 ;
        RECT  8.415000 14.780000  8.615000 14.980000 ;
        RECT  8.415000 15.220000  8.615000 15.420000 ;
        RECT  8.415000 15.660000  8.615000 15.860000 ;
        RECT  8.415000 16.100000  8.615000 16.300000 ;
        RECT  8.820000 13.020000  9.020000 13.220000 ;
        RECT  8.820000 13.460000  9.020000 13.660000 ;
        RECT  8.820000 13.900000  9.020000 14.100000 ;
        RECT  8.820000 14.340000  9.020000 14.540000 ;
        RECT  8.820000 14.780000  9.020000 14.980000 ;
        RECT  8.820000 15.220000  9.020000 15.420000 ;
        RECT  8.820000 15.660000  9.020000 15.860000 ;
        RECT  8.820000 16.100000  9.020000 16.300000 ;
        RECT  9.225000 13.020000  9.425000 13.220000 ;
        RECT  9.225000 13.460000  9.425000 13.660000 ;
        RECT  9.225000 13.900000  9.425000 14.100000 ;
        RECT  9.225000 14.340000  9.425000 14.540000 ;
        RECT  9.225000 14.780000  9.425000 14.980000 ;
        RECT  9.225000 15.220000  9.425000 15.420000 ;
        RECT  9.225000 15.660000  9.425000 15.860000 ;
        RECT  9.225000 16.100000  9.425000 16.300000 ;
        RECT  9.630000 13.020000  9.830000 13.220000 ;
        RECT  9.630000 13.460000  9.830000 13.660000 ;
        RECT  9.630000 13.900000  9.830000 14.100000 ;
        RECT  9.630000 14.340000  9.830000 14.540000 ;
        RECT  9.630000 14.780000  9.830000 14.980000 ;
        RECT  9.630000 15.220000  9.830000 15.420000 ;
        RECT  9.630000 15.660000  9.830000 15.860000 ;
        RECT  9.630000 16.100000  9.830000 16.300000 ;
        RECT 10.035000 13.020000 10.235000 13.220000 ;
        RECT 10.035000 13.460000 10.235000 13.660000 ;
        RECT 10.035000 13.900000 10.235000 14.100000 ;
        RECT 10.035000 14.340000 10.235000 14.540000 ;
        RECT 10.035000 14.780000 10.235000 14.980000 ;
        RECT 10.035000 15.220000 10.235000 15.420000 ;
        RECT 10.035000 15.660000 10.235000 15.860000 ;
        RECT 10.035000 16.100000 10.235000 16.300000 ;
        RECT 10.440000 13.020000 10.640000 13.220000 ;
        RECT 10.440000 13.460000 10.640000 13.660000 ;
        RECT 10.440000 13.900000 10.640000 14.100000 ;
        RECT 10.440000 14.340000 10.640000 14.540000 ;
        RECT 10.440000 14.780000 10.640000 14.980000 ;
        RECT 10.440000 15.220000 10.640000 15.420000 ;
        RECT 10.440000 15.660000 10.640000 15.860000 ;
        RECT 10.440000 16.100000 10.640000 16.300000 ;
        RECT 10.845000 13.020000 11.045000 13.220000 ;
        RECT 10.845000 13.460000 11.045000 13.660000 ;
        RECT 10.845000 13.900000 11.045000 14.100000 ;
        RECT 10.845000 14.340000 11.045000 14.540000 ;
        RECT 10.845000 14.780000 11.045000 14.980000 ;
        RECT 10.845000 15.220000 11.045000 15.420000 ;
        RECT 10.845000 15.660000 11.045000 15.860000 ;
        RECT 10.845000 16.100000 11.045000 16.300000 ;
        RECT 11.250000 13.020000 11.450000 13.220000 ;
        RECT 11.250000 13.460000 11.450000 13.660000 ;
        RECT 11.250000 13.900000 11.450000 14.100000 ;
        RECT 11.250000 14.340000 11.450000 14.540000 ;
        RECT 11.250000 14.780000 11.450000 14.980000 ;
        RECT 11.250000 15.220000 11.450000 15.420000 ;
        RECT 11.250000 15.660000 11.450000 15.860000 ;
        RECT 11.250000 16.100000 11.450000 16.300000 ;
        RECT 11.655000 13.020000 11.855000 13.220000 ;
        RECT 11.655000 13.460000 11.855000 13.660000 ;
        RECT 11.655000 13.900000 11.855000 14.100000 ;
        RECT 11.655000 14.340000 11.855000 14.540000 ;
        RECT 11.655000 14.780000 11.855000 14.980000 ;
        RECT 11.655000 15.220000 11.855000 15.420000 ;
        RECT 11.655000 15.660000 11.855000 15.860000 ;
        RECT 11.655000 16.100000 11.855000 16.300000 ;
        RECT 12.060000 13.020000 12.260000 13.220000 ;
        RECT 12.060000 13.460000 12.260000 13.660000 ;
        RECT 12.060000 13.900000 12.260000 14.100000 ;
        RECT 12.060000 14.340000 12.260000 14.540000 ;
        RECT 12.060000 14.780000 12.260000 14.980000 ;
        RECT 12.060000 15.220000 12.260000 15.420000 ;
        RECT 12.060000 15.660000 12.260000 15.860000 ;
        RECT 12.060000 16.100000 12.260000 16.300000 ;
        RECT 12.465000 13.020000 12.665000 13.220000 ;
        RECT 12.465000 13.460000 12.665000 13.660000 ;
        RECT 12.465000 13.900000 12.665000 14.100000 ;
        RECT 12.465000 14.340000 12.665000 14.540000 ;
        RECT 12.465000 14.780000 12.665000 14.980000 ;
        RECT 12.465000 15.220000 12.665000 15.420000 ;
        RECT 12.465000 15.660000 12.665000 15.860000 ;
        RECT 12.465000 16.100000 12.665000 16.300000 ;
        RECT 12.870000 13.020000 13.070000 13.220000 ;
        RECT 12.870000 13.460000 13.070000 13.660000 ;
        RECT 12.870000 13.900000 13.070000 14.100000 ;
        RECT 12.870000 14.340000 13.070000 14.540000 ;
        RECT 12.870000 14.780000 13.070000 14.980000 ;
        RECT 12.870000 15.220000 13.070000 15.420000 ;
        RECT 12.870000 15.660000 13.070000 15.860000 ;
        RECT 12.870000 16.100000 13.070000 16.300000 ;
        RECT 13.275000 13.020000 13.475000 13.220000 ;
        RECT 13.275000 13.460000 13.475000 13.660000 ;
        RECT 13.275000 13.900000 13.475000 14.100000 ;
        RECT 13.275000 14.340000 13.475000 14.540000 ;
        RECT 13.275000 14.780000 13.475000 14.980000 ;
        RECT 13.275000 15.220000 13.475000 15.420000 ;
        RECT 13.275000 15.660000 13.475000 15.860000 ;
        RECT 13.275000 16.100000 13.475000 16.300000 ;
        RECT 13.680000 13.020000 13.880000 13.220000 ;
        RECT 13.680000 13.460000 13.880000 13.660000 ;
        RECT 13.680000 13.900000 13.880000 14.100000 ;
        RECT 13.680000 14.340000 13.880000 14.540000 ;
        RECT 13.680000 14.780000 13.880000 14.980000 ;
        RECT 13.680000 15.220000 13.880000 15.420000 ;
        RECT 13.680000 15.660000 13.880000 15.860000 ;
        RECT 13.680000 16.100000 13.880000 16.300000 ;
        RECT 14.085000 13.020000 14.285000 13.220000 ;
        RECT 14.085000 13.460000 14.285000 13.660000 ;
        RECT 14.085000 13.900000 14.285000 14.100000 ;
        RECT 14.085000 14.340000 14.285000 14.540000 ;
        RECT 14.085000 14.780000 14.285000 14.980000 ;
        RECT 14.085000 15.220000 14.285000 15.420000 ;
        RECT 14.085000 15.660000 14.285000 15.860000 ;
        RECT 14.085000 16.100000 14.285000 16.300000 ;
        RECT 14.490000 13.020000 14.690000 13.220000 ;
        RECT 14.490000 13.460000 14.690000 13.660000 ;
        RECT 14.490000 13.900000 14.690000 14.100000 ;
        RECT 14.490000 14.340000 14.690000 14.540000 ;
        RECT 14.490000 14.780000 14.690000 14.980000 ;
        RECT 14.490000 15.220000 14.690000 15.420000 ;
        RECT 14.490000 15.660000 14.690000 15.860000 ;
        RECT 14.490000 16.100000 14.690000 16.300000 ;
        RECT 14.895000 13.020000 15.095000 13.220000 ;
        RECT 14.895000 13.460000 15.095000 13.660000 ;
        RECT 14.895000 13.900000 15.095000 14.100000 ;
        RECT 14.895000 14.340000 15.095000 14.540000 ;
        RECT 14.895000 14.780000 15.095000 14.980000 ;
        RECT 14.895000 15.220000 15.095000 15.420000 ;
        RECT 14.895000 15.660000 15.095000 15.860000 ;
        RECT 14.895000 16.100000 15.095000 16.300000 ;
        RECT 15.300000 13.020000 15.500000 13.220000 ;
        RECT 15.300000 13.460000 15.500000 13.660000 ;
        RECT 15.300000 13.900000 15.500000 14.100000 ;
        RECT 15.300000 14.340000 15.500000 14.540000 ;
        RECT 15.300000 14.780000 15.500000 14.980000 ;
        RECT 15.300000 15.220000 15.500000 15.420000 ;
        RECT 15.300000 15.660000 15.500000 15.860000 ;
        RECT 15.300000 16.100000 15.500000 16.300000 ;
        RECT 15.705000 13.020000 15.905000 13.220000 ;
        RECT 15.705000 13.460000 15.905000 13.660000 ;
        RECT 15.705000 13.900000 15.905000 14.100000 ;
        RECT 15.705000 14.340000 15.905000 14.540000 ;
        RECT 15.705000 14.780000 15.905000 14.980000 ;
        RECT 15.705000 15.220000 15.905000 15.420000 ;
        RECT 15.705000 15.660000 15.905000 15.860000 ;
        RECT 15.705000 16.100000 15.905000 16.300000 ;
        RECT 16.110000 13.020000 16.310000 13.220000 ;
        RECT 16.110000 13.460000 16.310000 13.660000 ;
        RECT 16.110000 13.900000 16.310000 14.100000 ;
        RECT 16.110000 14.340000 16.310000 14.540000 ;
        RECT 16.110000 14.780000 16.310000 14.980000 ;
        RECT 16.110000 15.220000 16.310000 15.420000 ;
        RECT 16.110000 15.660000 16.310000 15.860000 ;
        RECT 16.110000 16.100000 16.310000 16.300000 ;
        RECT 16.515000 13.020000 16.715000 13.220000 ;
        RECT 16.515000 13.460000 16.715000 13.660000 ;
        RECT 16.515000 13.900000 16.715000 14.100000 ;
        RECT 16.515000 14.340000 16.715000 14.540000 ;
        RECT 16.515000 14.780000 16.715000 14.980000 ;
        RECT 16.515000 15.220000 16.715000 15.420000 ;
        RECT 16.515000 15.660000 16.715000 15.860000 ;
        RECT 16.515000 16.100000 16.715000 16.300000 ;
        RECT 16.920000 13.020000 17.120000 13.220000 ;
        RECT 16.920000 13.460000 17.120000 13.660000 ;
        RECT 16.920000 13.900000 17.120000 14.100000 ;
        RECT 16.920000 14.340000 17.120000 14.540000 ;
        RECT 16.920000 14.780000 17.120000 14.980000 ;
        RECT 16.920000 15.220000 17.120000 15.420000 ;
        RECT 16.920000 15.660000 17.120000 15.860000 ;
        RECT 16.920000 16.100000 17.120000 16.300000 ;
        RECT 17.325000 13.020000 17.525000 13.220000 ;
        RECT 17.325000 13.460000 17.525000 13.660000 ;
        RECT 17.325000 13.900000 17.525000 14.100000 ;
        RECT 17.325000 14.340000 17.525000 14.540000 ;
        RECT 17.325000 14.780000 17.525000 14.980000 ;
        RECT 17.325000 15.220000 17.525000 15.420000 ;
        RECT 17.325000 15.660000 17.525000 15.860000 ;
        RECT 17.325000 16.100000 17.525000 16.300000 ;
        RECT 17.730000 13.020000 17.930000 13.220000 ;
        RECT 17.730000 13.460000 17.930000 13.660000 ;
        RECT 17.730000 13.900000 17.930000 14.100000 ;
        RECT 17.730000 14.340000 17.930000 14.540000 ;
        RECT 17.730000 14.780000 17.930000 14.980000 ;
        RECT 17.730000 15.220000 17.930000 15.420000 ;
        RECT 17.730000 15.660000 17.930000 15.860000 ;
        RECT 17.730000 16.100000 17.930000 16.300000 ;
        RECT 18.135000 13.020000 18.335000 13.220000 ;
        RECT 18.135000 13.460000 18.335000 13.660000 ;
        RECT 18.135000 13.900000 18.335000 14.100000 ;
        RECT 18.135000 14.340000 18.335000 14.540000 ;
        RECT 18.135000 14.780000 18.335000 14.980000 ;
        RECT 18.135000 15.220000 18.335000 15.420000 ;
        RECT 18.135000 15.660000 18.335000 15.860000 ;
        RECT 18.135000 16.100000 18.335000 16.300000 ;
        RECT 18.540000 13.020000 18.740000 13.220000 ;
        RECT 18.540000 13.460000 18.740000 13.660000 ;
        RECT 18.540000 13.900000 18.740000 14.100000 ;
        RECT 18.540000 14.340000 18.740000 14.540000 ;
        RECT 18.540000 14.780000 18.740000 14.980000 ;
        RECT 18.540000 15.220000 18.740000 15.420000 ;
        RECT 18.540000 15.660000 18.740000 15.860000 ;
        RECT 18.540000 16.100000 18.740000 16.300000 ;
        RECT 18.945000 13.020000 19.145000 13.220000 ;
        RECT 18.945000 13.460000 19.145000 13.660000 ;
        RECT 18.945000 13.900000 19.145000 14.100000 ;
        RECT 18.945000 14.340000 19.145000 14.540000 ;
        RECT 18.945000 14.780000 19.145000 14.980000 ;
        RECT 18.945000 15.220000 19.145000 15.420000 ;
        RECT 18.945000 15.660000 19.145000 15.860000 ;
        RECT 18.945000 16.100000 19.145000 16.300000 ;
        RECT 19.350000 13.020000 19.550000 13.220000 ;
        RECT 19.350000 13.460000 19.550000 13.660000 ;
        RECT 19.350000 13.900000 19.550000 14.100000 ;
        RECT 19.350000 14.340000 19.550000 14.540000 ;
        RECT 19.350000 14.780000 19.550000 14.980000 ;
        RECT 19.350000 15.220000 19.550000 15.420000 ;
        RECT 19.350000 15.660000 19.550000 15.860000 ;
        RECT 19.350000 16.100000 19.550000 16.300000 ;
        RECT 19.755000 13.020000 19.955000 13.220000 ;
        RECT 19.755000 13.460000 19.955000 13.660000 ;
        RECT 19.755000 13.900000 19.955000 14.100000 ;
        RECT 19.755000 14.340000 19.955000 14.540000 ;
        RECT 19.755000 14.780000 19.955000 14.980000 ;
        RECT 19.755000 15.220000 19.955000 15.420000 ;
        RECT 19.755000 15.660000 19.955000 15.860000 ;
        RECT 19.755000 16.100000 19.955000 16.300000 ;
        RECT 20.160000 13.020000 20.360000 13.220000 ;
        RECT 20.160000 13.460000 20.360000 13.660000 ;
        RECT 20.160000 13.900000 20.360000 14.100000 ;
        RECT 20.160000 14.340000 20.360000 14.540000 ;
        RECT 20.160000 14.780000 20.360000 14.980000 ;
        RECT 20.160000 15.220000 20.360000 15.420000 ;
        RECT 20.160000 15.660000 20.360000 15.860000 ;
        RECT 20.160000 16.100000 20.360000 16.300000 ;
        RECT 20.565000 13.020000 20.765000 13.220000 ;
        RECT 20.565000 13.460000 20.765000 13.660000 ;
        RECT 20.565000 13.900000 20.765000 14.100000 ;
        RECT 20.565000 14.340000 20.765000 14.540000 ;
        RECT 20.565000 14.780000 20.765000 14.980000 ;
        RECT 20.565000 15.220000 20.765000 15.420000 ;
        RECT 20.565000 15.660000 20.765000 15.860000 ;
        RECT 20.565000 16.100000 20.765000 16.300000 ;
        RECT 20.970000 13.020000 21.170000 13.220000 ;
        RECT 20.970000 13.460000 21.170000 13.660000 ;
        RECT 20.970000 13.900000 21.170000 14.100000 ;
        RECT 20.970000 14.340000 21.170000 14.540000 ;
        RECT 20.970000 14.780000 21.170000 14.980000 ;
        RECT 20.970000 15.220000 21.170000 15.420000 ;
        RECT 20.970000 15.660000 21.170000 15.860000 ;
        RECT 20.970000 16.100000 21.170000 16.300000 ;
        RECT 21.375000 13.020000 21.575000 13.220000 ;
        RECT 21.375000 13.460000 21.575000 13.660000 ;
        RECT 21.375000 13.900000 21.575000 14.100000 ;
        RECT 21.375000 14.340000 21.575000 14.540000 ;
        RECT 21.375000 14.780000 21.575000 14.980000 ;
        RECT 21.375000 15.220000 21.575000 15.420000 ;
        RECT 21.375000 15.660000 21.575000 15.860000 ;
        RECT 21.375000 16.100000 21.575000 16.300000 ;
        RECT 21.780000 13.020000 21.980000 13.220000 ;
        RECT 21.780000 13.460000 21.980000 13.660000 ;
        RECT 21.780000 13.900000 21.980000 14.100000 ;
        RECT 21.780000 14.340000 21.980000 14.540000 ;
        RECT 21.780000 14.780000 21.980000 14.980000 ;
        RECT 21.780000 15.220000 21.980000 15.420000 ;
        RECT 21.780000 15.660000 21.980000 15.860000 ;
        RECT 21.780000 16.100000 21.980000 16.300000 ;
        RECT 22.185000 13.020000 22.385000 13.220000 ;
        RECT 22.185000 13.460000 22.385000 13.660000 ;
        RECT 22.185000 13.900000 22.385000 14.100000 ;
        RECT 22.185000 14.340000 22.385000 14.540000 ;
        RECT 22.185000 14.780000 22.385000 14.980000 ;
        RECT 22.185000 15.220000 22.385000 15.420000 ;
        RECT 22.185000 15.660000 22.385000 15.860000 ;
        RECT 22.185000 16.100000 22.385000 16.300000 ;
        RECT 22.590000 13.020000 22.790000 13.220000 ;
        RECT 22.590000 13.460000 22.790000 13.660000 ;
        RECT 22.590000 13.900000 22.790000 14.100000 ;
        RECT 22.590000 14.340000 22.790000 14.540000 ;
        RECT 22.590000 14.780000 22.790000 14.980000 ;
        RECT 22.590000 15.220000 22.790000 15.420000 ;
        RECT 22.590000 15.660000 22.790000 15.860000 ;
        RECT 22.590000 16.100000 22.790000 16.300000 ;
        RECT 22.995000 13.020000 23.195000 13.220000 ;
        RECT 22.995000 13.460000 23.195000 13.660000 ;
        RECT 22.995000 13.900000 23.195000 14.100000 ;
        RECT 22.995000 14.340000 23.195000 14.540000 ;
        RECT 22.995000 14.780000 23.195000 14.980000 ;
        RECT 22.995000 15.220000 23.195000 15.420000 ;
        RECT 22.995000 15.660000 23.195000 15.860000 ;
        RECT 22.995000 16.100000 23.195000 16.300000 ;
        RECT 23.400000 13.020000 23.600000 13.220000 ;
        RECT 23.400000 13.460000 23.600000 13.660000 ;
        RECT 23.400000 13.900000 23.600000 14.100000 ;
        RECT 23.400000 14.340000 23.600000 14.540000 ;
        RECT 23.400000 14.780000 23.600000 14.980000 ;
        RECT 23.400000 15.220000 23.600000 15.420000 ;
        RECT 23.400000 15.660000 23.600000 15.860000 ;
        RECT 23.400000 16.100000 23.600000 16.300000 ;
        RECT 23.805000 13.020000 24.005000 13.220000 ;
        RECT 23.805000 13.460000 24.005000 13.660000 ;
        RECT 23.805000 13.900000 24.005000 14.100000 ;
        RECT 23.805000 14.340000 24.005000 14.540000 ;
        RECT 23.805000 14.780000 24.005000 14.980000 ;
        RECT 23.805000 15.220000 24.005000 15.420000 ;
        RECT 23.805000 15.660000 24.005000 15.860000 ;
        RECT 23.805000 16.100000 24.005000 16.300000 ;
        RECT 24.210000 13.020000 24.410000 13.220000 ;
        RECT 24.210000 13.460000 24.410000 13.660000 ;
        RECT 24.210000 13.900000 24.410000 14.100000 ;
        RECT 24.210000 14.340000 24.410000 14.540000 ;
        RECT 24.210000 14.780000 24.410000 14.980000 ;
        RECT 24.210000 15.220000 24.410000 15.420000 ;
        RECT 24.210000 15.660000 24.410000 15.860000 ;
        RECT 24.210000 16.100000 24.410000 16.300000 ;
        RECT 50.845000 13.020000 51.045000 13.220000 ;
        RECT 50.845000 13.460000 51.045000 13.660000 ;
        RECT 50.845000 13.900000 51.045000 14.100000 ;
        RECT 50.845000 14.340000 51.045000 14.540000 ;
        RECT 50.845000 14.780000 51.045000 14.980000 ;
        RECT 50.845000 15.220000 51.045000 15.420000 ;
        RECT 50.845000 15.660000 51.045000 15.860000 ;
        RECT 50.845000 16.100000 51.045000 16.300000 ;
        RECT 51.255000 13.020000 51.455000 13.220000 ;
        RECT 51.255000 13.460000 51.455000 13.660000 ;
        RECT 51.255000 13.900000 51.455000 14.100000 ;
        RECT 51.255000 14.340000 51.455000 14.540000 ;
        RECT 51.255000 14.780000 51.455000 14.980000 ;
        RECT 51.255000 15.220000 51.455000 15.420000 ;
        RECT 51.255000 15.660000 51.455000 15.860000 ;
        RECT 51.255000 16.100000 51.455000 16.300000 ;
        RECT 51.665000 13.020000 51.865000 13.220000 ;
        RECT 51.665000 13.460000 51.865000 13.660000 ;
        RECT 51.665000 13.900000 51.865000 14.100000 ;
        RECT 51.665000 14.340000 51.865000 14.540000 ;
        RECT 51.665000 14.780000 51.865000 14.980000 ;
        RECT 51.665000 15.220000 51.865000 15.420000 ;
        RECT 51.665000 15.660000 51.865000 15.860000 ;
        RECT 51.665000 16.100000 51.865000 16.300000 ;
        RECT 52.075000 13.020000 52.275000 13.220000 ;
        RECT 52.075000 13.460000 52.275000 13.660000 ;
        RECT 52.075000 13.900000 52.275000 14.100000 ;
        RECT 52.075000 14.340000 52.275000 14.540000 ;
        RECT 52.075000 14.780000 52.275000 14.980000 ;
        RECT 52.075000 15.220000 52.275000 15.420000 ;
        RECT 52.075000 15.660000 52.275000 15.860000 ;
        RECT 52.075000 16.100000 52.275000 16.300000 ;
        RECT 52.485000 13.020000 52.685000 13.220000 ;
        RECT 52.485000 13.460000 52.685000 13.660000 ;
        RECT 52.485000 13.900000 52.685000 14.100000 ;
        RECT 52.485000 14.340000 52.685000 14.540000 ;
        RECT 52.485000 14.780000 52.685000 14.980000 ;
        RECT 52.485000 15.220000 52.685000 15.420000 ;
        RECT 52.485000 15.660000 52.685000 15.860000 ;
        RECT 52.485000 16.100000 52.685000 16.300000 ;
        RECT 52.895000 13.020000 53.095000 13.220000 ;
        RECT 52.895000 13.460000 53.095000 13.660000 ;
        RECT 52.895000 13.900000 53.095000 14.100000 ;
        RECT 52.895000 14.340000 53.095000 14.540000 ;
        RECT 52.895000 14.780000 53.095000 14.980000 ;
        RECT 52.895000 15.220000 53.095000 15.420000 ;
        RECT 52.895000 15.660000 53.095000 15.860000 ;
        RECT 52.895000 16.100000 53.095000 16.300000 ;
        RECT 53.305000 13.020000 53.505000 13.220000 ;
        RECT 53.305000 13.460000 53.505000 13.660000 ;
        RECT 53.305000 13.900000 53.505000 14.100000 ;
        RECT 53.305000 14.340000 53.505000 14.540000 ;
        RECT 53.305000 14.780000 53.505000 14.980000 ;
        RECT 53.305000 15.220000 53.505000 15.420000 ;
        RECT 53.305000 15.660000 53.505000 15.860000 ;
        RECT 53.305000 16.100000 53.505000 16.300000 ;
        RECT 53.710000 13.020000 53.910000 13.220000 ;
        RECT 53.710000 13.460000 53.910000 13.660000 ;
        RECT 53.710000 13.900000 53.910000 14.100000 ;
        RECT 53.710000 14.340000 53.910000 14.540000 ;
        RECT 53.710000 14.780000 53.910000 14.980000 ;
        RECT 53.710000 15.220000 53.910000 15.420000 ;
        RECT 53.710000 15.660000 53.910000 15.860000 ;
        RECT 53.710000 16.100000 53.910000 16.300000 ;
        RECT 54.115000 13.020000 54.315000 13.220000 ;
        RECT 54.115000 13.460000 54.315000 13.660000 ;
        RECT 54.115000 13.900000 54.315000 14.100000 ;
        RECT 54.115000 14.340000 54.315000 14.540000 ;
        RECT 54.115000 14.780000 54.315000 14.980000 ;
        RECT 54.115000 15.220000 54.315000 15.420000 ;
        RECT 54.115000 15.660000 54.315000 15.860000 ;
        RECT 54.115000 16.100000 54.315000 16.300000 ;
        RECT 54.520000 13.020000 54.720000 13.220000 ;
        RECT 54.520000 13.460000 54.720000 13.660000 ;
        RECT 54.520000 13.900000 54.720000 14.100000 ;
        RECT 54.520000 14.340000 54.720000 14.540000 ;
        RECT 54.520000 14.780000 54.720000 14.980000 ;
        RECT 54.520000 15.220000 54.720000 15.420000 ;
        RECT 54.520000 15.660000 54.720000 15.860000 ;
        RECT 54.520000 16.100000 54.720000 16.300000 ;
        RECT 54.925000 13.020000 55.125000 13.220000 ;
        RECT 54.925000 13.460000 55.125000 13.660000 ;
        RECT 54.925000 13.900000 55.125000 14.100000 ;
        RECT 54.925000 14.340000 55.125000 14.540000 ;
        RECT 54.925000 14.780000 55.125000 14.980000 ;
        RECT 54.925000 15.220000 55.125000 15.420000 ;
        RECT 54.925000 15.660000 55.125000 15.860000 ;
        RECT 54.925000 16.100000 55.125000 16.300000 ;
        RECT 55.330000 13.020000 55.530000 13.220000 ;
        RECT 55.330000 13.460000 55.530000 13.660000 ;
        RECT 55.330000 13.900000 55.530000 14.100000 ;
        RECT 55.330000 14.340000 55.530000 14.540000 ;
        RECT 55.330000 14.780000 55.530000 14.980000 ;
        RECT 55.330000 15.220000 55.530000 15.420000 ;
        RECT 55.330000 15.660000 55.530000 15.860000 ;
        RECT 55.330000 16.100000 55.530000 16.300000 ;
        RECT 55.735000 13.020000 55.935000 13.220000 ;
        RECT 55.735000 13.460000 55.935000 13.660000 ;
        RECT 55.735000 13.900000 55.935000 14.100000 ;
        RECT 55.735000 14.340000 55.935000 14.540000 ;
        RECT 55.735000 14.780000 55.935000 14.980000 ;
        RECT 55.735000 15.220000 55.935000 15.420000 ;
        RECT 55.735000 15.660000 55.935000 15.860000 ;
        RECT 55.735000 16.100000 55.935000 16.300000 ;
        RECT 56.140000 13.020000 56.340000 13.220000 ;
        RECT 56.140000 13.460000 56.340000 13.660000 ;
        RECT 56.140000 13.900000 56.340000 14.100000 ;
        RECT 56.140000 14.340000 56.340000 14.540000 ;
        RECT 56.140000 14.780000 56.340000 14.980000 ;
        RECT 56.140000 15.220000 56.340000 15.420000 ;
        RECT 56.140000 15.660000 56.340000 15.860000 ;
        RECT 56.140000 16.100000 56.340000 16.300000 ;
        RECT 56.545000 13.020000 56.745000 13.220000 ;
        RECT 56.545000 13.460000 56.745000 13.660000 ;
        RECT 56.545000 13.900000 56.745000 14.100000 ;
        RECT 56.545000 14.340000 56.745000 14.540000 ;
        RECT 56.545000 14.780000 56.745000 14.980000 ;
        RECT 56.545000 15.220000 56.745000 15.420000 ;
        RECT 56.545000 15.660000 56.745000 15.860000 ;
        RECT 56.545000 16.100000 56.745000 16.300000 ;
        RECT 56.950000 13.020000 57.150000 13.220000 ;
        RECT 56.950000 13.460000 57.150000 13.660000 ;
        RECT 56.950000 13.900000 57.150000 14.100000 ;
        RECT 56.950000 14.340000 57.150000 14.540000 ;
        RECT 56.950000 14.780000 57.150000 14.980000 ;
        RECT 56.950000 15.220000 57.150000 15.420000 ;
        RECT 56.950000 15.660000 57.150000 15.860000 ;
        RECT 56.950000 16.100000 57.150000 16.300000 ;
        RECT 57.355000 13.020000 57.555000 13.220000 ;
        RECT 57.355000 13.460000 57.555000 13.660000 ;
        RECT 57.355000 13.900000 57.555000 14.100000 ;
        RECT 57.355000 14.340000 57.555000 14.540000 ;
        RECT 57.355000 14.780000 57.555000 14.980000 ;
        RECT 57.355000 15.220000 57.555000 15.420000 ;
        RECT 57.355000 15.660000 57.555000 15.860000 ;
        RECT 57.355000 16.100000 57.555000 16.300000 ;
        RECT 57.760000 13.020000 57.960000 13.220000 ;
        RECT 57.760000 13.460000 57.960000 13.660000 ;
        RECT 57.760000 13.900000 57.960000 14.100000 ;
        RECT 57.760000 14.340000 57.960000 14.540000 ;
        RECT 57.760000 14.780000 57.960000 14.980000 ;
        RECT 57.760000 15.220000 57.960000 15.420000 ;
        RECT 57.760000 15.660000 57.960000 15.860000 ;
        RECT 57.760000 16.100000 57.960000 16.300000 ;
        RECT 58.165000 13.020000 58.365000 13.220000 ;
        RECT 58.165000 13.460000 58.365000 13.660000 ;
        RECT 58.165000 13.900000 58.365000 14.100000 ;
        RECT 58.165000 14.340000 58.365000 14.540000 ;
        RECT 58.165000 14.780000 58.365000 14.980000 ;
        RECT 58.165000 15.220000 58.365000 15.420000 ;
        RECT 58.165000 15.660000 58.365000 15.860000 ;
        RECT 58.165000 16.100000 58.365000 16.300000 ;
        RECT 58.570000 13.020000 58.770000 13.220000 ;
        RECT 58.570000 13.460000 58.770000 13.660000 ;
        RECT 58.570000 13.900000 58.770000 14.100000 ;
        RECT 58.570000 14.340000 58.770000 14.540000 ;
        RECT 58.570000 14.780000 58.770000 14.980000 ;
        RECT 58.570000 15.220000 58.770000 15.420000 ;
        RECT 58.570000 15.660000 58.770000 15.860000 ;
        RECT 58.570000 16.100000 58.770000 16.300000 ;
        RECT 58.975000 13.020000 59.175000 13.220000 ;
        RECT 58.975000 13.460000 59.175000 13.660000 ;
        RECT 58.975000 13.900000 59.175000 14.100000 ;
        RECT 58.975000 14.340000 59.175000 14.540000 ;
        RECT 58.975000 14.780000 59.175000 14.980000 ;
        RECT 58.975000 15.220000 59.175000 15.420000 ;
        RECT 58.975000 15.660000 59.175000 15.860000 ;
        RECT 58.975000 16.100000 59.175000 16.300000 ;
        RECT 59.380000 13.020000 59.580000 13.220000 ;
        RECT 59.380000 13.460000 59.580000 13.660000 ;
        RECT 59.380000 13.900000 59.580000 14.100000 ;
        RECT 59.380000 14.340000 59.580000 14.540000 ;
        RECT 59.380000 14.780000 59.580000 14.980000 ;
        RECT 59.380000 15.220000 59.580000 15.420000 ;
        RECT 59.380000 15.660000 59.580000 15.860000 ;
        RECT 59.380000 16.100000 59.580000 16.300000 ;
        RECT 59.785000 13.020000 59.985000 13.220000 ;
        RECT 59.785000 13.460000 59.985000 13.660000 ;
        RECT 59.785000 13.900000 59.985000 14.100000 ;
        RECT 59.785000 14.340000 59.985000 14.540000 ;
        RECT 59.785000 14.780000 59.985000 14.980000 ;
        RECT 59.785000 15.220000 59.985000 15.420000 ;
        RECT 59.785000 15.660000 59.985000 15.860000 ;
        RECT 59.785000 16.100000 59.985000 16.300000 ;
        RECT 60.190000 13.020000 60.390000 13.220000 ;
        RECT 60.190000 13.460000 60.390000 13.660000 ;
        RECT 60.190000 13.900000 60.390000 14.100000 ;
        RECT 60.190000 14.340000 60.390000 14.540000 ;
        RECT 60.190000 14.780000 60.390000 14.980000 ;
        RECT 60.190000 15.220000 60.390000 15.420000 ;
        RECT 60.190000 15.660000 60.390000 15.860000 ;
        RECT 60.190000 16.100000 60.390000 16.300000 ;
        RECT 60.595000 13.020000 60.795000 13.220000 ;
        RECT 60.595000 13.460000 60.795000 13.660000 ;
        RECT 60.595000 13.900000 60.795000 14.100000 ;
        RECT 60.595000 14.340000 60.795000 14.540000 ;
        RECT 60.595000 14.780000 60.795000 14.980000 ;
        RECT 60.595000 15.220000 60.795000 15.420000 ;
        RECT 60.595000 15.660000 60.795000 15.860000 ;
        RECT 60.595000 16.100000 60.795000 16.300000 ;
        RECT 61.000000 13.020000 61.200000 13.220000 ;
        RECT 61.000000 13.460000 61.200000 13.660000 ;
        RECT 61.000000 13.900000 61.200000 14.100000 ;
        RECT 61.000000 14.340000 61.200000 14.540000 ;
        RECT 61.000000 14.780000 61.200000 14.980000 ;
        RECT 61.000000 15.220000 61.200000 15.420000 ;
        RECT 61.000000 15.660000 61.200000 15.860000 ;
        RECT 61.000000 16.100000 61.200000 16.300000 ;
        RECT 61.405000 13.020000 61.605000 13.220000 ;
        RECT 61.405000 13.460000 61.605000 13.660000 ;
        RECT 61.405000 13.900000 61.605000 14.100000 ;
        RECT 61.405000 14.340000 61.605000 14.540000 ;
        RECT 61.405000 14.780000 61.605000 14.980000 ;
        RECT 61.405000 15.220000 61.605000 15.420000 ;
        RECT 61.405000 15.660000 61.605000 15.860000 ;
        RECT 61.405000 16.100000 61.605000 16.300000 ;
        RECT 61.810000 13.020000 62.010000 13.220000 ;
        RECT 61.810000 13.460000 62.010000 13.660000 ;
        RECT 61.810000 13.900000 62.010000 14.100000 ;
        RECT 61.810000 14.340000 62.010000 14.540000 ;
        RECT 61.810000 14.780000 62.010000 14.980000 ;
        RECT 61.810000 15.220000 62.010000 15.420000 ;
        RECT 61.810000 15.660000 62.010000 15.860000 ;
        RECT 61.810000 16.100000 62.010000 16.300000 ;
        RECT 62.215000 13.020000 62.415000 13.220000 ;
        RECT 62.215000 13.460000 62.415000 13.660000 ;
        RECT 62.215000 13.900000 62.415000 14.100000 ;
        RECT 62.215000 14.340000 62.415000 14.540000 ;
        RECT 62.215000 14.780000 62.415000 14.980000 ;
        RECT 62.215000 15.220000 62.415000 15.420000 ;
        RECT 62.215000 15.660000 62.415000 15.860000 ;
        RECT 62.215000 16.100000 62.415000 16.300000 ;
        RECT 62.620000 13.020000 62.820000 13.220000 ;
        RECT 62.620000 13.460000 62.820000 13.660000 ;
        RECT 62.620000 13.900000 62.820000 14.100000 ;
        RECT 62.620000 14.340000 62.820000 14.540000 ;
        RECT 62.620000 14.780000 62.820000 14.980000 ;
        RECT 62.620000 15.220000 62.820000 15.420000 ;
        RECT 62.620000 15.660000 62.820000 15.860000 ;
        RECT 62.620000 16.100000 62.820000 16.300000 ;
        RECT 63.025000 13.020000 63.225000 13.220000 ;
        RECT 63.025000 13.460000 63.225000 13.660000 ;
        RECT 63.025000 13.900000 63.225000 14.100000 ;
        RECT 63.025000 14.340000 63.225000 14.540000 ;
        RECT 63.025000 14.780000 63.225000 14.980000 ;
        RECT 63.025000 15.220000 63.225000 15.420000 ;
        RECT 63.025000 15.660000 63.225000 15.860000 ;
        RECT 63.025000 16.100000 63.225000 16.300000 ;
        RECT 63.430000 13.020000 63.630000 13.220000 ;
        RECT 63.430000 13.460000 63.630000 13.660000 ;
        RECT 63.430000 13.900000 63.630000 14.100000 ;
        RECT 63.430000 14.340000 63.630000 14.540000 ;
        RECT 63.430000 14.780000 63.630000 14.980000 ;
        RECT 63.430000 15.220000 63.630000 15.420000 ;
        RECT 63.430000 15.660000 63.630000 15.860000 ;
        RECT 63.430000 16.100000 63.630000 16.300000 ;
        RECT 63.835000 13.020000 64.035000 13.220000 ;
        RECT 63.835000 13.460000 64.035000 13.660000 ;
        RECT 63.835000 13.900000 64.035000 14.100000 ;
        RECT 63.835000 14.340000 64.035000 14.540000 ;
        RECT 63.835000 14.780000 64.035000 14.980000 ;
        RECT 63.835000 15.220000 64.035000 15.420000 ;
        RECT 63.835000 15.660000 64.035000 15.860000 ;
        RECT 63.835000 16.100000 64.035000 16.300000 ;
        RECT 64.240000 13.020000 64.440000 13.220000 ;
        RECT 64.240000 13.460000 64.440000 13.660000 ;
        RECT 64.240000 13.900000 64.440000 14.100000 ;
        RECT 64.240000 14.340000 64.440000 14.540000 ;
        RECT 64.240000 14.780000 64.440000 14.980000 ;
        RECT 64.240000 15.220000 64.440000 15.420000 ;
        RECT 64.240000 15.660000 64.440000 15.860000 ;
        RECT 64.240000 16.100000 64.440000 16.300000 ;
        RECT 64.645000 13.020000 64.845000 13.220000 ;
        RECT 64.645000 13.460000 64.845000 13.660000 ;
        RECT 64.645000 13.900000 64.845000 14.100000 ;
        RECT 64.645000 14.340000 64.845000 14.540000 ;
        RECT 64.645000 14.780000 64.845000 14.980000 ;
        RECT 64.645000 15.220000 64.845000 15.420000 ;
        RECT 64.645000 15.660000 64.845000 15.860000 ;
        RECT 64.645000 16.100000 64.845000 16.300000 ;
        RECT 65.050000 13.020000 65.250000 13.220000 ;
        RECT 65.050000 13.460000 65.250000 13.660000 ;
        RECT 65.050000 13.900000 65.250000 14.100000 ;
        RECT 65.050000 14.340000 65.250000 14.540000 ;
        RECT 65.050000 14.780000 65.250000 14.980000 ;
        RECT 65.050000 15.220000 65.250000 15.420000 ;
        RECT 65.050000 15.660000 65.250000 15.860000 ;
        RECT 65.050000 16.100000 65.250000 16.300000 ;
        RECT 65.455000 13.020000 65.655000 13.220000 ;
        RECT 65.455000 13.460000 65.655000 13.660000 ;
        RECT 65.455000 13.900000 65.655000 14.100000 ;
        RECT 65.455000 14.340000 65.655000 14.540000 ;
        RECT 65.455000 14.780000 65.655000 14.980000 ;
        RECT 65.455000 15.220000 65.655000 15.420000 ;
        RECT 65.455000 15.660000 65.655000 15.860000 ;
        RECT 65.455000 16.100000 65.655000 16.300000 ;
        RECT 65.860000 13.020000 66.060000 13.220000 ;
        RECT 65.860000 13.460000 66.060000 13.660000 ;
        RECT 65.860000 13.900000 66.060000 14.100000 ;
        RECT 65.860000 14.340000 66.060000 14.540000 ;
        RECT 65.860000 14.780000 66.060000 14.980000 ;
        RECT 65.860000 15.220000 66.060000 15.420000 ;
        RECT 65.860000 15.660000 66.060000 15.860000 ;
        RECT 65.860000 16.100000 66.060000 16.300000 ;
        RECT 66.265000 13.020000 66.465000 13.220000 ;
        RECT 66.265000 13.460000 66.465000 13.660000 ;
        RECT 66.265000 13.900000 66.465000 14.100000 ;
        RECT 66.265000 14.340000 66.465000 14.540000 ;
        RECT 66.265000 14.780000 66.465000 14.980000 ;
        RECT 66.265000 15.220000 66.465000 15.420000 ;
        RECT 66.265000 15.660000 66.465000 15.860000 ;
        RECT 66.265000 16.100000 66.465000 16.300000 ;
        RECT 66.670000 13.020000 66.870000 13.220000 ;
        RECT 66.670000 13.460000 66.870000 13.660000 ;
        RECT 66.670000 13.900000 66.870000 14.100000 ;
        RECT 66.670000 14.340000 66.870000 14.540000 ;
        RECT 66.670000 14.780000 66.870000 14.980000 ;
        RECT 66.670000 15.220000 66.870000 15.420000 ;
        RECT 66.670000 15.660000 66.870000 15.860000 ;
        RECT 66.670000 16.100000 66.870000 16.300000 ;
        RECT 67.075000 13.020000 67.275000 13.220000 ;
        RECT 67.075000 13.460000 67.275000 13.660000 ;
        RECT 67.075000 13.900000 67.275000 14.100000 ;
        RECT 67.075000 14.340000 67.275000 14.540000 ;
        RECT 67.075000 14.780000 67.275000 14.980000 ;
        RECT 67.075000 15.220000 67.275000 15.420000 ;
        RECT 67.075000 15.660000 67.275000 15.860000 ;
        RECT 67.075000 16.100000 67.275000 16.300000 ;
        RECT 67.480000 13.020000 67.680000 13.220000 ;
        RECT 67.480000 13.460000 67.680000 13.660000 ;
        RECT 67.480000 13.900000 67.680000 14.100000 ;
        RECT 67.480000 14.340000 67.680000 14.540000 ;
        RECT 67.480000 14.780000 67.680000 14.980000 ;
        RECT 67.480000 15.220000 67.680000 15.420000 ;
        RECT 67.480000 15.660000 67.680000 15.860000 ;
        RECT 67.480000 16.100000 67.680000 16.300000 ;
        RECT 67.885000 13.020000 68.085000 13.220000 ;
        RECT 67.885000 13.460000 68.085000 13.660000 ;
        RECT 67.885000 13.900000 68.085000 14.100000 ;
        RECT 67.885000 14.340000 68.085000 14.540000 ;
        RECT 67.885000 14.780000 68.085000 14.980000 ;
        RECT 67.885000 15.220000 68.085000 15.420000 ;
        RECT 67.885000 15.660000 68.085000 15.860000 ;
        RECT 67.885000 16.100000 68.085000 16.300000 ;
        RECT 68.290000 13.020000 68.490000 13.220000 ;
        RECT 68.290000 13.460000 68.490000 13.660000 ;
        RECT 68.290000 13.900000 68.490000 14.100000 ;
        RECT 68.290000 14.340000 68.490000 14.540000 ;
        RECT 68.290000 14.780000 68.490000 14.980000 ;
        RECT 68.290000 15.220000 68.490000 15.420000 ;
        RECT 68.290000 15.660000 68.490000 15.860000 ;
        RECT 68.290000 16.100000 68.490000 16.300000 ;
        RECT 68.695000 13.020000 68.895000 13.220000 ;
        RECT 68.695000 13.460000 68.895000 13.660000 ;
        RECT 68.695000 13.900000 68.895000 14.100000 ;
        RECT 68.695000 14.340000 68.895000 14.540000 ;
        RECT 68.695000 14.780000 68.895000 14.980000 ;
        RECT 68.695000 15.220000 68.895000 15.420000 ;
        RECT 68.695000 15.660000 68.895000 15.860000 ;
        RECT 68.695000 16.100000 68.895000 16.300000 ;
        RECT 69.100000 13.020000 69.300000 13.220000 ;
        RECT 69.100000 13.460000 69.300000 13.660000 ;
        RECT 69.100000 13.900000 69.300000 14.100000 ;
        RECT 69.100000 14.340000 69.300000 14.540000 ;
        RECT 69.100000 14.780000 69.300000 14.980000 ;
        RECT 69.100000 15.220000 69.300000 15.420000 ;
        RECT 69.100000 15.660000 69.300000 15.860000 ;
        RECT 69.100000 16.100000 69.300000 16.300000 ;
        RECT 69.505000 13.020000 69.705000 13.220000 ;
        RECT 69.505000 13.460000 69.705000 13.660000 ;
        RECT 69.505000 13.900000 69.705000 14.100000 ;
        RECT 69.505000 14.340000 69.705000 14.540000 ;
        RECT 69.505000 14.780000 69.705000 14.980000 ;
        RECT 69.505000 15.220000 69.705000 15.420000 ;
        RECT 69.505000 15.660000 69.705000 15.860000 ;
        RECT 69.505000 16.100000 69.705000 16.300000 ;
        RECT 69.910000 13.020000 70.110000 13.220000 ;
        RECT 69.910000 13.460000 70.110000 13.660000 ;
        RECT 69.910000 13.900000 70.110000 14.100000 ;
        RECT 69.910000 14.340000 70.110000 14.540000 ;
        RECT 69.910000 14.780000 70.110000 14.980000 ;
        RECT 69.910000 15.220000 70.110000 15.420000 ;
        RECT 69.910000 15.660000 70.110000 15.860000 ;
        RECT 69.910000 16.100000 70.110000 16.300000 ;
        RECT 70.315000 13.020000 70.515000 13.220000 ;
        RECT 70.315000 13.460000 70.515000 13.660000 ;
        RECT 70.315000 13.900000 70.515000 14.100000 ;
        RECT 70.315000 14.340000 70.515000 14.540000 ;
        RECT 70.315000 14.780000 70.515000 14.980000 ;
        RECT 70.315000 15.220000 70.515000 15.420000 ;
        RECT 70.315000 15.660000 70.515000 15.860000 ;
        RECT 70.315000 16.100000 70.515000 16.300000 ;
        RECT 70.720000 13.020000 70.920000 13.220000 ;
        RECT 70.720000 13.460000 70.920000 13.660000 ;
        RECT 70.720000 13.900000 70.920000 14.100000 ;
        RECT 70.720000 14.340000 70.920000 14.540000 ;
        RECT 70.720000 14.780000 70.920000 14.980000 ;
        RECT 70.720000 15.220000 70.920000 15.420000 ;
        RECT 70.720000 15.660000 70.920000 15.860000 ;
        RECT 70.720000 16.100000 70.920000 16.300000 ;
        RECT 71.125000 13.020000 71.325000 13.220000 ;
        RECT 71.125000 13.460000 71.325000 13.660000 ;
        RECT 71.125000 13.900000 71.325000 14.100000 ;
        RECT 71.125000 14.340000 71.325000 14.540000 ;
        RECT 71.125000 14.780000 71.325000 14.980000 ;
        RECT 71.125000 15.220000 71.325000 15.420000 ;
        RECT 71.125000 15.660000 71.325000 15.860000 ;
        RECT 71.125000 16.100000 71.325000 16.300000 ;
        RECT 71.530000 13.020000 71.730000 13.220000 ;
        RECT 71.530000 13.460000 71.730000 13.660000 ;
        RECT 71.530000 13.900000 71.730000 14.100000 ;
        RECT 71.530000 14.340000 71.730000 14.540000 ;
        RECT 71.530000 14.780000 71.730000 14.980000 ;
        RECT 71.530000 15.220000 71.730000 15.420000 ;
        RECT 71.530000 15.660000 71.730000 15.860000 ;
        RECT 71.530000 16.100000 71.730000 16.300000 ;
        RECT 71.935000 13.020000 72.135000 13.220000 ;
        RECT 71.935000 13.460000 72.135000 13.660000 ;
        RECT 71.935000 13.900000 72.135000 14.100000 ;
        RECT 71.935000 14.340000 72.135000 14.540000 ;
        RECT 71.935000 14.780000 72.135000 14.980000 ;
        RECT 71.935000 15.220000 72.135000 15.420000 ;
        RECT 71.935000 15.660000 72.135000 15.860000 ;
        RECT 71.935000 16.100000 72.135000 16.300000 ;
        RECT 72.340000 13.020000 72.540000 13.220000 ;
        RECT 72.340000 13.460000 72.540000 13.660000 ;
        RECT 72.340000 13.900000 72.540000 14.100000 ;
        RECT 72.340000 14.340000 72.540000 14.540000 ;
        RECT 72.340000 14.780000 72.540000 14.980000 ;
        RECT 72.340000 15.220000 72.540000 15.420000 ;
        RECT 72.340000 15.660000 72.540000 15.860000 ;
        RECT 72.340000 16.100000 72.540000 16.300000 ;
        RECT 72.745000 13.020000 72.945000 13.220000 ;
        RECT 72.745000 13.460000 72.945000 13.660000 ;
        RECT 72.745000 13.900000 72.945000 14.100000 ;
        RECT 72.745000 14.340000 72.945000 14.540000 ;
        RECT 72.745000 14.780000 72.945000 14.980000 ;
        RECT 72.745000 15.220000 72.945000 15.420000 ;
        RECT 72.745000 15.660000 72.945000 15.860000 ;
        RECT 72.745000 16.100000 72.945000 16.300000 ;
        RECT 73.150000 13.020000 73.350000 13.220000 ;
        RECT 73.150000 13.460000 73.350000 13.660000 ;
        RECT 73.150000 13.900000 73.350000 14.100000 ;
        RECT 73.150000 14.340000 73.350000 14.540000 ;
        RECT 73.150000 14.780000 73.350000 14.980000 ;
        RECT 73.150000 15.220000 73.350000 15.420000 ;
        RECT 73.150000 15.660000 73.350000 15.860000 ;
        RECT 73.150000 16.100000 73.350000 16.300000 ;
        RECT 73.555000 13.020000 73.755000 13.220000 ;
        RECT 73.555000 13.460000 73.755000 13.660000 ;
        RECT 73.555000 13.900000 73.755000 14.100000 ;
        RECT 73.555000 14.340000 73.755000 14.540000 ;
        RECT 73.555000 14.780000 73.755000 14.980000 ;
        RECT 73.555000 15.220000 73.755000 15.420000 ;
        RECT 73.555000 15.660000 73.755000 15.860000 ;
        RECT 73.555000 16.100000 73.755000 16.300000 ;
        RECT 73.960000 13.020000 74.160000 13.220000 ;
        RECT 73.960000 13.460000 74.160000 13.660000 ;
        RECT 73.960000 13.900000 74.160000 14.100000 ;
        RECT 73.960000 14.340000 74.160000 14.540000 ;
        RECT 73.960000 14.780000 74.160000 14.980000 ;
        RECT 73.960000 15.220000 74.160000 15.420000 ;
        RECT 73.960000 15.660000 74.160000 15.860000 ;
        RECT 73.960000 16.100000 74.160000 16.300000 ;
        RECT 74.365000 13.020000 74.565000 13.220000 ;
        RECT 74.365000 13.460000 74.565000 13.660000 ;
        RECT 74.365000 13.900000 74.565000 14.100000 ;
        RECT 74.365000 14.340000 74.565000 14.540000 ;
        RECT 74.365000 14.780000 74.565000 14.980000 ;
        RECT 74.365000 15.220000 74.565000 15.420000 ;
        RECT 74.365000 15.660000 74.565000 15.860000 ;
        RECT 74.365000 16.100000 74.565000 16.300000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 17.785000 1.270000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 68.035000 1.270000 93.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 17.785000 75.000000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 68.035000 75.000000 93.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 17.885000 1.270000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 68.035000 1.270000 92.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 17.885000 75.000000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 62.085000 1.270000 66.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 62.085000 75.000000 66.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 62.185000 1.270000 66.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 34.735000 1.270000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 45.735000 1.270000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 49.645000 1.270000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 54.405000 1.270000 54.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 34.735000 75.000000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 45.735000 75.000000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 49.645000 75.000000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 54.405000 75.000000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 34.840000 1.270000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 45.735000 1.270000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 34.840000 75.000000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 39.585000 1.270000 44.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 39.585000 75.000000 44.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 39.685000 1.270000 44.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 23.835000 1.270000 28.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 23.835000 75.000000 28.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 23.935000 1.270000 28.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 56.235000 1.270000 60.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.235000 75.000000 60.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 56.335000 1.270000 60.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 29.885000 1.270000 33.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 29.885000 75.000000 33.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 29.985000 1.270000 33.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 198.000000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 75.000000 198.000000 ;
    LAYER met3 ;
      RECT  0.000000  0.000000 75.000000  12.540000 ;
      RECT  0.000000 16.780000 75.000000 198.000000 ;
      RECT 24.900000 12.540000 50.355000  16.780000 ;
    LAYER met4 ;
      RECT  0.000000   5.885000  1.670000   6.485000 ;
      RECT  0.000000  11.935000  1.670000  12.535000 ;
      RECT  0.000000  16.785000  1.670000  17.385000 ;
      RECT  0.000000  22.835000  1.670000  23.435000 ;
      RECT  0.000000  28.885000  1.670000  29.485000 ;
      RECT  0.000000  33.735000  1.670000  34.335000 ;
      RECT  0.000000  38.585000  1.670000  39.185000 ;
      RECT  0.000000  44.635000  1.670000  45.335000 ;
      RECT  0.000000  55.135000  1.670000  55.835000 ;
      RECT  0.000000  61.085000  1.670000  61.685000 ;
      RECT  0.000000  66.935000  1.670000  67.635000 ;
      RECT  0.000000  93.400000 75.000000 173.385000 ;
      RECT  1.670000   0.000000 73.330000  12.535000 ;
      RECT  1.670000  16.785000 73.330000  93.400000 ;
      RECT  1.670000 173.385000 73.330000 198.000000 ;
      RECT 24.875000  12.535000 50.380000  16.785000 ;
      RECT 73.330000   5.885000 75.000000   6.485000 ;
      RECT 73.330000  11.935000 75.000000  12.535000 ;
      RECT 73.330000  16.785000 75.000000  17.385000 ;
      RECT 73.330000  22.835000 75.000000  23.435000 ;
      RECT 73.330000  28.885000 75.000000  29.485000 ;
      RECT 73.330000  33.735000 75.000000  34.335000 ;
      RECT 73.330000  38.585000 75.000000  39.185000 ;
      RECT 73.330000  44.635000 75.000000  45.335000 ;
      RECT 73.330000  55.135000 75.000000  55.835000 ;
      RECT 73.330000  61.085000 75.000000  61.685000 ;
      RECT 73.330000  66.935000 75.000000  67.635000 ;
    LAYER met5 ;
      RECT 0.000000  93.785000 75.000000 172.985000 ;
      RECT 1.765000  12.235000 73.235000  17.085000 ;
      RECT 2.070000   0.000000 72.930000  12.235000 ;
      RECT 2.070000  17.085000 72.930000  93.785000 ;
      RECT 2.070000 172.985000 72.930000 198.000000 ;
  END
END sky130_fd_io__overlay_vdda_lvc
END LIBRARY
