# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sky130_fd_io__top_hvclamp
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 75 BY 200 ;
  SYMMETRY R90 ;

  PIN ogc_hvc
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 25.895 0 27.895 1.92 ;
    END
  END ogc_hvc

  PIN src_bdy_hvc
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 25.895 0 36.895 90.39 ;
        RECT 25.895 90.39 36.895 90.54 ;
        RECT 25.745 90.54 36.895 90.69 ;
        RECT 25.595 90.69 36.895 90.84 ;
        RECT 25.445 90.84 36.895 90.99 ;
        RECT 25.295 90.99 36.895 91.14 ;
        RECT 25.145 91.14 36.895 91.29 ;
        RECT 24.995 91.29 36.895 91.44 ;
        RECT 24.845 91.44 36.895 91.59 ;
        RECT 24.695 91.59 36.895 91.74 ;
        RECT 24.545 91.74 36.895 91.89 ;
        RECT 24.395 91.89 36.895 92.04 ;
        RECT 24.245 92.04 36.895 92.19 ;
        RECT 24.095 92.19 36.895 92.34 ;
        RECT 23.945 92.34 36.895 92.39 ;
        RECT 31.385 92.39 36.895 92.54 ;
        RECT 31.535 92.54 36.895 92.69 ;
        RECT 31.685 92.69 36.895 92.84 ;
        RECT 31.835 92.84 36.895 92.99 ;
        RECT 31.945 92.99 36.895 93.1 ;
        RECT 23.895 92.39 30.16 92.465 ;
        RECT 23.82 92.465 30.085 92.54 ;
        RECT 31.945 93.1 36.895 96.375 ;
        RECT 23.745 92.54 29.935 92.69 ;
        RECT 23.745 92.69 29.785 92.84 ;
        RECT 23.745 92.84 29.635 92.99 ;
        RECT 23.745 92.99 29.525 93.1 ;
        RECT 31.945 96.375 36.895 96.525 ;
        RECT 31.795 96.525 36.895 96.675 ;
        RECT 31.645 96.675 36.895 96.825 ;
        RECT 31.495 96.825 36.895 96.975 ;
        RECT 31.345 96.975 36.895 97.125 ;
        RECT 31.195 97.125 36.895 97.275 ;
        RECT 31.045 97.275 36.895 97.425 ;
        RECT 30.895 97.425 36.895 97.575 ;
        RECT 30.745 97.575 36.895 97.725 ;
        RECT 30.595 97.725 36.895 97.875 ;
        RECT 30.445 97.875 36.895 98.025 ;
        RECT 30.295 98.025 36.895 98.175 ;
        RECT 30.145 98.175 36.895 98.325 ;
        RECT 29.995 98.325 36.895 98.475 ;
        RECT 29.845 98.475 36.895 98.625 ;
        RECT 29.695 98.625 36.895 98.775 ;
        RECT 29.545 98.775 36.895 98.925 ;
        RECT 29.395 98.925 36.895 99.075 ;
        RECT 29.245 99.075 36.895 99.225 ;
        RECT 29.095 99.225 36.895 99.375 ;
        RECT 28.945 99.375 36.895 99.525 ;
        RECT 28.795 99.525 36.895 99.675 ;
        RECT 28.645 99.675 36.895 99.825 ;
        RECT 28.495 99.825 36.895 99.895 ;
        RECT 23.745 93.1 29.525 93.955 ;
        RECT 28.425 99.895 36.745 100.045 ;
        RECT 28.275 100.045 36.595 100.195 ;
        RECT 28.125 100.195 36.445 100.345 ;
        RECT 27.975 100.345 36.295 100.495 ;
        RECT 27.825 100.495 36.145 100.645 ;
        RECT 27.675 100.645 35.995 100.795 ;
        RECT 27.525 100.795 35.845 100.945 ;
        RECT 27.375 100.945 35.695 101.095 ;
        RECT 27.225 101.095 35.545 101.245 ;
        RECT 27.075 101.245 35.395 101.395 ;
        RECT 26.925 101.395 35.245 101.545 ;
        RECT 26.775 101.545 35.095 101.695 ;
        RECT 26.625 101.695 34.945 101.845 ;
        RECT 26.475 101.845 34.795 101.995 ;
        RECT 26.325 101.995 34.645 102.145 ;
        RECT 26.175 102.145 34.495 102.295 ;
        RECT 26.025 102.295 34.4 102.39 ;
        RECT 23.745 93.955 29.525 94.105 ;
        RECT 23.595 94.105 29.525 94.255 ;
        RECT 23.445 94.255 29.525 94.405 ;
        RECT 23.295 94.405 29.525 94.555 ;
        RECT 23.145 94.555 29.525 94.705 ;
        RECT 22.995 94.705 29.525 94.855 ;
        RECT 22.845 94.855 29.525 95.005 ;
        RECT 22.695 95.005 29.525 95.155 ;
        RECT 22.545 95.155 29.525 95.305 ;
        RECT 22.395 95.305 29.525 95.455 ;
        RECT 22.245 95.455 29.525 95.605 ;
        RECT 22.095 95.605 29.525 95.755 ;
        RECT 21.945 95.755 29.525 95.905 ;
        RECT 21.795 95.905 29.525 96.055 ;
        RECT 21.645 96.055 29.525 96.205 ;
        RECT 21.495 96.205 29.525 96.355 ;
        RECT 21.345 96.355 29.525 96.505 ;
        RECT 21.195 96.505 29.525 96.655 ;
        RECT 25.93 102.39 34.25 102.54 ;
        RECT 25.93 102.54 34.1 102.69 ;
        RECT 25.93 102.69 33.95 102.84 ;
        RECT 25.93 102.84 33.8 102.99 ;
        RECT 25.93 102.99 33.65 103.14 ;
        RECT 25.93 103.14 33.5 103.29 ;
        RECT 25.93 103.29 33.35 103.44 ;
        RECT 25.93 103.44 33.2 103.59 ;
        RECT 25.93 103.59 33.05 103.74 ;
        RECT 25.93 103.74 32.9 103.89 ;
        RECT 25.93 103.89 32.75 104.04 ;
        RECT 25.93 104.04 32.6 104.19 ;
        RECT 25.93 104.19 32.45 104.34 ;
        RECT 25.93 104.34 32.3 104.49 ;
        RECT 25.93 104.49 32.15 104.64 ;
        RECT 25.93 104.64 32 104.79 ;
        RECT 25.93 104.79 31.93 104.86 ;
        RECT 21.045 96.655 29.375 96.805 ;
        RECT 20.895 96.805 29.225 96.955 ;
        RECT 20.745 96.955 29.075 97.105 ;
        RECT 20.595 97.105 28.925 97.255 ;
        RECT 20.445 97.255 28.775 97.405 ;
        RECT 20.295 97.405 28.625 97.555 ;
        RECT 20.145 97.555 28.475 97.705 ;
        RECT 19.995 97.705 28.325 97.855 ;
        RECT 19.845 97.855 28.175 98.005 ;
        RECT 19.695 98.005 28.025 98.155 ;
        RECT 19.545 98.155 27.875 98.305 ;
        RECT 19.395 98.305 27.725 98.455 ;
        RECT 19.245 98.455 27.575 98.605 ;
        RECT 19.095 98.605 27.425 98.755 ;
        RECT 18.945 98.755 27.275 98.905 ;
        RECT 18.795 98.905 27.125 99.055 ;
        RECT 18.645 99.055 26.975 99.205 ;
        RECT 18.495 99.205 26.825 99.355 ;
        RECT 18.345 99.355 26.675 99.505 ;
        RECT 18.195 99.505 26.525 99.655 ;
        RECT 18.045 99.655 26.375 99.805 ;
        RECT 17.895 99.805 26.225 99.955 ;
        RECT 17.745 99.955 26.075 100.105 ;
        RECT 17.595 100.105 25.925 100.255 ;
        RECT 17.445 100.255 25.775 100.405 ;
        RECT 17.295 100.405 25.625 100.555 ;
        RECT 17.145 100.555 25.475 100.705 ;
        RECT 16.995 100.705 25.325 100.855 ;
        RECT 16.845 100.855 25.175 101.005 ;
        RECT 16.695 101.005 25.025 101.155 ;
        RECT 16.545 101.155 24.875 101.305 ;
        RECT 16.395 101.305 24.725 101.455 ;
        RECT 16.245 101.455 24.575 101.605 ;
        RECT 16.095 101.605 24.425 101.755 ;
        RECT 15.945 101.755 24.275 101.905 ;
        RECT 15.795 101.905 24.125 102.055 ;
        RECT 15.645 102.055 23.98 102.2 ;
        RECT 25.93 104.86 31.93 170.46 ;
        RECT 15.5 102.2 23.83 102.35 ;
        RECT 15.5 102.35 23.68 102.5 ;
        RECT 15.5 102.5 23.53 102.65 ;
        RECT 15.5 102.65 23.38 102.8 ;
        RECT 15.5 102.8 23.23 102.95 ;
        RECT 15.5 102.95 23.08 103.1 ;
        RECT 15.5 103.1 22.93 103.25 ;
        RECT 15.5 103.25 22.78 103.4 ;
        RECT 15.5 103.4 22.63 103.55 ;
        RECT 15.5 103.55 22.48 103.7 ;
        RECT 15.5 103.7 22.33 103.85 ;
        RECT 15.5 103.85 22.18 104 ;
        RECT 15.5 104 22.03 104.15 ;
        RECT 15.5 104.15 21.88 104.3 ;
        RECT 15.5 104.3 21.73 104.45 ;
        RECT 15.5 104.45 21.58 104.6 ;
        RECT 15.5 104.6 21.5 104.68 ;
        RECT 25.93 170.46 31.93 170.61 ;
        RECT 25.93 170.61 32.08 170.76 ;
        RECT 25.93 170.76 32.23 170.91 ;
        RECT 25.93 170.91 32.38 171.06 ;
        RECT 25.93 171.06 32.53 171.21 ;
        RECT 25.93 171.21 32.68 171.36 ;
        RECT 25.93 171.36 32.83 171.51 ;
        RECT 25.93 171.51 32.98 171.66 ;
        RECT 25.93 171.66 33.13 171.81 ;
        RECT 25.93 171.81 33.28 171.96 ;
        RECT 25.93 171.96 33.43 172.11 ;
        RECT 25.93 172.11 33.58 172.26 ;
        RECT 25.93 172.26 33.73 172.41 ;
        RECT 25.93 172.41 33.88 172.56 ;
        RECT 25.93 172.56 34.03 172.71 ;
        RECT 25.93 172.71 34.18 172.86 ;
        RECT 25.93 172.86 34.33 173.01 ;
        RECT 25.93 173.01 34.48 173.16 ;
        RECT 25.93 173.16 34.63 173.31 ;
        RECT 25.93 173.31 34.78 173.46 ;
        RECT 25.93 173.46 34.93 173.61 ;
        RECT 25.93 173.61 35.08 173.76 ;
        RECT 25.93 173.76 35.23 173.91 ;
        RECT 25.93 173.91 35.38 174.06 ;
        RECT 25.93 174.06 35.53 174.21 ;
        RECT 25.93 174.21 35.68 174.36 ;
        RECT 25.93 174.36 35.83 174.51 ;
        RECT 25.93 174.51 35.98 174.66 ;
        RECT 25.93 174.66 36.13 174.81 ;
        RECT 25.93 174.81 36.28 174.96 ;
        RECT 25.93 174.96 36.43 175.11 ;
        RECT 25.93 175.11 36.58 175.26 ;
        RECT 25.93 175.26 36.73 175.35 ;
        RECT 15.5 104.68 21.5 169.13 ;
        RECT 25.93 175.35 36.82 195.075 ;
        RECT 15.5 169.13 21.5 169.28 ;
        RECT 15.5 169.28 21.65 169.43 ;
        RECT 15.5 169.43 21.8 169.58 ;
        RECT 15.5 169.58 21.95 169.73 ;
        RECT 15.5 169.73 22.1 169.88 ;
        RECT 15.5 169.88 22.25 170.03 ;
        RECT 15.5 170.03 22.4 170.18 ;
        RECT 15.5 170.18 22.55 170.33 ;
        RECT 15.5 170.33 22.7 170.48 ;
        RECT 15.5 170.48 22.85 170.63 ;
        RECT 15.5 170.63 23 170.78 ;
        RECT 15.5 170.78 23.15 170.93 ;
        RECT 15.5 170.93 23.3 171.08 ;
        RECT 15.5 171.08 23.45 171.23 ;
        RECT 15.5 171.23 23.6 171.38 ;
        RECT 15.5 171.38 23.75 171.53 ;
        RECT 15.5 171.53 23.9 171.68 ;
        RECT 15.5 171.68 24.05 171.83 ;
        RECT 15.5 171.83 24.2 171.98 ;
        RECT 15.5 171.98 24.35 172.13 ;
        RECT 15.5 172.13 24.5 172.28 ;
        RECT 15.5 172.28 24.65 172.43 ;
        RECT 15.5 172.43 24.8 172.58 ;
        RECT 15.5 172.58 24.95 172.64 ;
        RECT 15.5 173.02 25.01 173.17 ;
        RECT 15.35 173.17 25.01 173.32 ;
        RECT 15.2 173.32 25.01 173.47 ;
        RECT 15.05 173.47 25.01 173.62 ;
        RECT 14.9 173.62 25.01 173.77 ;
        RECT 14.75 173.77 25.01 173.92 ;
        RECT 14.6 173.92 25.01 174.07 ;
        RECT 14.45 174.07 25.01 174.22 ;
        RECT 14.3 174.22 25.01 174.37 ;
        RECT 14.15 174.37 25.01 174.52 ;
        RECT 14 174.52 25.01 174.67 ;
        RECT 13.85 174.67 25.01 174.82 ;
        RECT 13.7 174.82 25.01 174.97 ;
        RECT 13.55 174.97 25.01 175.12 ;
        RECT 13.4 175.12 25.01 175.27 ;
        RECT 13.25 175.27 25.01 175.42 ;
        RECT 13.1 175.42 25.01 175.57 ;
        RECT 12.95 175.57 25.01 175.72 ;
        RECT 12.8 175.72 25.01 175.87 ;
        RECT 12.65 175.87 25.01 175.895 ;
        RECT 12.625 175.895 25.01 195.075 ;
        RECT 15.5 172.64 25.01 173.02 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.935 190.56 67.2 195.075 ;
        RECT 0.935 189.585 14.12 189.655 ;
        RECT 0.935 189.655 14.19 189.725 ;
        RECT 0.935 189.725 14.26 189.795 ;
        RECT 0.935 189.795 14.33 189.865 ;
        RECT 0.935 189.865 14.4 189.935 ;
        RECT 0.935 189.935 14.47 190.005 ;
        RECT 0.935 190.005 14.54 190.075 ;
        RECT 0.935 190.075 14.61 190.145 ;
        RECT 0.935 190.145 14.68 190.215 ;
        RECT 0.935 190.215 14.75 190.285 ;
        RECT 0.935 190.285 14.82 190.355 ;
        RECT 0.935 190.355 14.89 190.425 ;
        RECT 0.935 190.425 14.96 190.495 ;
        RECT 0.935 190.495 15.03 190.56 ;
        RECT 0.935 185.055 14.12 189.585 ;
        RECT 0.935 183.905 15.2 183.975 ;
        RECT 0.935 183.975 15.13 184.045 ;
        RECT 0.935 184.045 15.06 184.115 ;
        RECT 0.935 184.115 14.99 184.185 ;
        RECT 0.935 184.185 14.92 184.255 ;
        RECT 0.935 184.255 14.85 184.325 ;
        RECT 0.935 184.325 14.78 184.395 ;
        RECT 0.935 184.395 14.71 184.465 ;
        RECT 0.935 184.465 14.64 184.535 ;
        RECT 0.935 184.535 14.57 184.605 ;
        RECT 0.935 184.605 14.5 184.675 ;
        RECT 0.935 184.675 14.43 184.745 ;
        RECT 0.935 184.745 14.36 184.815 ;
        RECT 0.935 184.815 14.29 184.885 ;
        RECT 0.935 184.885 14.22 184.955 ;
        RECT 0.935 184.955 14.15 185.025 ;
        RECT 0.935 185.025 14.12 185.055 ;
        RECT 0.935 183.855 15.32 183.905 ;
        RECT 0.935 181.48 17.625 181.55 ;
        RECT 0.935 181.55 17.555 181.62 ;
        RECT 0.935 181.62 17.485 181.69 ;
        RECT 0.935 181.69 17.415 181.76 ;
        RECT 0.935 181.76 17.345 181.83 ;
        RECT 0.935 181.83 17.275 181.9 ;
        RECT 0.935 181.9 17.205 181.97 ;
        RECT 0.935 181.97 17.135 182.04 ;
        RECT 0.935 182.04 17.065 182.11 ;
        RECT 0.935 182.11 16.995 182.18 ;
        RECT 0.935 182.18 16.925 182.25 ;
        RECT 0.935 182.25 16.855 182.32 ;
        RECT 0.935 182.32 16.785 182.39 ;
        RECT 0.935 182.39 16.715 182.46 ;
        RECT 0.935 182.46 16.645 182.53 ;
        RECT 0.935 182.53 16.575 182.6 ;
        RECT 0.935 182.6 16.505 182.67 ;
        RECT 0.935 182.67 16.435 182.74 ;
        RECT 0.935 182.74 16.365 182.81 ;
        RECT 0.935 182.81 16.295 182.88 ;
        RECT 0.935 182.88 16.225 182.95 ;
        RECT 0.935 182.95 16.155 183.02 ;
        RECT 0.935 183.02 16.085 183.09 ;
        RECT 0.935 183.09 16.015 183.16 ;
        RECT 0.935 183.16 15.945 183.23 ;
        RECT 0.935 183.23 15.875 183.3 ;
        RECT 0.935 183.3 15.805 183.37 ;
        RECT 0.935 183.37 15.735 183.44 ;
        RECT 0.935 183.44 15.665 183.51 ;
        RECT 0.935 183.51 15.595 183.58 ;
        RECT 0.935 183.58 15.525 183.65 ;
        RECT 0.935 183.65 15.455 183.72 ;
        RECT 0.935 183.72 15.385 183.79 ;
        RECT 0.935 183.79 15.32 183.855 ;
        RECT 0.935 172.78 57.96 181.48 ;
        RECT 0.935 169.22 14.12 169.29 ;
        RECT 0.935 169.29 14.19 169.36 ;
        RECT 0.935 169.36 14.26 169.43 ;
        RECT 0.935 169.43 14.33 169.5 ;
        RECT 0.935 169.5 14.4 169.57 ;
        RECT 0.935 169.57 14.47 169.64 ;
        RECT 0.935 169.64 14.54 169.71 ;
        RECT 0.935 169.71 14.61 169.78 ;
        RECT 0.935 169.78 14.68 169.85 ;
        RECT 0.935 169.85 14.75 169.92 ;
        RECT 0.935 169.92 14.82 169.99 ;
        RECT 0.935 169.99 14.89 170.06 ;
        RECT 0.935 170.06 14.96 170.13 ;
        RECT 0.935 170.13 15.03 170.2 ;
        RECT 0.935 170.2 15.1 170.27 ;
        RECT 0.935 170.27 15.17 170.34 ;
        RECT 0.935 170.34 15.24 170.41 ;
        RECT 0.935 170.41 15.31 170.48 ;
        RECT 0.935 170.48 15.38 170.55 ;
        RECT 0.935 170.55 15.45 170.62 ;
        RECT 0.935 170.62 15.52 170.69 ;
        RECT 0.935 170.69 15.59 170.76 ;
        RECT 0.935 170.76 15.66 170.83 ;
        RECT 0.935 170.83 15.73 170.9 ;
        RECT 0.935 170.9 15.8 170.97 ;
        RECT 0.935 170.97 15.87 171.04 ;
        RECT 0.935 171.04 15.94 171.11 ;
        RECT 0.935 171.11 16.01 171.18 ;
        RECT 0.935 171.18 16.08 171.25 ;
        RECT 0.935 171.25 16.15 171.32 ;
        RECT 0.935 171.32 16.22 171.39 ;
        RECT 0.935 171.39 16.29 171.46 ;
        RECT 0.935 171.46 16.36 171.53 ;
        RECT 0.935 171.53 16.43 171.6 ;
        RECT 0.935 171.6 16.5 171.67 ;
        RECT 0.935 171.67 16.57 171.74 ;
        RECT 0.935 171.74 16.64 171.81 ;
        RECT 0.935 171.81 16.71 171.88 ;
        RECT 0.935 171.88 16.78 171.95 ;
        RECT 0.935 171.95 16.85 172.02 ;
        RECT 0.935 172.02 16.92 172.09 ;
        RECT 0.935 172.09 16.99 172.16 ;
        RECT 0.935 172.16 17.06 172.23 ;
        RECT 0.935 172.23 17.13 172.3 ;
        RECT 0.935 172.3 17.2 172.37 ;
        RECT 0.935 172.37 17.27 172.44 ;
        RECT 0.935 172.44 17.34 172.51 ;
        RECT 0.935 172.51 17.41 172.58 ;
        RECT 0.935 172.58 17.48 172.65 ;
        RECT 0.935 172.65 17.55 172.72 ;
        RECT 0.935 172.72 17.62 172.78 ;
        RECT 0.935 162.08 14.12 169.22 ;
        RECT 0.935 158.48 17.65 158.55 ;
        RECT 0.935 158.55 17.58 158.62 ;
        RECT 0.935 158.62 17.51 158.69 ;
        RECT 0.935 158.69 17.44 158.76 ;
        RECT 0.935 158.76 17.37 158.83 ;
        RECT 0.935 158.83 17.3 158.9 ;
        RECT 0.935 158.9 17.23 158.97 ;
        RECT 0.935 158.97 17.16 159.04 ;
        RECT 0.935 159.04 17.09 159.11 ;
        RECT 0.935 159.11 17.02 159.18 ;
        RECT 0.935 159.18 16.95 159.25 ;
        RECT 0.935 159.25 16.88 159.32 ;
        RECT 0.935 159.32 16.81 159.39 ;
        RECT 0.935 159.39 16.74 159.46 ;
        RECT 0.935 159.46 16.67 159.53 ;
        RECT 0.935 159.53 16.6 159.6 ;
        RECT 0.935 159.6 16.53 159.67 ;
        RECT 0.935 159.67 16.46 159.74 ;
        RECT 0.935 159.74 16.39 159.81 ;
        RECT 0.935 159.81 16.32 159.88 ;
        RECT 0.935 159.88 16.25 159.95 ;
        RECT 0.935 159.95 16.18 160.02 ;
        RECT 0.935 160.02 16.11 160.09 ;
        RECT 0.935 160.09 16.04 160.16 ;
        RECT 0.935 160.16 15.97 160.23 ;
        RECT 0.935 160.23 15.9 160.3 ;
        RECT 0.935 160.3 15.83 160.37 ;
        RECT 0.935 160.37 15.76 160.44 ;
        RECT 0.935 160.44 15.69 160.51 ;
        RECT 0.935 160.51 15.62 160.58 ;
        RECT 0.935 160.58 15.55 160.65 ;
        RECT 0.935 160.65 15.48 160.72 ;
        RECT 0.935 160.72 15.41 160.79 ;
        RECT 0.935 160.79 15.34 160.86 ;
        RECT 0.935 160.86 15.27 160.93 ;
        RECT 0.935 160.93 15.2 161 ;
        RECT 0.935 161 15.13 161.07 ;
        RECT 0.935 161.07 15.06 161.14 ;
        RECT 0.935 161.14 14.99 161.21 ;
        RECT 0.935 161.21 14.92 161.28 ;
        RECT 0.935 161.28 14.85 161.35 ;
        RECT 0.935 161.35 14.78 161.42 ;
        RECT 0.935 161.42 14.71 161.49 ;
        RECT 0.935 161.49 14.64 161.56 ;
        RECT 0.935 161.56 14.57 161.63 ;
        RECT 0.935 161.63 14.5 161.7 ;
        RECT 0.935 161.7 14.43 161.77 ;
        RECT 0.935 161.77 14.36 161.84 ;
        RECT 0.935 161.84 14.29 161.91 ;
        RECT 0.935 161.91 14.22 161.98 ;
        RECT 0.935 161.98 14.15 162.05 ;
        RECT 0.935 162.05 14.12 162.08 ;
        RECT 0.935 149.78 56.705 158.48 ;
        RECT 0.935 146.215 14.12 146.285 ;
        RECT 0.935 146.285 14.19 146.355 ;
        RECT 0.935 146.355 14.26 146.425 ;
        RECT 0.935 146.425 14.33 146.495 ;
        RECT 0.935 146.495 14.4 146.565 ;
        RECT 0.935 146.565 14.47 146.635 ;
        RECT 0.935 146.635 14.54 146.705 ;
        RECT 0.935 146.705 14.61 146.775 ;
        RECT 0.935 146.775 14.68 146.845 ;
        RECT 0.935 146.845 14.75 146.915 ;
        RECT 0.935 146.915 14.82 146.985 ;
        RECT 0.935 146.985 14.89 147.055 ;
        RECT 0.935 147.055 14.96 147.125 ;
        RECT 0.935 147.125 15.03 147.195 ;
        RECT 0.935 147.195 15.1 147.265 ;
        RECT 0.935 147.265 15.17 147.335 ;
        RECT 0.935 147.335 15.24 147.405 ;
        RECT 0.935 147.405 15.31 147.475 ;
        RECT 0.935 147.475 15.38 147.545 ;
        RECT 0.935 147.545 15.45 147.615 ;
        RECT 0.935 147.615 15.52 147.685 ;
        RECT 0.935 147.685 15.59 147.755 ;
        RECT 0.935 147.755 15.66 147.825 ;
        RECT 0.935 147.825 15.73 147.895 ;
        RECT 0.935 147.895 15.8 147.965 ;
        RECT 0.935 147.965 15.87 148.035 ;
        RECT 0.935 148.035 15.94 148.105 ;
        RECT 0.935 148.105 16.01 148.175 ;
        RECT 0.935 148.175 16.08 148.245 ;
        RECT 0.935 148.245 16.15 148.315 ;
        RECT 0.935 148.315 16.22 148.385 ;
        RECT 0.935 148.385 16.29 148.455 ;
        RECT 0.935 148.455 16.36 148.525 ;
        RECT 0.935 148.525 16.43 148.595 ;
        RECT 0.935 148.595 16.5 148.665 ;
        RECT 0.935 148.665 16.57 148.735 ;
        RECT 0.935 148.735 16.64 148.805 ;
        RECT 0.935 148.805 16.71 148.875 ;
        RECT 0.935 148.875 16.78 148.945 ;
        RECT 0.935 148.945 16.85 149.015 ;
        RECT 0.935 149.015 16.92 149.085 ;
        RECT 0.935 149.085 16.99 149.155 ;
        RECT 0.935 149.155 17.06 149.225 ;
        RECT 0.935 149.225 17.13 149.295 ;
        RECT 0.935 149.295 17.2 149.365 ;
        RECT 0.935 149.365 17.27 149.435 ;
        RECT 0.935 149.435 17.34 149.505 ;
        RECT 0.935 149.505 17.41 149.575 ;
        RECT 0.935 149.575 17.48 149.645 ;
        RECT 0.935 149.645 17.55 149.715 ;
        RECT 0.935 149.715 17.62 149.78 ;
        RECT 0.935 139.17 14.12 146.215 ;
        RECT 0.935 135.48 17.74 135.55 ;
        RECT 0.935 135.55 17.67 135.62 ;
        RECT 0.935 135.62 17.6 135.69 ;
        RECT 0.935 135.69 17.53 135.76 ;
        RECT 0.935 135.76 17.46 135.83 ;
        RECT 0.935 135.83 17.39 135.9 ;
        RECT 0.935 135.9 17.32 135.97 ;
        RECT 0.935 135.97 17.25 136.04 ;
        RECT 0.935 136.04 17.18 136.11 ;
        RECT 0.935 136.11 17.11 136.18 ;
        RECT 0.935 136.18 17.04 136.25 ;
        RECT 0.935 136.25 16.97 136.32 ;
        RECT 0.935 136.32 16.9 136.39 ;
        RECT 0.935 136.39 16.83 136.46 ;
        RECT 0.935 136.46 16.76 136.53 ;
        RECT 0.935 136.53 16.69 136.6 ;
        RECT 0.935 136.6 16.62 136.67 ;
        RECT 0.935 136.67 16.55 136.74 ;
        RECT 0.935 136.74 16.48 136.81 ;
        RECT 0.935 136.81 16.41 136.88 ;
        RECT 0.935 136.88 16.34 136.95 ;
        RECT 0.935 136.95 16.27 137.02 ;
        RECT 0.935 137.02 16.2 137.09 ;
        RECT 0.935 137.09 16.13 137.16 ;
        RECT 0.935 137.16 16.06 137.23 ;
        RECT 0.935 137.23 15.99 137.3 ;
        RECT 0.935 137.3 15.92 137.37 ;
        RECT 0.935 137.37 15.85 137.44 ;
        RECT 0.935 137.44 15.78 137.51 ;
        RECT 0.935 137.51 15.71 137.58 ;
        RECT 0.935 137.58 15.64 137.65 ;
        RECT 0.935 137.65 15.57 137.72 ;
        RECT 0.935 137.72 15.5 137.79 ;
        RECT 0.935 137.79 15.43 137.86 ;
        RECT 0.935 137.86 15.36 137.93 ;
        RECT 0.935 137.93 15.29 138 ;
        RECT 0.935 138 15.22 138.07 ;
        RECT 0.935 138.07 15.15 138.14 ;
        RECT 0.935 138.14 15.08 138.21 ;
        RECT 0.935 138.21 15.01 138.28 ;
        RECT 0.935 138.28 14.94 138.35 ;
        RECT 0.935 138.35 14.87 138.42 ;
        RECT 0.935 138.42 14.8 138.49 ;
        RECT 0.935 138.49 14.73 138.56 ;
        RECT 0.935 138.56 14.66 138.63 ;
        RECT 0.935 138.63 14.59 138.7 ;
        RECT 0.935 138.7 14.52 138.77 ;
        RECT 0.935 138.77 14.45 138.84 ;
        RECT 0.935 138.84 14.38 138.91 ;
        RECT 0.935 138.91 14.31 138.98 ;
        RECT 0.935 138.98 14.24 139.05 ;
        RECT 0.935 139.05 14.17 139.12 ;
        RECT 0.935 139.12 14.12 139.17 ;
        RECT 0.935 126.78 56.705 135.48 ;
        RECT 0.935 123.145 14.12 123.215 ;
        RECT 0.935 123.215 14.19 123.285 ;
        RECT 0.935 123.285 14.26 123.355 ;
        RECT 0.935 123.355 14.33 123.425 ;
        RECT 0.935 123.425 14.4 123.495 ;
        RECT 0.935 123.495 14.47 123.565 ;
        RECT 0.935 123.565 14.54 123.635 ;
        RECT 0.935 123.635 14.61 123.705 ;
        RECT 0.935 123.705 14.68 123.775 ;
        RECT 0.935 123.775 14.75 123.845 ;
        RECT 0.935 123.845 14.82 123.915 ;
        RECT 0.935 123.915 14.89 123.985 ;
        RECT 0.935 123.985 14.96 124.055 ;
        RECT 0.935 124.055 15.03 124.125 ;
        RECT 0.935 124.125 15.1 124.195 ;
        RECT 0.935 124.195 15.17 124.265 ;
        RECT 0.935 124.265 15.24 124.335 ;
        RECT 0.935 124.335 15.31 124.405 ;
        RECT 0.935 124.405 15.38 124.475 ;
        RECT 0.935 124.475 15.45 124.545 ;
        RECT 0.935 124.545 15.52 124.615 ;
        RECT 0.935 124.615 15.59 124.685 ;
        RECT 0.935 124.685 15.66 124.755 ;
        RECT 0.935 124.755 15.73 124.825 ;
        RECT 0.935 124.825 15.8 124.895 ;
        RECT 0.935 124.895 15.87 124.965 ;
        RECT 0.935 124.965 15.94 125.035 ;
        RECT 0.935 125.035 16.01 125.105 ;
        RECT 0.935 125.105 16.08 125.175 ;
        RECT 0.935 125.175 16.15 125.245 ;
        RECT 0.935 125.245 16.22 125.315 ;
        RECT 0.935 125.315 16.29 125.385 ;
        RECT 0.935 125.385 16.36 125.455 ;
        RECT 0.935 125.455 16.43 125.525 ;
        RECT 0.935 125.525 16.5 125.595 ;
        RECT 0.935 125.595 16.57 125.665 ;
        RECT 0.935 125.665 16.64 125.735 ;
        RECT 0.935 125.735 16.71 125.805 ;
        RECT 0.935 125.805 16.78 125.875 ;
        RECT 0.935 125.875 16.85 125.945 ;
        RECT 0.935 125.945 16.92 126.015 ;
        RECT 0.935 126.015 16.99 126.085 ;
        RECT 0.935 126.085 17.06 126.155 ;
        RECT 0.935 126.155 17.13 126.225 ;
        RECT 0.935 126.225 17.2 126.295 ;
        RECT 0.935 126.295 17.27 126.365 ;
        RECT 0.935 126.365 17.34 126.435 ;
        RECT 0.935 126.435 17.41 126.505 ;
        RECT 0.935 126.505 17.48 126.575 ;
        RECT 0.935 126.575 17.55 126.645 ;
        RECT 0.935 126.645 17.62 126.715 ;
        RECT 0.935 126.715 17.69 126.78 ;
        RECT 0.935 116.065 14.12 123.145 ;
        RECT 0.935 112.48 17.635 112.55 ;
        RECT 0.935 112.55 17.565 112.62 ;
        RECT 0.935 112.62 17.495 112.69 ;
        RECT 0.935 112.69 17.425 112.76 ;
        RECT 0.935 112.76 17.355 112.83 ;
        RECT 0.935 112.83 17.285 112.9 ;
        RECT 0.935 112.9 17.215 112.97 ;
        RECT 0.935 112.97 17.145 113.04 ;
        RECT 0.935 113.04 17.075 113.11 ;
        RECT 0.935 113.11 17.005 113.18 ;
        RECT 0.935 113.18 16.935 113.25 ;
        RECT 0.935 113.25 16.865 113.32 ;
        RECT 0.935 113.32 16.795 113.39 ;
        RECT 0.935 113.39 16.725 113.46 ;
        RECT 0.935 113.46 16.655 113.53 ;
        RECT 0.935 113.53 16.585 113.6 ;
        RECT 0.935 113.6 16.515 113.67 ;
        RECT 0.935 113.67 16.445 113.74 ;
        RECT 0.935 113.74 16.375 113.81 ;
        RECT 0.935 113.81 16.305 113.88 ;
        RECT 0.935 113.88 16.235 113.95 ;
        RECT 0.935 113.95 16.165 114.02 ;
        RECT 0.935 114.02 16.095 114.09 ;
        RECT 0.935 114.09 16.025 114.16 ;
        RECT 0.935 114.16 15.955 114.23 ;
        RECT 0.935 114.23 15.885 114.3 ;
        RECT 0.935 114.3 15.815 114.37 ;
        RECT 0.935 114.37 15.745 114.44 ;
        RECT 0.935 114.44 15.675 114.51 ;
        RECT 0.935 114.51 15.605 114.58 ;
        RECT 0.935 114.58 15.535 114.65 ;
        RECT 0.935 114.65 15.465 114.72 ;
        RECT 0.935 114.72 15.395 114.79 ;
        RECT 0.935 114.79 15.325 114.86 ;
        RECT 0.935 114.86 15.255 114.93 ;
        RECT 0.935 114.93 15.185 115 ;
        RECT 0.935 115 15.115 115.07 ;
        RECT 0.935 115.07 15.045 115.14 ;
        RECT 0.935 115.14 14.975 115.21 ;
        RECT 0.935 115.21 14.905 115.28 ;
        RECT 0.935 115.28 14.835 115.35 ;
        RECT 0.935 115.35 14.765 115.42 ;
        RECT 0.935 115.42 14.695 115.49 ;
        RECT 0.935 115.49 14.625 115.56 ;
        RECT 0.935 115.56 14.555 115.63 ;
        RECT 0.935 115.63 14.485 115.7 ;
        RECT 0.935 115.7 14.415 115.77 ;
        RECT 0.935 115.77 14.345 115.84 ;
        RECT 0.935 115.84 14.275 115.91 ;
        RECT 0.935 115.91 14.205 115.98 ;
        RECT 0.935 115.98 14.135 116.05 ;
        RECT 0.935 116.05 14.12 116.065 ;
        RECT 0.935 103.78 56.705 112.48 ;
        RECT 0.935 100.24 14.12 100.31 ;
        RECT 0.935 100.31 14.19 100.38 ;
        RECT 0.935 100.38 14.26 100.45 ;
        RECT 0.935 100.45 14.33 100.52 ;
        RECT 0.935 100.52 14.4 100.59 ;
        RECT 0.935 100.59 14.47 100.66 ;
        RECT 0.935 100.66 14.54 100.73 ;
        RECT 0.935 100.73 14.61 100.8 ;
        RECT 0.935 100.8 14.68 100.87 ;
        RECT 0.935 100.87 14.75 100.94 ;
        RECT 0.935 100.94 14.82 101.01 ;
        RECT 0.935 101.01 14.89 101.08 ;
        RECT 0.935 101.08 14.96 101.15 ;
        RECT 0.935 101.15 15.03 101.22 ;
        RECT 0.935 101.22 15.1 101.29 ;
        RECT 0.935 101.29 15.17 101.36 ;
        RECT 0.935 101.36 15.24 101.43 ;
        RECT 0.935 101.43 15.31 101.5 ;
        RECT 0.935 101.5 15.38 101.57 ;
        RECT 0.935 101.57 15.45 101.64 ;
        RECT 0.935 101.64 15.52 101.71 ;
        RECT 0.935 101.71 15.59 101.78 ;
        RECT 0.935 101.78 15.66 101.85 ;
        RECT 0.935 101.85 15.73 101.92 ;
        RECT 0.935 101.92 15.8 101.99 ;
        RECT 0.935 101.99 15.87 102.06 ;
        RECT 0.935 102.06 15.94 102.13 ;
        RECT 0.935 102.13 16.01 102.2 ;
        RECT 0.935 102.2 16.08 102.27 ;
        RECT 0.935 102.27 16.15 102.34 ;
        RECT 0.935 102.34 16.22 102.41 ;
        RECT 0.935 102.41 16.29 102.48 ;
        RECT 0.935 102.48 16.36 102.55 ;
        RECT 0.935 102.55 16.43 102.62 ;
        RECT 0.935 102.62 16.5 102.69 ;
        RECT 0.935 102.69 16.57 102.76 ;
        RECT 0.935 102.76 16.64 102.83 ;
        RECT 0.935 102.83 16.71 102.9 ;
        RECT 0.935 102.9 16.78 102.97 ;
        RECT 0.935 102.97 16.85 103.04 ;
        RECT 0.935 103.04 16.92 103.11 ;
        RECT 0.935 103.11 16.99 103.18 ;
        RECT 0.935 103.18 17.06 103.25 ;
        RECT 0.935 103.25 17.13 103.32 ;
        RECT 0.935 103.32 17.2 103.39 ;
        RECT 0.935 103.39 17.27 103.46 ;
        RECT 0.935 103.46 17.34 103.53 ;
        RECT 0.935 103.53 17.41 103.6 ;
        RECT 0.935 103.6 17.48 103.67 ;
        RECT 0.935 103.67 17.55 103.74 ;
        RECT 0.935 103.74 17.62 103.78 ;
        RECT 0.935 93.025 14.12 100.24 ;
        RECT 0.935 89.48 17.595 89.55 ;
        RECT 0.935 89.55 17.525 89.62 ;
        RECT 0.935 89.62 17.455 89.69 ;
        RECT 0.935 89.69 17.385 89.76 ;
        RECT 0.935 89.76 17.315 89.83 ;
        RECT 0.935 89.83 17.245 89.9 ;
        RECT 0.935 89.9 17.175 89.97 ;
        RECT 0.935 89.97 17.105 90.04 ;
        RECT 0.935 90.04 17.035 90.11 ;
        RECT 0.935 90.11 16.965 90.18 ;
        RECT 0.935 90.18 16.895 90.25 ;
        RECT 0.935 90.25 16.825 90.32 ;
        RECT 0.935 90.32 16.755 90.39 ;
        RECT 0.935 90.39 16.685 90.46 ;
        RECT 0.935 90.46 16.615 90.53 ;
        RECT 0.935 90.53 16.545 90.6 ;
        RECT 0.935 90.6 16.475 90.67 ;
        RECT 0.935 90.67 16.405 90.74 ;
        RECT 0.935 90.74 16.335 90.81 ;
        RECT 0.935 90.81 16.265 90.88 ;
        RECT 0.935 90.88 16.195 90.95 ;
        RECT 0.935 90.95 16.125 91.02 ;
        RECT 0.935 91.02 16.055 91.09 ;
        RECT 0.935 91.09 15.985 91.16 ;
        RECT 0.935 91.16 15.915 91.23 ;
        RECT 0.935 91.23 15.845 91.3 ;
        RECT 0.935 91.3 15.775 91.37 ;
        RECT 0.935 91.37 15.705 91.44 ;
        RECT 0.935 91.44 15.635 91.51 ;
        RECT 0.935 91.51 15.565 91.58 ;
        RECT 0.935 91.58 15.495 91.65 ;
        RECT 0.935 91.65 15.425 91.72 ;
        RECT 0.935 91.72 15.355 91.79 ;
        RECT 0.935 91.79 15.285 91.86 ;
        RECT 0.935 91.86 15.215 91.93 ;
        RECT 0.935 91.93 15.145 92 ;
        RECT 0.935 92 15.075 92.07 ;
        RECT 0.935 92.07 15.005 92.14 ;
        RECT 0.935 92.14 14.935 92.21 ;
        RECT 0.935 92.21 14.865 92.28 ;
        RECT 0.935 92.28 14.795 92.35 ;
        RECT 0.935 92.35 14.725 92.42 ;
        RECT 0.935 92.42 14.655 92.49 ;
        RECT 0.935 92.49 14.585 92.56 ;
        RECT 0.935 92.56 14.515 92.63 ;
        RECT 0.935 92.63 14.445 92.7 ;
        RECT 0.935 92.7 14.375 92.77 ;
        RECT 0.935 92.77 14.305 92.84 ;
        RECT 0.935 92.84 14.235 92.91 ;
        RECT 0.935 92.91 14.165 92.98 ;
        RECT 0.935 92.98 14.12 93.025 ;
        RECT 0.935 80.78 56.705 89.48 ;
        RECT 0.935 77.24 14.12 77.31 ;
        RECT 0.935 77.31 14.19 77.38 ;
        RECT 0.935 77.38 14.26 77.45 ;
        RECT 0.935 77.45 14.33 77.52 ;
        RECT 0.935 77.52 14.4 77.59 ;
        RECT 0.935 77.59 14.47 77.66 ;
        RECT 0.935 77.66 14.54 77.73 ;
        RECT 0.935 77.73 14.61 77.8 ;
        RECT 0.935 77.8 14.68 77.87 ;
        RECT 0.935 77.87 14.75 77.94 ;
        RECT 0.935 77.94 14.82 78.01 ;
        RECT 0.935 78.01 14.89 78.08 ;
        RECT 0.935 78.08 14.96 78.15 ;
        RECT 0.935 78.15 15.03 78.22 ;
        RECT 0.935 78.22 15.1 78.29 ;
        RECT 0.935 78.29 15.17 78.36 ;
        RECT 0.935 78.36 15.24 78.43 ;
        RECT 0.935 78.43 15.31 78.5 ;
        RECT 0.935 78.5 15.38 78.57 ;
        RECT 0.935 78.57 15.45 78.64 ;
        RECT 0.935 78.64 15.52 78.71 ;
        RECT 0.935 78.71 15.59 78.78 ;
        RECT 0.935 78.78 15.66 78.85 ;
        RECT 0.935 78.85 15.73 78.92 ;
        RECT 0.935 78.92 15.8 78.99 ;
        RECT 0.935 78.99 15.87 79.06 ;
        RECT 0.935 79.06 15.94 79.13 ;
        RECT 0.935 79.13 16.01 79.2 ;
        RECT 0.935 79.2 16.08 79.27 ;
        RECT 0.935 79.27 16.15 79.34 ;
        RECT 0.935 79.34 16.22 79.41 ;
        RECT 0.935 79.41 16.29 79.48 ;
        RECT 0.935 79.48 16.36 79.55 ;
        RECT 0.935 79.55 16.43 79.62 ;
        RECT 0.935 79.62 16.5 79.69 ;
        RECT 0.935 79.69 16.57 79.76 ;
        RECT 0.935 79.76 16.64 79.83 ;
        RECT 0.935 79.83 16.71 79.9 ;
        RECT 0.935 79.9 16.78 79.97 ;
        RECT 0.935 79.97 16.85 80.04 ;
        RECT 0.935 80.04 16.92 80.11 ;
        RECT 0.935 80.11 16.99 80.18 ;
        RECT 0.935 80.18 17.06 80.25 ;
        RECT 0.935 80.25 17.13 80.32 ;
        RECT 0.935 80.32 17.2 80.39 ;
        RECT 0.935 80.39 17.27 80.46 ;
        RECT 0.935 80.46 17.34 80.53 ;
        RECT 0.935 80.53 17.41 80.6 ;
        RECT 0.935 80.6 17.48 80.67 ;
        RECT 0.935 80.67 17.55 80.74 ;
        RECT 0.935 80.74 17.62 80.78 ;
        RECT 0.935 70.025 14.12 77.24 ;
        RECT 0.935 66.48 17.595 66.55 ;
        RECT 0.935 66.55 17.525 66.62 ;
        RECT 0.935 66.62 17.455 66.69 ;
        RECT 0.935 66.69 17.385 66.76 ;
        RECT 0.935 66.76 17.315 66.83 ;
        RECT 0.935 66.83 17.245 66.9 ;
        RECT 0.935 66.9 17.175 66.97 ;
        RECT 0.935 66.97 17.105 67.04 ;
        RECT 0.935 67.04 17.035 67.11 ;
        RECT 0.935 67.11 16.965 67.18 ;
        RECT 0.935 67.18 16.895 67.25 ;
        RECT 0.935 67.25 16.825 67.32 ;
        RECT 0.935 67.32 16.755 67.39 ;
        RECT 0.935 67.39 16.685 67.46 ;
        RECT 0.935 67.46 16.615 67.53 ;
        RECT 0.935 67.53 16.545 67.6 ;
        RECT 0.935 67.6 16.475 67.67 ;
        RECT 0.935 67.67 16.405 67.74 ;
        RECT 0.935 67.74 16.335 67.81 ;
        RECT 0.935 67.81 16.265 67.88 ;
        RECT 0.935 67.88 16.195 67.95 ;
        RECT 0.935 67.95 16.125 68.02 ;
        RECT 0.935 68.02 16.055 68.09 ;
        RECT 0.935 68.09 15.985 68.16 ;
        RECT 0.935 68.16 15.915 68.23 ;
        RECT 0.935 68.23 15.845 68.3 ;
        RECT 0.935 68.3 15.775 68.37 ;
        RECT 0.935 68.37 15.705 68.44 ;
        RECT 0.935 68.44 15.635 68.51 ;
        RECT 0.935 68.51 15.565 68.58 ;
        RECT 0.935 68.58 15.495 68.65 ;
        RECT 0.935 68.65 15.425 68.72 ;
        RECT 0.935 68.72 15.355 68.79 ;
        RECT 0.935 68.79 15.285 68.86 ;
        RECT 0.935 68.86 15.215 68.93 ;
        RECT 0.935 68.93 15.145 69 ;
        RECT 0.935 69 15.075 69.07 ;
        RECT 0.935 69.07 15.005 69.14 ;
        RECT 0.935 69.14 14.935 69.21 ;
        RECT 0.935 69.21 14.865 69.28 ;
        RECT 0.935 69.28 14.795 69.35 ;
        RECT 0.935 69.35 14.725 69.42 ;
        RECT 0.935 69.42 14.655 69.49 ;
        RECT 0.935 69.49 14.585 69.56 ;
        RECT 0.935 69.56 14.515 69.63 ;
        RECT 0.935 69.63 14.445 69.7 ;
        RECT 0.935 69.7 14.375 69.77 ;
        RECT 0.935 69.77 14.305 69.84 ;
        RECT 0.935 69.84 14.235 69.91 ;
        RECT 0.935 69.91 14.165 69.98 ;
        RECT 0.935 69.98 14.12 70.025 ;
        RECT 0.935 57.78 56.71 66.48 ;
        RECT 0.935 54.215 14.12 54.285 ;
        RECT 0.935 54.285 14.19 54.355 ;
        RECT 0.935 54.355 14.26 54.425 ;
        RECT 0.935 54.425 14.33 54.495 ;
        RECT 0.935 54.495 14.4 54.565 ;
        RECT 0.935 54.565 14.47 54.635 ;
        RECT 0.935 54.635 14.54 54.705 ;
        RECT 0.935 54.705 14.61 54.775 ;
        RECT 0.935 54.775 14.68 54.845 ;
        RECT 0.935 54.845 14.75 54.915 ;
        RECT 0.935 54.915 14.82 54.985 ;
        RECT 0.935 54.985 14.89 55.055 ;
        RECT 0.935 55.055 14.96 55.125 ;
        RECT 0.935 55.125 15.03 55.195 ;
        RECT 0.935 55.195 15.1 55.265 ;
        RECT 0.935 55.265 15.17 55.335 ;
        RECT 0.935 55.335 15.24 55.405 ;
        RECT 0.935 55.405 15.31 55.475 ;
        RECT 0.935 55.475 15.38 55.545 ;
        RECT 0.935 55.545 15.45 55.615 ;
        RECT 0.935 55.615 15.52 55.685 ;
        RECT 0.935 55.685 15.59 55.755 ;
        RECT 0.935 55.755 15.66 55.825 ;
        RECT 0.935 55.825 15.73 55.895 ;
        RECT 0.935 55.895 15.8 55.965 ;
        RECT 0.935 55.965 15.87 56.035 ;
        RECT 0.935 56.035 15.94 56.105 ;
        RECT 0.935 56.105 16.01 56.175 ;
        RECT 0.935 56.175 16.08 56.245 ;
        RECT 0.935 56.245 16.15 56.315 ;
        RECT 0.935 56.315 16.22 56.385 ;
        RECT 0.935 56.385 16.29 56.455 ;
        RECT 0.935 56.455 16.36 56.525 ;
        RECT 0.935 56.525 16.43 56.595 ;
        RECT 0.935 56.595 16.5 56.665 ;
        RECT 0.935 56.665 16.57 56.735 ;
        RECT 0.935 56.735 16.64 56.805 ;
        RECT 0.935 56.805 16.71 56.875 ;
        RECT 0.935 56.875 16.78 56.945 ;
        RECT 0.935 56.945 16.85 57.015 ;
        RECT 0.935 57.015 16.92 57.085 ;
        RECT 0.935 57.085 16.99 57.155 ;
        RECT 0.935 57.155 17.06 57.225 ;
        RECT 0.935 57.225 17.13 57.295 ;
        RECT 0.935 57.295 17.2 57.365 ;
        RECT 0.935 57.365 17.27 57.435 ;
        RECT 0.935 57.435 17.34 57.505 ;
        RECT 0.935 57.505 17.41 57.575 ;
        RECT 0.935 57.575 17.48 57.645 ;
        RECT 0.935 57.645 17.55 57.715 ;
        RECT 0.935 57.715 17.62 57.78 ;
        RECT 0.935 45.315 14.12 54.215 ;
        RECT 0.935 42.38 16.985 42.45 ;
        RECT 0.935 42.45 16.915 42.52 ;
        RECT 0.935 42.52 16.845 42.59 ;
        RECT 0.935 42.59 16.775 42.66 ;
        RECT 0.935 42.66 16.705 42.73 ;
        RECT 0.935 42.73 16.635 42.8 ;
        RECT 0.935 42.8 16.565 42.87 ;
        RECT 0.935 42.87 16.495 42.94 ;
        RECT 0.935 42.94 16.425 43.01 ;
        RECT 0.935 43.01 16.355 43.08 ;
        RECT 0.935 43.08 16.285 43.15 ;
        RECT 0.935 43.15 16.215 43.22 ;
        RECT 0.935 43.22 16.145 43.29 ;
        RECT 0.935 43.29 16.075 43.36 ;
        RECT 0.935 43.36 16.005 43.43 ;
        RECT 0.935 43.43 15.935 43.5 ;
        RECT 0.935 43.5 15.865 43.57 ;
        RECT 0.935 43.57 15.795 43.64 ;
        RECT 0.935 43.64 15.725 43.71 ;
        RECT 0.935 43.71 15.655 43.78 ;
        RECT 0.935 43.78 15.585 43.85 ;
        RECT 0.935 43.85 15.515 43.92 ;
        RECT 0.935 43.92 15.445 43.99 ;
        RECT 0.935 43.99 15.375 44.06 ;
        RECT 0.935 44.06 15.305 44.13 ;
        RECT 0.935 44.13 15.235 44.2 ;
        RECT 0.935 44.2 15.165 44.27 ;
        RECT 0.935 44.27 15.095 44.34 ;
        RECT 0.935 44.34 15.025 44.41 ;
        RECT 0.935 44.41 14.955 44.48 ;
        RECT 0.935 44.48 14.885 44.55 ;
        RECT 0.935 44.55 14.815 44.62 ;
        RECT 0.935 44.62 14.745 44.69 ;
        RECT 0.935 44.69 14.675 44.76 ;
        RECT 0.935 44.76 14.605 44.83 ;
        RECT 0.935 44.83 14.535 44.9 ;
        RECT 0.935 44.9 14.465 44.97 ;
        RECT 0.935 44.97 14.395 45.04 ;
        RECT 0.935 45.04 14.325 45.11 ;
        RECT 0.935 45.11 14.255 45.18 ;
        RECT 0.935 45.18 14.185 45.25 ;
        RECT 0.935 45.25 14.12 45.315 ;
        RECT 0.935 40.35 56.16 40.42 ;
        RECT 0.935 40.42 56.09 40.49 ;
        RECT 0.935 40.49 56.02 40.56 ;
        RECT 0.935 40.56 55.95 40.63 ;
        RECT 0.935 40.63 55.88 40.7 ;
        RECT 0.935 40.7 55.81 40.77 ;
        RECT 0.935 40.77 55.74 40.84 ;
        RECT 0.935 40.84 55.67 40.91 ;
        RECT 0.935 40.91 55.6 40.98 ;
        RECT 0.935 40.98 55.53 41.05 ;
        RECT 0.935 41.05 55.46 41.12 ;
        RECT 0.935 41.12 55.39 41.19 ;
        RECT 0.935 41.19 55.32 41.26 ;
        RECT 0.935 41.26 55.25 41.33 ;
        RECT 0.935 41.33 55.18 41.4 ;
        RECT 0.935 41.4 55.11 41.47 ;
        RECT 0.935 41.47 55.04 41.54 ;
        RECT 0.935 41.54 54.97 41.61 ;
        RECT 0.935 41.61 54.9 41.68 ;
        RECT 0.935 41.68 54.83 41.75 ;
        RECT 0.935 41.75 54.76 41.82 ;
        RECT 0.935 41.82 54.69 41.89 ;
        RECT 0.935 41.89 54.62 41.96 ;
        RECT 0.935 41.96 54.55 42.03 ;
        RECT 0.935 42.03 54.48 42.1 ;
        RECT 0.935 42.1 54.41 42.17 ;
        RECT 0.935 42.17 54.34 42.24 ;
        RECT 0.935 42.24 54.27 42.31 ;
        RECT 0.935 42.31 54.2 42.38 ;
        RECT 53.26 39.665 56.845 39.735 ;
        RECT 53.19 39.735 56.775 39.805 ;
        RECT 53.12 39.805 56.705 39.875 ;
        RECT 53.05 39.875 56.635 39.945 ;
        RECT 52.98 39.945 56.565 40.015 ;
        RECT 52.91 40.015 56.495 40.085 ;
        RECT 52.84 40.085 56.425 40.155 ;
        RECT 52.77 40.155 56.355 40.225 ;
        RECT 52.7 40.225 56.285 40.295 ;
        RECT 52.63 40.295 56.23 40.35 ;
        RECT 54.67 38.255 56.915 38.325 ;
        RECT 54.6 38.325 56.915 38.395 ;
        RECT 54.53 38.395 56.915 38.465 ;
        RECT 54.46 38.465 56.915 38.535 ;
        RECT 54.39 38.535 56.915 38.605 ;
        RECT 54.32 38.605 56.915 38.675 ;
        RECT 54.25 38.675 56.915 38.745 ;
        RECT 54.18 38.745 56.915 38.815 ;
        RECT 54.11 38.815 56.915 38.885 ;
        RECT 54.04 38.885 56.915 38.955 ;
        RECT 53.97 38.955 56.915 39.025 ;
        RECT 53.9 39.025 56.915 39.095 ;
        RECT 53.83 39.095 56.915 39.165 ;
        RECT 53.76 39.165 56.915 39.235 ;
        RECT 53.69 39.235 56.915 39.305 ;
        RECT 53.62 39.305 56.915 39.375 ;
        RECT 53.55 39.375 56.915 39.445 ;
        RECT 53.48 39.445 56.915 39.515 ;
        RECT 53.41 39.515 56.915 39.585 ;
        RECT 53.34 39.585 56.915 39.655 ;
        RECT 53.27 39.655 56.915 39.665 ;
        RECT 54.67 36.115 56.915 38.255 ;
        RECT 0.935 40.285 19.825 40.35 ;
        RECT 0.935 40.215 19.755 40.285 ;
        RECT 0.935 40.145 19.685 40.215 ;
        RECT 0.935 40.075 19.615 40.145 ;
        RECT 0.935 40.005 19.545 40.075 ;
        RECT 0.935 39.935 19.475 40.005 ;
        RECT 0.935 39.865 19.405 39.935 ;
        RECT 0.935 39.795 19.335 39.865 ;
        RECT 0.935 39.725 19.265 39.795 ;
        RECT 0.935 39.655 19.195 39.725 ;
        RECT 0.935 39.585 19.125 39.655 ;
        RECT 0.935 39.515 19.055 39.585 ;
        RECT 0.935 39.445 18.985 39.515 ;
        RECT 0.935 39.375 18.915 39.445 ;
        RECT 0.935 39.305 18.845 39.375 ;
        RECT 0.935 39.235 18.775 39.305 ;
        RECT 0.935 39.165 18.705 39.235 ;
        RECT 0.935 39.095 18.635 39.165 ;
        RECT 0.935 39.025 18.565 39.095 ;
        RECT 0.935 38.955 18.495 39.025 ;
        RECT 0.935 38.885 18.425 38.955 ;
        RECT 0.935 38.815 18.355 38.885 ;
        RECT 0.935 38.745 18.285 38.815 ;
        RECT 0.935 38.675 18.215 38.745 ;
        RECT 0.935 38.605 18.145 38.675 ;
        RECT 0.935 38.535 18.075 38.605 ;
        RECT 0.935 38.465 18.005 38.535 ;
        RECT 0.935 38.395 17.935 38.465 ;
        RECT 0.935 38.325 17.865 38.395 ;
        RECT 0.935 38.255 17.795 38.325 ;
        RECT 0.935 38.185 17.725 38.255 ;
        RECT 0.935 38.115 17.655 38.185 ;
        RECT 0.935 38.045 17.585 38.115 ;
        RECT 0.935 37.975 17.515 38.045 ;
        RECT 0.935 37.905 17.445 37.975 ;
        RECT 0.935 37.835 17.375 37.905 ;
        RECT 0.935 37.765 17.305 37.835 ;
        RECT 0.935 37.695 17.235 37.765 ;
        RECT 0.935 37.625 17.165 37.695 ;
        RECT 0.935 37.555 17.095 37.625 ;
        RECT 0.935 37.485 17.025 37.555 ;
        RECT 0.935 37.415 16.955 37.485 ;
        RECT 0.935 37.345 16.885 37.415 ;
        RECT 0.935 37.275 16.815 37.345 ;
        RECT 0.935 37.205 16.745 37.275 ;
        RECT 0.935 37.135 16.675 37.205 ;
        RECT 0.935 37.065 16.605 37.135 ;
        RECT 0.935 36.995 16.535 37.065 ;
        RECT 0.935 36.925 16.465 36.995 ;
        RECT 0.935 36.855 16.395 36.925 ;
        RECT 0.935 36.785 16.325 36.855 ;
        RECT 0.935 36.715 16.255 36.785 ;
        RECT 0.935 36.645 16.185 36.715 ;
        RECT 0.935 36.575 16.115 36.645 ;
        RECT 0.935 36.505 16.045 36.575 ;
        RECT 0.935 36.435 15.975 36.505 ;
        RECT 0.935 36.365 15.905 36.435 ;
        RECT 0.935 36.295 15.835 36.365 ;
        RECT 0.935 36.225 15.765 36.295 ;
        RECT 0.935 36.155 15.695 36.225 ;
        RECT 0.935 36.085 15.625 36.155 ;
        RECT 0.935 36.015 15.555 36.085 ;
        RECT 0.935 35.945 15.485 36.015 ;
        RECT 0.935 35.875 15.415 35.945 ;
        RECT 0.935 35.805 15.345 35.875 ;
        RECT 0.935 35.735 15.275 35.805 ;
        RECT 0.935 35.665 15.205 35.735 ;
        RECT 0.935 29.315 15.205 35.665 ;
        RECT 0.935 25.7 18.75 25.77 ;
        RECT 0.935 25.77 18.68 25.84 ;
        RECT 0.935 25.84 18.61 25.91 ;
        RECT 0.935 25.91 18.54 25.98 ;
        RECT 0.935 25.98 18.47 26.05 ;
        RECT 0.935 26.05 18.4 26.12 ;
        RECT 0.935 26.12 18.33 26.19 ;
        RECT 0.935 26.19 18.26 26.26 ;
        RECT 0.935 26.26 18.19 26.33 ;
        RECT 0.935 26.33 18.12 26.4 ;
        RECT 0.935 26.4 18.05 26.47 ;
        RECT 0.935 26.47 17.98 26.54 ;
        RECT 0.935 26.54 17.91 26.61 ;
        RECT 0.935 26.61 17.84 26.68 ;
        RECT 0.935 26.68 17.77 26.75 ;
        RECT 0.935 26.75 17.7 26.82 ;
        RECT 0.935 26.82 17.63 26.89 ;
        RECT 0.935 26.89 17.56 26.96 ;
        RECT 0.935 26.96 17.49 27.03 ;
        RECT 0.935 27.03 17.42 27.1 ;
        RECT 0.935 27.1 17.35 27.17 ;
        RECT 0.935 27.17 17.28 27.24 ;
        RECT 0.935 27.24 17.21 27.31 ;
        RECT 0.935 27.31 17.14 27.38 ;
        RECT 0.935 27.38 17.07 27.45 ;
        RECT 0.935 27.45 17 27.52 ;
        RECT 0.935 27.52 16.93 27.59 ;
        RECT 0.935 27.59 16.86 27.66 ;
        RECT 0.935 27.66 16.79 27.73 ;
        RECT 0.935 27.73 16.72 27.8 ;
        RECT 0.935 27.8 16.65 27.87 ;
        RECT 0.935 27.87 16.58 27.94 ;
        RECT 0.935 27.94 16.51 28.01 ;
        RECT 0.935 28.01 16.44 28.08 ;
        RECT 0.935 28.08 16.37 28.15 ;
        RECT 0.935 28.15 16.3 28.22 ;
        RECT 0.935 28.22 16.23 28.29 ;
        RECT 0.935 28.29 16.16 28.36 ;
        RECT 0.935 28.36 16.09 28.43 ;
        RECT 0.935 28.43 16.02 28.5 ;
        RECT 0.935 28.5 15.95 28.57 ;
        RECT 0.935 28.57 15.88 28.64 ;
        RECT 0.935 28.64 15.81 28.71 ;
        RECT 0.935 28.71 15.74 28.78 ;
        RECT 0.935 28.78 15.67 28.85 ;
        RECT 0.935 28.85 15.6 28.92 ;
        RECT 0.935 28.92 15.53 28.99 ;
        RECT 0.935 28.99 15.46 29.06 ;
        RECT 0.935 29.06 15.39 29.13 ;
        RECT 0.935 29.13 15.32 29.2 ;
        RECT 0.935 29.2 15.25 29.27 ;
        RECT 0.935 29.27 15.205 29.315 ;
        RECT 0.935 12.4 36.895 25.7 ;
        RECT 0.935 8.595 24.395 8.665 ;
        RECT 0.935 8.665 24.465 8.735 ;
        RECT 0.935 8.735 24.535 8.805 ;
        RECT 0.935 8.805 24.605 8.875 ;
        RECT 0.935 8.875 24.675 8.945 ;
        RECT 0.935 8.945 24.745 9.015 ;
        RECT 0.935 9.015 24.815 9.085 ;
        RECT 0.935 9.085 24.885 9.155 ;
        RECT 0.935 9.155 24.955 9.225 ;
        RECT 0.935 9.225 25.025 9.295 ;
        RECT 0.935 9.295 25.095 9.365 ;
        RECT 0.935 9.365 25.165 9.435 ;
        RECT 0.935 9.435 25.235 9.505 ;
        RECT 0.935 9.505 25.305 9.575 ;
        RECT 0.935 9.575 25.375 9.645 ;
        RECT 0.935 9.645 25.445 9.715 ;
        RECT 0.935 9.715 25.515 9.785 ;
        RECT 0.935 9.785 25.585 9.855 ;
        RECT 0.935 9.855 25.655 9.925 ;
        RECT 0.935 9.925 25.725 9.995 ;
        RECT 0.935 9.995 25.795 10.065 ;
        RECT 0.935 10.065 25.865 10.135 ;
        RECT 0.935 10.135 25.935 10.205 ;
        RECT 0.935 10.205 26.005 10.275 ;
        RECT 0.935 10.275 26.075 10.345 ;
        RECT 0.935 10.345 26.145 10.415 ;
        RECT 0.935 10.415 26.215 10.485 ;
        RECT 0.935 10.485 26.285 10.555 ;
        RECT 0.935 10.555 26.355 10.625 ;
        RECT 0.935 10.625 26.425 10.695 ;
        RECT 0.935 10.695 26.495 10.765 ;
        RECT 0.935 10.765 26.565 10.835 ;
        RECT 0.935 10.835 26.635 10.905 ;
        RECT 0.935 10.905 26.705 10.975 ;
        RECT 0.935 10.975 26.775 11.045 ;
        RECT 0.935 11.045 26.845 11.115 ;
        RECT 0.935 11.115 26.915 11.185 ;
        RECT 0.935 11.185 26.985 11.255 ;
        RECT 0.935 11.255 27.055 11.325 ;
        RECT 0.935 11.325 27.125 11.395 ;
        RECT 0.935 11.395 27.195 11.465 ;
        RECT 0.935 11.465 27.265 11.535 ;
        RECT 0.935 11.535 27.335 11.605 ;
        RECT 0.935 11.605 27.405 11.675 ;
        RECT 0.935 11.675 27.475 11.745 ;
        RECT 0.935 11.745 27.545 11.815 ;
        RECT 0.935 11.815 27.615 11.885 ;
        RECT 0.935 11.885 27.685 11.955 ;
        RECT 0.935 11.955 27.755 12.025 ;
        RECT 0.935 12.025 27.825 12.095 ;
        RECT 0.935 12.095 27.895 12.165 ;
        RECT 0.935 12.165 27.965 12.235 ;
        RECT 0.935 12.235 28.035 12.305 ;
        RECT 0.935 12.305 28.105 12.375 ;
        RECT 0.935 12.375 28.175 12.4 ;
        RECT 0.935 2.495 24.395 8.595 ;
        RECT 0.565 2.055 24.395 2.125 ;
        RECT 0.635 2.125 24.395 2.195 ;
        RECT 0.705 2.195 24.395 2.265 ;
        RECT 0.775 2.265 24.395 2.335 ;
        RECT 0.845 2.335 24.395 2.405 ;
        RECT 0.915 2.405 24.395 2.475 ;
        RECT 0.935 2.475 24.395 2.495 ;
        RECT 0.495 0 24.395 2.055 ;
    END
  END src_bdy_hvc

  PIN drn_hvc
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 37.89 0 48.89 96.15 ;
        RECT 37.89 96.15 48.89 96.3 ;
        RECT 37.89 96.3 49.04 96.45 ;
        RECT 37.89 96.45 49.19 96.6 ;
        RECT 37.89 96.6 49.34 96.75 ;
        RECT 37.89 96.75 49.49 96.9 ;
        RECT 37.89 96.9 49.64 97.05 ;
        RECT 37.89 97.05 49.79 97.2 ;
        RECT 37.89 97.2 49.94 97.35 ;
        RECT 37.89 97.35 50.09 97.5 ;
        RECT 37.89 97.5 50.24 97.65 ;
        RECT 37.89 97.65 50.39 97.8 ;
        RECT 37.89 97.8 50.54 97.95 ;
        RECT 37.89 97.95 50.69 98.1 ;
        RECT 37.89 98.1 50.84 98.25 ;
        RECT 37.89 98.25 50.99 98.3 ;
        RECT 37.89 98.3 51.04 99.505 ;
        RECT 44.73 99.505 51.04 99.61 ;
        RECT 44.835 99.61 51.04 99.715 ;
        RECT 45.35 100.23 51.555 100.38 ;
        RECT 45.35 100.38 51.705 100.53 ;
        RECT 45.35 100.53 51.855 100.68 ;
        RECT 45.35 100.68 52.005 100.83 ;
        RECT 45.35 100.83 52.155 100.98 ;
        RECT 45.35 100.98 52.305 101.13 ;
        RECT 45.35 101.13 52.455 101.28 ;
        RECT 45.35 101.28 52.605 101.43 ;
        RECT 45.35 101.43 52.755 101.58 ;
        RECT 45.35 101.58 52.905 101.73 ;
        RECT 45.35 101.73 53.055 101.88 ;
        RECT 45.35 101.88 53.205 102.03 ;
        RECT 45.35 102.03 53.355 102.18 ;
        RECT 45.35 102.18 53.505 102.33 ;
        RECT 45.35 102.33 53.655 102.48 ;
        RECT 45.35 102.48 53.805 102.505 ;
        RECT 44.985 99.715 51.04 99.865 ;
        RECT 45.135 99.865 51.19 100.015 ;
        RECT 45.285 100.015 51.34 100.165 ;
        RECT 45.35 100.165 51.49 100.23 ;
        RECT 37.89 99.505 43.47 99.655 ;
        RECT 37.89 99.655 43.32 99.805 ;
        RECT 37.89 99.805 43.17 99.955 ;
        RECT 37.89 99.955 43.02 100.105 ;
        RECT 37.89 100.105 42.87 100.255 ;
        RECT 37.89 100.255 42.84 100.285 ;
        RECT 37.89 100.285 42.84 102.135 ;
        RECT 37.89 102.135 42.84 102.285 ;
        RECT 37.89 102.285 42.99 102.435 ;
        RECT 37.89 102.435 43.14 102.585 ;
        RECT 37.89 102.585 43.29 102.735 ;
        RECT 37.89 102.735 43.44 102.885 ;
        RECT 37.89 102.885 43.59 103.035 ;
        RECT 37.89 103.035 43.74 103.185 ;
        RECT 37.89 103.185 43.89 103.335 ;
        RECT 37.89 103.335 44.04 103.485 ;
        RECT 37.89 103.485 44.19 103.635 ;
        RECT 37.89 103.635 44.34 103.785 ;
        RECT 37.89 103.785 44.49 103.935 ;
        RECT 37.89 103.935 44.64 104.085 ;
        RECT 37.89 104.085 44.79 104.235 ;
        RECT 37.89 104.235 44.94 104.385 ;
        RECT 37.89 104.385 45.09 104.535 ;
        RECT 37.89 104.535 45.24 104.685 ;
        RECT 37.89 104.685 45.39 104.835 ;
        RECT 37.89 104.835 45.54 104.985 ;
        RECT 37.89 104.985 45.69 105.135 ;
        RECT 37.89 105.135 45.84 105.285 ;
        RECT 37.89 105.285 45.99 105.435 ;
        RECT 37.89 105.435 46.14 105.585 ;
        RECT 37.89 105.585 46.29 105.655 ;
        RECT 45.5 102.505 53.83 102.655 ;
        RECT 45.65 102.655 53.98 102.805 ;
        RECT 45.8 102.805 54.13 102.955 ;
        RECT 45.95 102.955 54.28 103.105 ;
        RECT 46.1 103.105 54.43 103.255 ;
        RECT 46.25 103.255 54.58 103.405 ;
        RECT 46.4 103.405 54.73 103.555 ;
        RECT 46.55 103.555 54.88 103.705 ;
        RECT 46.7 103.705 55.03 103.855 ;
        RECT 46.85 103.855 55.18 104.005 ;
        RECT 47 104.005 55.33 104.155 ;
        RECT 47.15 104.155 55.48 104.305 ;
        RECT 47.3 104.305 55.63 104.455 ;
        RECT 47.45 104.455 55.78 104.605 ;
        RECT 47.6 104.605 55.93 104.755 ;
        RECT 47.75 104.755 56.08 104.905 ;
        RECT 47.9 104.905 56.23 105.055 ;
        RECT 48.05 105.055 56.38 105.205 ;
        RECT 48.2 105.205 56.53 105.355 ;
        RECT 48.35 105.355 56.68 105.505 ;
        RECT 48.5 105.505 56.83 105.655 ;
        RECT 48.65 105.655 56.98 105.805 ;
        RECT 48.8 105.805 57.13 105.955 ;
        RECT 48.95 105.955 57.28 106.105 ;
        RECT 49.1 106.105 57.43 106.255 ;
        RECT 49.25 106.255 57.58 106.405 ;
        RECT 49.4 106.405 57.73 106.555 ;
        RECT 49.55 106.555 57.88 106.705 ;
        RECT 49.7 106.705 58.03 106.855 ;
        RECT 49.85 106.855 58.18 107.005 ;
        RECT 50 107.005 58.33 107.155 ;
        RECT 50.15 107.155 58.48 107.305 ;
        RECT 50.3 107.305 58.63 107.455 ;
        RECT 50.45 107.455 58.78 107.605 ;
        RECT 50.6 107.605 58.93 107.755 ;
        RECT 50.75 107.755 59.08 107.905 ;
        RECT 50.805 107.905 59.23 107.96 ;
        RECT 38.04 105.655 46.36 105.805 ;
        RECT 38.19 105.805 46.51 105.955 ;
        RECT 38.34 105.955 46.66 106.105 ;
        RECT 38.49 106.105 46.81 106.255 ;
        RECT 38.64 106.255 46.96 106.405 ;
        RECT 38.79 106.405 47.11 106.555 ;
        RECT 38.94 106.555 47.26 106.705 ;
        RECT 39.09 106.705 47.41 106.855 ;
        RECT 39.24 106.855 47.56 107.005 ;
        RECT 39.39 107.005 47.71 107.155 ;
        RECT 39.54 107.155 47.86 107.305 ;
        RECT 39.69 107.305 48.01 107.455 ;
        RECT 39.84 107.455 48.16 107.605 ;
        RECT 39.99 107.605 48.31 107.755 ;
        RECT 40.14 107.755 48.46 107.905 ;
        RECT 40.29 107.905 48.61 108.055 ;
        RECT 40.385 108.055 48.76 108.15 ;
        RECT 50.955 107.96 59.285 108.11 ;
        RECT 51.105 108.11 59.285 108.26 ;
        RECT 51.255 108.26 59.285 108.41 ;
        RECT 51.405 108.41 59.285 108.56 ;
        RECT 51.555 108.56 59.285 108.71 ;
        RECT 51.705 108.71 59.285 108.86 ;
        RECT 51.855 108.86 59.285 109.01 ;
        RECT 52.005 109.01 59.285 109.16 ;
        RECT 52.155 109.16 59.285 109.31 ;
        RECT 52.305 109.31 59.285 109.46 ;
        RECT 52.455 109.46 59.285 109.61 ;
        RECT 52.605 109.61 59.285 109.76 ;
        RECT 52.755 109.76 59.285 109.91 ;
        RECT 52.905 109.91 59.285 110.06 ;
        RECT 53.055 110.06 59.285 110.21 ;
        RECT 53.205 110.21 59.285 110.36 ;
        RECT 53.285 110.36 59.285 110.44 ;
        RECT 40.535 108.15 48.855 108.3 ;
        RECT 40.685 108.3 48.855 108.45 ;
        RECT 40.835 108.45 48.855 108.6 ;
        RECT 40.985 108.6 48.855 108.75 ;
        RECT 41.135 108.75 48.855 108.9 ;
        RECT 41.285 108.9 48.855 109.05 ;
        RECT 41.435 109.05 48.855 109.2 ;
        RECT 41.585 109.2 48.855 109.35 ;
        RECT 41.735 109.35 48.855 109.5 ;
        RECT 41.885 109.5 48.855 109.65 ;
        RECT 42.035 109.65 48.855 109.8 ;
        RECT 42.185 109.8 48.855 109.95 ;
        RECT 42.335 109.95 48.855 110.1 ;
        RECT 42.485 110.1 48.855 110.25 ;
        RECT 42.635 110.25 48.855 110.4 ;
        RECT 42.785 110.4 48.855 110.55 ;
        RECT 42.855 110.55 48.855 110.62 ;
        RECT 53.285 169.135 59.285 169.285 ;
        RECT 53.135 169.285 59.285 169.435 ;
        RECT 52.985 169.435 59.285 169.585 ;
        RECT 52.835 169.585 59.285 169.735 ;
        RECT 52.685 169.735 59.285 169.885 ;
        RECT 52.535 169.885 59.285 170.035 ;
        RECT 52.385 170.035 59.285 170.185 ;
        RECT 52.235 170.185 59.285 170.335 ;
        RECT 52.085 170.335 59.285 170.485 ;
        RECT 51.935 170.485 59.285 170.635 ;
        RECT 51.785 170.635 59.285 170.785 ;
        RECT 51.635 170.785 59.285 170.935 ;
        RECT 51.485 170.935 59.285 171.085 ;
        RECT 51.335 171.085 59.285 171.235 ;
        RECT 51.185 171.235 59.285 171.385 ;
        RECT 51.035 171.385 59.285 171.535 ;
        RECT 50.885 171.535 59.285 171.685 ;
        RECT 50.735 171.685 59.285 171.835 ;
        RECT 50.585 171.835 59.285 171.985 ;
        RECT 50.435 171.985 59.285 172.135 ;
        RECT 50.285 172.135 59.285 172.285 ;
        RECT 50.135 172.285 59.285 172.435 ;
        RECT 49.985 172.435 59.285 172.585 ;
        RECT 49.835 172.585 59.285 172.645 ;
        RECT 42.855 170.46 48.855 170.61 ;
        RECT 42.705 170.61 48.855 170.76 ;
        RECT 42.555 170.76 48.855 170.91 ;
        RECT 42.405 170.91 48.855 171.06 ;
        RECT 42.255 171.06 48.855 171.21 ;
        RECT 42.105 171.21 48.855 171.36 ;
        RECT 41.955 171.36 48.855 171.51 ;
        RECT 41.805 171.51 48.855 171.66 ;
        RECT 41.655 171.66 48.855 171.81 ;
        RECT 41.505 171.81 48.855 171.96 ;
        RECT 41.355 171.96 48.855 172.11 ;
        RECT 41.205 172.11 48.855 172.26 ;
        RECT 41.055 172.26 48.855 172.41 ;
        RECT 40.905 172.41 48.855 172.56 ;
        RECT 40.755 172.56 48.855 172.71 ;
        RECT 40.605 172.71 48.855 172.86 ;
        RECT 40.455 172.86 48.855 173.01 ;
        RECT 40.305 173.01 48.855 173.16 ;
        RECT 40.155 173.16 48.855 173.31 ;
        RECT 40.005 173.31 48.855 173.46 ;
        RECT 39.855 173.46 48.855 173.61 ;
        RECT 39.705 173.61 48.855 173.76 ;
        RECT 39.555 173.76 48.855 173.91 ;
        RECT 39.405 173.91 48.855 174.06 ;
        RECT 39.255 174.06 48.855 174.21 ;
        RECT 39.105 174.21 48.855 174.36 ;
        RECT 38.955 174.36 48.855 174.51 ;
        RECT 38.805 174.51 48.855 174.66 ;
        RECT 38.655 174.66 48.855 174.81 ;
        RECT 38.505 174.81 48.855 174.96 ;
        RECT 38.355 174.96 48.855 175.11 ;
        RECT 38.205 175.11 48.855 175.26 ;
        RECT 38.055 175.26 48.855 175.35 ;
        RECT 49.775 172.645 59.285 173.02 ;
        RECT 37.965 175.35 48.855 190.02 ;
        RECT 49.775 173.02 59.285 173.17 ;
        RECT 49.775 173.17 59.435 173.32 ;
        RECT 49.775 173.32 59.585 173.47 ;
        RECT 49.775 173.47 59.735 173.62 ;
        RECT 49.775 173.62 59.885 173.77 ;
        RECT 49.775 173.77 60.035 173.92 ;
        RECT 49.775 173.92 60.185 174.07 ;
        RECT 49.775 174.07 60.335 174.22 ;
        RECT 49.775 174.22 60.485 174.37 ;
        RECT 49.775 174.37 60.635 174.52 ;
        RECT 49.775 174.52 60.785 174.67 ;
        RECT 49.775 174.67 60.935 174.82 ;
        RECT 49.775 174.82 61.085 174.97 ;
        RECT 49.775 174.97 61.235 175.12 ;
        RECT 49.775 175.12 61.385 175.225 ;
        RECT 49.775 175.225 61.49 190.04 ;
        RECT 53.285 110.44 59.285 169.135 ;
        RECT 42.855 110.62 48.855 170.46 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.62 185.295 74.29 190.015 ;
        RECT 61.11 182.88 74.29 182.95 ;
        RECT 61.04 182.95 74.29 183.02 ;
        RECT 60.97 183.02 74.29 183.09 ;
        RECT 60.9 183.09 74.29 183.16 ;
        RECT 60.83 183.16 74.29 183.23 ;
        RECT 60.76 183.23 74.29 183.3 ;
        RECT 60.69 183.3 74.29 183.37 ;
        RECT 60.62 183.37 74.29 183.44 ;
        RECT 60.55 183.44 74.29 183.51 ;
        RECT 60.48 183.51 74.29 183.58 ;
        RECT 60.41 183.58 74.29 183.65 ;
        RECT 60.34 183.65 74.29 183.72 ;
        RECT 60.27 183.72 74.29 183.79 ;
        RECT 60.2 183.79 74.29 183.86 ;
        RECT 60.13 183.86 74.29 183.93 ;
        RECT 60.06 183.93 74.29 184 ;
        RECT 59.99 184 74.29 184.07 ;
        RECT 59.92 184.07 74.29 184.14 ;
        RECT 59.85 184.14 74.29 184.21 ;
        RECT 59.78 184.21 74.29 184.28 ;
        RECT 59.71 184.28 74.29 184.35 ;
        RECT 59.64 184.35 74.29 184.42 ;
        RECT 59.57 184.42 74.29 184.49 ;
        RECT 59.5 184.49 74.29 184.56 ;
        RECT 59.43 184.56 74.29 184.63 ;
        RECT 59.36 184.63 74.29 184.7 ;
        RECT 59.29 184.7 74.29 184.77 ;
        RECT 59.22 184.77 74.29 184.84 ;
        RECT 59.15 184.84 74.29 184.91 ;
        RECT 59.08 184.91 74.29 184.98 ;
        RECT 59.01 184.98 74.29 185.05 ;
        RECT 58.94 185.05 74.29 185.12 ;
        RECT 58.87 185.12 74.29 185.19 ;
        RECT 58.8 185.19 74.29 185.26 ;
        RECT 58.73 185.26 74.29 185.295 ;
        RECT 61.11 174.7 74.29 182.88 ;
        RECT 57.635 171.155 74.29 171.225 ;
        RECT 57.705 171.225 74.29 171.295 ;
        RECT 57.775 171.295 74.29 171.365 ;
        RECT 57.845 171.365 74.29 171.435 ;
        RECT 57.915 171.435 74.29 171.505 ;
        RECT 57.985 171.505 74.29 171.575 ;
        RECT 58.055 171.575 74.29 171.645 ;
        RECT 58.125 171.645 74.29 171.715 ;
        RECT 58.195 171.715 74.29 171.785 ;
        RECT 58.265 171.785 74.29 171.855 ;
        RECT 58.335 171.855 74.29 171.925 ;
        RECT 58.405 171.925 74.29 171.995 ;
        RECT 58.475 171.995 74.29 172.065 ;
        RECT 58.545 172.065 74.29 172.135 ;
        RECT 58.615 172.135 74.29 172.205 ;
        RECT 58.685 172.205 74.29 172.275 ;
        RECT 58.755 172.275 74.29 172.345 ;
        RECT 58.825 172.345 74.29 172.415 ;
        RECT 58.895 172.415 74.29 172.485 ;
        RECT 58.965 172.485 74.29 172.555 ;
        RECT 59.035 172.555 74.29 172.625 ;
        RECT 59.105 172.625 74.29 172.695 ;
        RECT 59.175 172.695 74.29 172.765 ;
        RECT 59.245 172.765 74.29 172.835 ;
        RECT 59.315 172.835 74.29 172.905 ;
        RECT 59.385 172.905 74.29 172.975 ;
        RECT 59.455 172.975 74.29 173.045 ;
        RECT 59.525 173.045 74.29 173.115 ;
        RECT 59.595 173.115 74.29 173.185 ;
        RECT 59.665 173.185 74.29 173.255 ;
        RECT 59.735 173.255 74.29 173.325 ;
        RECT 59.805 173.325 74.29 173.395 ;
        RECT 59.875 173.395 74.29 173.465 ;
        RECT 59.945 173.465 74.29 173.535 ;
        RECT 60.015 173.535 74.29 173.605 ;
        RECT 60.085 173.605 74.29 173.675 ;
        RECT 60.155 173.675 74.29 173.745 ;
        RECT 60.225 173.745 74.29 173.815 ;
        RECT 60.295 173.815 74.29 173.885 ;
        RECT 60.365 173.885 74.29 173.955 ;
        RECT 60.435 173.955 74.29 174.025 ;
        RECT 60.505 174.025 74.29 174.095 ;
        RECT 60.575 174.095 74.29 174.165 ;
        RECT 60.645 174.165 74.29 174.235 ;
        RECT 60.715 174.235 74.29 174.305 ;
        RECT 60.785 174.305 74.29 174.375 ;
        RECT 60.855 174.375 74.29 174.445 ;
        RECT 60.925 174.445 74.29 174.515 ;
        RECT 60.995 174.515 74.29 174.585 ;
        RECT 61.065 174.585 74.29 174.655 ;
        RECT 61.11 174.655 74.29 174.7 ;
        RECT 16.805 162.455 74.29 171.155 ;
        RECT 61.11 158.87 74.29 158.94 ;
        RECT 61.04 158.94 74.29 159.01 ;
        RECT 60.97 159.01 74.29 159.08 ;
        RECT 60.9 159.08 74.29 159.15 ;
        RECT 60.83 159.15 74.29 159.22 ;
        RECT 60.76 159.22 74.29 159.29 ;
        RECT 60.69 159.29 74.29 159.36 ;
        RECT 60.62 159.36 74.29 159.43 ;
        RECT 60.55 159.43 74.29 159.5 ;
        RECT 60.48 159.5 74.29 159.57 ;
        RECT 60.41 159.57 74.29 159.64 ;
        RECT 60.34 159.64 74.29 159.71 ;
        RECT 60.27 159.71 74.29 159.78 ;
        RECT 60.2 159.78 74.29 159.85 ;
        RECT 60.13 159.85 74.29 159.92 ;
        RECT 60.06 159.92 74.29 159.99 ;
        RECT 59.99 159.99 74.29 160.06 ;
        RECT 59.92 160.06 74.29 160.13 ;
        RECT 59.85 160.13 74.29 160.2 ;
        RECT 59.78 160.2 74.29 160.27 ;
        RECT 59.71 160.27 74.29 160.34 ;
        RECT 59.64 160.34 74.29 160.41 ;
        RECT 59.57 160.41 74.29 160.48 ;
        RECT 59.5 160.48 74.29 160.55 ;
        RECT 59.43 160.55 74.29 160.62 ;
        RECT 59.36 160.62 74.29 160.69 ;
        RECT 59.29 160.69 74.29 160.76 ;
        RECT 59.22 160.76 74.29 160.83 ;
        RECT 59.15 160.83 74.29 160.9 ;
        RECT 59.08 160.9 74.29 160.97 ;
        RECT 59.01 160.97 74.29 161.04 ;
        RECT 58.94 161.04 74.29 161.11 ;
        RECT 58.87 161.11 74.29 161.18 ;
        RECT 58.8 161.18 74.29 161.25 ;
        RECT 58.73 161.25 74.29 161.32 ;
        RECT 58.66 161.32 74.29 161.39 ;
        RECT 58.59 161.39 74.29 161.46 ;
        RECT 58.52 161.46 74.29 161.53 ;
        RECT 58.45 161.53 74.29 161.6 ;
        RECT 58.38 161.6 74.29 161.67 ;
        RECT 58.31 161.67 74.29 161.74 ;
        RECT 58.24 161.74 74.29 161.81 ;
        RECT 58.17 161.81 74.29 161.88 ;
        RECT 58.1 161.88 74.29 161.95 ;
        RECT 58.03 161.95 74.29 162.02 ;
        RECT 57.96 162.02 74.29 162.09 ;
        RECT 57.89 162.09 74.29 162.16 ;
        RECT 57.82 162.16 74.29 162.23 ;
        RECT 57.75 162.23 74.29 162.3 ;
        RECT 57.68 162.3 74.29 162.37 ;
        RECT 57.61 162.37 74.29 162.44 ;
        RECT 57.54 162.44 74.29 162.455 ;
        RECT 61.11 151.78 74.29 158.87 ;
        RECT 57.555 148.155 74.29 148.225 ;
        RECT 57.625 148.225 74.29 148.295 ;
        RECT 57.695 148.295 74.29 148.365 ;
        RECT 57.765 148.365 74.29 148.435 ;
        RECT 57.835 148.435 74.29 148.505 ;
        RECT 57.905 148.505 74.29 148.575 ;
        RECT 57.975 148.575 74.29 148.645 ;
        RECT 58.045 148.645 74.29 148.715 ;
        RECT 58.115 148.715 74.29 148.785 ;
        RECT 58.185 148.785 74.29 148.855 ;
        RECT 58.255 148.855 74.29 148.925 ;
        RECT 58.325 148.925 74.29 148.995 ;
        RECT 58.395 148.995 74.29 149.065 ;
        RECT 58.465 149.065 74.29 149.135 ;
        RECT 58.535 149.135 74.29 149.205 ;
        RECT 58.605 149.205 74.29 149.275 ;
        RECT 58.675 149.275 74.29 149.345 ;
        RECT 58.745 149.345 74.29 149.415 ;
        RECT 58.815 149.415 74.29 149.485 ;
        RECT 58.885 149.485 74.29 149.555 ;
        RECT 58.955 149.555 74.29 149.625 ;
        RECT 59.025 149.625 74.29 149.695 ;
        RECT 59.095 149.695 74.29 149.765 ;
        RECT 59.165 149.765 74.29 149.835 ;
        RECT 59.235 149.835 74.29 149.905 ;
        RECT 59.305 149.905 74.29 149.975 ;
        RECT 59.375 149.975 74.29 150.045 ;
        RECT 59.445 150.045 74.29 150.115 ;
        RECT 59.515 150.115 74.29 150.185 ;
        RECT 59.585 150.185 74.29 150.255 ;
        RECT 59.655 150.255 74.29 150.325 ;
        RECT 59.725 150.325 74.29 150.395 ;
        RECT 59.795 150.395 74.29 150.465 ;
        RECT 59.865 150.465 74.29 150.535 ;
        RECT 59.935 150.535 74.29 150.605 ;
        RECT 60.005 150.605 74.29 150.675 ;
        RECT 60.075 150.675 74.29 150.745 ;
        RECT 60.145 150.745 74.29 150.815 ;
        RECT 60.215 150.815 74.29 150.885 ;
        RECT 60.285 150.885 74.29 150.955 ;
        RECT 60.355 150.955 74.29 151.025 ;
        RECT 60.425 151.025 74.29 151.095 ;
        RECT 60.495 151.095 74.29 151.165 ;
        RECT 60.565 151.165 74.29 151.235 ;
        RECT 60.635 151.235 74.29 151.305 ;
        RECT 60.705 151.305 74.29 151.375 ;
        RECT 60.775 151.375 74.29 151.445 ;
        RECT 60.845 151.445 74.29 151.515 ;
        RECT 60.915 151.515 74.29 151.585 ;
        RECT 60.985 151.585 74.29 151.655 ;
        RECT 61.055 151.655 74.29 151.725 ;
        RECT 61.11 151.725 74.29 151.78 ;
        RECT 16.875 146.71 74.29 146.78 ;
        RECT 16.945 146.78 74.29 146.85 ;
        RECT 17.015 146.85 74.29 146.92 ;
        RECT 17.085 146.92 74.29 146.99 ;
        RECT 17.155 146.99 74.29 147.06 ;
        RECT 17.225 147.06 74.29 147.13 ;
        RECT 17.295 147.13 74.29 147.2 ;
        RECT 17.365 147.2 74.29 147.27 ;
        RECT 17.435 147.27 74.29 147.34 ;
        RECT 17.505 147.34 74.29 147.41 ;
        RECT 17.575 147.41 74.29 147.48 ;
        RECT 17.645 147.48 74.29 147.55 ;
        RECT 17.715 147.55 74.29 147.62 ;
        RECT 17.785 147.62 74.29 147.69 ;
        RECT 17.855 147.69 74.29 147.76 ;
        RECT 17.925 147.76 74.29 147.83 ;
        RECT 17.995 147.83 74.29 147.9 ;
        RECT 18.065 147.9 74.29 147.97 ;
        RECT 18.135 147.97 74.29 148.04 ;
        RECT 18.205 148.04 74.29 148.11 ;
        RECT 18.25 148.11 74.29 148.155 ;
        RECT 16.805 139.455 74.29 146.71 ;
        RECT 61.11 135.855 74.29 135.925 ;
        RECT 61.04 135.925 74.29 135.995 ;
        RECT 60.97 135.995 74.29 136.065 ;
        RECT 60.9 136.065 74.29 136.135 ;
        RECT 60.83 136.135 74.29 136.205 ;
        RECT 60.76 136.205 74.29 136.275 ;
        RECT 60.69 136.275 74.29 136.345 ;
        RECT 60.62 136.345 74.29 136.415 ;
        RECT 60.55 136.415 74.29 136.485 ;
        RECT 60.48 136.485 74.29 136.555 ;
        RECT 60.41 136.555 74.29 136.625 ;
        RECT 60.34 136.625 74.29 136.695 ;
        RECT 60.27 136.695 74.29 136.765 ;
        RECT 60.2 136.765 74.29 136.835 ;
        RECT 60.13 136.835 74.29 136.905 ;
        RECT 60.06 136.905 74.29 136.975 ;
        RECT 59.99 136.975 74.29 137.045 ;
        RECT 59.92 137.045 74.29 137.115 ;
        RECT 59.85 137.115 74.29 137.185 ;
        RECT 59.78 137.185 74.29 137.255 ;
        RECT 59.71 137.255 74.29 137.325 ;
        RECT 59.64 137.325 74.29 137.395 ;
        RECT 59.57 137.395 74.29 137.465 ;
        RECT 59.5 137.465 74.29 137.535 ;
        RECT 59.43 137.535 74.29 137.605 ;
        RECT 59.36 137.605 74.29 137.675 ;
        RECT 59.29 137.675 74.29 137.745 ;
        RECT 59.22 137.745 74.29 137.815 ;
        RECT 59.15 137.815 74.29 137.885 ;
        RECT 59.08 137.885 74.29 137.955 ;
        RECT 59.01 137.955 74.29 138.025 ;
        RECT 58.94 138.025 74.29 138.095 ;
        RECT 58.87 138.095 74.29 138.165 ;
        RECT 58.8 138.165 74.29 138.235 ;
        RECT 58.73 138.235 74.29 138.305 ;
        RECT 58.66 138.305 74.29 138.375 ;
        RECT 58.59 138.375 74.29 138.445 ;
        RECT 58.52 138.445 74.29 138.515 ;
        RECT 58.45 138.515 74.29 138.585 ;
        RECT 58.38 138.585 74.29 138.655 ;
        RECT 58.31 138.655 74.29 138.725 ;
        RECT 58.24 138.725 74.29 138.795 ;
        RECT 58.17 138.795 74.29 138.865 ;
        RECT 58.1 138.865 74.29 138.935 ;
        RECT 58.03 138.935 74.29 139.005 ;
        RECT 57.96 139.005 74.29 139.075 ;
        RECT 57.89 139.075 74.29 139.145 ;
        RECT 57.82 139.145 74.29 139.215 ;
        RECT 57.75 139.215 74.29 139.285 ;
        RECT 57.68 139.285 74.29 139.355 ;
        RECT 57.61 139.355 74.29 139.425 ;
        RECT 57.54 139.425 74.29 139.455 ;
        RECT 61.11 128.71 74.29 135.855 ;
        RECT 57.625 125.155 74.29 125.225 ;
        RECT 57.695 125.225 74.29 125.295 ;
        RECT 57.765 125.295 74.29 125.365 ;
        RECT 57.835 125.365 74.29 125.435 ;
        RECT 57.905 125.435 74.29 125.505 ;
        RECT 57.975 125.505 74.29 125.575 ;
        RECT 58.045 125.575 74.29 125.645 ;
        RECT 58.115 125.645 74.29 125.715 ;
        RECT 58.185 125.715 74.29 125.785 ;
        RECT 58.255 125.785 74.29 125.855 ;
        RECT 58.325 125.855 74.29 125.925 ;
        RECT 58.395 125.925 74.29 125.995 ;
        RECT 58.465 125.995 74.29 126.065 ;
        RECT 58.535 126.065 74.29 126.135 ;
        RECT 58.605 126.135 74.29 126.205 ;
        RECT 58.675 126.205 74.29 126.275 ;
        RECT 58.745 126.275 74.29 126.345 ;
        RECT 58.815 126.345 74.29 126.415 ;
        RECT 58.885 126.415 74.29 126.485 ;
        RECT 58.955 126.485 74.29 126.555 ;
        RECT 59.025 126.555 74.29 126.625 ;
        RECT 59.095 126.625 74.29 126.695 ;
        RECT 59.165 126.695 74.29 126.765 ;
        RECT 59.235 126.765 74.29 126.835 ;
        RECT 59.305 126.835 74.29 126.905 ;
        RECT 59.375 126.905 74.29 126.975 ;
        RECT 59.445 126.975 74.29 127.045 ;
        RECT 59.515 127.045 74.29 127.115 ;
        RECT 59.585 127.115 74.29 127.185 ;
        RECT 59.655 127.185 74.29 127.255 ;
        RECT 59.725 127.255 74.29 127.325 ;
        RECT 59.795 127.325 74.29 127.395 ;
        RECT 59.865 127.395 74.29 127.465 ;
        RECT 59.935 127.465 74.29 127.535 ;
        RECT 60.005 127.535 74.29 127.605 ;
        RECT 60.075 127.605 74.29 127.675 ;
        RECT 60.145 127.675 74.29 127.745 ;
        RECT 60.215 127.745 74.29 127.815 ;
        RECT 60.285 127.815 74.29 127.885 ;
        RECT 60.355 127.885 74.29 127.955 ;
        RECT 60.425 127.955 74.29 128.025 ;
        RECT 60.495 128.025 74.29 128.095 ;
        RECT 60.565 128.095 74.29 128.165 ;
        RECT 60.635 128.165 74.29 128.235 ;
        RECT 60.705 128.235 74.29 128.305 ;
        RECT 60.775 128.305 74.29 128.375 ;
        RECT 60.845 128.375 74.29 128.445 ;
        RECT 60.915 128.445 74.29 128.515 ;
        RECT 60.985 128.515 74.29 128.585 ;
        RECT 61.055 128.585 74.29 128.655 ;
        RECT 61.11 128.655 74.29 128.71 ;
        RECT 24.82 116.455 74.29 125.155 ;
        RECT 61.11 112.82 74.29 112.89 ;
        RECT 61.04 112.89 74.29 112.96 ;
        RECT 60.97 112.96 74.29 113.03 ;
        RECT 60.9 113.03 74.29 113.1 ;
        RECT 60.83 113.1 74.29 113.17 ;
        RECT 60.76 113.17 74.29 113.24 ;
        RECT 60.69 113.24 74.29 113.31 ;
        RECT 60.62 113.31 74.29 113.38 ;
        RECT 60.55 113.38 74.29 113.45 ;
        RECT 60.48 113.45 74.29 113.52 ;
        RECT 60.41 113.52 74.29 113.59 ;
        RECT 60.34 113.59 74.29 113.66 ;
        RECT 60.27 113.66 74.29 113.73 ;
        RECT 60.2 113.73 74.29 113.8 ;
        RECT 60.13 113.8 74.29 113.87 ;
        RECT 60.06 113.87 74.29 113.94 ;
        RECT 59.99 113.94 74.29 114.01 ;
        RECT 59.92 114.01 74.29 114.08 ;
        RECT 59.85 114.08 74.29 114.15 ;
        RECT 59.78 114.15 74.29 114.22 ;
        RECT 59.71 114.22 74.29 114.29 ;
        RECT 59.64 114.29 74.29 114.36 ;
        RECT 59.57 114.36 74.29 114.43 ;
        RECT 59.5 114.43 74.29 114.5 ;
        RECT 59.43 114.5 74.29 114.57 ;
        RECT 59.36 114.57 74.29 114.64 ;
        RECT 59.29 114.64 74.29 114.71 ;
        RECT 59.22 114.71 74.29 114.78 ;
        RECT 59.15 114.78 74.29 114.85 ;
        RECT 59.08 114.85 74.29 114.92 ;
        RECT 59.01 114.92 74.29 114.99 ;
        RECT 58.94 114.99 74.29 115.06 ;
        RECT 58.87 115.06 74.29 115.13 ;
        RECT 58.8 115.13 74.29 115.2 ;
        RECT 58.73 115.2 74.29 115.27 ;
        RECT 58.66 115.27 74.29 115.34 ;
        RECT 58.59 115.34 74.29 115.41 ;
        RECT 58.52 115.41 74.29 115.48 ;
        RECT 58.45 115.48 74.29 115.55 ;
        RECT 58.38 115.55 74.29 115.62 ;
        RECT 58.31 115.62 74.29 115.69 ;
        RECT 58.24 115.69 74.29 115.76 ;
        RECT 58.17 115.76 74.29 115.83 ;
        RECT 58.1 115.83 74.29 115.9 ;
        RECT 58.03 115.9 74.29 115.97 ;
        RECT 57.96 115.97 74.29 116.04 ;
        RECT 57.89 116.04 74.29 116.11 ;
        RECT 57.82 116.11 74.29 116.18 ;
        RECT 57.75 116.18 74.29 116.25 ;
        RECT 57.68 116.25 74.29 116.32 ;
        RECT 57.61 116.32 74.29 116.39 ;
        RECT 57.54 116.39 74.29 116.455 ;
        RECT 61.11 105.71 74.29 112.82 ;
        RECT 57.625 102.155 74.29 102.225 ;
        RECT 57.695 102.225 74.29 102.295 ;
        RECT 57.765 102.295 74.29 102.365 ;
        RECT 57.835 102.365 74.29 102.435 ;
        RECT 57.905 102.435 74.29 102.505 ;
        RECT 57.975 102.505 74.29 102.575 ;
        RECT 58.045 102.575 74.29 102.645 ;
        RECT 58.115 102.645 74.29 102.715 ;
        RECT 58.185 102.715 74.29 102.785 ;
        RECT 58.255 102.785 74.29 102.855 ;
        RECT 58.325 102.855 74.29 102.925 ;
        RECT 58.395 102.925 74.29 102.995 ;
        RECT 58.465 102.995 74.29 103.065 ;
        RECT 58.535 103.065 74.29 103.135 ;
        RECT 58.605 103.135 74.29 103.205 ;
        RECT 58.675 103.205 74.29 103.275 ;
        RECT 58.745 103.275 74.29 103.345 ;
        RECT 58.815 103.345 74.29 103.415 ;
        RECT 58.885 103.415 74.29 103.485 ;
        RECT 58.955 103.485 74.29 103.555 ;
        RECT 59.025 103.555 74.29 103.625 ;
        RECT 59.095 103.625 74.29 103.695 ;
        RECT 59.165 103.695 74.29 103.765 ;
        RECT 59.235 103.765 74.29 103.835 ;
        RECT 59.305 103.835 74.29 103.905 ;
        RECT 59.375 103.905 74.29 103.975 ;
        RECT 59.445 103.975 74.29 104.045 ;
        RECT 59.515 104.045 74.29 104.115 ;
        RECT 59.585 104.115 74.29 104.185 ;
        RECT 59.655 104.185 74.29 104.255 ;
        RECT 59.725 104.255 74.29 104.325 ;
        RECT 59.795 104.325 74.29 104.395 ;
        RECT 59.865 104.395 74.29 104.465 ;
        RECT 59.935 104.465 74.29 104.535 ;
        RECT 60.005 104.535 74.29 104.605 ;
        RECT 60.075 104.605 74.29 104.675 ;
        RECT 60.145 104.675 74.29 104.745 ;
        RECT 60.215 104.745 74.29 104.815 ;
        RECT 60.285 104.815 74.29 104.885 ;
        RECT 60.355 104.885 74.29 104.955 ;
        RECT 60.425 104.955 74.29 105.025 ;
        RECT 60.495 105.025 74.29 105.095 ;
        RECT 60.565 105.095 74.29 105.165 ;
        RECT 60.635 105.165 74.29 105.235 ;
        RECT 60.705 105.235 74.29 105.305 ;
        RECT 60.775 105.305 74.29 105.375 ;
        RECT 60.845 105.375 74.29 105.445 ;
        RECT 60.915 105.445 74.29 105.515 ;
        RECT 60.985 105.515 74.29 105.585 ;
        RECT 61.055 105.585 74.29 105.655 ;
        RECT 61.11 105.655 74.29 105.71 ;
        RECT 24.82 93.455 74.29 102.155 ;
        RECT 61.11 89.91 74.29 89.98 ;
        RECT 61.04 89.98 74.29 90.05 ;
        RECT 60.97 90.05 74.29 90.12 ;
        RECT 60.9 90.12 74.29 90.19 ;
        RECT 60.83 90.19 74.29 90.26 ;
        RECT 60.76 90.26 74.29 90.33 ;
        RECT 60.69 90.33 74.29 90.4 ;
        RECT 60.62 90.4 74.29 90.47 ;
        RECT 60.55 90.47 74.29 90.54 ;
        RECT 60.48 90.54 74.29 90.61 ;
        RECT 60.41 90.61 74.29 90.68 ;
        RECT 60.34 90.68 74.29 90.75 ;
        RECT 60.27 90.75 74.29 90.82 ;
        RECT 60.2 90.82 74.29 90.89 ;
        RECT 60.13 90.89 74.29 90.96 ;
        RECT 60.06 90.96 74.29 91.03 ;
        RECT 59.99 91.03 74.29 91.1 ;
        RECT 59.92 91.1 74.29 91.17 ;
        RECT 59.85 91.17 74.29 91.24 ;
        RECT 59.78 91.24 74.29 91.31 ;
        RECT 59.71 91.31 74.29 91.38 ;
        RECT 59.64 91.38 74.29 91.45 ;
        RECT 59.57 91.45 74.29 91.52 ;
        RECT 59.5 91.52 74.29 91.59 ;
        RECT 59.43 91.59 74.29 91.66 ;
        RECT 59.36 91.66 74.29 91.73 ;
        RECT 59.29 91.73 74.29 91.8 ;
        RECT 59.22 91.8 74.29 91.87 ;
        RECT 59.15 91.87 74.29 91.94 ;
        RECT 59.08 91.94 74.29 92.01 ;
        RECT 59.01 92.01 74.29 92.08 ;
        RECT 58.94 92.08 74.29 92.15 ;
        RECT 58.87 92.15 74.29 92.22 ;
        RECT 58.8 92.22 74.29 92.29 ;
        RECT 58.73 92.29 74.29 92.36 ;
        RECT 58.66 92.36 74.29 92.43 ;
        RECT 58.59 92.43 74.29 92.5 ;
        RECT 58.52 92.5 74.29 92.57 ;
        RECT 58.45 92.57 74.29 92.64 ;
        RECT 58.38 92.64 74.29 92.71 ;
        RECT 58.31 92.71 74.29 92.78 ;
        RECT 58.24 92.78 74.29 92.85 ;
        RECT 58.17 92.85 74.29 92.92 ;
        RECT 58.1 92.92 74.29 92.99 ;
        RECT 58.03 92.99 74.29 93.06 ;
        RECT 57.96 93.06 74.29 93.13 ;
        RECT 57.89 93.13 74.29 93.2 ;
        RECT 57.82 93.2 74.29 93.27 ;
        RECT 57.75 93.27 74.29 93.34 ;
        RECT 57.68 93.34 74.29 93.41 ;
        RECT 57.61 93.41 74.29 93.455 ;
        RECT 61.11 82.71 74.29 89.91 ;
        RECT 57.625 79.155 74.29 79.225 ;
        RECT 57.695 79.225 74.29 79.295 ;
        RECT 57.765 79.295 74.29 79.365 ;
        RECT 57.835 79.365 74.29 79.435 ;
        RECT 57.905 79.435 74.29 79.505 ;
        RECT 57.975 79.505 74.29 79.575 ;
        RECT 58.045 79.575 74.29 79.645 ;
        RECT 58.115 79.645 74.29 79.715 ;
        RECT 58.185 79.715 74.29 79.785 ;
        RECT 58.255 79.785 74.29 79.855 ;
        RECT 58.325 79.855 74.29 79.925 ;
        RECT 58.395 79.925 74.29 79.995 ;
        RECT 58.465 79.995 74.29 80.065 ;
        RECT 58.535 80.065 74.29 80.135 ;
        RECT 58.605 80.135 74.29 80.205 ;
        RECT 58.675 80.205 74.29 80.275 ;
        RECT 58.745 80.275 74.29 80.345 ;
        RECT 58.815 80.345 74.29 80.415 ;
        RECT 58.885 80.415 74.29 80.485 ;
        RECT 58.955 80.485 74.29 80.555 ;
        RECT 59.025 80.555 74.29 80.625 ;
        RECT 59.095 80.625 74.29 80.695 ;
        RECT 59.165 80.695 74.29 80.765 ;
        RECT 59.235 80.765 74.29 80.835 ;
        RECT 59.305 80.835 74.29 80.905 ;
        RECT 59.375 80.905 74.29 80.975 ;
        RECT 59.445 80.975 74.29 81.045 ;
        RECT 59.515 81.045 74.29 81.115 ;
        RECT 59.585 81.115 74.29 81.185 ;
        RECT 59.655 81.185 74.29 81.255 ;
        RECT 59.725 81.255 74.29 81.325 ;
        RECT 59.795 81.325 74.29 81.395 ;
        RECT 59.865 81.395 74.29 81.465 ;
        RECT 59.935 81.465 74.29 81.535 ;
        RECT 60.005 81.535 74.29 81.605 ;
        RECT 60.075 81.605 74.29 81.675 ;
        RECT 60.145 81.675 74.29 81.745 ;
        RECT 60.215 81.745 74.29 81.815 ;
        RECT 60.285 81.815 74.29 81.885 ;
        RECT 60.355 81.885 74.29 81.955 ;
        RECT 60.425 81.955 74.29 82.025 ;
        RECT 60.495 82.025 74.29 82.095 ;
        RECT 60.565 82.095 74.29 82.165 ;
        RECT 60.635 82.165 74.29 82.235 ;
        RECT 60.705 82.235 74.29 82.305 ;
        RECT 60.775 82.305 74.29 82.375 ;
        RECT 60.845 82.375 74.29 82.445 ;
        RECT 60.915 82.445 74.29 82.515 ;
        RECT 60.985 82.515 74.29 82.585 ;
        RECT 61.055 82.585 74.29 82.655 ;
        RECT 61.11 82.655 74.29 82.71 ;
        RECT 24.82 75.615 74.29 79.155 ;
        RECT 23.69 74.415 74.29 74.485 ;
        RECT 23.76 74.485 74.29 74.555 ;
        RECT 23.83 74.555 74.29 74.625 ;
        RECT 23.9 74.625 74.29 74.695 ;
        RECT 23.97 74.695 74.29 74.765 ;
        RECT 24.04 74.765 74.29 74.835 ;
        RECT 24.11 74.835 74.29 74.905 ;
        RECT 24.18 74.905 74.29 74.975 ;
        RECT 24.25 74.975 74.29 75.045 ;
        RECT 24.32 75.045 74.29 75.115 ;
        RECT 24.39 75.115 74.29 75.185 ;
        RECT 24.46 75.185 74.29 75.255 ;
        RECT 24.53 75.255 74.29 75.325 ;
        RECT 24.6 75.325 74.29 75.395 ;
        RECT 24.67 75.395 74.29 75.465 ;
        RECT 24.74 75.465 74.29 75.535 ;
        RECT 24.81 75.535 74.29 75.605 ;
        RECT 24.82 75.605 74.29 75.615 ;
        RECT 18.41 74.155 74.29 74.415 ;
        RECT 24.82 72.985 74.29 73.055 ;
        RECT 24.75 73.055 74.29 73.125 ;
        RECT 24.68 73.125 74.29 73.195 ;
        RECT 24.61 73.195 74.29 73.265 ;
        RECT 24.54 73.265 74.29 73.335 ;
        RECT 24.47 73.335 74.29 73.405 ;
        RECT 24.4 73.405 74.29 73.475 ;
        RECT 24.33 73.475 74.29 73.545 ;
        RECT 24.26 73.545 74.29 73.615 ;
        RECT 24.19 73.615 74.29 73.685 ;
        RECT 24.12 73.685 74.29 73.755 ;
        RECT 24.05 73.755 74.29 73.825 ;
        RECT 23.98 73.825 74.29 73.895 ;
        RECT 23.91 73.895 74.29 73.965 ;
        RECT 23.84 73.965 74.29 74.035 ;
        RECT 23.77 74.035 74.29 74.105 ;
        RECT 23.7 74.105 74.29 74.155 ;
        RECT 24.82 70.455 74.29 72.985 ;
        RECT 61.11 66.85 74.29 66.92 ;
        RECT 61.04 66.92 74.29 66.99 ;
        RECT 60.97 66.99 74.29 67.06 ;
        RECT 60.9 67.06 74.29 67.13 ;
        RECT 60.83 67.13 74.29 67.2 ;
        RECT 60.76 67.2 74.29 67.27 ;
        RECT 60.69 67.27 74.29 67.34 ;
        RECT 60.62 67.34 74.29 67.41 ;
        RECT 60.55 67.41 74.29 67.48 ;
        RECT 60.48 67.48 74.29 67.55 ;
        RECT 60.41 67.55 74.29 67.62 ;
        RECT 60.34 67.62 74.29 67.69 ;
        RECT 60.27 67.69 74.29 67.76 ;
        RECT 60.2 67.76 74.29 67.83 ;
        RECT 60.13 67.83 74.29 67.9 ;
        RECT 60.06 67.9 74.29 67.97 ;
        RECT 59.99 67.97 74.29 68.04 ;
        RECT 59.92 68.04 74.29 68.11 ;
        RECT 59.85 68.11 74.29 68.18 ;
        RECT 59.78 68.18 74.29 68.25 ;
        RECT 59.71 68.25 74.29 68.32 ;
        RECT 59.64 68.32 74.29 68.39 ;
        RECT 59.57 68.39 74.29 68.46 ;
        RECT 59.5 68.46 74.29 68.53 ;
        RECT 59.43 68.53 74.29 68.6 ;
        RECT 59.36 68.6 74.29 68.67 ;
        RECT 59.29 68.67 74.29 68.74 ;
        RECT 59.22 68.74 74.29 68.81 ;
        RECT 59.15 68.81 74.29 68.88 ;
        RECT 59.08 68.88 74.29 68.95 ;
        RECT 59.01 68.95 74.29 69.02 ;
        RECT 58.94 69.02 74.29 69.09 ;
        RECT 58.87 69.09 74.29 69.16 ;
        RECT 58.8 69.16 74.29 69.23 ;
        RECT 58.73 69.23 74.29 69.3 ;
        RECT 58.66 69.3 74.29 69.37 ;
        RECT 58.59 69.37 74.29 69.44 ;
        RECT 58.52 69.44 74.29 69.51 ;
        RECT 58.45 69.51 74.29 69.58 ;
        RECT 58.38 69.58 74.29 69.65 ;
        RECT 58.31 69.65 74.29 69.72 ;
        RECT 58.24 69.72 74.29 69.79 ;
        RECT 58.17 69.79 74.29 69.86 ;
        RECT 58.1 69.86 74.29 69.93 ;
        RECT 58.03 69.93 74.29 70 ;
        RECT 57.96 70 74.29 70.07 ;
        RECT 57.89 70.07 74.29 70.14 ;
        RECT 57.82 70.14 74.29 70.21 ;
        RECT 57.75 70.21 74.29 70.28 ;
        RECT 57.68 70.28 74.29 70.35 ;
        RECT 57.61 70.35 74.29 70.42 ;
        RECT 57.54 70.42 74.29 70.455 ;
        RECT 61.11 59.74 74.29 66.85 ;
        RECT 57.595 56.155 74.29 56.225 ;
        RECT 57.665 56.225 74.29 56.295 ;
        RECT 57.735 56.295 74.29 56.365 ;
        RECT 57.805 56.365 74.29 56.435 ;
        RECT 57.875 56.435 74.29 56.505 ;
        RECT 57.945 56.505 74.29 56.575 ;
        RECT 58.015 56.575 74.29 56.645 ;
        RECT 58.085 56.645 74.29 56.715 ;
        RECT 58.155 56.715 74.29 56.785 ;
        RECT 58.225 56.785 74.29 56.855 ;
        RECT 58.295 56.855 74.29 56.925 ;
        RECT 58.365 56.925 74.29 56.995 ;
        RECT 58.435 56.995 74.29 57.065 ;
        RECT 58.505 57.065 74.29 57.135 ;
        RECT 58.575 57.135 74.29 57.205 ;
        RECT 58.645 57.205 74.29 57.275 ;
        RECT 58.715 57.275 74.29 57.345 ;
        RECT 58.785 57.345 74.29 57.415 ;
        RECT 58.855 57.415 74.29 57.485 ;
        RECT 58.925 57.485 74.29 57.555 ;
        RECT 58.995 57.555 74.29 57.625 ;
        RECT 59.065 57.625 74.29 57.695 ;
        RECT 59.135 57.695 74.29 57.765 ;
        RECT 59.205 57.765 74.29 57.835 ;
        RECT 59.275 57.835 74.29 57.905 ;
        RECT 59.345 57.905 74.29 57.975 ;
        RECT 59.415 57.975 74.29 58.045 ;
        RECT 59.485 58.045 74.29 58.115 ;
        RECT 59.555 58.115 74.29 58.185 ;
        RECT 59.625 58.185 74.29 58.255 ;
        RECT 59.695 58.255 74.29 58.325 ;
        RECT 59.765 58.325 74.29 58.395 ;
        RECT 59.835 58.395 74.29 58.465 ;
        RECT 59.905 58.465 74.29 58.535 ;
        RECT 59.975 58.535 74.29 58.605 ;
        RECT 60.045 58.605 74.29 58.675 ;
        RECT 60.115 58.675 74.29 58.745 ;
        RECT 60.185 58.745 74.29 58.815 ;
        RECT 60.255 58.815 74.29 58.885 ;
        RECT 60.325 58.885 74.29 58.955 ;
        RECT 60.395 58.955 74.29 59.025 ;
        RECT 60.465 59.025 74.29 59.095 ;
        RECT 60.535 59.095 74.29 59.165 ;
        RECT 60.605 59.165 74.29 59.235 ;
        RECT 60.675 59.235 74.29 59.305 ;
        RECT 60.745 59.305 74.29 59.375 ;
        RECT 60.815 59.375 74.29 59.445 ;
        RECT 60.885 59.445 74.29 59.515 ;
        RECT 60.955 59.515 74.29 59.585 ;
        RECT 61.025 59.585 74.29 59.655 ;
        RECT 61.095 59.655 74.29 59.725 ;
        RECT 61.11 59.725 74.29 59.74 ;
        RECT 17.53 54.765 74.29 54.835 ;
        RECT 17.6 54.835 74.29 54.905 ;
        RECT 17.67 54.905 74.29 54.975 ;
        RECT 17.74 54.975 74.29 55.045 ;
        RECT 17.81 55.045 74.29 55.115 ;
        RECT 17.88 55.115 74.29 55.185 ;
        RECT 17.95 55.185 74.29 55.255 ;
        RECT 18.02 55.255 74.29 55.325 ;
        RECT 18.09 55.325 74.29 55.395 ;
        RECT 18.16 55.395 74.29 55.465 ;
        RECT 18.23 55.465 74.29 55.535 ;
        RECT 18.3 55.535 74.29 55.605 ;
        RECT 18.37 55.605 74.29 55.675 ;
        RECT 18.44 55.675 74.29 55.745 ;
        RECT 18.51 55.745 74.29 55.815 ;
        RECT 18.58 55.815 74.29 55.885 ;
        RECT 18.65 55.885 74.29 55.955 ;
        RECT 18.72 55.955 74.29 56.025 ;
        RECT 18.79 56.025 74.29 56.095 ;
        RECT 18.85 56.095 74.29 56.155 ;
        RECT 16.805 47.455 74.29 54.765 ;
        RECT 61.11 43.82 74.29 43.89 ;
        RECT 61.04 43.89 74.29 43.96 ;
        RECT 60.97 43.96 74.29 44.03 ;
        RECT 60.9 44.03 74.29 44.1 ;
        RECT 60.83 44.1 74.29 44.17 ;
        RECT 60.76 44.17 74.29 44.24 ;
        RECT 60.69 44.24 74.29 44.31 ;
        RECT 60.62 44.31 74.29 44.38 ;
        RECT 60.55 44.38 74.29 44.45 ;
        RECT 60.48 44.45 74.29 44.52 ;
        RECT 60.41 44.52 74.29 44.59 ;
        RECT 60.34 44.59 74.29 44.66 ;
        RECT 60.27 44.66 74.29 44.73 ;
        RECT 60.2 44.73 74.29 44.8 ;
        RECT 60.13 44.8 74.29 44.87 ;
        RECT 60.06 44.87 74.29 44.94 ;
        RECT 59.99 44.94 74.29 45.01 ;
        RECT 59.92 45.01 74.29 45.08 ;
        RECT 59.85 45.08 74.29 45.15 ;
        RECT 59.78 45.15 74.29 45.22 ;
        RECT 59.71 45.22 74.29 45.29 ;
        RECT 59.64 45.29 74.29 45.36 ;
        RECT 59.57 45.36 74.29 45.43 ;
        RECT 59.5 45.43 74.29 45.5 ;
        RECT 59.43 45.5 74.29 45.57 ;
        RECT 59.36 45.57 74.29 45.64 ;
        RECT 59.29 45.64 74.29 45.71 ;
        RECT 59.22 45.71 74.29 45.78 ;
        RECT 59.15 45.78 74.29 45.85 ;
        RECT 59.08 45.85 74.29 45.92 ;
        RECT 59.01 45.92 74.29 45.99 ;
        RECT 58.94 45.99 74.29 46.06 ;
        RECT 58.87 46.06 74.29 46.13 ;
        RECT 58.8 46.13 74.29 46.2 ;
        RECT 58.73 46.2 74.29 46.27 ;
        RECT 58.66 46.27 74.29 46.34 ;
        RECT 58.59 46.34 74.29 46.41 ;
        RECT 58.52 46.41 74.29 46.48 ;
        RECT 58.45 46.48 74.29 46.55 ;
        RECT 58.38 46.55 74.29 46.62 ;
        RECT 58.31 46.62 74.29 46.69 ;
        RECT 58.24 46.69 74.29 46.76 ;
        RECT 58.17 46.76 74.29 46.83 ;
        RECT 58.1 46.83 74.29 46.9 ;
        RECT 58.03 46.9 74.29 46.97 ;
        RECT 57.96 46.97 74.29 47.04 ;
        RECT 57.89 47.04 74.29 47.11 ;
        RECT 57.82 47.11 74.29 47.18 ;
        RECT 57.75 47.18 74.29 47.25 ;
        RECT 57.68 47.25 74.29 47.32 ;
        RECT 57.61 47.32 74.29 47.39 ;
        RECT 57.54 47.39 74.29 47.455 ;
        RECT 61.11 30.955 74.29 43.82 ;
        RECT 61.11 30.91 74.29 30.955 ;
        RECT 61.065 30.84 74.29 30.91 ;
        RECT 60.995 30.77 74.29 30.84 ;
        RECT 60.925 30.7 74.29 30.77 ;
        RECT 60.855 30.63 74.29 30.7 ;
        RECT 60.785 30.56 74.29 30.63 ;
        RECT 60.715 30.49 74.29 30.56 ;
        RECT 60.645 30.42 74.29 30.49 ;
        RECT 60.575 30.35 74.29 30.42 ;
        RECT 60.505 30.28 74.29 30.35 ;
        RECT 60.435 30.21 74.29 30.28 ;
        RECT 60.365 30.14 74.29 30.21 ;
        RECT 60.295 30.07 74.29 30.14 ;
        RECT 60.225 30 74.29 30.07 ;
        RECT 60.155 29.93 74.29 30 ;
        RECT 60.085 29.86 74.29 29.93 ;
        RECT 60.015 29.79 74.29 29.86 ;
        RECT 59.945 29.72 74.29 29.79 ;
        RECT 59.875 29.65 74.29 29.72 ;
        RECT 59.805 29.58 74.29 29.65 ;
        RECT 59.735 29.51 74.29 29.58 ;
        RECT 59.665 29.44 74.29 29.51 ;
        RECT 59.595 29.37 74.29 29.44 ;
        RECT 59.525 29.3 74.29 29.37 ;
        RECT 59.455 29.23 74.29 29.3 ;
        RECT 59.385 29.16 74.29 29.23 ;
        RECT 59.315 29.09 74.29 29.16 ;
        RECT 59.245 29.02 74.29 29.09 ;
        RECT 59.175 28.95 74.29 29.02 ;
        RECT 59.105 28.88 74.29 28.95 ;
        RECT 59.035 28.81 74.29 28.88 ;
        RECT 58.965 28.74 74.29 28.81 ;
        RECT 58.895 28.67 74.29 28.74 ;
        RECT 58.825 28.6 74.29 28.67 ;
        RECT 58.755 28.53 74.29 28.6 ;
        RECT 58.685 28.46 74.29 28.53 ;
        RECT 58.615 28.39 74.29 28.46 ;
        RECT 58.545 28.32 74.29 28.39 ;
        RECT 58.475 28.25 74.29 28.32 ;
        RECT 58.405 28.18 74.29 28.25 ;
        RECT 58.335 28.11 74.29 28.18 ;
        RECT 58.265 28.04 74.29 28.11 ;
        RECT 58.195 27.97 74.29 28.04 ;
        RECT 58.125 27.9 74.29 27.97 ;
        RECT 58.055 27.83 74.29 27.9 ;
        RECT 57.985 27.76 74.29 27.83 ;
        RECT 57.915 27.69 74.29 27.76 ;
        RECT 57.845 27.62 74.29 27.69 ;
        RECT 57.775 27.55 74.29 27.62 ;
        RECT 57.705 27.48 74.29 27.55 ;
        RECT 57.635 27.41 74.29 27.48 ;
        RECT 57.565 27.34 74.29 27.41 ;
        RECT 57.495 27.27 74.29 27.34 ;
        RECT 57.425 27.2 74.29 27.27 ;
        RECT 57.355 27.13 74.29 27.2 ;
        RECT 57.285 27.06 74.29 27.13 ;
        RECT 57.215 26.99 74.29 27.06 ;
        RECT 57.145 26.92 74.29 26.99 ;
        RECT 57.075 26.85 74.29 26.92 ;
        RECT 57.005 26.78 74.29 26.85 ;
        RECT 56.935 26.71 74.29 26.78 ;
        RECT 56.865 26.64 74.29 26.71 ;
        RECT 56.795 26.57 74.29 26.64 ;
        RECT 56.725 26.5 74.29 26.57 ;
        RECT 56.655 26.43 74.29 26.5 ;
        RECT 56.585 26.36 74.29 26.43 ;
        RECT 56.515 26.29 74.29 26.36 ;
        RECT 56.445 26.22 74.29 26.29 ;
        RECT 56.375 26.15 74.29 26.22 ;
        RECT 56.305 26.08 74.29 26.15 ;
        RECT 56.235 26.01 74.29 26.08 ;
        RECT 56.165 25.94 74.29 26.01 ;
        RECT 56.095 25.87 74.29 25.94 ;
        RECT 56.025 25.8 74.29 25.87 ;
        RECT 55.955 25.73 74.29 25.8 ;
        RECT 55.885 25.66 74.29 25.73 ;
        RECT 37.89 12.295 74.29 25.66 ;
        RECT 50.39 8.625 74.29 8.695 ;
        RECT 50.32 8.695 74.29 8.765 ;
        RECT 50.25 8.765 74.29 8.835 ;
        RECT 50.18 8.835 74.29 8.905 ;
        RECT 50.11 8.905 74.29 8.975 ;
        RECT 50.04 8.975 74.29 9.045 ;
        RECT 49.97 9.045 74.29 9.115 ;
        RECT 49.9 9.115 74.29 9.185 ;
        RECT 49.83 9.185 74.29 9.255 ;
        RECT 49.76 9.255 74.29 9.325 ;
        RECT 49.69 9.325 74.29 9.395 ;
        RECT 49.62 9.395 74.29 9.465 ;
        RECT 49.55 9.465 74.29 9.535 ;
        RECT 49.48 9.535 74.29 9.605 ;
        RECT 49.41 9.605 74.29 9.675 ;
        RECT 49.34 9.675 74.29 9.745 ;
        RECT 49.27 9.745 74.29 9.815 ;
        RECT 49.2 9.815 74.29 9.885 ;
        RECT 49.13 9.885 74.29 9.955 ;
        RECT 49.06 9.955 74.29 10.025 ;
        RECT 48.99 10.025 74.29 10.095 ;
        RECT 48.92 10.095 74.29 10.165 ;
        RECT 48.85 10.165 74.29 10.235 ;
        RECT 48.78 10.235 74.29 10.305 ;
        RECT 48.71 10.305 74.29 10.375 ;
        RECT 48.64 10.375 74.29 10.445 ;
        RECT 48.57 10.445 74.29 10.515 ;
        RECT 48.5 10.515 74.29 10.585 ;
        RECT 48.43 10.585 74.29 10.655 ;
        RECT 48.36 10.655 74.29 10.725 ;
        RECT 48.29 10.725 74.29 10.795 ;
        RECT 48.22 10.795 74.29 10.865 ;
        RECT 48.15 10.865 74.29 10.935 ;
        RECT 48.08 10.935 74.29 11.005 ;
        RECT 48.01 11.005 74.29 11.075 ;
        RECT 47.94 11.075 74.29 11.145 ;
        RECT 47.87 11.145 74.29 11.215 ;
        RECT 47.8 11.215 74.29 11.285 ;
        RECT 47.73 11.285 74.29 11.355 ;
        RECT 47.66 11.355 74.29 11.425 ;
        RECT 47.59 11.425 74.29 11.495 ;
        RECT 47.52 11.495 74.29 11.565 ;
        RECT 47.45 11.565 74.29 11.635 ;
        RECT 47.38 11.635 74.29 11.705 ;
        RECT 47.31 11.705 74.29 11.775 ;
        RECT 47.24 11.775 74.29 11.845 ;
        RECT 47.17 11.845 74.29 11.915 ;
        RECT 47.1 11.915 74.29 11.985 ;
        RECT 47.03 11.985 74.29 12.055 ;
        RECT 46.96 12.055 74.29 12.125 ;
        RECT 46.89 12.125 74.29 12.195 ;
        RECT 46.82 12.195 74.29 12.265 ;
        RECT 46.75 12.265 74.29 12.295 ;
        RECT 50.39 0 74.29 8.625 ;
    END
  END drn_hvc
  OBS
    LAYER met2 ;
      RECT 14.4 74.015 18.27 74.555 ;
      RECT 14.4 72.925 23.59 74.015 ;
      RECT 14.4 70.315 24.68 72.925 ;
      RECT 14.4 70.14 57.445 70.315 ;
      RECT 17.75 66.79 57.62 70.14 ;
      RECT 17.78 66.76 60.97 66.79 ;
      RECT 56.99 59.8 60.97 66.76 ;
      RECT 56.99 57.5 60.97 59.8 ;
      RECT 16.595 56.295 58.67 57.5 ;
      RECT 15.205 54.905 18.79 56.295 ;
      RECT 14.4 54.1 16.665 54.905 ;
      RECT 14.4 47.315 16.665 54.1 ;
      RECT 14.4 45.43 57.415 47.315 ;
      RECT 16.07 43.76 59.3 45.43 ;
      RECT 17.17 42.66 60.97 43.76 ;
      RECT 22.85 42.52 60.97 42.66 ;
      RECT 20.4 40.07 52.515 40.21 ;
      RECT 57.055 39.725 60.97 42.52 ;
      RECT 18.13 38.195 52.655 40.07 ;
      RECT 57.055 35.975 60.97 39.725 ;
      RECT 15.91 35.975 54.53 38.195 ;
      RECT 15.485 35.55 60.97 35.975 ;
      RECT 15.485 31.015 60.97 35.55 ;
      RECT 15.485 29.43 60.97 31.015 ;
      RECT 18.935 25.98 59.39 29.43 ;
      RECT 37.175 25.8 55.935 25.98 ;
      RECT 37.175 12.155 37.75 25.8 ;
      RECT 37.175 12.12 46.66 12.155 ;
      RECT 24.765 8.565 46.695 12.12 ;
      RECT 24.675 8.48 50.25 8.565 ;
      RECT 0 2.61 0.655 195.355 ;
      RECT 74.43 0 75 190.155 ;
      RECT 24.675 2.06 50.25 8.48 ;
      RECT 0 2.17 0.655 2.61 ;
      RECT 0 0 0.215 2.17 ;
      RECT 28.035 0 50.25 2.06 ;
      RECT 24.675 0 25.755 2.06 ;
      RECT 0 195.355 75 200 ;
      RECT 67.48 190.28 75 195.355 ;
      RECT 15.085 190.155 75 190.28 ;
      RECT 14.4 189.47 15.48 190.155 ;
      RECT 14.4 185.17 15.48 189.47 ;
      RECT 14.415 185.155 15.48 185.17 ;
      RECT 15.385 184.185 58.635 185.155 ;
      RECT 15.6 183.97 59.605 184.185 ;
      RECT 16.75 182.82 59.82 183.97 ;
      RECT 17.81 181.76 60.97 182.82 ;
      RECT 58.24 174.76 60.97 181.76 ;
      RECT 58.24 172.5 60.97 174.76 ;
      RECT 16.59 171.295 58.71 172.5 ;
      RECT 14.4 169.105 16.665 171.295 ;
      RECT 14.4 162.315 16.665 169.105 ;
      RECT 14.4 162.195 57.465 162.315 ;
      RECT 17.785 158.81 57.585 162.195 ;
      RECT 17.835 158.76 60.97 158.81 ;
      RECT 56.985 151.84 60.97 158.76 ;
      RECT 56.985 149.5 60.97 151.84 ;
      RECT 16.595 148.295 58.63 149.5 ;
      RECT 15.07 146.77 18.19 148.295 ;
      RECT 14.4 146.1 16.665 146.77 ;
      RECT 14.4 139.315 16.665 146.1 ;
      RECT 14.4 139.285 57.45 139.315 ;
      RECT 17.89 135.795 57.48 139.285 ;
      RECT 17.925 135.76 60.97 135.795 ;
      RECT 56.985 128.77 60.97 135.76 ;
      RECT 56.985 126.5 60.97 128.77 ;
      RECT 16.665 125.295 58.7 126.5 ;
      RECT 14.4 123.03 24.68 125.295 ;
      RECT 14.4 116.315 24.68 123.03 ;
      RECT 14.4 116.18 57.415 116.315 ;
      RECT 17.82 112.76 57.55 116.18 ;
      RECT 17.82 112.76 60.97 112.76 ;
      RECT 56.985 105.77 60.97 112.76 ;
      RECT 56.985 103.5 60.97 105.77 ;
      RECT 16.57 102.295 58.7 103.5 ;
      RECT 14.4 100.125 24.68 102.295 ;
      RECT 14.4 93.315 24.68 100.125 ;
      RECT 14.4 93.14 57.505 93.315 ;
      RECT 17.69 89.85 57.68 93.14 ;
      RECT 17.78 89.76 60.97 89.85 ;
      RECT 56.985 82.77 60.97 89.76 ;
      RECT 56.985 80.5 60.97 82.77 ;
      RECT 16.57 79.295 58.7 80.5 ;
      RECT 14.4 77.125 24.68 79.295 ;
      RECT 14.4 75.675 24.68 77.125 ;
      RECT 14.4 74.555 24.68 75.675 ;
      RECT 54.465 42.51 60.83 42.58 ;
      RECT 54.395 42.58 60.83 42.65 ;
      RECT 54.325 42.65 60.83 42.66 ;
      RECT 15.555 35.55 60.83 35.62 ;
      RECT 15.625 35.62 60.83 35.69 ;
      RECT 15.695 35.69 60.83 35.76 ;
      RECT 15.765 35.76 60.83 35.83 ;
      RECT 15.77 35.83 60.83 35.835 ;
      RECT 15.485 29.43 59.19 29.5 ;
      RECT 15.485 29.5 59.26 29.57 ;
      RECT 15.485 29.57 59.33 29.64 ;
      RECT 15.485 29.64 59.4 29.71 ;
      RECT 15.485 29.71 59.47 29.78 ;
      RECT 15.485 29.78 59.54 29.85 ;
      RECT 15.485 29.85 59.61 29.92 ;
      RECT 15.485 29.92 59.68 29.99 ;
      RECT 15.485 29.99 59.75 30.06 ;
      RECT 15.485 30.06 59.82 30.13 ;
      RECT 15.485 30.13 59.89 30.2 ;
      RECT 15.485 30.2 59.96 30.27 ;
      RECT 15.485 30.27 60.03 30.34 ;
      RECT 15.485 30.34 60.1 30.41 ;
      RECT 15.485 30.41 60.17 30.48 ;
      RECT 15.485 30.48 60.24 30.55 ;
      RECT 15.485 30.55 60.31 30.62 ;
      RECT 15.485 30.62 60.38 30.69 ;
      RECT 15.485 30.69 60.45 30.76 ;
      RECT 15.485 30.76 60.52 30.83 ;
      RECT 15.485 30.83 60.59 30.9 ;
      RECT 15.485 30.9 60.66 30.97 ;
      RECT 15.485 30.97 60.73 31.04 ;
      RECT 15.485 31.04 60.8 31.07 ;
      RECT 17.78 89.76 60.83 89.775 ;
      RECT 17.765 89.775 60.83 89.79 ;
      RECT 17.75 89.79 60.83 89.795 ;
      RECT 56.985 82.81 60.815 82.825 ;
      RECT 56.985 82.74 60.745 82.81 ;
      RECT 56.985 82.67 60.675 82.74 ;
      RECT 56.985 82.6 60.605 82.67 ;
      RECT 56.985 82.53 60.535 82.6 ;
      RECT 56.985 82.46 60.465 82.53 ;
      RECT 56.985 82.39 60.395 82.46 ;
      RECT 56.985 82.32 60.325 82.39 ;
      RECT 56.985 82.25 60.255 82.32 ;
      RECT 56.985 82.18 60.185 82.25 ;
      RECT 56.985 82.11 60.115 82.18 ;
      RECT 56.985 82.04 60.045 82.11 ;
      RECT 56.985 81.97 59.975 82.04 ;
      RECT 56.985 81.9 59.905 81.97 ;
      RECT 56.985 81.83 59.835 81.9 ;
      RECT 56.985 81.76 59.765 81.83 ;
      RECT 56.985 81.69 59.695 81.76 ;
      RECT 56.985 81.62 59.625 81.69 ;
      RECT 56.985 81.55 59.555 81.62 ;
      RECT 56.985 81.48 59.485 81.55 ;
      RECT 56.985 81.41 59.415 81.48 ;
      RECT 56.985 81.34 59.345 81.41 ;
      RECT 56.985 81.27 59.275 81.34 ;
      RECT 56.985 81.2 59.205 81.27 ;
      RECT 56.985 81.13 59.135 81.2 ;
      RECT 56.985 81.06 59.065 81.13 ;
      RECT 56.985 80.99 58.995 81.06 ;
      RECT 56.985 80.92 58.925 80.99 ;
      RECT 56.985 80.85 58.855 80.92 ;
      RECT 56.985 80.78 58.785 80.85 ;
      RECT 56.985 80.71 58.715 80.78 ;
      RECT 56.985 80.64 58.645 80.71 ;
      RECT 56.985 80.57 58.575 80.64 ;
      RECT 56.985 80.5 58.505 80.57 ;
      RECT 24.69 8.48 50.11 8.495 ;
      RECT 24.705 8.495 50.11 8.51 ;
      RECT 15.52 78.175 24.54 78.245 ;
      RECT 15.59 78.245 24.54 78.315 ;
      RECT 15.66 78.315 24.54 78.385 ;
      RECT 15.73 78.385 24.54 78.455 ;
      RECT 15.8 78.455 24.54 78.525 ;
      RECT 15.87 78.525 24.54 78.595 ;
      RECT 15.94 78.595 24.54 78.665 ;
      RECT 16.01 78.665 24.54 78.735 ;
      RECT 16.08 78.735 24.54 78.805 ;
      RECT 16.15 78.805 24.54 78.875 ;
      RECT 16.22 78.875 24.54 78.945 ;
      RECT 16.29 78.945 24.54 79.015 ;
      RECT 16.36 79.015 24.54 79.085 ;
      RECT 16.43 79.085 24.54 79.155 ;
      RECT 16.5 79.155 24.54 79.225 ;
      RECT 16.57 79.225 24.54 79.295 ;
      RECT 16.64 79.295 24.54 79.365 ;
      RECT 16.71 79.365 24.54 79.435 ;
      RECT 14.4 74.695 23.505 74.765 ;
      RECT 14.4 74.765 23.575 74.835 ;
      RECT 14.4 74.835 23.645 74.905 ;
      RECT 14.4 74.905 23.715 74.975 ;
      RECT 14.4 74.975 23.785 75.045 ;
      RECT 14.4 75.045 23.855 75.115 ;
      RECT 14.4 75.115 23.925 75.185 ;
      RECT 14.4 75.185 23.995 75.255 ;
      RECT 14.4 75.255 24.065 75.325 ;
      RECT 14.4 75.325 24.135 75.395 ;
      RECT 14.4 75.395 24.205 75.465 ;
      RECT 14.4 75.465 24.275 75.535 ;
      RECT 14.4 75.535 24.345 75.605 ;
      RECT 14.4 75.605 24.415 75.675 ;
      RECT 14.4 75.675 24.485 75.73 ;
      RECT 14.4 72.87 24.47 72.94 ;
      RECT 14.4 72.94 24.4 73.01 ;
      RECT 14.4 73.01 24.33 73.08 ;
      RECT 14.4 73.08 24.26 73.15 ;
      RECT 14.4 73.15 24.19 73.22 ;
      RECT 14.4 73.22 24.12 73.29 ;
      RECT 14.4 73.29 24.05 73.36 ;
      RECT 14.4 73.36 23.98 73.43 ;
      RECT 14.4 73.43 23.91 73.5 ;
      RECT 14.4 73.5 23.84 73.57 ;
      RECT 14.4 73.57 23.77 73.64 ;
      RECT 14.4 73.64 23.7 73.71 ;
      RECT 14.4 73.71 23.63 73.78 ;
      RECT 14.4 73.78 23.56 73.85 ;
      RECT 14.4 73.85 23.535 73.875 ;
      RECT 14.4 70.14 57.405 70.16 ;
      RECT 14.4 70.16 57.39 70.175 ;
      RECT 56.99 66.735 60.82 66.745 ;
      RECT 56.99 66.745 60.805 66.76 ;
      RECT 56.99 59.81 60.785 59.855 ;
      RECT 56.99 59.74 60.715 59.81 ;
      RECT 56.99 59.67 60.645 59.74 ;
      RECT 56.99 59.6 60.575 59.67 ;
      RECT 56.99 59.53 60.505 59.6 ;
      RECT 56.99 59.46 60.435 59.53 ;
      RECT 56.99 59.39 60.365 59.46 ;
      RECT 56.99 59.32 60.295 59.39 ;
      RECT 56.99 59.25 60.225 59.32 ;
      RECT 56.99 59.18 60.155 59.25 ;
      RECT 56.99 59.11 60.085 59.18 ;
      RECT 56.99 59.04 60.015 59.11 ;
      RECT 56.99 58.97 59.945 59.04 ;
      RECT 56.99 58.9 59.875 58.97 ;
      RECT 56.99 58.83 59.805 58.9 ;
      RECT 56.99 58.76 59.735 58.83 ;
      RECT 56.99 58.69 59.665 58.76 ;
      RECT 56.99 58.62 59.595 58.69 ;
      RECT 56.99 58.55 59.525 58.62 ;
      RECT 56.99 58.48 59.455 58.55 ;
      RECT 56.99 58.41 59.385 58.48 ;
      RECT 56.99 58.34 59.315 58.41 ;
      RECT 56.99 58.27 59.245 58.34 ;
      RECT 56.99 58.2 59.175 58.27 ;
      RECT 56.99 58.13 59.105 58.2 ;
      RECT 56.99 58.06 59.035 58.13 ;
      RECT 56.99 57.99 58.965 58.06 ;
      RECT 56.99 57.92 58.895 57.99 ;
      RECT 56.99 57.85 58.825 57.92 ;
      RECT 56.99 57.78 58.755 57.85 ;
      RECT 56.99 57.71 58.685 57.78 ;
      RECT 56.99 57.64 58.615 57.71 ;
      RECT 56.99 57.57 58.545 57.64 ;
      RECT 56.99 57.5 58.475 57.57 ;
      RECT 57.195 39.78 60.83 39.85 ;
      RECT 57.125 39.85 60.83 39.92 ;
      RECT 57.055 39.92 60.83 39.99 ;
      RECT 56.985 39.99 60.83 40.06 ;
      RECT 56.915 40.06 60.83 40.13 ;
      RECT 56.845 40.13 60.83 40.2 ;
      RECT 56.775 40.2 60.83 40.27 ;
      RECT 56.705 40.27 60.83 40.34 ;
      RECT 56.635 40.34 60.83 40.41 ;
      RECT 56.565 40.41 60.83 40.48 ;
      RECT 56.495 40.48 60.83 40.55 ;
      RECT 56.425 40.55 60.83 40.62 ;
      RECT 56.355 40.62 60.83 40.69 ;
      RECT 56.285 40.69 60.83 40.76 ;
      RECT 56.215 40.76 60.83 40.83 ;
      RECT 56.145 40.83 60.83 40.9 ;
      RECT 56.075 40.9 60.83 40.97 ;
      RECT 56.005 40.97 60.83 41.04 ;
      RECT 55.935 41.04 60.83 41.11 ;
      RECT 55.865 41.11 60.83 41.18 ;
      RECT 55.795 41.18 60.83 41.25 ;
      RECT 55.725 41.25 60.83 41.32 ;
      RECT 55.655 41.32 60.83 41.39 ;
      RECT 55.585 41.39 60.83 41.46 ;
      RECT 55.515 41.46 60.83 41.53 ;
      RECT 55.445 41.53 60.83 41.6 ;
      RECT 55.375 41.6 60.83 41.67 ;
      RECT 55.305 41.67 60.83 41.74 ;
      RECT 55.235 41.74 60.83 41.81 ;
      RECT 55.165 41.81 60.83 41.88 ;
      RECT 55.095 41.88 60.83 41.95 ;
      RECT 55.025 41.95 60.83 42.02 ;
      RECT 54.955 42.02 60.83 42.09 ;
      RECT 54.885 42.09 60.83 42.16 ;
      RECT 54.815 42.16 60.83 42.23 ;
      RECT 54.745 42.23 60.83 42.3 ;
      RECT 54.675 42.3 60.83 42.37 ;
      RECT 54.605 42.37 60.83 42.44 ;
      RECT 54.535 42.44 60.83 42.51 ;
      RECT 56.985 126.64 58.645 126.71 ;
      RECT 56.985 126.57 58.575 126.64 ;
      RECT 56.985 126.5 58.505 126.57 ;
      RECT 14.47 123.03 24.54 123.1 ;
      RECT 14.54 123.1 24.54 123.17 ;
      RECT 14.61 123.17 24.54 123.24 ;
      RECT 14.68 123.24 24.54 123.31 ;
      RECT 14.75 123.31 24.54 123.38 ;
      RECT 14.82 123.38 24.54 123.45 ;
      RECT 14.89 123.45 24.54 123.52 ;
      RECT 14.96 123.52 24.54 123.59 ;
      RECT 15.03 123.59 24.54 123.66 ;
      RECT 15.1 123.66 24.54 123.73 ;
      RECT 15.17 123.73 24.54 123.8 ;
      RECT 15.24 123.8 24.54 123.87 ;
      RECT 15.31 123.87 24.54 123.94 ;
      RECT 15.38 123.94 24.54 124.01 ;
      RECT 15.45 124.01 24.54 124.08 ;
      RECT 15.52 124.08 24.54 124.15 ;
      RECT 15.59 124.15 24.54 124.22 ;
      RECT 15.66 124.22 24.54 124.29 ;
      RECT 15.73 124.29 24.54 124.36 ;
      RECT 15.8 124.36 24.54 124.43 ;
      RECT 15.87 124.43 24.54 124.5 ;
      RECT 15.94 124.5 24.54 124.57 ;
      RECT 16.01 124.57 24.54 124.64 ;
      RECT 16.08 124.64 24.54 124.71 ;
      RECT 16.15 124.71 24.54 124.78 ;
      RECT 16.22 124.78 24.54 124.85 ;
      RECT 16.29 124.85 24.54 124.92 ;
      RECT 16.36 124.92 24.54 124.99 ;
      RECT 16.43 124.99 24.54 125.06 ;
      RECT 16.5 125.06 24.54 125.13 ;
      RECT 16.57 125.13 24.54 125.2 ;
      RECT 16.64 125.2 24.54 125.27 ;
      RECT 16.71 125.27 24.54 125.34 ;
      RECT 16.78 125.34 24.54 125.41 ;
      RECT 16.805 125.41 24.54 125.435 ;
      RECT 14.405 116.175 24.54 116.18 ;
      RECT 56.985 112.705 60.805 112.73 ;
      RECT 56.985 112.73 60.775 112.76 ;
      RECT 56.985 105.81 60.815 105.825 ;
      RECT 56.985 105.74 60.745 105.81 ;
      RECT 56.985 105.67 60.675 105.74 ;
      RECT 56.985 105.6 60.605 105.67 ;
      RECT 56.985 105.53 60.535 105.6 ;
      RECT 56.985 105.46 60.465 105.53 ;
      RECT 56.985 105.39 60.395 105.46 ;
      RECT 56.985 105.32 60.325 105.39 ;
      RECT 56.985 105.25 60.255 105.32 ;
      RECT 56.985 105.18 60.185 105.25 ;
      RECT 56.985 105.11 60.115 105.18 ;
      RECT 56.985 105.04 60.045 105.11 ;
      RECT 56.985 104.97 59.975 105.04 ;
      RECT 56.985 104.9 59.905 104.97 ;
      RECT 56.985 104.83 59.835 104.9 ;
      RECT 56.985 104.76 59.765 104.83 ;
      RECT 56.985 104.69 59.695 104.76 ;
      RECT 56.985 104.62 59.625 104.69 ;
      RECT 56.985 104.55 59.555 104.62 ;
      RECT 56.985 104.48 59.485 104.55 ;
      RECT 56.985 104.41 59.415 104.48 ;
      RECT 56.985 104.34 59.345 104.41 ;
      RECT 56.985 104.27 59.275 104.34 ;
      RECT 56.985 104.2 59.205 104.27 ;
      RECT 56.985 104.13 59.135 104.2 ;
      RECT 56.985 104.06 59.065 104.13 ;
      RECT 56.985 103.99 58.995 104.06 ;
      RECT 56.985 103.92 58.925 103.99 ;
      RECT 56.985 103.85 58.855 103.92 ;
      RECT 56.985 103.78 58.785 103.85 ;
      RECT 56.985 103.71 58.715 103.78 ;
      RECT 56.985 103.64 58.645 103.71 ;
      RECT 56.985 103.57 58.575 103.64 ;
      RECT 56.985 103.5 58.505 103.57 ;
      RECT 14.47 100.125 24.54 100.195 ;
      RECT 14.54 100.195 24.54 100.265 ;
      RECT 14.61 100.265 24.54 100.335 ;
      RECT 14.68 100.335 24.54 100.405 ;
      RECT 14.75 100.405 24.54 100.475 ;
      RECT 14.82 100.475 24.54 100.545 ;
      RECT 14.89 100.545 24.54 100.615 ;
      RECT 14.96 100.615 24.54 100.685 ;
      RECT 15.03 100.685 24.54 100.755 ;
      RECT 15.1 100.755 24.54 100.825 ;
      RECT 15.17 100.825 24.54 100.895 ;
      RECT 15.24 100.895 24.54 100.965 ;
      RECT 15.31 100.965 24.54 101.035 ;
      RECT 15.38 101.035 24.54 101.105 ;
      RECT 15.45 101.105 24.54 101.175 ;
      RECT 15.52 101.175 24.54 101.245 ;
      RECT 15.59 101.245 24.54 101.315 ;
      RECT 15.66 101.315 24.54 101.385 ;
      RECT 15.73 101.385 24.54 101.455 ;
      RECT 15.8 101.455 24.54 101.525 ;
      RECT 15.87 101.525 24.54 101.595 ;
      RECT 15.94 101.595 24.54 101.665 ;
      RECT 16.01 101.665 24.54 101.735 ;
      RECT 16.08 101.735 24.54 101.805 ;
      RECT 16.15 101.805 24.54 101.875 ;
      RECT 16.22 101.875 24.54 101.945 ;
      RECT 16.29 101.945 24.54 102.015 ;
      RECT 16.36 102.015 24.54 102.085 ;
      RECT 16.43 102.085 24.54 102.155 ;
      RECT 16.5 102.155 24.54 102.225 ;
      RECT 16.57 102.225 24.54 102.295 ;
      RECT 16.64 102.295 24.54 102.365 ;
      RECT 16.71 102.365 24.54 102.435 ;
      RECT 14.4 93.14 57.465 93.16 ;
      RECT 14.4 93.16 57.45 93.175 ;
      RECT 14.47 77.125 24.54 77.195 ;
      RECT 14.54 77.195 24.54 77.265 ;
      RECT 14.61 77.265 24.54 77.335 ;
      RECT 14.68 77.335 24.54 77.405 ;
      RECT 14.75 77.405 24.54 77.475 ;
      RECT 14.82 77.475 24.54 77.545 ;
      RECT 14.89 77.545 24.54 77.615 ;
      RECT 14.96 77.615 24.54 77.685 ;
      RECT 15.03 77.685 24.54 77.755 ;
      RECT 15.1 77.755 24.54 77.825 ;
      RECT 15.17 77.825 24.54 77.895 ;
      RECT 15.24 77.895 24.54 77.965 ;
      RECT 15.31 77.965 24.54 78.035 ;
      RECT 15.38 78.035 24.54 78.105 ;
      RECT 15.45 78.105 24.54 78.175 ;
      RECT 26.525 10.26 48.29 10.33 ;
      RECT 26.595 10.33 48.22 10.4 ;
      RECT 26.665 10.4 48.15 10.47 ;
      RECT 26.735 10.47 48.08 10.54 ;
      RECT 26.805 10.54 48.01 10.61 ;
      RECT 26.875 10.61 47.94 10.68 ;
      RECT 26.945 10.68 47.87 10.75 ;
      RECT 27.015 10.75 47.8 10.82 ;
      RECT 27.085 10.82 47.73 10.89 ;
      RECT 27.155 10.89 47.66 10.96 ;
      RECT 27.225 10.96 47.59 11.03 ;
      RECT 27.295 11.03 47.52 11.1 ;
      RECT 27.365 11.1 47.45 11.17 ;
      RECT 27.435 11.17 47.38 11.24 ;
      RECT 27.505 11.24 47.31 11.31 ;
      RECT 27.575 11.31 47.24 11.38 ;
      RECT 27.645 11.38 47.17 11.45 ;
      RECT 27.715 11.45 47.1 11.52 ;
      RECT 27.785 11.52 47.03 11.59 ;
      RECT 27.855 11.59 46.96 11.66 ;
      RECT 27.925 11.66 46.89 11.73 ;
      RECT 27.995 11.73 46.82 11.8 ;
      RECT 28.065 11.8 46.75 11.87 ;
      RECT 28.135 11.87 46.68 11.94 ;
      RECT 28.205 11.94 46.61 12.01 ;
      RECT 28.21 12.01 46.605 12.015 ;
      RECT 14.4 45.43 59.035 45.5 ;
      RECT 14.4 45.5 58.965 45.57 ;
      RECT 14.4 45.57 58.895 45.64 ;
      RECT 14.4 45.64 58.825 45.71 ;
      RECT 14.4 45.71 58.755 45.78 ;
      RECT 14.4 45.78 58.685 45.85 ;
      RECT 14.4 45.85 58.615 45.92 ;
      RECT 14.4 45.92 58.545 45.99 ;
      RECT 14.4 45.99 58.475 46.06 ;
      RECT 14.4 46.06 58.405 46.13 ;
      RECT 14.4 46.13 58.335 46.2 ;
      RECT 14.4 46.2 58.265 46.27 ;
      RECT 14.4 46.27 58.195 46.34 ;
      RECT 14.4 46.34 58.125 46.41 ;
      RECT 14.4 46.41 58.055 46.48 ;
      RECT 14.4 46.48 57.985 46.55 ;
      RECT 14.4 46.55 57.915 46.62 ;
      RECT 14.4 46.62 57.845 46.69 ;
      RECT 14.4 46.69 57.775 46.76 ;
      RECT 14.4 46.76 57.705 46.83 ;
      RECT 14.4 46.83 57.635 46.9 ;
      RECT 14.4 46.9 57.565 46.97 ;
      RECT 14.4 46.97 57.495 47.04 ;
      RECT 14.4 47.04 57.425 47.11 ;
      RECT 14.4 47.11 57.36 47.175 ;
      RECT 28.26 12.015 37.61 12.065 ;
      RECT 28.31 12.065 37.61 12.115 ;
      RECT 28.315 12.115 37.61 12.12 ;
      RECT 37.175 25.94 55.7 25.96 ;
      RECT 37.175 25.96 55.72 25.98 ;
      RECT 56.985 158.755 60.825 158.76 ;
      RECT 56.985 151.88 60.815 151.895 ;
      RECT 56.985 151.81 60.745 151.88 ;
      RECT 56.985 151.74 60.675 151.81 ;
      RECT 56.985 151.67 60.605 151.74 ;
      RECT 56.985 151.6 60.535 151.67 ;
      RECT 56.985 151.53 60.465 151.6 ;
      RECT 56.985 151.46 60.395 151.53 ;
      RECT 56.985 151.39 60.325 151.46 ;
      RECT 56.985 151.32 60.255 151.39 ;
      RECT 56.985 151.25 60.185 151.32 ;
      RECT 56.985 151.18 60.115 151.25 ;
      RECT 56.985 151.11 60.045 151.18 ;
      RECT 56.985 151.04 59.975 151.11 ;
      RECT 56.985 150.97 59.905 151.04 ;
      RECT 56.985 150.9 59.835 150.97 ;
      RECT 56.985 150.83 59.765 150.9 ;
      RECT 56.985 150.76 59.695 150.83 ;
      RECT 56.985 150.69 59.625 150.76 ;
      RECT 56.985 150.62 59.555 150.69 ;
      RECT 56.985 150.55 59.485 150.62 ;
      RECT 56.985 150.48 59.415 150.55 ;
      RECT 56.985 150.41 59.345 150.48 ;
      RECT 56.985 150.34 59.275 150.41 ;
      RECT 56.985 150.27 59.205 150.34 ;
      RECT 56.985 150.2 59.135 150.27 ;
      RECT 56.985 150.13 59.065 150.2 ;
      RECT 56.985 150.06 58.995 150.13 ;
      RECT 56.985 149.99 58.925 150.06 ;
      RECT 56.985 149.92 58.855 149.99 ;
      RECT 56.985 149.85 58.785 149.92 ;
      RECT 56.985 149.78 58.715 149.85 ;
      RECT 56.985 149.71 58.645 149.78 ;
      RECT 56.985 149.64 58.575 149.71 ;
      RECT 56.985 149.57 58.505 149.64 ;
      RECT 56.985 149.5 58.435 149.57 ;
      RECT 56.985 135.74 60.82 135.75 ;
      RECT 56.985 135.75 60.81 135.76 ;
      RECT 56.985 128.81 60.815 128.825 ;
      RECT 56.985 128.74 60.745 128.81 ;
      RECT 56.985 128.67 60.675 128.74 ;
      RECT 56.985 128.6 60.605 128.67 ;
      RECT 56.985 128.53 60.535 128.6 ;
      RECT 56.985 128.46 60.465 128.53 ;
      RECT 56.985 128.39 60.395 128.46 ;
      RECT 56.985 128.32 60.325 128.39 ;
      RECT 56.985 128.25 60.255 128.32 ;
      RECT 56.985 128.18 60.185 128.25 ;
      RECT 56.985 128.11 60.115 128.18 ;
      RECT 56.985 128.04 60.045 128.11 ;
      RECT 56.985 127.97 59.975 128.04 ;
      RECT 56.985 127.9 59.905 127.97 ;
      RECT 56.985 127.83 59.835 127.9 ;
      RECT 56.985 127.76 59.765 127.83 ;
      RECT 56.985 127.69 59.695 127.76 ;
      RECT 56.985 127.62 59.625 127.69 ;
      RECT 56.985 127.55 59.555 127.62 ;
      RECT 56.985 127.48 59.485 127.55 ;
      RECT 56.985 127.41 59.415 127.48 ;
      RECT 56.985 127.34 59.345 127.41 ;
      RECT 56.985 127.27 59.275 127.34 ;
      RECT 56.985 127.2 59.205 127.27 ;
      RECT 56.985 127.13 59.135 127.2 ;
      RECT 56.985 127.06 59.065 127.13 ;
      RECT 56.985 126.99 58.995 127.06 ;
      RECT 56.985 126.92 58.925 126.99 ;
      RECT 56.985 126.85 58.855 126.92 ;
      RECT 56.985 126.78 58.785 126.85 ;
      RECT 56.985 126.71 58.715 126.78 ;
      RECT 18.845 38.84 53.62 38.91 ;
      RECT 18.915 38.91 53.55 38.98 ;
      RECT 18.985 38.98 53.48 39.05 ;
      RECT 19.055 39.05 53.41 39.12 ;
      RECT 19.125 39.12 53.34 39.19 ;
      RECT 19.195 39.19 53.27 39.26 ;
      RECT 19.265 39.26 53.2 39.33 ;
      RECT 19.335 39.33 53.13 39.4 ;
      RECT 19.405 39.4 53.06 39.47 ;
      RECT 19.475 39.47 52.99 39.54 ;
      RECT 19.545 39.54 52.92 39.61 ;
      RECT 19.615 39.61 52.85 39.68 ;
      RECT 19.685 39.68 52.78 39.75 ;
      RECT 19.755 39.75 52.71 39.82 ;
      RECT 19.825 39.82 52.64 39.89 ;
      RECT 19.895 39.89 52.57 39.96 ;
      RECT 19.965 39.96 52.5 40.03 ;
      RECT 20.005 40.03 52.46 40.07 ;
      RECT 15.84 35.835 54.39 35.905 ;
      RECT 15.91 35.905 54.39 35.975 ;
      RECT 15.98 35.975 54.39 36.045 ;
      RECT 16.05 36.045 54.39 36.115 ;
      RECT 16.12 36.115 54.39 36.185 ;
      RECT 16.19 36.185 54.39 36.255 ;
      RECT 16.26 36.255 54.39 36.325 ;
      RECT 16.33 36.325 54.39 36.395 ;
      RECT 16.4 36.395 54.39 36.465 ;
      RECT 16.47 36.465 54.39 36.535 ;
      RECT 16.54 36.535 54.39 36.605 ;
      RECT 16.61 36.605 54.39 36.675 ;
      RECT 16.68 36.675 54.39 36.745 ;
      RECT 16.75 36.745 54.39 36.815 ;
      RECT 16.82 36.815 54.39 36.885 ;
      RECT 16.89 36.885 54.39 36.955 ;
      RECT 16.96 36.955 54.39 37.025 ;
      RECT 17.03 37.025 54.39 37.095 ;
      RECT 17.1 37.095 54.39 37.165 ;
      RECT 17.17 37.165 54.39 37.235 ;
      RECT 17.24 37.235 54.39 37.305 ;
      RECT 17.31 37.305 54.39 37.375 ;
      RECT 17.38 37.375 54.39 37.445 ;
      RECT 17.45 37.445 54.39 37.515 ;
      RECT 17.52 37.515 54.39 37.585 ;
      RECT 17.59 37.585 54.39 37.655 ;
      RECT 17.66 37.655 54.39 37.725 ;
      RECT 17.73 37.725 54.39 37.795 ;
      RECT 17.8 37.795 54.39 37.865 ;
      RECT 17.87 37.865 54.39 37.935 ;
      RECT 17.94 37.935 54.39 38.005 ;
      RECT 18.01 38.005 54.39 38.075 ;
      RECT 18.075 38.075 54.39 38.14 ;
      RECT 15.505 29.41 59.17 29.43 ;
      RECT 15.575 29.34 59.1 29.41 ;
      RECT 15.645 29.27 59.03 29.34 ;
      RECT 15.715 29.2 58.96 29.27 ;
      RECT 15.785 29.13 58.89 29.2 ;
      RECT 15.855 29.06 58.82 29.13 ;
      RECT 15.925 28.99 58.75 29.06 ;
      RECT 15.995 28.92 58.68 28.99 ;
      RECT 16.065 28.85 58.61 28.92 ;
      RECT 16.135 28.78 58.54 28.85 ;
      RECT 16.205 28.71 58.47 28.78 ;
      RECT 16.275 28.64 58.4 28.71 ;
      RECT 16.345 28.57 58.33 28.64 ;
      RECT 16.415 28.5 58.26 28.57 ;
      RECT 16.485 28.43 58.19 28.5 ;
      RECT 16.555 28.36 58.12 28.43 ;
      RECT 16.625 28.29 58.05 28.36 ;
      RECT 16.695 28.22 57.98 28.29 ;
      RECT 16.765 28.15 57.91 28.22 ;
      RECT 16.835 28.08 57.84 28.15 ;
      RECT 16.905 28.01 57.77 28.08 ;
      RECT 16.975 27.94 57.7 28.01 ;
      RECT 17.045 27.87 57.63 27.94 ;
      RECT 17.115 27.8 57.56 27.87 ;
      RECT 17.185 27.73 57.49 27.8 ;
      RECT 17.255 27.66 57.42 27.73 ;
      RECT 17.325 27.59 57.35 27.66 ;
      RECT 17.395 27.52 57.28 27.59 ;
      RECT 17.465 27.45 57.21 27.52 ;
      RECT 17.535 27.38 57.14 27.45 ;
      RECT 17.605 27.31 57.07 27.38 ;
      RECT 17.675 27.24 57.0 27.31 ;
      RECT 17.745 27.17 56.93 27.24 ;
      RECT 17.815 27.1 56.86 27.17 ;
      RECT 17.885 27.03 56.79 27.1 ;
      RECT 17.955 26.96 56.72 27.03 ;
      RECT 18.025 26.89 56.65 26.96 ;
      RECT 18.095 26.82 56.58 26.89 ;
      RECT 18.165 26.75 56.51 26.82 ;
      RECT 18.235 26.68 56.44 26.75 ;
      RECT 18.305 26.61 56.37 26.68 ;
      RECT 18.375 26.54 56.3 26.61 ;
      RECT 18.445 26.47 56.23 26.54 ;
      RECT 18.515 26.4 56.16 26.47 ;
      RECT 18.585 26.33 56.09 26.4 ;
      RECT 18.655 26.26 56.02 26.33 ;
      RECT 18.725 26.19 55.95 26.26 ;
      RECT 18.795 26.12 55.88 26.19 ;
      RECT 18.865 26.05 55.81 26.12 ;
      RECT 18.935 25.98 55.74 26.05 ;
      RECT 24.775 8.51 50.04 8.58 ;
      RECT 24.845 8.58 49.97 8.65 ;
      RECT 24.915 8.65 49.9 8.72 ;
      RECT 24.985 8.72 49.83 8.79 ;
      RECT 25.055 8.79 49.76 8.86 ;
      RECT 25.125 8.86 49.69 8.93 ;
      RECT 25.195 8.93 49.62 9 ;
      RECT 25.265 9 49.55 9.07 ;
      RECT 25.335 9.07 49.48 9.14 ;
      RECT 25.405 9.14 49.41 9.21 ;
      RECT 25.475 9.21 49.34 9.28 ;
      RECT 25.545 9.28 49.27 9.35 ;
      RECT 25.615 9.35 49.2 9.42 ;
      RECT 25.685 9.42 49.13 9.49 ;
      RECT 25.755 9.49 49.06 9.56 ;
      RECT 25.825 9.56 48.99 9.63 ;
      RECT 25.895 9.63 48.92 9.7 ;
      RECT 25.965 9.7 48.85 9.77 ;
      RECT 26.035 9.77 48.78 9.84 ;
      RECT 26.105 9.84 48.71 9.91 ;
      RECT 26.175 9.91 48.64 9.98 ;
      RECT 26.245 9.98 48.57 10.05 ;
      RECT 26.315 10.05 48.5 10.12 ;
      RECT 26.385 10.12 48.43 10.19 ;
      RECT 26.455 10.19 48.36 10.26 ;
      RECT 17.2 79.855 24.54 79.925 ;
      RECT 17.27 79.925 24.54 79.995 ;
      RECT 17.34 79.995 24.54 80.065 ;
      RECT 17.41 80.065 24.54 80.135 ;
      RECT 17.48 80.135 24.54 80.205 ;
      RECT 17.55 80.205 24.54 80.275 ;
      RECT 17.62 80.275 24.54 80.345 ;
      RECT 17.69 80.345 24.54 80.415 ;
      RECT 17.76 80.415 24.54 80.485 ;
      RECT 17.775 80.485 24.54 80.5 ;
      RECT 14.42 70.12 57.425 70.14 ;
      RECT 14.49 70.05 57.445 70.12 ;
      RECT 14.56 69.98 57.515 70.05 ;
      RECT 14.63 69.91 57.585 69.98 ;
      RECT 14.7 69.84 57.655 69.91 ;
      RECT 14.77 69.77 57.725 69.84 ;
      RECT 14.84 69.7 57.795 69.77 ;
      RECT 14.91 69.63 57.865 69.7 ;
      RECT 14.98 69.56 57.935 69.63 ;
      RECT 15.05 69.49 58.005 69.56 ;
      RECT 15.12 69.42 58.075 69.49 ;
      RECT 15.19 69.35 58.145 69.42 ;
      RECT 15.26 69.28 58.215 69.35 ;
      RECT 15.33 69.21 58.285 69.28 ;
      RECT 15.4 69.14 58.355 69.21 ;
      RECT 15.47 69.07 58.425 69.14 ;
      RECT 15.54 69 58.495 69.07 ;
      RECT 15.61 68.93 58.565 69 ;
      RECT 15.68 68.86 58.635 68.93 ;
      RECT 15.75 68.79 58.705 68.86 ;
      RECT 15.82 68.72 58.775 68.79 ;
      RECT 15.89 68.65 58.845 68.72 ;
      RECT 15.96 68.58 58.915 68.65 ;
      RECT 16.03 68.51 58.985 68.58 ;
      RECT 16.1 68.44 59.055 68.51 ;
      RECT 16.17 68.37 59.125 68.44 ;
      RECT 16.24 68.3 59.195 68.37 ;
      RECT 16.31 68.23 59.265 68.3 ;
      RECT 16.38 68.16 59.335 68.23 ;
      RECT 16.45 68.09 59.405 68.16 ;
      RECT 16.52 68.02 59.475 68.09 ;
      RECT 16.59 67.95 59.545 68.02 ;
      RECT 16.66 67.88 59.615 67.95 ;
      RECT 16.73 67.81 59.685 67.88 ;
      RECT 16.8 67.74 59.755 67.81 ;
      RECT 16.87 67.67 59.825 67.74 ;
      RECT 16.94 67.6 59.895 67.67 ;
      RECT 17.01 67.53 59.965 67.6 ;
      RECT 17.08 67.46 60.035 67.53 ;
      RECT 17.15 67.39 60.105 67.46 ;
      RECT 17.22 67.32 60.175 67.39 ;
      RECT 17.29 67.25 60.245 67.32 ;
      RECT 17.36 67.18 60.315 67.25 ;
      RECT 17.43 67.11 60.385 67.18 ;
      RECT 17.5 67.04 60.455 67.11 ;
      RECT 17.57 66.97 60.525 67.04 ;
      RECT 17.64 66.9 60.595 66.97 ;
      RECT 17.71 66.83 60.665 66.9 ;
      RECT 17.78 66.76 60.735 66.83 ;
      RECT 56.99 56.435 57.41 56.505 ;
      RECT 56.99 56.505 57.48 56.575 ;
      RECT 56.99 56.575 57.55 56.645 ;
      RECT 56.99 56.645 57.62 56.715 ;
      RECT 56.99 56.715 57.69 56.785 ;
      RECT 56.99 56.785 57.76 56.855 ;
      RECT 56.99 56.855 57.83 56.925 ;
      RECT 56.99 56.925 57.9 56.995 ;
      RECT 56.99 56.995 57.97 57.065 ;
      RECT 56.99 57.065 58.04 57.135 ;
      RECT 56.99 57.135 58.11 57.205 ;
      RECT 56.99 57.205 58.18 57.275 ;
      RECT 56.99 57.275 58.25 57.345 ;
      RECT 56.99 57.345 58.32 57.415 ;
      RECT 56.99 57.415 58.39 57.485 ;
      RECT 56.99 57.485 58.46 57.5 ;
      RECT 16.125 43.705 60.76 43.775 ;
      RECT 16.055 43.775 60.69 43.845 ;
      RECT 15.985 43.845 60.62 43.915 ;
      RECT 15.915 43.915 60.55 43.985 ;
      RECT 15.845 43.985 60.48 44.055 ;
      RECT 15.775 44.055 60.41 44.125 ;
      RECT 15.705 44.125 60.34 44.195 ;
      RECT 15.635 44.195 60.27 44.265 ;
      RECT 15.565 44.265 60.2 44.335 ;
      RECT 15.495 44.335 60.13 44.405 ;
      RECT 15.425 44.405 60.06 44.475 ;
      RECT 15.355 44.475 59.99 44.545 ;
      RECT 15.285 44.545 59.92 44.615 ;
      RECT 15.215 44.615 59.85 44.685 ;
      RECT 15.145 44.685 59.78 44.755 ;
      RECT 15.075 44.755 59.71 44.825 ;
      RECT 15.005 44.825 59.64 44.895 ;
      RECT 14.935 44.895 59.57 44.965 ;
      RECT 14.865 44.965 59.5 45.035 ;
      RECT 14.795 45.035 59.43 45.105 ;
      RECT 14.725 45.105 59.36 45.175 ;
      RECT 14.655 45.175 59.29 45.245 ;
      RECT 14.585 45.245 59.22 45.315 ;
      RECT 14.515 45.315 59.15 45.385 ;
      RECT 14.445 45.385 59.105 45.43 ;
      RECT 17.17 42.66 60.83 42.73 ;
      RECT 17.1 42.73 60.83 42.8 ;
      RECT 17.03 42.8 60.83 42.87 ;
      RECT 16.96 42.87 60.83 42.94 ;
      RECT 16.89 42.94 60.83 43.01 ;
      RECT 16.82 43.01 60.83 43.08 ;
      RECT 16.75 43.08 60.83 43.15 ;
      RECT 16.68 43.15 60.83 43.22 ;
      RECT 16.61 43.22 60.83 43.29 ;
      RECT 16.54 43.29 60.83 43.36 ;
      RECT 16.47 43.36 60.83 43.43 ;
      RECT 16.4 43.43 60.83 43.5 ;
      RECT 16.33 43.5 60.83 43.57 ;
      RECT 16.26 43.57 60.83 43.64 ;
      RECT 16.19 43.64 60.83 43.705 ;
      RECT 18.145 38.14 54.32 38.21 ;
      RECT 18.215 38.21 54.25 38.28 ;
      RECT 18.285 38.28 54.18 38.35 ;
      RECT 18.355 38.35 54.11 38.42 ;
      RECT 18.425 38.42 54.04 38.49 ;
      RECT 18.495 38.49 53.97 38.56 ;
      RECT 18.565 38.56 53.9 38.63 ;
      RECT 18.635 38.63 53.83 38.7 ;
      RECT 18.705 38.7 53.76 38.77 ;
      RECT 18.775 38.77 53.69 38.84 ;
      RECT 16.07 114.51 58.955 114.58 ;
      RECT 16.0 114.58 58.885 114.65 ;
      RECT 15.93 114.65 58.815 114.72 ;
      RECT 15.86 114.72 58.745 114.79 ;
      RECT 15.79 114.79 58.675 114.86 ;
      RECT 15.72 114.86 58.605 114.93 ;
      RECT 15.65 114.93 58.535 115 ;
      RECT 15.58 115 58.465 115.07 ;
      RECT 15.51 115.07 58.395 115.14 ;
      RECT 15.44 115.14 58.325 115.21 ;
      RECT 15.37 115.21 58.255 115.28 ;
      RECT 15.3 115.28 58.185 115.35 ;
      RECT 15.23 115.35 58.115 115.42 ;
      RECT 15.16 115.42 58.045 115.49 ;
      RECT 15.09 115.49 57.975 115.56 ;
      RECT 15.02 115.56 57.905 115.63 ;
      RECT 14.95 115.63 57.835 115.7 ;
      RECT 14.88 115.7 57.765 115.77 ;
      RECT 14.81 115.77 57.695 115.84 ;
      RECT 14.74 115.84 57.625 115.91 ;
      RECT 14.67 115.91 57.555 115.98 ;
      RECT 14.6 115.98 57.485 116.05 ;
      RECT 14.53 116.05 57.415 116.12 ;
      RECT 14.46 116.12 57.36 116.175 ;
      RECT 56.985 102.435 57.44 102.505 ;
      RECT 56.985 102.505 57.51 102.575 ;
      RECT 56.985 102.575 57.58 102.645 ;
      RECT 56.985 102.645 57.65 102.715 ;
      RECT 56.985 102.715 57.72 102.785 ;
      RECT 56.985 102.785 57.79 102.855 ;
      RECT 56.985 102.855 57.86 102.925 ;
      RECT 56.985 102.925 57.93 102.995 ;
      RECT 56.985 102.995 58.0 103.065 ;
      RECT 56.985 103.065 58.07 103.135 ;
      RECT 56.985 103.135 58.14 103.205 ;
      RECT 56.985 103.205 58.21 103.275 ;
      RECT 56.985 103.275 58.28 103.345 ;
      RECT 56.985 103.345 58.35 103.415 ;
      RECT 56.985 103.415 58.42 103.485 ;
      RECT 56.985 103.485 58.49 103.5 ;
      RECT 16.78 102.435 24.54 102.505 ;
      RECT 16.85 102.505 24.54 102.575 ;
      RECT 16.92 102.575 24.54 102.645 ;
      RECT 16.99 102.645 24.54 102.715 ;
      RECT 17.06 102.715 24.54 102.785 ;
      RECT 17.13 102.785 24.54 102.855 ;
      RECT 17.2 102.855 24.54 102.925 ;
      RECT 17.27 102.925 24.54 102.995 ;
      RECT 17.34 102.995 24.54 103.065 ;
      RECT 17.41 103.065 24.54 103.135 ;
      RECT 17.48 103.135 24.54 103.205 ;
      RECT 17.55 103.205 24.54 103.275 ;
      RECT 17.62 103.275 24.54 103.345 ;
      RECT 17.69 103.345 24.54 103.415 ;
      RECT 17.76 103.415 24.54 103.485 ;
      RECT 17.775 103.485 24.54 103.5 ;
      RECT 14.455 93.085 57.485 93.14 ;
      RECT 14.525 93.015 57.54 93.085 ;
      RECT 14.595 92.945 57.61 93.015 ;
      RECT 14.665 92.875 57.68 92.945 ;
      RECT 14.735 92.805 57.75 92.875 ;
      RECT 14.805 92.735 57.82 92.805 ;
      RECT 14.875 92.665 57.89 92.735 ;
      RECT 14.945 92.595 57.96 92.665 ;
      RECT 15.015 92.525 58.03 92.595 ;
      RECT 15.085 92.455 58.1 92.525 ;
      RECT 15.155 92.385 58.17 92.455 ;
      RECT 15.225 92.315 58.24 92.385 ;
      RECT 15.295 92.245 58.31 92.315 ;
      RECT 15.365 92.175 58.38 92.245 ;
      RECT 15.435 92.105 58.45 92.175 ;
      RECT 15.505 92.035 58.52 92.105 ;
      RECT 15.575 91.965 58.59 92.035 ;
      RECT 15.645 91.895 58.66 91.965 ;
      RECT 15.715 91.825 58.73 91.895 ;
      RECT 15.785 91.755 58.8 91.825 ;
      RECT 15.855 91.685 58.87 91.755 ;
      RECT 15.925 91.615 58.94 91.685 ;
      RECT 15.995 91.545 59.01 91.615 ;
      RECT 16.065 91.475 59.08 91.545 ;
      RECT 16.135 91.405 59.15 91.475 ;
      RECT 16.205 91.335 59.22 91.405 ;
      RECT 16.275 91.265 59.29 91.335 ;
      RECT 16.345 91.195 59.36 91.265 ;
      RECT 16.415 91.125 59.43 91.195 ;
      RECT 16.485 91.055 59.5 91.125 ;
      RECT 16.555 90.985 59.57 91.055 ;
      RECT 16.625 90.915 59.64 90.985 ;
      RECT 16.695 90.845 59.71 90.915 ;
      RECT 16.765 90.775 59.78 90.845 ;
      RECT 16.835 90.705 59.85 90.775 ;
      RECT 16.905 90.635 59.92 90.705 ;
      RECT 16.975 90.565 59.99 90.635 ;
      RECT 17.045 90.495 60.06 90.565 ;
      RECT 17.115 90.425 60.13 90.495 ;
      RECT 17.185 90.355 60.2 90.425 ;
      RECT 17.255 90.285 60.27 90.355 ;
      RECT 17.325 90.215 60.34 90.285 ;
      RECT 17.395 90.145 60.41 90.215 ;
      RECT 17.465 90.075 60.48 90.145 ;
      RECT 17.535 90.005 60.55 90.075 ;
      RECT 17.605 89.935 60.62 90.005 ;
      RECT 17.675 89.865 60.69 89.935 ;
      RECT 17.745 89.795 60.76 89.865 ;
      RECT 56.985 79.435 57.44 79.505 ;
      RECT 56.985 79.505 57.51 79.575 ;
      RECT 56.985 79.575 57.58 79.645 ;
      RECT 56.985 79.645 57.65 79.715 ;
      RECT 56.985 79.715 57.72 79.785 ;
      RECT 56.985 79.785 57.79 79.855 ;
      RECT 56.985 79.855 57.86 79.925 ;
      RECT 56.985 79.925 57.93 79.995 ;
      RECT 56.985 79.995 58.0 80.065 ;
      RECT 56.985 80.065 58.07 80.135 ;
      RECT 56.985 80.135 58.14 80.205 ;
      RECT 56.985 80.205 58.21 80.275 ;
      RECT 56.985 80.275 58.28 80.345 ;
      RECT 56.985 80.345 58.35 80.415 ;
      RECT 56.985 80.415 58.42 80.485 ;
      RECT 56.985 80.485 58.49 80.5 ;
      RECT 16.78 79.435 24.54 79.505 ;
      RECT 16.85 79.505 24.54 79.575 ;
      RECT 16.92 79.575 24.54 79.645 ;
      RECT 16.99 79.645 24.54 79.715 ;
      RECT 17.06 79.715 24.54 79.785 ;
      RECT 17.13 79.785 24.54 79.855 ;
      RECT 14.755 161.84 57.675 161.91 ;
      RECT 14.685 161.91 57.605 161.98 ;
      RECT 14.615 161.98 57.535 162.05 ;
      RECT 14.545 162.05 57.465 162.12 ;
      RECT 14.475 162.12 57.41 162.175 ;
      RECT 56.985 148.435 57.37 148.505 ;
      RECT 56.985 148.505 57.44 148.575 ;
      RECT 56.985 148.575 57.51 148.645 ;
      RECT 56.985 148.645 57.58 148.715 ;
      RECT 56.985 148.715 57.65 148.785 ;
      RECT 56.985 148.785 57.72 148.855 ;
      RECT 56.985 148.855 57.79 148.925 ;
      RECT 56.985 148.925 57.86 148.995 ;
      RECT 56.985 148.995 57.93 149.065 ;
      RECT 56.985 149.065 58.0 149.135 ;
      RECT 56.985 149.135 58.07 149.205 ;
      RECT 56.985 149.205 58.14 149.275 ;
      RECT 56.985 149.275 58.21 149.345 ;
      RECT 56.985 149.345 58.28 149.415 ;
      RECT 56.985 149.415 58.35 149.485 ;
      RECT 56.985 149.485 58.42 149.5 ;
      RECT 17.925 135.76 60.74 135.83 ;
      RECT 17.855 135.83 60.67 135.9 ;
      RECT 17.785 135.9 60.6 135.97 ;
      RECT 17.715 135.97 60.53 136.04 ;
      RECT 17.645 136.04 60.46 136.11 ;
      RECT 17.575 136.11 60.39 136.18 ;
      RECT 17.505 136.18 60.32 136.25 ;
      RECT 17.435 136.25 60.25 136.32 ;
      RECT 17.365 136.32 60.18 136.39 ;
      RECT 17.295 136.39 60.11 136.46 ;
      RECT 17.225 136.46 60.04 136.53 ;
      RECT 17.155 136.53 59.97 136.6 ;
      RECT 17.085 136.6 59.9 136.67 ;
      RECT 17.015 136.67 59.83 136.74 ;
      RECT 16.945 136.74 59.76 136.81 ;
      RECT 16.875 136.81 59.69 136.88 ;
      RECT 16.805 136.88 59.62 136.95 ;
      RECT 16.735 136.95 59.55 137.02 ;
      RECT 16.665 137.02 59.48 137.09 ;
      RECT 16.595 137.09 59.41 137.16 ;
      RECT 16.525 137.16 59.34 137.23 ;
      RECT 16.455 137.23 59.27 137.3 ;
      RECT 16.385 137.3 59.2 137.37 ;
      RECT 16.315 137.37 59.13 137.44 ;
      RECT 16.245 137.44 59.06 137.51 ;
      RECT 16.175 137.51 58.99 137.58 ;
      RECT 16.105 137.58 58.92 137.65 ;
      RECT 16.035 137.65 58.85 137.72 ;
      RECT 15.965 137.72 58.78 137.79 ;
      RECT 15.895 137.79 58.71 137.86 ;
      RECT 15.825 137.86 58.64 137.93 ;
      RECT 15.755 137.93 58.57 138 ;
      RECT 15.685 138 58.5 138.07 ;
      RECT 15.615 138.07 58.43 138.14 ;
      RECT 15.545 138.14 58.36 138.21 ;
      RECT 15.475 138.21 58.29 138.28 ;
      RECT 15.405 138.28 58.22 138.35 ;
      RECT 15.335 138.35 58.15 138.42 ;
      RECT 15.265 138.42 58.08 138.49 ;
      RECT 15.195 138.49 58.01 138.56 ;
      RECT 15.125 138.56 57.94 138.63 ;
      RECT 15.055 138.63 57.87 138.7 ;
      RECT 14.985 138.7 57.8 138.77 ;
      RECT 14.915 138.77 57.73 138.84 ;
      RECT 14.845 138.84 57.66 138.91 ;
      RECT 14.775 138.91 57.59 138.98 ;
      RECT 14.705 138.98 57.52 139.05 ;
      RECT 14.635 139.05 57.45 139.12 ;
      RECT 14.565 139.12 57.395 139.175 ;
      RECT 56.985 125.435 57.44 125.505 ;
      RECT 56.985 125.505 57.51 125.575 ;
      RECT 56.985 125.575 57.58 125.645 ;
      RECT 56.985 125.645 57.65 125.715 ;
      RECT 56.985 125.715 57.72 125.785 ;
      RECT 56.985 125.785 57.79 125.855 ;
      RECT 56.985 125.855 57.86 125.925 ;
      RECT 56.985 125.925 57.93 125.995 ;
      RECT 56.985 125.995 58.0 126.065 ;
      RECT 56.985 126.065 58.07 126.135 ;
      RECT 56.985 126.135 58.14 126.205 ;
      RECT 56.985 126.205 58.21 126.275 ;
      RECT 56.985 126.275 58.28 126.345 ;
      RECT 56.985 126.345 58.35 126.415 ;
      RECT 56.985 126.415 58.42 126.485 ;
      RECT 56.985 126.485 58.49 126.5 ;
      RECT 16.875 125.435 24.54 125.505 ;
      RECT 16.945 125.505 24.54 125.575 ;
      RECT 17.015 125.575 24.54 125.645 ;
      RECT 17.085 125.645 24.54 125.715 ;
      RECT 17.155 125.715 24.54 125.785 ;
      RECT 17.225 125.785 24.54 125.855 ;
      RECT 17.295 125.855 24.54 125.925 ;
      RECT 17.365 125.925 24.54 125.995 ;
      RECT 17.435 125.995 24.54 126.065 ;
      RECT 17.505 126.065 24.54 126.135 ;
      RECT 17.575 126.135 24.54 126.205 ;
      RECT 17.645 126.205 24.54 126.275 ;
      RECT 17.715 126.275 24.54 126.345 ;
      RECT 17.785 126.345 24.54 126.415 ;
      RECT 17.855 126.415 24.54 126.485 ;
      RECT 17.87 126.485 24.54 126.5 ;
      RECT 17.82 112.76 60.705 112.83 ;
      RECT 17.75 112.83 60.635 112.9 ;
      RECT 17.68 112.9 60.565 112.97 ;
      RECT 17.61 112.97 60.495 113.04 ;
      RECT 17.54 113.04 60.425 113.11 ;
      RECT 17.47 113.11 60.355 113.18 ;
      RECT 17.4 113.18 60.285 113.25 ;
      RECT 17.33 113.25 60.215 113.32 ;
      RECT 17.26 113.32 60.145 113.39 ;
      RECT 17.19 113.39 60.075 113.46 ;
      RECT 17.12 113.46 60.005 113.53 ;
      RECT 17.05 113.53 59.935 113.6 ;
      RECT 16.98 113.6 59.865 113.67 ;
      RECT 16.91 113.67 59.795 113.74 ;
      RECT 16.84 113.74 59.725 113.81 ;
      RECT 16.77 113.81 59.655 113.88 ;
      RECT 16.7 113.88 59.585 113.95 ;
      RECT 16.63 113.95 59.515 114.02 ;
      RECT 16.56 114.02 59.445 114.09 ;
      RECT 16.49 114.09 59.375 114.16 ;
      RECT 16.42 114.16 59.305 114.23 ;
      RECT 16.35 114.23 59.235 114.3 ;
      RECT 16.28 114.3 59.165 114.37 ;
      RECT 16.21 114.37 59.095 114.44 ;
      RECT 16.14 114.44 59.025 114.51 ;
      RECT 17.745 27.17 56.93 27.24 ;
      RECT 17.815 27.1 56.86 27.17 ;
      RECT 17.885 27.03 56.79 27.1 ;
      RECT 17.955 26.96 56.72 27.03 ;
      RECT 18.025 26.89 56.65 26.96 ;
      RECT 18.095 26.82 56.58 26.89 ;
      RECT 18.165 26.75 56.51 26.82 ;
      RECT 18.235 26.68 56.44 26.75 ;
      RECT 18.305 26.61 56.37 26.68 ;
      RECT 18.375 26.54 56.3 26.61 ;
      RECT 18.445 26.47 56.23 26.54 ;
      RECT 18.515 26.4 56.16 26.47 ;
      RECT 18.585 26.33 56.09 26.4 ;
      RECT 18.655 26.26 56.02 26.33 ;
      RECT 18.725 26.19 55.95 26.26 ;
      RECT 18.795 26.12 55.88 26.19 ;
      RECT 18.865 26.05 55.81 26.12 ;
      RECT 18.935 25.98 55.74 26.05 ;
      RECT 37.175 25.94 55.7 25.96 ;
      RECT 37.175 25.96 55.72 25.98 ;
      RECT 28.26 12.015 37.61 12.065 ;
      RECT 28.31 12.065 37.61 12.115 ;
      RECT 28.315 12.115 37.61 12.12 ;
      RECT 24.775 8.51 50.04 8.58 ;
      RECT 24.845 8.58 49.97 8.65 ;
      RECT 24.915 8.65 49.9 8.72 ;
      RECT 24.985 8.72 49.83 8.79 ;
      RECT 25.055 8.79 49.76 8.86 ;
      RECT 25.125 8.86 49.69 8.93 ;
      RECT 25.195 8.93 49.62 9 ;
      RECT 25.265 9 49.55 9.07 ;
      RECT 25.335 9.07 49.48 9.14 ;
      RECT 25.405 9.14 49.41 9.21 ;
      RECT 25.475 9.21 49.34 9.28 ;
      RECT 25.545 9.28 49.27 9.35 ;
      RECT 25.615 9.35 49.2 9.42 ;
      RECT 25.685 9.42 49.13 9.49 ;
      RECT 25.755 9.49 49.06 9.56 ;
      RECT 25.825 9.56 48.99 9.63 ;
      RECT 25.895 9.63 48.92 9.7 ;
      RECT 25.965 9.7 48.85 9.77 ;
      RECT 26.035 9.77 48.78 9.84 ;
      RECT 26.105 9.84 48.71 9.91 ;
      RECT 26.175 9.91 48.64 9.98 ;
      RECT 26.245 9.98 48.57 10.05 ;
      RECT 26.315 10.05 48.5 10.12 ;
      RECT 26.385 10.12 48.43 10.19 ;
      RECT 26.455 10.19 48.36 10.26 ;
      RECT 26.525 10.26 48.29 10.33 ;
      RECT 26.595 10.33 48.22 10.4 ;
      RECT 26.665 10.4 48.15 10.47 ;
      RECT 26.735 10.47 48.08 10.54 ;
      RECT 26.805 10.54 48.01 10.61 ;
      RECT 26.875 10.61 47.94 10.68 ;
      RECT 26.945 10.68 47.87 10.75 ;
      RECT 27.015 10.75 47.8 10.82 ;
      RECT 27.085 10.82 47.73 10.89 ;
      RECT 27.155 10.89 47.66 10.96 ;
      RECT 27.225 10.96 47.59 11.03 ;
      RECT 27.295 11.03 47.52 11.1 ;
      RECT 27.365 11.1 47.45 11.17 ;
      RECT 27.435 11.17 47.38 11.24 ;
      RECT 27.505 11.24 47.31 11.31 ;
      RECT 27.575 11.31 47.24 11.38 ;
      RECT 27.645 11.38 47.17 11.45 ;
      RECT 27.715 11.45 47.1 11.52 ;
      RECT 27.785 11.52 47.03 11.59 ;
      RECT 27.855 11.59 46.96 11.66 ;
      RECT 27.925 11.66 46.89 11.73 ;
      RECT 27.995 11.73 46.82 11.8 ;
      RECT 28.065 11.8 46.75 11.87 ;
      RECT 28.135 11.87 46.68 11.94 ;
      RECT 28.205 11.94 46.61 12.01 ;
      RECT 28.21 12.01 46.605 12.015 ;
      RECT 24.69 8.48 50.11 8.495 ;
      RECT 24.705 8.495 50.11 8.51 ;
      RECT 56.985 158.755 60.825 158.76 ;
      RECT 56.985 135.74 60.82 135.75 ;
      RECT 56.985 135.75 60.81 135.76 ;
      RECT 56.985 112.705 60.805 112.73 ;
      RECT 56.985 112.73 60.775 112.76 ;
      RECT 56.99 66.735 60.82 66.745 ;
      RECT 56.99 66.745 60.805 66.76 ;
      RECT 17.835 158.76 60.755 158.83 ;
      RECT 17.765 158.83 60.685 158.9 ;
      RECT 17.695 158.9 60.615 158.97 ;
      RECT 17.625 158.97 60.545 159.04 ;
      RECT 17.555 159.04 60.475 159.11 ;
      RECT 17.485 159.11 60.405 159.18 ;
      RECT 17.415 159.18 60.335 159.25 ;
      RECT 17.345 159.25 60.265 159.32 ;
      RECT 17.275 159.32 60.195 159.39 ;
      RECT 17.205 159.39 60.125 159.46 ;
      RECT 17.135 159.46 60.055 159.53 ;
      RECT 17.065 159.53 59.985 159.6 ;
      RECT 16.995 159.6 59.915 159.67 ;
      RECT 16.925 159.67 59.845 159.74 ;
      RECT 16.855 159.74 59.775 159.81 ;
      RECT 16.785 159.81 59.705 159.88 ;
      RECT 16.715 159.88 59.635 159.95 ;
      RECT 16.645 159.95 59.565 160.02 ;
      RECT 16.575 160.02 59.495 160.09 ;
      RECT 16.505 160.09 59.425 160.16 ;
      RECT 16.435 160.16 59.355 160.23 ;
      RECT 16.365 160.23 59.285 160.3 ;
      RECT 16.295 160.3 59.215 160.37 ;
      RECT 16.225 160.37 59.145 160.44 ;
      RECT 16.155 160.44 59.075 160.51 ;
      RECT 16.085 160.51 59.005 160.58 ;
      RECT 16.015 160.58 58.935 160.65 ;
      RECT 15.945 160.65 58.865 160.72 ;
      RECT 15.875 160.72 58.795 160.79 ;
      RECT 15.805 160.79 58.725 160.86 ;
      RECT 15.735 160.86 58.655 160.93 ;
      RECT 15.665 160.93 58.585 161 ;
      RECT 15.595 161 58.515 161.07 ;
      RECT 15.525 161.07 58.445 161.14 ;
      RECT 15.455 161.14 58.375 161.21 ;
      RECT 15.385 161.21 58.305 161.28 ;
      RECT 15.315 161.28 58.235 161.35 ;
      RECT 15.245 161.35 58.165 161.42 ;
      RECT 15.175 161.42 58.095 161.49 ;
      RECT 15.105 161.49 58.025 161.56 ;
      RECT 15.035 161.56 57.955 161.63 ;
      RECT 14.965 161.63 57.885 161.7 ;
      RECT 14.895 161.7 57.815 161.77 ;
      RECT 14.825 161.77 57.745 161.84 ;
      RECT 54.465 42.51 60.83 42.58 ;
      RECT 54.395 42.58 60.83 42.65 ;
      RECT 54.325 42.65 60.83 42.66 ;
      RECT 18.145 38.14 54.32 38.21 ;
      RECT 18.215 38.21 54.25 38.28 ;
      RECT 18.285 38.28 54.18 38.35 ;
      RECT 18.355 38.35 54.11 38.42 ;
      RECT 18.425 38.42 54.04 38.49 ;
      RECT 18.495 38.49 53.97 38.56 ;
      RECT 18.565 38.56 53.9 38.63 ;
      RECT 18.635 38.63 53.83 38.7 ;
      RECT 18.705 38.7 53.76 38.77 ;
      RECT 18.775 38.77 53.69 38.84 ;
      RECT 18.845 38.84 53.62 38.91 ;
      RECT 18.915 38.91 53.55 38.98 ;
      RECT 18.985 38.98 53.48 39.05 ;
      RECT 19.055 39.05 53.41 39.12 ;
      RECT 19.125 39.12 53.34 39.19 ;
      RECT 19.195 39.19 53.27 39.26 ;
      RECT 19.265 39.26 53.2 39.33 ;
      RECT 19.335 39.33 53.13 39.4 ;
      RECT 19.405 39.4 53.06 39.47 ;
      RECT 19.475 39.47 52.99 39.54 ;
      RECT 19.545 39.54 52.92 39.61 ;
      RECT 19.615 39.61 52.85 39.68 ;
      RECT 19.685 39.68 52.78 39.75 ;
      RECT 19.755 39.75 52.71 39.82 ;
      RECT 19.825 39.82 52.64 39.89 ;
      RECT 19.895 39.89 52.57 39.96 ;
      RECT 19.965 39.96 52.5 40.03 ;
      RECT 20.005 40.03 52.46 40.07 ;
      RECT 15.84 35.835 54.39 35.905 ;
      RECT 15.91 35.905 54.39 35.975 ;
      RECT 15.98 35.975 54.39 36.045 ;
      RECT 16.05 36.045 54.39 36.115 ;
      RECT 16.12 36.115 54.39 36.185 ;
      RECT 16.19 36.185 54.39 36.255 ;
      RECT 16.26 36.255 54.39 36.325 ;
      RECT 16.33 36.325 54.39 36.395 ;
      RECT 16.4 36.395 54.39 36.465 ;
      RECT 16.47 36.465 54.39 36.535 ;
      RECT 16.54 36.535 54.39 36.605 ;
      RECT 16.61 36.605 54.39 36.675 ;
      RECT 16.68 36.675 54.39 36.745 ;
      RECT 16.75 36.745 54.39 36.815 ;
      RECT 16.82 36.815 54.39 36.885 ;
      RECT 16.89 36.885 54.39 36.955 ;
      RECT 16.96 36.955 54.39 37.025 ;
      RECT 17.03 37.025 54.39 37.095 ;
      RECT 17.1 37.095 54.39 37.165 ;
      RECT 17.17 37.165 54.39 37.235 ;
      RECT 17.24 37.235 54.39 37.305 ;
      RECT 17.31 37.305 54.39 37.375 ;
      RECT 17.38 37.375 54.39 37.445 ;
      RECT 17.45 37.445 54.39 37.515 ;
      RECT 17.52 37.515 54.39 37.585 ;
      RECT 17.59 37.585 54.39 37.655 ;
      RECT 17.66 37.655 54.39 37.725 ;
      RECT 17.73 37.725 54.39 37.795 ;
      RECT 17.8 37.795 54.39 37.865 ;
      RECT 17.87 37.865 54.39 37.935 ;
      RECT 17.94 37.935 54.39 38.005 ;
      RECT 18.01 38.005 54.39 38.075 ;
      RECT 18.075 38.075 54.39 38.14 ;
      RECT 15.555 35.55 60.83 35.62 ;
      RECT 15.625 35.62 60.83 35.69 ;
      RECT 15.695 35.69 60.83 35.76 ;
      RECT 15.765 35.76 60.83 35.83 ;
      RECT 15.77 35.83 60.83 35.835 ;
      RECT 15.485 29.43 59.19 29.5 ;
      RECT 15.485 29.5 59.26 29.57 ;
      RECT 15.485 29.57 59.33 29.64 ;
      RECT 15.485 29.64 59.4 29.71 ;
      RECT 15.485 29.71 59.47 29.78 ;
      RECT 15.485 29.78 59.54 29.85 ;
      RECT 15.485 29.85 59.61 29.92 ;
      RECT 15.485 29.92 59.68 29.99 ;
      RECT 15.485 29.99 59.75 30.06 ;
      RECT 15.485 30.06 59.82 30.13 ;
      RECT 15.485 30.13 59.89 30.2 ;
      RECT 15.485 30.2 59.96 30.27 ;
      RECT 15.485 30.27 60.03 30.34 ;
      RECT 15.485 30.34 60.1 30.41 ;
      RECT 15.485 30.41 60.17 30.48 ;
      RECT 15.485 30.48 60.24 30.55 ;
      RECT 15.485 30.55 60.31 30.62 ;
      RECT 15.485 30.62 60.38 30.69 ;
      RECT 15.485 30.69 60.45 30.76 ;
      RECT 15.485 30.76 60.52 30.83 ;
      RECT 15.485 30.83 60.59 30.9 ;
      RECT 15.485 30.9 60.66 30.97 ;
      RECT 15.485 30.97 60.73 31.04 ;
      RECT 15.485 31.04 60.8 31.07 ;
      RECT 15.505 29.41 59.17 29.43 ;
      RECT 15.575 29.34 59.1 29.41 ;
      RECT 15.645 29.27 59.03 29.34 ;
      RECT 15.715 29.2 58.96 29.27 ;
      RECT 15.785 29.13 58.89 29.2 ;
      RECT 15.855 29.06 58.82 29.13 ;
      RECT 15.925 28.99 58.75 29.06 ;
      RECT 15.995 28.92 58.68 28.99 ;
      RECT 16.065 28.85 58.61 28.92 ;
      RECT 16.135 28.78 58.54 28.85 ;
      RECT 16.205 28.71 58.47 28.78 ;
      RECT 16.275 28.64 58.4 28.71 ;
      RECT 16.345 28.57 58.33 28.64 ;
      RECT 16.415 28.5 58.26 28.57 ;
      RECT 16.485 28.43 58.19 28.5 ;
      RECT 16.555 28.36 58.12 28.43 ;
      RECT 16.625 28.29 58.05 28.36 ;
      RECT 16.695 28.22 57.98 28.29 ;
      RECT 16.765 28.15 57.91 28.22 ;
      RECT 16.835 28.08 57.84 28.15 ;
      RECT 16.905 28.01 57.77 28.08 ;
      RECT 16.975 27.94 57.7 28.01 ;
      RECT 17.045 27.87 57.63 27.94 ;
      RECT 17.115 27.8 57.56 27.87 ;
      RECT 17.185 27.73 57.49 27.8 ;
      RECT 17.255 27.66 57.42 27.73 ;
      RECT 17.325 27.59 57.35 27.66 ;
      RECT 17.395 27.52 57.28 27.59 ;
      RECT 17.465 27.45 57.21 27.52 ;
      RECT 17.535 27.38 57.14 27.45 ;
      RECT 17.605 27.31 57.07 27.38 ;
      RECT 17.675 27.24 57.0 27.31 ;
      RECT 56.99 57.85 58.825 57.92 ;
      RECT 56.99 57.78 58.755 57.85 ;
      RECT 56.99 57.71 58.685 57.78 ;
      RECT 56.99 57.64 58.615 57.71 ;
      RECT 56.99 57.57 58.545 57.64 ;
      RECT 56.99 57.5 58.475 57.57 ;
      RECT 56.99 56.435 57.41 56.505 ;
      RECT 56.99 56.505 57.48 56.575 ;
      RECT 56.99 56.575 57.55 56.645 ;
      RECT 56.99 56.645 57.62 56.715 ;
      RECT 56.99 56.715 57.69 56.785 ;
      RECT 56.99 56.785 57.76 56.855 ;
      RECT 56.99 56.855 57.83 56.925 ;
      RECT 56.99 56.925 57.9 56.995 ;
      RECT 56.99 56.995 57.97 57.065 ;
      RECT 56.99 57.065 58.04 57.135 ;
      RECT 56.99 57.135 58.11 57.205 ;
      RECT 56.99 57.205 58.18 57.275 ;
      RECT 56.99 57.275 58.25 57.345 ;
      RECT 56.99 57.345 58.32 57.415 ;
      RECT 56.99 57.415 58.39 57.485 ;
      RECT 56.99 57.485 58.46 57.5 ;
      RECT 14.4 45.43 59.035 45.5 ;
      RECT 14.4 45.5 58.965 45.57 ;
      RECT 14.4 45.57 58.895 45.64 ;
      RECT 14.4 45.64 58.825 45.71 ;
      RECT 14.4 45.71 58.755 45.78 ;
      RECT 14.4 45.78 58.685 45.85 ;
      RECT 14.4 45.85 58.615 45.92 ;
      RECT 14.4 45.92 58.545 45.99 ;
      RECT 14.4 45.99 58.475 46.06 ;
      RECT 14.4 46.06 58.405 46.13 ;
      RECT 14.4 46.13 58.335 46.2 ;
      RECT 14.4 46.2 58.265 46.27 ;
      RECT 14.4 46.27 58.195 46.34 ;
      RECT 14.4 46.34 58.125 46.41 ;
      RECT 14.4 46.41 58.055 46.48 ;
      RECT 14.4 46.48 57.985 46.55 ;
      RECT 14.4 46.55 57.915 46.62 ;
      RECT 14.4 46.62 57.845 46.69 ;
      RECT 14.4 46.69 57.775 46.76 ;
      RECT 14.4 46.76 57.705 46.83 ;
      RECT 14.4 46.83 57.635 46.9 ;
      RECT 14.4 46.9 57.565 46.97 ;
      RECT 14.4 46.97 57.495 47.04 ;
      RECT 14.4 47.04 57.425 47.11 ;
      RECT 14.4 47.11 57.36 47.175 ;
      RECT 16.125 43.705 60.76 43.775 ;
      RECT 16.055 43.775 60.69 43.845 ;
      RECT 15.985 43.845 60.62 43.915 ;
      RECT 15.915 43.915 60.55 43.985 ;
      RECT 15.845 43.985 60.48 44.055 ;
      RECT 15.775 44.055 60.41 44.125 ;
      RECT 15.705 44.125 60.34 44.195 ;
      RECT 15.635 44.195 60.27 44.265 ;
      RECT 15.565 44.265 60.2 44.335 ;
      RECT 15.495 44.335 60.13 44.405 ;
      RECT 15.425 44.405 60.06 44.475 ;
      RECT 15.355 44.475 59.99 44.545 ;
      RECT 15.285 44.545 59.92 44.615 ;
      RECT 15.215 44.615 59.85 44.685 ;
      RECT 15.145 44.685 59.78 44.755 ;
      RECT 15.075 44.755 59.71 44.825 ;
      RECT 15.005 44.825 59.64 44.895 ;
      RECT 14.935 44.895 59.57 44.965 ;
      RECT 14.865 44.965 59.5 45.035 ;
      RECT 14.795 45.035 59.43 45.105 ;
      RECT 14.725 45.105 59.36 45.175 ;
      RECT 14.655 45.175 59.29 45.245 ;
      RECT 14.585 45.245 59.22 45.315 ;
      RECT 14.515 45.315 59.15 45.385 ;
      RECT 14.445 45.385 59.105 45.43 ;
      RECT 17.17 42.66 60.83 42.73 ;
      RECT 17.1 42.73 60.83 42.8 ;
      RECT 17.03 42.8 60.83 42.87 ;
      RECT 16.96 42.87 60.83 42.94 ;
      RECT 16.89 42.94 60.83 43.01 ;
      RECT 16.82 43.01 60.83 43.08 ;
      RECT 16.75 43.08 60.83 43.15 ;
      RECT 16.68 43.15 60.83 43.22 ;
      RECT 16.61 43.22 60.83 43.29 ;
      RECT 16.54 43.29 60.83 43.36 ;
      RECT 16.47 43.36 60.83 43.43 ;
      RECT 16.4 43.43 60.83 43.5 ;
      RECT 16.33 43.5 60.83 43.57 ;
      RECT 16.26 43.57 60.83 43.64 ;
      RECT 16.19 43.64 60.83 43.705 ;
      RECT 57.195 39.78 60.83 39.85 ;
      RECT 57.125 39.85 60.83 39.92 ;
      RECT 57.055 39.92 60.83 39.99 ;
      RECT 56.985 39.99 60.83 40.06 ;
      RECT 56.915 40.06 60.83 40.13 ;
      RECT 56.845 40.13 60.83 40.2 ;
      RECT 56.775 40.2 60.83 40.27 ;
      RECT 56.705 40.27 60.83 40.34 ;
      RECT 56.635 40.34 60.83 40.41 ;
      RECT 56.565 40.41 60.83 40.48 ;
      RECT 56.495 40.48 60.83 40.55 ;
      RECT 56.425 40.55 60.83 40.62 ;
      RECT 56.355 40.62 60.83 40.69 ;
      RECT 56.285 40.69 60.83 40.76 ;
      RECT 56.215 40.76 60.83 40.83 ;
      RECT 56.145 40.83 60.83 40.9 ;
      RECT 56.075 40.9 60.83 40.97 ;
      RECT 56.005 40.97 60.83 41.04 ;
      RECT 55.935 41.04 60.83 41.11 ;
      RECT 55.865 41.11 60.83 41.18 ;
      RECT 55.795 41.18 60.83 41.25 ;
      RECT 55.725 41.25 60.83 41.32 ;
      RECT 55.655 41.32 60.83 41.39 ;
      RECT 55.585 41.39 60.83 41.46 ;
      RECT 55.515 41.46 60.83 41.53 ;
      RECT 55.445 41.53 60.83 41.6 ;
      RECT 55.375 41.6 60.83 41.67 ;
      RECT 55.305 41.67 60.83 41.74 ;
      RECT 55.235 41.74 60.83 41.81 ;
      RECT 55.165 41.81 60.83 41.88 ;
      RECT 55.095 41.88 60.83 41.95 ;
      RECT 55.025 41.95 60.83 42.02 ;
      RECT 54.955 42.02 60.83 42.09 ;
      RECT 54.885 42.09 60.83 42.16 ;
      RECT 54.815 42.16 60.83 42.23 ;
      RECT 54.745 42.23 60.83 42.3 ;
      RECT 54.675 42.3 60.83 42.37 ;
      RECT 54.605 42.37 60.83 42.44 ;
      RECT 54.535 42.44 60.83 42.51 ;
      RECT 15.73 78.385 24.54 78.455 ;
      RECT 15.8 78.455 24.54 78.525 ;
      RECT 15.87 78.525 24.54 78.595 ;
      RECT 15.94 78.595 24.54 78.665 ;
      RECT 16.01 78.665 24.54 78.735 ;
      RECT 16.08 78.735 24.54 78.805 ;
      RECT 16.15 78.805 24.54 78.875 ;
      RECT 16.22 78.875 24.54 78.945 ;
      RECT 16.29 78.945 24.54 79.015 ;
      RECT 16.36 79.015 24.54 79.085 ;
      RECT 16.43 79.085 24.54 79.155 ;
      RECT 16.5 79.155 24.54 79.225 ;
      RECT 16.57 79.225 24.54 79.295 ;
      RECT 16.64 79.295 24.54 79.365 ;
      RECT 16.71 79.365 24.54 79.435 ;
      RECT 14.4 74.695 23.505 74.765 ;
      RECT 14.4 74.765 23.575 74.835 ;
      RECT 14.4 74.835 23.645 74.905 ;
      RECT 14.4 74.905 23.715 74.975 ;
      RECT 14.4 74.975 23.785 75.045 ;
      RECT 14.4 75.045 23.855 75.115 ;
      RECT 14.4 75.115 23.925 75.185 ;
      RECT 14.4 75.185 23.995 75.255 ;
      RECT 14.4 75.255 24.065 75.325 ;
      RECT 14.4 75.325 24.135 75.395 ;
      RECT 14.4 75.395 24.205 75.465 ;
      RECT 14.4 75.465 24.275 75.535 ;
      RECT 14.4 75.535 24.345 75.605 ;
      RECT 14.4 75.605 24.415 75.675 ;
      RECT 14.4 75.675 24.485 75.73 ;
      RECT 14.4 72.87 24.47 72.94 ;
      RECT 14.4 72.94 24.4 73.01 ;
      RECT 14.4 73.01 24.33 73.08 ;
      RECT 14.4 73.08 24.26 73.15 ;
      RECT 14.4 73.15 24.19 73.22 ;
      RECT 14.4 73.22 24.12 73.29 ;
      RECT 14.4 73.29 24.05 73.36 ;
      RECT 14.4 73.36 23.98 73.43 ;
      RECT 14.4 73.43 23.91 73.5 ;
      RECT 14.4 73.5 23.84 73.57 ;
      RECT 14.4 73.57 23.77 73.64 ;
      RECT 14.4 73.64 23.7 73.71 ;
      RECT 14.4 73.71 23.63 73.78 ;
      RECT 14.4 73.78 23.56 73.85 ;
      RECT 14.4 73.85 23.535 73.875 ;
      RECT 14.4 70.14 57.405 70.16 ;
      RECT 14.4 70.16 57.39 70.175 ;
      RECT 14.42 70.12 57.425 70.14 ;
      RECT 14.49 70.05 57.445 70.12 ;
      RECT 14.56 69.98 57.515 70.05 ;
      RECT 14.63 69.91 57.585 69.98 ;
      RECT 14.7 69.84 57.655 69.91 ;
      RECT 14.77 69.77 57.725 69.84 ;
      RECT 14.84 69.7 57.795 69.77 ;
      RECT 14.91 69.63 57.865 69.7 ;
      RECT 14.98 69.56 57.935 69.63 ;
      RECT 15.05 69.49 58.005 69.56 ;
      RECT 15.12 69.42 58.075 69.49 ;
      RECT 15.19 69.35 58.145 69.42 ;
      RECT 15.26 69.28 58.215 69.35 ;
      RECT 15.33 69.21 58.285 69.28 ;
      RECT 15.4 69.14 58.355 69.21 ;
      RECT 15.47 69.07 58.425 69.14 ;
      RECT 15.54 69 58.495 69.07 ;
      RECT 15.61 68.93 58.565 69 ;
      RECT 15.68 68.86 58.635 68.93 ;
      RECT 15.75 68.79 58.705 68.86 ;
      RECT 15.82 68.72 58.775 68.79 ;
      RECT 15.89 68.65 58.845 68.72 ;
      RECT 15.96 68.58 58.915 68.65 ;
      RECT 16.03 68.51 58.985 68.58 ;
      RECT 16.1 68.44 59.055 68.51 ;
      RECT 16.17 68.37 59.125 68.44 ;
      RECT 16.24 68.3 59.195 68.37 ;
      RECT 16.31 68.23 59.265 68.3 ;
      RECT 16.38 68.16 59.335 68.23 ;
      RECT 16.45 68.09 59.405 68.16 ;
      RECT 16.52 68.02 59.475 68.09 ;
      RECT 16.59 67.95 59.545 68.02 ;
      RECT 16.66 67.88 59.615 67.95 ;
      RECT 16.73 67.81 59.685 67.88 ;
      RECT 16.8 67.74 59.755 67.81 ;
      RECT 16.87 67.67 59.825 67.74 ;
      RECT 16.94 67.6 59.895 67.67 ;
      RECT 17.01 67.53 59.965 67.6 ;
      RECT 17.08 67.46 60.035 67.53 ;
      RECT 17.15 67.39 60.105 67.46 ;
      RECT 17.22 67.32 60.175 67.39 ;
      RECT 17.29 67.25 60.245 67.32 ;
      RECT 17.36 67.18 60.315 67.25 ;
      RECT 17.43 67.11 60.385 67.18 ;
      RECT 17.5 67.04 60.455 67.11 ;
      RECT 17.57 66.97 60.525 67.04 ;
      RECT 17.64 66.9 60.595 66.97 ;
      RECT 17.71 66.83 60.665 66.9 ;
      RECT 17.78 66.76 60.735 66.83 ;
      RECT 56.99 59.81 60.785 59.855 ;
      RECT 56.99 59.74 60.715 59.81 ;
      RECT 56.99 59.67 60.645 59.74 ;
      RECT 56.99 59.6 60.575 59.67 ;
      RECT 56.99 59.53 60.505 59.6 ;
      RECT 56.99 59.46 60.435 59.53 ;
      RECT 56.99 59.39 60.365 59.46 ;
      RECT 56.99 59.32 60.295 59.39 ;
      RECT 56.99 59.25 60.225 59.32 ;
      RECT 56.99 59.18 60.155 59.25 ;
      RECT 56.99 59.11 60.085 59.18 ;
      RECT 56.99 59.04 60.015 59.11 ;
      RECT 56.99 58.97 59.945 59.04 ;
      RECT 56.99 58.9 59.875 58.97 ;
      RECT 56.99 58.83 59.805 58.9 ;
      RECT 56.99 58.76 59.735 58.83 ;
      RECT 56.99 58.69 59.665 58.76 ;
      RECT 56.99 58.62 59.595 58.69 ;
      RECT 56.99 58.55 59.525 58.62 ;
      RECT 56.99 58.48 59.455 58.55 ;
      RECT 56.99 58.41 59.385 58.48 ;
      RECT 56.99 58.34 59.315 58.41 ;
      RECT 56.99 58.27 59.245 58.34 ;
      RECT 56.99 58.2 59.175 58.27 ;
      RECT 56.99 58.13 59.105 58.2 ;
      RECT 56.99 58.06 59.035 58.13 ;
      RECT 56.99 57.99 58.965 58.06 ;
      RECT 56.99 57.92 58.895 57.99 ;
      RECT 15.085 92.455 58.1 92.525 ;
      RECT 15.155 92.385 58.17 92.455 ;
      RECT 15.225 92.315 58.24 92.385 ;
      RECT 15.295 92.245 58.31 92.315 ;
      RECT 15.365 92.175 58.38 92.245 ;
      RECT 15.435 92.105 58.45 92.175 ;
      RECT 15.505 92.035 58.52 92.105 ;
      RECT 15.575 91.965 58.59 92.035 ;
      RECT 15.645 91.895 58.66 91.965 ;
      RECT 15.715 91.825 58.73 91.895 ;
      RECT 15.785 91.755 58.8 91.825 ;
      RECT 15.855 91.685 58.87 91.755 ;
      RECT 15.925 91.615 58.94 91.685 ;
      RECT 15.995 91.545 59.01 91.615 ;
      RECT 16.065 91.475 59.08 91.545 ;
      RECT 16.135 91.405 59.15 91.475 ;
      RECT 16.205 91.335 59.22 91.405 ;
      RECT 16.275 91.265 59.29 91.335 ;
      RECT 16.345 91.195 59.36 91.265 ;
      RECT 16.415 91.125 59.43 91.195 ;
      RECT 16.485 91.055 59.5 91.125 ;
      RECT 16.555 90.985 59.57 91.055 ;
      RECT 16.625 90.915 59.64 90.985 ;
      RECT 16.695 90.845 59.71 90.915 ;
      RECT 16.765 90.775 59.78 90.845 ;
      RECT 16.835 90.705 59.85 90.775 ;
      RECT 16.905 90.635 59.92 90.705 ;
      RECT 16.975 90.565 59.99 90.635 ;
      RECT 17.045 90.495 60.06 90.565 ;
      RECT 17.115 90.425 60.13 90.495 ;
      RECT 17.185 90.355 60.2 90.425 ;
      RECT 17.255 90.285 60.27 90.355 ;
      RECT 17.325 90.215 60.34 90.285 ;
      RECT 17.395 90.145 60.41 90.215 ;
      RECT 17.465 90.075 60.48 90.145 ;
      RECT 17.535 90.005 60.55 90.075 ;
      RECT 17.605 89.935 60.62 90.005 ;
      RECT 17.675 89.865 60.69 89.935 ;
      RECT 17.745 89.795 60.76 89.865 ;
      RECT 17.78 89.76 60.83 89.775 ;
      RECT 17.765 89.775 60.83 89.79 ;
      RECT 17.75 89.79 60.83 89.795 ;
      RECT 56.985 82.81 60.815 82.825 ;
      RECT 56.985 82.74 60.745 82.81 ;
      RECT 56.985 82.67 60.675 82.74 ;
      RECT 56.985 82.6 60.605 82.67 ;
      RECT 56.985 82.53 60.535 82.6 ;
      RECT 56.985 82.46 60.465 82.53 ;
      RECT 56.985 82.39 60.395 82.46 ;
      RECT 56.985 82.32 60.325 82.39 ;
      RECT 56.985 82.25 60.255 82.32 ;
      RECT 56.985 82.18 60.185 82.25 ;
      RECT 56.985 82.11 60.115 82.18 ;
      RECT 56.985 82.04 60.045 82.11 ;
      RECT 56.985 81.97 59.975 82.04 ;
      RECT 56.985 81.9 59.905 81.97 ;
      RECT 56.985 81.83 59.835 81.9 ;
      RECT 56.985 81.76 59.765 81.83 ;
      RECT 56.985 81.69 59.695 81.76 ;
      RECT 56.985 81.62 59.625 81.69 ;
      RECT 56.985 81.55 59.555 81.62 ;
      RECT 56.985 81.48 59.485 81.55 ;
      RECT 56.985 81.41 59.415 81.48 ;
      RECT 56.985 81.34 59.345 81.41 ;
      RECT 56.985 81.27 59.275 81.34 ;
      RECT 56.985 81.2 59.205 81.27 ;
      RECT 56.985 81.13 59.135 81.2 ;
      RECT 56.985 81.06 59.065 81.13 ;
      RECT 56.985 80.99 58.995 81.06 ;
      RECT 56.985 80.92 58.925 80.99 ;
      RECT 56.985 80.85 58.855 80.92 ;
      RECT 56.985 80.78 58.785 80.85 ;
      RECT 56.985 80.71 58.715 80.78 ;
      RECT 56.985 80.64 58.645 80.71 ;
      RECT 56.985 80.57 58.575 80.64 ;
      RECT 56.985 80.5 58.505 80.57 ;
      RECT 56.985 79.435 57.44 79.505 ;
      RECT 56.985 79.505 57.51 79.575 ;
      RECT 56.985 79.575 57.58 79.645 ;
      RECT 56.985 79.645 57.65 79.715 ;
      RECT 56.985 79.715 57.72 79.785 ;
      RECT 56.985 79.785 57.79 79.855 ;
      RECT 56.985 79.855 57.86 79.925 ;
      RECT 56.985 79.925 57.93 79.995 ;
      RECT 56.985 79.995 58.0 80.065 ;
      RECT 56.985 80.065 58.07 80.135 ;
      RECT 56.985 80.135 58.14 80.205 ;
      RECT 56.985 80.205 58.21 80.275 ;
      RECT 56.985 80.275 58.28 80.345 ;
      RECT 56.985 80.345 58.35 80.415 ;
      RECT 56.985 80.415 58.42 80.485 ;
      RECT 56.985 80.485 58.49 80.5 ;
      RECT 16.78 79.435 24.54 79.505 ;
      RECT 16.85 79.505 24.54 79.575 ;
      RECT 16.92 79.575 24.54 79.645 ;
      RECT 16.99 79.645 24.54 79.715 ;
      RECT 17.06 79.715 24.54 79.785 ;
      RECT 17.13 79.785 24.54 79.855 ;
      RECT 17.2 79.855 24.54 79.925 ;
      RECT 17.27 79.925 24.54 79.995 ;
      RECT 17.34 79.995 24.54 80.065 ;
      RECT 17.41 80.065 24.54 80.135 ;
      RECT 17.48 80.135 24.54 80.205 ;
      RECT 17.55 80.205 24.54 80.275 ;
      RECT 17.62 80.275 24.54 80.345 ;
      RECT 17.69 80.345 24.54 80.415 ;
      RECT 17.76 80.415 24.54 80.485 ;
      RECT 17.775 80.485 24.54 80.5 ;
      RECT 14.47 77.125 24.54 77.195 ;
      RECT 14.54 77.195 24.54 77.265 ;
      RECT 14.61 77.265 24.54 77.335 ;
      RECT 14.68 77.335 24.54 77.405 ;
      RECT 14.75 77.405 24.54 77.475 ;
      RECT 14.82 77.475 24.54 77.545 ;
      RECT 14.89 77.545 24.54 77.615 ;
      RECT 14.96 77.615 24.54 77.685 ;
      RECT 15.03 77.685 24.54 77.755 ;
      RECT 15.1 77.755 24.54 77.825 ;
      RECT 15.17 77.825 24.54 77.895 ;
      RECT 15.24 77.895 24.54 77.965 ;
      RECT 15.31 77.965 24.54 78.035 ;
      RECT 15.38 78.035 24.54 78.105 ;
      RECT 15.45 78.105 24.54 78.175 ;
      RECT 15.52 78.175 24.54 78.245 ;
      RECT 15.59 78.245 24.54 78.315 ;
      RECT 15.66 78.315 24.54 78.385 ;
      RECT 15.44 115.14 58.325 115.21 ;
      RECT 15.37 115.21 58.255 115.28 ;
      RECT 15.3 115.28 58.185 115.35 ;
      RECT 15.23 115.35 58.115 115.42 ;
      RECT 15.16 115.42 58.045 115.49 ;
      RECT 15.09 115.49 57.975 115.56 ;
      RECT 15.02 115.56 57.905 115.63 ;
      RECT 14.95 115.63 57.835 115.7 ;
      RECT 14.88 115.7 57.765 115.77 ;
      RECT 14.81 115.77 57.695 115.84 ;
      RECT 14.74 115.84 57.625 115.91 ;
      RECT 14.67 115.91 57.555 115.98 ;
      RECT 14.6 115.98 57.485 116.05 ;
      RECT 14.53 116.05 57.415 116.12 ;
      RECT 14.46 116.12 57.36 116.175 ;
      RECT 56.985 105.81 60.815 105.825 ;
      RECT 56.985 105.74 60.745 105.81 ;
      RECT 56.985 105.67 60.675 105.74 ;
      RECT 56.985 105.6 60.605 105.67 ;
      RECT 56.985 105.53 60.535 105.6 ;
      RECT 56.985 105.46 60.465 105.53 ;
      RECT 56.985 105.39 60.395 105.46 ;
      RECT 56.985 105.32 60.325 105.39 ;
      RECT 56.985 105.25 60.255 105.32 ;
      RECT 56.985 105.18 60.185 105.25 ;
      RECT 56.985 105.11 60.115 105.18 ;
      RECT 56.985 105.04 60.045 105.11 ;
      RECT 56.985 104.97 59.975 105.04 ;
      RECT 56.985 104.9 59.905 104.97 ;
      RECT 56.985 104.83 59.835 104.9 ;
      RECT 56.985 104.76 59.765 104.83 ;
      RECT 56.985 104.69 59.695 104.76 ;
      RECT 56.985 104.62 59.625 104.69 ;
      RECT 56.985 104.55 59.555 104.62 ;
      RECT 56.985 104.48 59.485 104.55 ;
      RECT 56.985 104.41 59.415 104.48 ;
      RECT 56.985 104.34 59.345 104.41 ;
      RECT 56.985 104.27 59.275 104.34 ;
      RECT 56.985 104.2 59.205 104.27 ;
      RECT 56.985 104.13 59.135 104.2 ;
      RECT 56.985 104.06 59.065 104.13 ;
      RECT 56.985 103.99 58.995 104.06 ;
      RECT 56.985 103.92 58.925 103.99 ;
      RECT 56.985 103.85 58.855 103.92 ;
      RECT 56.985 103.78 58.785 103.85 ;
      RECT 56.985 103.71 58.715 103.78 ;
      RECT 56.985 103.64 58.645 103.71 ;
      RECT 56.985 103.57 58.575 103.64 ;
      RECT 56.985 103.5 58.505 103.57 ;
      RECT 56.985 102.435 57.44 102.505 ;
      RECT 56.985 102.505 57.51 102.575 ;
      RECT 56.985 102.575 57.58 102.645 ;
      RECT 56.985 102.645 57.65 102.715 ;
      RECT 56.985 102.715 57.72 102.785 ;
      RECT 56.985 102.785 57.79 102.855 ;
      RECT 56.985 102.855 57.86 102.925 ;
      RECT 56.985 102.925 57.93 102.995 ;
      RECT 56.985 102.995 58.0 103.065 ;
      RECT 56.985 103.065 58.07 103.135 ;
      RECT 56.985 103.135 58.14 103.205 ;
      RECT 56.985 103.205 58.21 103.275 ;
      RECT 56.985 103.275 58.28 103.345 ;
      RECT 56.985 103.345 58.35 103.415 ;
      RECT 56.985 103.415 58.42 103.485 ;
      RECT 56.985 103.485 58.49 103.5 ;
      RECT 16.78 102.435 24.54 102.505 ;
      RECT 16.85 102.505 24.54 102.575 ;
      RECT 16.92 102.575 24.54 102.645 ;
      RECT 16.99 102.645 24.54 102.715 ;
      RECT 17.06 102.715 24.54 102.785 ;
      RECT 17.13 102.785 24.54 102.855 ;
      RECT 17.2 102.855 24.54 102.925 ;
      RECT 17.27 102.925 24.54 102.995 ;
      RECT 17.34 102.995 24.54 103.065 ;
      RECT 17.41 103.065 24.54 103.135 ;
      RECT 17.48 103.135 24.54 103.205 ;
      RECT 17.55 103.205 24.54 103.275 ;
      RECT 17.62 103.275 24.54 103.345 ;
      RECT 17.69 103.345 24.54 103.415 ;
      RECT 17.76 103.415 24.54 103.485 ;
      RECT 17.775 103.485 24.54 103.5 ;
      RECT 14.47 100.125 24.54 100.195 ;
      RECT 14.54 100.195 24.54 100.265 ;
      RECT 14.61 100.265 24.54 100.335 ;
      RECT 14.68 100.335 24.54 100.405 ;
      RECT 14.75 100.405 24.54 100.475 ;
      RECT 14.82 100.475 24.54 100.545 ;
      RECT 14.89 100.545 24.54 100.615 ;
      RECT 14.96 100.615 24.54 100.685 ;
      RECT 15.03 100.685 24.54 100.755 ;
      RECT 15.1 100.755 24.54 100.825 ;
      RECT 15.17 100.825 24.54 100.895 ;
      RECT 15.24 100.895 24.54 100.965 ;
      RECT 15.31 100.965 24.54 101.035 ;
      RECT 15.38 101.035 24.54 101.105 ;
      RECT 15.45 101.105 24.54 101.175 ;
      RECT 15.52 101.175 24.54 101.245 ;
      RECT 15.59 101.245 24.54 101.315 ;
      RECT 15.66 101.315 24.54 101.385 ;
      RECT 15.73 101.385 24.54 101.455 ;
      RECT 15.8 101.455 24.54 101.525 ;
      RECT 15.87 101.525 24.54 101.595 ;
      RECT 15.94 101.595 24.54 101.665 ;
      RECT 16.01 101.665 24.54 101.735 ;
      RECT 16.08 101.735 24.54 101.805 ;
      RECT 16.15 101.805 24.54 101.875 ;
      RECT 16.22 101.875 24.54 101.945 ;
      RECT 16.29 101.945 24.54 102.015 ;
      RECT 16.36 102.015 24.54 102.085 ;
      RECT 16.43 102.085 24.54 102.155 ;
      RECT 16.5 102.155 24.54 102.225 ;
      RECT 16.57 102.225 24.54 102.295 ;
      RECT 16.64 102.295 24.54 102.365 ;
      RECT 16.71 102.365 24.54 102.435 ;
      RECT 14.4 93.14 57.465 93.16 ;
      RECT 14.4 93.16 57.45 93.175 ;
      RECT 14.455 93.085 57.485 93.14 ;
      RECT 14.525 93.015 57.54 93.085 ;
      RECT 14.595 92.945 57.61 93.015 ;
      RECT 14.665 92.875 57.68 92.945 ;
      RECT 14.735 92.805 57.75 92.875 ;
      RECT 14.805 92.735 57.82 92.805 ;
      RECT 14.875 92.665 57.89 92.735 ;
      RECT 14.945 92.595 57.96 92.665 ;
      RECT 15.015 92.525 58.03 92.595 ;
      RECT 56.985 128.11 60.115 128.18 ;
      RECT 56.985 128.04 60.045 128.11 ;
      RECT 56.985 127.97 59.975 128.04 ;
      RECT 56.985 127.9 59.905 127.97 ;
      RECT 56.985 127.83 59.835 127.9 ;
      RECT 56.985 127.76 59.765 127.83 ;
      RECT 56.985 127.69 59.695 127.76 ;
      RECT 56.985 127.62 59.625 127.69 ;
      RECT 56.985 127.55 59.555 127.62 ;
      RECT 56.985 127.48 59.485 127.55 ;
      RECT 56.985 127.41 59.415 127.48 ;
      RECT 56.985 127.34 59.345 127.41 ;
      RECT 56.985 127.27 59.275 127.34 ;
      RECT 56.985 127.2 59.205 127.27 ;
      RECT 56.985 127.13 59.135 127.2 ;
      RECT 56.985 127.06 59.065 127.13 ;
      RECT 56.985 126.99 58.995 127.06 ;
      RECT 56.985 126.92 58.925 126.99 ;
      RECT 56.985 126.85 58.855 126.92 ;
      RECT 56.985 126.78 58.785 126.85 ;
      RECT 56.985 126.71 58.715 126.78 ;
      RECT 56.985 126.64 58.645 126.71 ;
      RECT 56.985 126.57 58.575 126.64 ;
      RECT 56.985 126.5 58.505 126.57 ;
      RECT 56.985 125.435 57.44 125.505 ;
      RECT 56.985 125.505 57.51 125.575 ;
      RECT 56.985 125.575 57.58 125.645 ;
      RECT 56.985 125.645 57.65 125.715 ;
      RECT 56.985 125.715 57.72 125.785 ;
      RECT 56.985 125.785 57.79 125.855 ;
      RECT 56.985 125.855 57.86 125.925 ;
      RECT 56.985 125.925 57.93 125.995 ;
      RECT 56.985 125.995 58.0 126.065 ;
      RECT 56.985 126.065 58.07 126.135 ;
      RECT 56.985 126.135 58.14 126.205 ;
      RECT 56.985 126.205 58.21 126.275 ;
      RECT 56.985 126.275 58.28 126.345 ;
      RECT 56.985 126.345 58.35 126.415 ;
      RECT 56.985 126.415 58.42 126.485 ;
      RECT 56.985 126.485 58.49 126.5 ;
      RECT 16.875 125.435 24.54 125.505 ;
      RECT 16.945 125.505 24.54 125.575 ;
      RECT 17.015 125.575 24.54 125.645 ;
      RECT 17.085 125.645 24.54 125.715 ;
      RECT 17.155 125.715 24.54 125.785 ;
      RECT 17.225 125.785 24.54 125.855 ;
      RECT 17.295 125.855 24.54 125.925 ;
      RECT 17.365 125.925 24.54 125.995 ;
      RECT 17.435 125.995 24.54 126.065 ;
      RECT 17.505 126.065 24.54 126.135 ;
      RECT 17.575 126.135 24.54 126.205 ;
      RECT 17.645 126.205 24.54 126.275 ;
      RECT 17.715 126.275 24.54 126.345 ;
      RECT 17.785 126.345 24.54 126.415 ;
      RECT 17.855 126.415 24.54 126.485 ;
      RECT 17.87 126.485 24.54 126.5 ;
      RECT 14.47 123.03 24.54 123.1 ;
      RECT 14.54 123.1 24.54 123.17 ;
      RECT 14.61 123.17 24.54 123.24 ;
      RECT 14.68 123.24 24.54 123.31 ;
      RECT 14.75 123.31 24.54 123.38 ;
      RECT 14.82 123.38 24.54 123.45 ;
      RECT 14.89 123.45 24.54 123.52 ;
      RECT 14.96 123.52 24.54 123.59 ;
      RECT 15.03 123.59 24.54 123.66 ;
      RECT 15.1 123.66 24.54 123.73 ;
      RECT 15.17 123.73 24.54 123.8 ;
      RECT 15.24 123.8 24.54 123.87 ;
      RECT 15.31 123.87 24.54 123.94 ;
      RECT 15.38 123.94 24.54 124.01 ;
      RECT 15.45 124.01 24.54 124.08 ;
      RECT 15.52 124.08 24.54 124.15 ;
      RECT 15.59 124.15 24.54 124.22 ;
      RECT 15.66 124.22 24.54 124.29 ;
      RECT 15.73 124.29 24.54 124.36 ;
      RECT 15.8 124.36 24.54 124.43 ;
      RECT 15.87 124.43 24.54 124.5 ;
      RECT 15.94 124.5 24.54 124.57 ;
      RECT 16.01 124.57 24.54 124.64 ;
      RECT 16.08 124.64 24.54 124.71 ;
      RECT 16.15 124.71 24.54 124.78 ;
      RECT 16.22 124.78 24.54 124.85 ;
      RECT 16.29 124.85 24.54 124.92 ;
      RECT 16.36 124.92 24.54 124.99 ;
      RECT 16.43 124.99 24.54 125.06 ;
      RECT 16.5 125.06 24.54 125.13 ;
      RECT 16.57 125.13 24.54 125.2 ;
      RECT 16.64 125.2 24.54 125.27 ;
      RECT 16.71 125.27 24.54 125.34 ;
      RECT 16.78 125.34 24.54 125.41 ;
      RECT 16.805 125.41 24.54 125.435 ;
      RECT 14.405 116.175 24.54 116.18 ;
      RECT 17.82 112.76 60.705 112.83 ;
      RECT 17.75 112.83 60.635 112.9 ;
      RECT 17.68 112.9 60.565 112.97 ;
      RECT 17.61 112.97 60.495 113.04 ;
      RECT 17.54 113.04 60.425 113.11 ;
      RECT 17.47 113.11 60.355 113.18 ;
      RECT 17.4 113.18 60.285 113.25 ;
      RECT 17.33 113.25 60.215 113.32 ;
      RECT 17.26 113.32 60.145 113.39 ;
      RECT 17.19 113.39 60.075 113.46 ;
      RECT 17.12 113.46 60.005 113.53 ;
      RECT 17.05 113.53 59.935 113.6 ;
      RECT 16.98 113.6 59.865 113.67 ;
      RECT 16.91 113.67 59.795 113.74 ;
      RECT 16.84 113.74 59.725 113.81 ;
      RECT 16.77 113.81 59.655 113.88 ;
      RECT 16.7 113.88 59.585 113.95 ;
      RECT 16.63 113.95 59.515 114.02 ;
      RECT 16.56 114.02 59.445 114.09 ;
      RECT 16.49 114.09 59.375 114.16 ;
      RECT 16.42 114.16 59.305 114.23 ;
      RECT 16.35 114.23 59.235 114.3 ;
      RECT 16.28 114.3 59.165 114.37 ;
      RECT 16.21 114.37 59.095 114.44 ;
      RECT 16.14 114.44 59.025 114.51 ;
      RECT 16.07 114.51 58.955 114.58 ;
      RECT 16.0 114.58 58.885 114.65 ;
      RECT 15.93 114.65 58.815 114.72 ;
      RECT 15.86 114.72 58.745 114.79 ;
      RECT 15.79 114.79 58.675 114.86 ;
      RECT 15.72 114.86 58.605 114.93 ;
      RECT 15.65 114.93 58.535 115 ;
      RECT 15.58 115 58.465 115.07 ;
      RECT 15.51 115.07 58.395 115.14 ;
      RECT 15.455 161.14 58.375 161.21 ;
      RECT 15.385 161.21 58.305 161.28 ;
      RECT 15.315 161.28 58.235 161.35 ;
      RECT 15.245 161.35 58.165 161.42 ;
      RECT 15.175 161.42 58.095 161.49 ;
      RECT 15.105 161.49 58.025 161.56 ;
      RECT 15.035 161.56 57.955 161.63 ;
      RECT 14.965 161.63 57.885 161.7 ;
      RECT 14.895 161.7 57.815 161.77 ;
      RECT 14.825 161.77 57.745 161.84 ;
      RECT 14.755 161.84 57.675 161.91 ;
      RECT 14.685 161.91 57.605 161.98 ;
      RECT 14.615 161.98 57.535 162.05 ;
      RECT 14.545 162.05 57.465 162.12 ;
      RECT 14.475 162.12 57.41 162.175 ;
      RECT 56.985 151.88 60.815 151.895 ;
      RECT 56.985 151.81 60.745 151.88 ;
      RECT 56.985 151.74 60.675 151.81 ;
      RECT 56.985 151.67 60.605 151.74 ;
      RECT 56.985 151.6 60.535 151.67 ;
      RECT 56.985 151.53 60.465 151.6 ;
      RECT 56.985 151.46 60.395 151.53 ;
      RECT 56.985 151.39 60.325 151.46 ;
      RECT 56.985 151.32 60.255 151.39 ;
      RECT 56.985 151.25 60.185 151.32 ;
      RECT 56.985 151.18 60.115 151.25 ;
      RECT 56.985 151.11 60.045 151.18 ;
      RECT 56.985 151.04 59.975 151.11 ;
      RECT 56.985 150.97 59.905 151.04 ;
      RECT 56.985 150.9 59.835 150.97 ;
      RECT 56.985 150.83 59.765 150.9 ;
      RECT 56.985 150.76 59.695 150.83 ;
      RECT 56.985 150.69 59.625 150.76 ;
      RECT 56.985 150.62 59.555 150.69 ;
      RECT 56.985 150.55 59.485 150.62 ;
      RECT 56.985 150.48 59.415 150.55 ;
      RECT 56.985 150.41 59.345 150.48 ;
      RECT 56.985 150.34 59.275 150.41 ;
      RECT 56.985 150.27 59.205 150.34 ;
      RECT 56.985 150.2 59.135 150.27 ;
      RECT 56.985 150.13 59.065 150.2 ;
      RECT 56.985 150.06 58.995 150.13 ;
      RECT 56.985 149.99 58.925 150.06 ;
      RECT 56.985 149.92 58.855 149.99 ;
      RECT 56.985 149.85 58.785 149.92 ;
      RECT 56.985 149.78 58.715 149.85 ;
      RECT 56.985 149.71 58.645 149.78 ;
      RECT 56.985 149.64 58.575 149.71 ;
      RECT 56.985 149.57 58.505 149.64 ;
      RECT 56.985 149.5 58.435 149.57 ;
      RECT 56.985 148.435 57.37 148.505 ;
      RECT 56.985 148.505 57.44 148.575 ;
      RECT 56.985 148.575 57.51 148.645 ;
      RECT 56.985 148.645 57.58 148.715 ;
      RECT 56.985 148.715 57.65 148.785 ;
      RECT 56.985 148.785 57.72 148.855 ;
      RECT 56.985 148.855 57.79 148.925 ;
      RECT 56.985 148.925 57.86 148.995 ;
      RECT 56.985 148.995 57.93 149.065 ;
      RECT 56.985 149.065 58.0 149.135 ;
      RECT 56.985 149.135 58.07 149.205 ;
      RECT 56.985 149.205 58.14 149.275 ;
      RECT 56.985 149.275 58.21 149.345 ;
      RECT 56.985 149.345 58.28 149.415 ;
      RECT 56.985 149.415 58.35 149.485 ;
      RECT 56.985 149.485 58.42 149.5 ;
      RECT 17.925 135.76 60.74 135.83 ;
      RECT 17.855 135.83 60.67 135.9 ;
      RECT 17.785 135.9 60.6 135.97 ;
      RECT 17.715 135.97 60.53 136.04 ;
      RECT 17.645 136.04 60.46 136.11 ;
      RECT 17.575 136.11 60.39 136.18 ;
      RECT 17.505 136.18 60.32 136.25 ;
      RECT 17.435 136.25 60.25 136.32 ;
      RECT 17.365 136.32 60.18 136.39 ;
      RECT 17.295 136.39 60.11 136.46 ;
      RECT 17.225 136.46 60.04 136.53 ;
      RECT 17.155 136.53 59.97 136.6 ;
      RECT 17.085 136.6 59.9 136.67 ;
      RECT 17.015 136.67 59.83 136.74 ;
      RECT 16.945 136.74 59.76 136.81 ;
      RECT 16.875 136.81 59.69 136.88 ;
      RECT 16.805 136.88 59.62 136.95 ;
      RECT 16.735 136.95 59.55 137.02 ;
      RECT 16.665 137.02 59.48 137.09 ;
      RECT 16.595 137.09 59.41 137.16 ;
      RECT 16.525 137.16 59.34 137.23 ;
      RECT 16.455 137.23 59.27 137.3 ;
      RECT 16.385 137.3 59.2 137.37 ;
      RECT 16.315 137.37 59.13 137.44 ;
      RECT 16.245 137.44 59.06 137.51 ;
      RECT 16.175 137.51 58.99 137.58 ;
      RECT 16.105 137.58 58.92 137.65 ;
      RECT 16.035 137.65 58.85 137.72 ;
      RECT 15.965 137.72 58.78 137.79 ;
      RECT 15.895 137.79 58.71 137.86 ;
      RECT 15.825 137.86 58.64 137.93 ;
      RECT 15.755 137.93 58.57 138 ;
      RECT 15.685 138 58.5 138.07 ;
      RECT 15.615 138.07 58.43 138.14 ;
      RECT 15.545 138.14 58.36 138.21 ;
      RECT 15.475 138.21 58.29 138.28 ;
      RECT 15.405 138.28 58.22 138.35 ;
      RECT 15.335 138.35 58.15 138.42 ;
      RECT 15.265 138.42 58.08 138.49 ;
      RECT 15.195 138.49 58.01 138.56 ;
      RECT 15.125 138.56 57.94 138.63 ;
      RECT 15.055 138.63 57.87 138.7 ;
      RECT 14.985 138.7 57.8 138.77 ;
      RECT 14.915 138.77 57.73 138.84 ;
      RECT 14.845 138.84 57.66 138.91 ;
      RECT 14.775 138.91 57.59 138.98 ;
      RECT 14.705 138.98 57.52 139.05 ;
      RECT 14.635 139.05 57.45 139.12 ;
      RECT 14.565 139.12 57.395 139.175 ;
      RECT 56.985 128.81 60.815 128.825 ;
      RECT 56.985 128.74 60.745 128.81 ;
      RECT 56.985 128.67 60.675 128.74 ;
      RECT 56.985 128.6 60.605 128.67 ;
      RECT 56.985 128.53 60.535 128.6 ;
      RECT 56.985 128.46 60.465 128.53 ;
      RECT 56.985 128.39 60.395 128.46 ;
      RECT 56.985 128.32 60.325 128.39 ;
      RECT 56.985 128.25 60.255 128.32 ;
      RECT 56.985 128.18 60.185 128.25 ;
      RECT 15.905 55.535 17.835 55.605 ;
      RECT 15.975 55.605 17.905 55.675 ;
      RECT 16.045 55.675 17.975 55.745 ;
      RECT 16.115 55.745 18.045 55.815 ;
      RECT 16.185 55.815 18.115 55.885 ;
      RECT 16.255 55.885 18.185 55.955 ;
      RECT 16.325 55.955 18.255 56.025 ;
      RECT 16.395 56.025 18.325 56.095 ;
      RECT 16.465 56.095 18.395 56.165 ;
      RECT 16.535 56.165 18.465 56.235 ;
      RECT 16.605 56.235 18.535 56.305 ;
      RECT 16.675 56.305 18.605 56.375 ;
      RECT 16.735 56.375 18.675 56.435 ;
      RECT 16.78 79.435 57.44 79.505 ;
      RECT 16.85 79.505 57.51 79.575 ;
      RECT 16.92 79.575 57.58 79.645 ;
      RECT 16.99 79.645 57.65 79.715 ;
      RECT 17.06 79.715 57.72 79.785 ;
      RECT 17.13 79.785 57.79 79.855 ;
      RECT 17.2 79.855 57.86 79.925 ;
      RECT 17.27 79.925 57.93 79.995 ;
      RECT 17.34 79.995 58.0 80.065 ;
      RECT 17.41 80.065 58.07 80.135 ;
      RECT 17.48 80.135 58.14 80.205 ;
      RECT 17.55 80.205 58.21 80.275 ;
      RECT 17.62 80.275 58.28 80.345 ;
      RECT 17.69 80.345 58.35 80.415 ;
      RECT 17.76 80.415 58.42 80.485 ;
      RECT 17.775 80.485 58.49 80.5 ;
      RECT 16.78 102.435 57.44 102.505 ;
      RECT 16.85 102.505 57.51 102.575 ;
      RECT 16.92 102.575 57.58 102.645 ;
      RECT 16.99 102.645 57.65 102.715 ;
      RECT 17.06 102.715 57.72 102.785 ;
      RECT 17.13 102.785 57.79 102.855 ;
      RECT 17.2 102.855 57.86 102.925 ;
      RECT 17.27 102.925 57.93 102.995 ;
      RECT 17.34 102.995 58.0 103.065 ;
      RECT 17.41 103.065 58.07 103.135 ;
      RECT 17.48 103.135 58.14 103.205 ;
      RECT 17.55 103.205 58.21 103.275 ;
      RECT 17.62 103.275 58.28 103.345 ;
      RECT 17.69 103.345 58.35 103.415 ;
      RECT 17.76 103.415 58.42 103.485 ;
      RECT 17.775 103.485 58.49 103.5 ;
      RECT 16.805 56.435 57.41 56.505 ;
      RECT 16.875 56.505 57.48 56.575 ;
      RECT 16.945 56.575 57.55 56.645 ;
      RECT 17.015 56.645 57.62 56.715 ;
      RECT 17.085 56.715 57.69 56.785 ;
      RECT 17.155 56.785 57.76 56.855 ;
      RECT 17.225 56.855 57.83 56.925 ;
      RECT 17.295 56.925 57.9 56.995 ;
      RECT 17.365 56.995 57.97 57.065 ;
      RECT 17.435 57.065 58.04 57.135 ;
      RECT 17.505 57.135 58.11 57.205 ;
      RECT 17.575 57.205 58.18 57.275 ;
      RECT 17.645 57.275 58.25 57.345 ;
      RECT 17.715 57.345 58.32 57.415 ;
      RECT 17.785 57.415 58.39 57.485 ;
      RECT 17.8 57.485 58.46 57.5 ;
      RECT 16.805 148.435 57.37 148.505 ;
      RECT 16.875 148.505 57.44 148.575 ;
      RECT 16.945 148.575 57.51 148.645 ;
      RECT 17.015 148.645 57.58 148.715 ;
      RECT 17.085 148.715 57.65 148.785 ;
      RECT 17.155 148.785 57.72 148.855 ;
      RECT 17.225 148.855 57.79 148.925 ;
      RECT 17.295 148.925 57.86 148.995 ;
      RECT 17.365 148.995 57.93 149.065 ;
      RECT 17.435 149.065 58.0 149.135 ;
      RECT 17.505 149.135 58.07 149.205 ;
      RECT 17.575 149.205 58.14 149.275 ;
      RECT 17.645 149.275 58.21 149.345 ;
      RECT 17.715 149.345 58.28 149.415 ;
      RECT 17.785 149.415 58.35 149.485 ;
      RECT 17.8 149.485 58.42 149.5 ;
      RECT 16.875 125.435 57.44 125.505 ;
      RECT 16.945 125.505 57.51 125.575 ;
      RECT 17.015 125.575 57.58 125.645 ;
      RECT 17.085 125.645 57.65 125.715 ;
      RECT 17.155 125.715 57.72 125.785 ;
      RECT 17.225 125.785 57.79 125.855 ;
      RECT 17.295 125.855 57.86 125.925 ;
      RECT 17.365 125.925 57.93 125.995 ;
      RECT 17.435 125.995 58.0 126.065 ;
      RECT 17.505 126.065 58.07 126.135 ;
      RECT 17.575 126.135 58.14 126.205 ;
      RECT 17.645 126.205 58.21 126.275 ;
      RECT 17.715 126.275 58.28 126.345 ;
      RECT 17.785 126.345 58.35 126.415 ;
      RECT 17.855 126.415 58.42 126.485 ;
      RECT 17.87 126.485 58.49 126.5 ;
      RECT 17.835 158.76 60.755 158.83 ;
      RECT 17.765 158.83 60.685 158.9 ;
      RECT 17.695 158.9 60.615 158.97 ;
      RECT 17.625 158.97 60.545 159.04 ;
      RECT 17.555 159.04 60.475 159.11 ;
      RECT 17.485 159.11 60.405 159.18 ;
      RECT 17.415 159.18 60.335 159.25 ;
      RECT 17.345 159.25 60.265 159.32 ;
      RECT 17.275 159.32 60.195 159.39 ;
      RECT 17.205 159.39 60.125 159.46 ;
      RECT 17.135 159.46 60.055 159.53 ;
      RECT 17.065 159.53 59.985 159.6 ;
      RECT 16.995 159.6 59.915 159.67 ;
      RECT 16.925 159.67 59.845 159.74 ;
      RECT 16.855 159.74 59.775 159.81 ;
      RECT 16.785 159.81 59.705 159.88 ;
      RECT 16.715 159.88 59.635 159.95 ;
      RECT 16.645 159.95 59.565 160.02 ;
      RECT 16.575 160.02 59.495 160.09 ;
      RECT 16.505 160.09 59.425 160.16 ;
      RECT 16.435 160.16 59.355 160.23 ;
      RECT 16.365 160.23 59.285 160.3 ;
      RECT 16.295 160.3 59.215 160.37 ;
      RECT 16.225 160.37 59.145 160.44 ;
      RECT 16.155 160.44 59.075 160.51 ;
      RECT 16.085 160.51 59.005 160.58 ;
      RECT 16.015 160.58 58.935 160.65 ;
      RECT 15.945 160.65 58.865 160.72 ;
      RECT 15.875 160.72 58.795 160.79 ;
      RECT 15.805 160.79 58.725 160.86 ;
      RECT 15.735 160.86 58.655 160.93 ;
      RECT 15.665 160.93 58.585 161 ;
      RECT 15.595 161 58.515 161.07 ;
      RECT 15.525 161.07 58.445 161.14 ;
      RECT 16.87 171.505 57.52 171.575 ;
      RECT 16.94 171.575 57.59 171.645 ;
      RECT 17.01 171.645 57.66 171.715 ;
      RECT 17.08 171.715 57.73 171.785 ;
      RECT 17.15 171.785 57.8 171.855 ;
      RECT 17.22 171.855 57.87 171.925 ;
      RECT 17.29 171.925 57.94 171.995 ;
      RECT 17.36 171.995 58.01 172.065 ;
      RECT 17.43 172.065 58.08 172.135 ;
      RECT 17.5 172.135 58.15 172.205 ;
      RECT 17.57 172.205 58.22 172.275 ;
      RECT 17.64 172.275 58.29 172.345 ;
      RECT 17.71 172.345 58.36 172.415 ;
      RECT 17.78 172.415 58.43 172.485 ;
      RECT 17.795 172.485 58.5 172.5 ;
      RECT 14.4 47.175 16.525 54.1 ;
      RECT 14.4 162.195 16.525 169.105 ;
      RECT 14.4 139.285 16.525 146.1 ;
      RECT 24.675 0 25.615 2.2 ;
      RECT 37.175 12.12 37.61 25.94 ;
      RECT 56.985 151.895 60.83 158.755 ;
      RECT 56.985 128.825 60.83 135.74 ;
      RECT 14.4 116.18 24.54 123.03 ;
      RECT 56.985 105.825 60.83 112.705 ;
      RECT 14.4 93.175 24.54 100.125 ;
      RECT 14.4 75.73 24.54 77.125 ;
      RECT 14.4 73.875 18.13 74.695 ;
      RECT 14.4 70.175 24.54 72.87 ;
      RECT 56.99 59.855 60.83 66.735 ;
      RECT 57.195 35.835 60.83 39.78 ;
      RECT 15.485 31.07 60.83 35.55 ;
      RECT 56.985 82.825 60.83 89.76 ;
      RECT 24.675 2.2 50.11 8.48 ;
      RECT 28.175 0 50.11 8.48 ;
      RECT 28.175 0 50.11 2.2 ;
      RECT 14.51 139.175 16.525 139.23 ;
      RECT 14.455 139.23 16.525 139.285 ;
      RECT 14.47 169.105 16.525 169.175 ;
      RECT 14.54 169.175 16.525 169.245 ;
      RECT 14.61 169.245 16.525 169.315 ;
      RECT 14.68 169.315 16.525 169.385 ;
      RECT 14.75 169.385 16.525 169.455 ;
      RECT 14.82 169.455 16.525 169.525 ;
      RECT 14.89 169.525 16.525 169.595 ;
      RECT 14.96 169.595 16.525 169.665 ;
      RECT 15.03 169.665 16.525 169.735 ;
      RECT 15.1 169.735 16.525 169.805 ;
      RECT 15.17 169.805 16.525 169.875 ;
      RECT 15.24 169.875 16.525 169.945 ;
      RECT 15.31 169.945 16.525 170.015 ;
      RECT 15.38 170.015 16.525 170.085 ;
      RECT 15.45 170.085 16.525 170.155 ;
      RECT 15.52 170.155 16.525 170.225 ;
      RECT 15.59 170.225 16.525 170.295 ;
      RECT 15.66 170.295 16.525 170.365 ;
      RECT 15.73 170.365 16.525 170.435 ;
      RECT 15.8 170.435 16.525 170.505 ;
      RECT 15.87 170.505 16.525 170.575 ;
      RECT 15.94 170.575 16.525 170.645 ;
      RECT 16.01 170.645 16.525 170.715 ;
      RECT 16.08 170.715 16.525 170.785 ;
      RECT 16.15 170.785 16.525 170.855 ;
      RECT 16.22 170.855 16.525 170.925 ;
      RECT 16.29 170.925 16.525 170.995 ;
      RECT 16.36 170.995 16.525 171.065 ;
      RECT 16.43 171.065 16.525 171.135 ;
      RECT 16.5 171.135 16.525 171.205 ;
      RECT 14.42 162.175 16.525 162.185 ;
      RECT 14.41 162.185 16.525 162.195 ;
      RECT 14.47 146.1 16.525 146.17 ;
      RECT 14.54 146.17 16.525 146.24 ;
      RECT 14.61 146.24 16.525 146.31 ;
      RECT 14.68 146.31 16.525 146.38 ;
      RECT 14.75 146.38 16.525 146.45 ;
      RECT 14.82 146.45 16.525 146.52 ;
      RECT 14.89 146.52 16.525 146.59 ;
      RECT 14.96 146.59 16.525 146.66 ;
      RECT 15.03 146.66 16.525 146.73 ;
      RECT 15.1 146.73 16.525 146.8 ;
      RECT 15.125 146.8 16.525 146.825 ;
      RECT 14.47 54.1 16.525 54.17 ;
      RECT 14.54 54.17 16.525 54.24 ;
      RECT 14.61 54.24 16.525 54.31 ;
      RECT 14.68 54.31 16.525 54.38 ;
      RECT 14.75 54.38 16.525 54.45 ;
      RECT 14.82 54.45 16.525 54.52 ;
      RECT 14.89 54.52 16.525 54.59 ;
      RECT 14.96 54.59 16.525 54.66 ;
      RECT 15.03 54.66 16.525 54.73 ;
      RECT 15.1 54.73 16.525 54.8 ;
      RECT 15.17 54.8 16.525 54.87 ;
      RECT 15.24 54.87 16.525 54.94 ;
      RECT 15.31 54.94 16.525 55.01 ;
      RECT 15.345 55.01 16.525 55.045 ;
      RECT 15.195 146.825 16.525 146.895 ;
      RECT 15.265 146.895 16.595 146.965 ;
      RECT 15.335 146.965 16.665 147.035 ;
      RECT 15.405 147.035 16.735 147.105 ;
      RECT 15.475 147.105 16.805 147.175 ;
      RECT 15.545 147.175 16.875 147.245 ;
      RECT 15.615 147.245 16.945 147.315 ;
      RECT 15.685 147.315 17.015 147.385 ;
      RECT 15.755 147.385 17.085 147.455 ;
      RECT 15.825 147.455 17.155 147.525 ;
      RECT 15.895 147.525 17.225 147.595 ;
      RECT 15.965 147.595 17.295 147.665 ;
      RECT 16.035 147.665 17.365 147.735 ;
      RECT 16.105 147.735 17.435 147.805 ;
      RECT 16.175 147.805 17.505 147.875 ;
      RECT 16.245 147.875 17.575 147.945 ;
      RECT 16.315 147.945 17.645 148.015 ;
      RECT 16.385 148.015 17.715 148.085 ;
      RECT 16.455 148.085 17.785 148.155 ;
      RECT 16.525 148.155 17.855 148.225 ;
      RECT 16.595 148.225 17.925 148.295 ;
      RECT 16.665 148.295 17.995 148.365 ;
      RECT 16.735 148.365 18.065 148.435 ;
      RECT 15.415 55.045 17.345 55.115 ;
      RECT 15.485 55.115 17.415 55.185 ;
      RECT 15.555 55.185 17.485 55.255 ;
      RECT 15.625 55.255 17.555 55.325 ;
      RECT 15.695 55.325 17.625 55.395 ;
      RECT 15.765 55.395 17.695 55.465 ;
      RECT 15.835 55.465 17.765 55.535 ;
      RECT 0 195.355 67.48 200 ;
      RECT 0 2.61 0.655 195.355 ;
      RECT 0 0 0.215 2.17 ;
      RECT 74.57 0 75 190.295 ;
      RECT 67.48 190.295 75 200 ;
      RECT 70.48 193.295 72.0 197.0 ;
      RECT 0 2.17 0.215 2.24 ;
      RECT 0 2.24 0.285 2.31 ;
      RECT 0 2.31 0.355 2.38 ;
      RECT 0 2.38 0.425 2.45 ;
      RECT 0 2.45 0.495 2.52 ;
      RECT 0 2.52 0.565 2.59 ;
      RECT 0 2.59 0.635 2.61 ;
      RECT 14.4 185.17 15.34 189.47 ;
      RECT 58.24 174.815 60.83 181.76 ;
      RECT 14.47 189.47 15.34 189.54 ;
      RECT 14.54 189.54 15.34 189.61 ;
      RECT 14.61 189.61 15.34 189.68 ;
      RECT 14.68 189.68 15.34 189.75 ;
      RECT 14.75 189.75 15.34 189.82 ;
      RECT 14.82 189.82 15.34 189.89 ;
      RECT 14.89 189.89 15.34 189.96 ;
      RECT 14.96 189.96 15.34 190.03 ;
      RECT 15.03 190.03 15.34 190.1 ;
      RECT 15.1 190.1 15.34 190.17 ;
      RECT 15.17 190.17 15.34 190.24 ;
      RECT 15.21 190.24 15.34 190.28 ;
      RECT 14.555 185.015 15.34 185.085 ;
      RECT 14.485 185.085 15.34 185.155 ;
      RECT 14.415 185.155 15.34 185.17 ;
      RECT 15.385 184.185 59.34 184.255 ;
      RECT 15.315 184.255 59.27 184.325 ;
      RECT 15.245 184.325 59.2 184.395 ;
      RECT 15.175 184.395 59.13 184.465 ;
      RECT 15.105 184.465 59.06 184.535 ;
      RECT 15.035 184.535 58.99 184.605 ;
      RECT 14.965 184.605 58.92 184.675 ;
      RECT 14.895 184.675 58.85 184.745 ;
      RECT 14.825 184.745 58.78 184.815 ;
      RECT 14.755 184.815 58.71 184.885 ;
      RECT 14.685 184.885 58.64 184.955 ;
      RECT 14.615 184.955 58.58 185.015 ;
      RECT 15.6 183.97 59.555 184.04 ;
      RECT 15.6 184.04 59.485 184.11 ;
      RECT 15.6 184.11 59.415 184.18 ;
      RECT 15.6 184.18 59.41 184.185 ;
      RECT 16.805 182.765 60.76 182.835 ;
      RECT 16.735 182.835 60.69 182.905 ;
      RECT 16.665 182.905 60.62 182.975 ;
      RECT 16.595 182.975 60.55 183.045 ;
      RECT 16.525 183.045 60.48 183.115 ;
      RECT 16.455 183.115 60.41 183.185 ;
      RECT 16.385 183.185 60.34 183.255 ;
      RECT 16.315 183.255 60.27 183.325 ;
      RECT 16.245 183.325 60.2 183.395 ;
      RECT 16.175 183.395 60.13 183.465 ;
      RECT 16.105 183.465 60.06 183.535 ;
      RECT 16.035 183.535 59.99 183.605 ;
      RECT 15.965 183.605 59.92 183.675 ;
      RECT 15.895 183.675 59.85 183.745 ;
      RECT 15.825 183.745 59.78 183.815 ;
      RECT 15.755 183.815 59.71 183.885 ;
      RECT 15.685 183.885 59.64 183.955 ;
      RECT 15.615 183.955 59.625 183.97 ;
      RECT 17.81 181.76 60.83 181.83 ;
      RECT 17.74 181.83 60.83 181.9 ;
      RECT 17.67 181.9 60.83 181.97 ;
      RECT 17.6 181.97 60.83 182.04 ;
      RECT 17.53 182.04 60.83 182.11 ;
      RECT 17.46 182.11 60.83 182.18 ;
      RECT 17.39 182.18 60.83 182.25 ;
      RECT 17.32 182.25 60.83 182.32 ;
      RECT 17.25 182.32 60.83 182.39 ;
      RECT 17.18 182.39 60.83 182.46 ;
      RECT 17.11 182.46 60.83 182.53 ;
      RECT 17.04 182.53 60.83 182.6 ;
      RECT 16.97 182.6 60.83 182.67 ;
      RECT 16.9 182.67 60.83 182.74 ;
      RECT 16.83 182.74 60.83 182.765 ;
      RECT 58.24 174.81 60.825 174.815 ;
      RECT 58.24 174.74 60.755 174.81 ;
      RECT 58.24 174.67 60.685 174.74 ;
      RECT 58.24 174.6 60.615 174.67 ;
      RECT 58.24 174.53 60.545 174.6 ;
      RECT 58.24 174.46 60.475 174.53 ;
      RECT 58.24 174.39 60.405 174.46 ;
      RECT 58.24 174.32 60.335 174.39 ;
      RECT 58.24 174.25 60.265 174.32 ;
      RECT 58.24 174.18 60.195 174.25 ;
      RECT 58.24 174.11 60.125 174.18 ;
      RECT 58.24 174.04 60.055 174.11 ;
      RECT 58.24 173.97 59.985 174.04 ;
      RECT 58.24 173.9 59.915 173.97 ;
      RECT 58.24 173.83 59.845 173.9 ;
      RECT 58.24 173.76 59.775 173.83 ;
      RECT 58.24 173.69 59.705 173.76 ;
      RECT 58.24 173.62 59.635 173.69 ;
      RECT 58.24 173.55 59.565 173.62 ;
      RECT 58.24 173.48 59.495 173.55 ;
      RECT 58.24 173.41 59.425 173.48 ;
      RECT 58.24 173.34 59.355 173.41 ;
      RECT 58.24 173.27 59.285 173.34 ;
      RECT 58.24 173.2 59.215 173.27 ;
      RECT 58.24 173.13 59.145 173.2 ;
      RECT 58.24 173.06 59.075 173.13 ;
      RECT 58.24 172.99 59.005 173.06 ;
      RECT 58.24 172.92 58.935 172.99 ;
      RECT 58.24 172.85 58.865 172.92 ;
      RECT 58.24 172.78 58.795 172.85 ;
      RECT 58.24 172.71 58.725 172.78 ;
      RECT 58.24 172.64 58.655 172.71 ;
      RECT 58.24 172.57 58.585 172.64 ;
      RECT 58.24 172.5 58.515 172.57 ;
      RECT 16.8 171.435 57.45 171.505 ;
    LAYER li1 ;
      RECT 61.78 195.37 62.49 195.54 ;
      RECT 62.865 162.525 63.395 180.695 ;
      RECT 62.885 180.695 63.395 182.035 ;
      RECT 62.885 162.325 63.395 162.525 ;
      RECT 60.245 185.16 61.435 195.01 ;
      RECT 60.385 195.01 61.275 195.14 ;
      RECT 60.245 162.16 61.435 181.87 ;
      RECT 72.245 199.21 72.775 199.38 ;
      RECT 72.345 199.38 72.675 199.42 ;
      RECT 59.575 3.075 67.575 3.305 ;
      RECT 49.815 3.075 57.815 3.305 ;
      RECT 40.055 3.075 48.055 3.305 ;
      RECT 30.295 3.075 38.295 3.305 ;
      RECT 20.535 3.075 28.535 3.305 ;
      RECT 59.575 9.295 67.575 9.525 ;
      RECT 49.815 9.295 57.815 9.525 ;
      RECT 40.055 9.295 48.055 9.525 ;
      RECT 30.295 9.295 38.295 9.525 ;
      RECT 20.535 9.295 28.535 9.525 ;
      RECT 59.575 15.515 67.575 15.745 ;
      RECT 49.815 15.515 57.815 15.745 ;
      RECT 40.055 15.515 48.055 15.745 ;
      RECT 30.295 15.515 38.295 15.745 ;
      RECT 20.535 15.515 28.535 15.745 ;
      RECT 54.94 39.77 66.335 39.94 ;
      RECT 6.34 36.97 45.06 37.23 ;
      RECT 53.685 139.325 54.195 139.525 ;
      RECT 53.665 116.525 54.195 134.695 ;
      RECT 53.685 134.695 54.195 136.035 ;
      RECT 53.685 116.325 54.195 116.525 ;
      RECT 58.265 116.525 58.795 134.695 ;
      RECT 58.285 134.695 58.795 136.035 ;
      RECT 58.285 116.325 58.795 116.525 ;
      RECT 55.645 116.16 56.835 135.87 ;
      RECT 55.645 139.16 56.835 158.87 ;
      RECT 64.845 116.16 65.875 135.93 ;
      RECT 64.845 139.16 65.875 158.93 ;
      RECT 62.865 139.525 63.395 157.695 ;
      RECT 62.885 157.695 63.395 159.035 ;
      RECT 62.885 139.325 63.395 139.525 ;
      RECT 62.865 116.525 63.395 134.695 ;
      RECT 62.885 134.695 63.395 136.035 ;
      RECT 62.885 116.325 63.395 116.525 ;
      RECT 60.245 116.16 61.435 135.87 ;
      RECT 60.245 139.16 61.435 158.87 ;
      RECT 14.385 162.16 15.435 181.93 ;
      RECT 14.385 185.16 15.435 195.185 ;
      RECT 16.865 185.525 17.395 195.055 ;
      RECT 16.885 185.325 17.395 185.525 ;
      RECT 17.79 195.37 18.5 195.54 ;
      RECT 15.78 195.37 16.49 195.54 ;
      RECT 16.865 162.525 17.395 180.695 ;
      RECT 16.885 180.695 17.395 182.035 ;
      RECT 16.885 162.325 17.395 162.525 ;
      RECT 18.845 185.16 20.035 195.01 ;
      RECT 18.985 195.01 19.875 195.075 ;
      RECT 18.845 162.16 20.035 181.87 ;
      RECT 15.78 159.34 64.5 159.555 ;
      RECT 12.4 159.555 64.5 161.99 ;
      RECT 15.78 182.34 66.685 182.57 ;
      RECT 12.83 182.57 66.685 184.99 ;
      RECT 21.465 185.525 21.995 195.055 ;
      RECT 21.485 185.325 21.995 185.525 ;
      RECT 22.39 195.37 23.1 195.54 ;
      RECT 24.98 195.37 25.69 195.54 ;
      RECT 20.38 195.37 21.09 195.54 ;
      RECT 21.465 162.525 21.995 180.695 ;
      RECT 21.485 180.695 21.995 182.035 ;
      RECT 21.485 162.325 21.995 162.525 ;
      RECT 23.445 185.16 24.635 195.01 ;
      RECT 23.585 195.01 24.475 195.03 ;
      RECT 23.445 162.16 24.635 181.87 ;
      RECT 26.065 185.525 26.595 195.055 ;
      RECT 26.085 185.325 26.595 185.525 ;
      RECT 30.665 185.525 31.195 195.055 ;
      RECT 30.685 185.325 31.195 185.525 ;
      RECT 26.99 195.37 27.7 195.54 ;
      RECT 31.59 195.37 32.3 195.54 ;
      RECT 29.58 195.37 30.29 195.54 ;
      RECT 30.665 162.525 31.195 180.695 ;
      RECT 30.685 180.695 31.195 182.035 ;
      RECT 30.685 162.325 31.195 162.525 ;
      RECT 26.065 162.525 26.595 180.695 ;
      RECT 26.085 180.695 26.595 182.035 ;
      RECT 26.085 162.325 26.595 162.525 ;
      RECT 28.045 185.16 29.235 195.01 ;
      RECT 28.185 195.01 29.075 195.03 ;
      RECT 28.045 162.16 29.235 181.87 ;
      RECT 35.265 185.525 35.795 195.055 ;
      RECT 35.285 185.325 35.795 185.525 ;
      RECT 36.19 195.37 36.9 195.54 ;
      RECT 38.78 195.37 39.49 195.54 ;
      RECT 34.18 195.37 34.89 195.54 ;
      RECT 35.265 162.525 35.795 180.695 ;
      RECT 35.285 180.695 35.795 182.035 ;
      RECT 35.285 162.325 35.795 162.525 ;
      RECT 37.245 185.16 38.435 195.01 ;
      RECT 37.385 195.01 38.275 195.03 ;
      RECT 32.645 185.16 33.835 195.01 ;
      RECT 32.785 195.01 33.675 195.03 ;
      RECT 37.245 162.16 38.435 181.87 ;
      RECT 32.645 162.16 33.835 181.87 ;
      RECT 39.865 185.525 40.395 195.055 ;
      RECT 39.885 185.325 40.395 185.525 ;
      RECT 44.465 185.525 44.995 195.055 ;
      RECT 44.485 185.325 44.995 185.525 ;
      RECT 40.79 195.37 41.5 195.54 ;
      RECT 45.39 195.37 46.1 195.54 ;
      RECT 43.38 195.37 44.09 195.54 ;
      RECT 44.465 162.525 44.995 180.695 ;
      RECT 44.485 180.695 44.995 182.035 ;
      RECT 44.485 162.325 44.995 162.525 ;
      RECT 39.865 162.525 40.395 180.695 ;
      RECT 39.885 180.695 40.395 182.035 ;
      RECT 39.885 162.325 40.395 162.525 ;
      RECT 41.845 185.16 43.035 195.01 ;
      RECT 41.985 195.01 42.875 195.03 ;
      RECT 41.845 162.16 43.035 181.87 ;
      RECT 49.065 185.525 49.595 195.055 ;
      RECT 49.085 185.325 49.595 185.525 ;
      RECT 49.99 195.37 50.7 195.54 ;
      RECT 47.98 195.37 48.69 195.54 ;
      RECT 49.065 162.525 49.595 180.695 ;
      RECT 49.085 180.695 49.595 182.035 ;
      RECT 49.085 162.325 49.595 162.525 ;
      RECT 51.045 185.16 52.235 195.01 ;
      RECT 51.185 195.01 52.075 195.03 ;
      RECT 46.445 185.16 47.635 195.01 ;
      RECT 46.585 195.01 47.475 195.03 ;
      RECT 51.045 162.16 52.235 181.87 ;
      RECT 46.445 162.16 47.635 181.87 ;
      RECT 52.58 195.37 53.29 195.54 ;
      RECT 53.665 185.525 54.195 195.055 ;
      RECT 53.685 185.325 54.195 185.525 ;
      RECT 58.265 185.525 58.795 195.055 ;
      RECT 58.285 185.325 58.795 185.525 ;
      RECT 54.59 195.37 55.3 195.54 ;
      RECT 59.19 195.37 59.9 195.54 ;
      RECT 57.18 195.37 57.89 195.54 ;
      RECT 58.265 162.525 58.795 180.695 ;
      RECT 58.285 180.695 58.795 182.035 ;
      RECT 58.285 162.325 58.795 162.525 ;
      RECT 53.665 162.525 54.195 180.695 ;
      RECT 53.685 180.695 54.195 182.035 ;
      RECT 53.685 162.325 54.195 162.525 ;
      RECT 55.645 185.16 56.835 195.01 ;
      RECT 55.785 195.01 56.675 195.14 ;
      RECT 55.645 162.16 56.835 181.87 ;
      RECT 64.845 162.16 65.875 181.93 ;
      RECT 64.845 185.16 65.875 195.18 ;
      RECT 62.865 185.525 63.395 195.055 ;
      RECT 62.885 185.325 63.395 185.525 ;
      RECT 63.79 195.37 64.5 195.54 ;
      RECT 60.93 39.29 61.1 39.35 ;
      RECT 60.93 32.56 61.1 36.19 ;
      RECT 60.145 32.62 60.32 35.77 ;
      RECT 60.15 35.77 60.32 39.35 ;
      RECT 60.15 32.56 60.32 32.62 ;
      RECT 59.37 36.19 59.545 39.29 ;
      RECT 59.37 39.29 59.54 39.35 ;
      RECT 59.37 32.56 59.54 36.19 ;
      RECT 60.245 47.16 61.435 66.87 ;
      RECT 66.385 32.62 66.56 35.77 ;
      RECT 66.39 35.77 66.56 39.35 ;
      RECT 66.39 32.56 66.56 32.62 ;
      RECT 70.725 42.99 71.055 43.015 ;
      RECT 70.725 42.735 71.055 42.82 ;
      RECT 70.47 42.82 71.055 42.99 ;
      RECT 9.405 74.18 9.935 74.35 ;
      RECT 9.5 74.35 9.83 74.355 ;
      RECT 18.41 74.2 19 74.37 ;
      RECT 18.41 74.37 18.74 74.385 ;
      RECT 18.41 74.185 18.74 74.2 ;
      RECT 23.585 93.16 24.635 112.93 ;
      RECT 23.055 113.34 64.5 115.99 ;
      RECT 23.025 90.495 64.5 92.99 ;
      RECT 24.98 90.37 64.5 90.495 ;
      RECT 25.67 90.34 64.5 90.37 ;
      RECT 26.065 93.525 26.595 111.695 ;
      RECT 26.085 111.695 26.595 113.035 ;
      RECT 26.085 93.325 26.595 93.525 ;
      RECT 30.665 93.525 31.195 111.695 ;
      RECT 30.685 111.695 31.195 113.035 ;
      RECT 30.685 93.325 31.195 93.525 ;
      RECT 28.045 93.16 29.235 112.87 ;
      RECT 35.265 93.525 35.795 111.695 ;
      RECT 35.285 111.695 35.795 113.035 ;
      RECT 35.285 93.325 35.795 93.525 ;
      RECT 37.245 93.16 38.435 112.87 ;
      RECT 32.645 93.16 33.835 112.87 ;
      RECT 39.865 93.525 40.395 111.695 ;
      RECT 39.885 111.695 40.395 113.035 ;
      RECT 39.885 93.325 40.395 93.525 ;
      RECT 44.465 93.525 44.995 111.695 ;
      RECT 44.485 111.695 44.995 113.035 ;
      RECT 44.485 93.325 44.995 93.525 ;
      RECT 41.845 93.16 43.035 112.87 ;
      RECT 49.065 93.525 49.595 111.695 ;
      RECT 49.085 111.695 49.595 113.035 ;
      RECT 49.085 93.325 49.595 93.525 ;
      RECT 51.045 93.16 52.235 112.87 ;
      RECT 46.445 93.16 47.635 112.87 ;
      RECT 53.665 93.525 54.195 111.695 ;
      RECT 53.685 111.695 54.195 113.035 ;
      RECT 53.685 93.325 54.195 93.525 ;
      RECT 58.265 93.525 58.795 111.695 ;
      RECT 58.285 111.695 58.795 113.035 ;
      RECT 58.285 93.325 58.795 93.525 ;
      RECT 55.645 93.16 56.835 112.87 ;
      RECT 64.845 93.16 65.875 112.935 ;
      RECT 62.865 93.525 63.395 111.695 ;
      RECT 62.885 111.695 63.395 113.035 ;
      RECT 62.885 93.325 63.395 93.525 ;
      RECT 60.245 93.16 61.435 112.87 ;
      RECT 14.385 139.16 15.435 158.93 ;
      RECT 16.865 139.525 17.395 157.695 ;
      RECT 16.885 157.695 17.395 159.035 ;
      RECT 16.885 139.325 17.395 139.525 ;
      RECT 18.845 139.16 20.035 158.87 ;
      RECT 15.78 136.54 64.5 138.99 ;
      RECT 25.67 136.34 64.5 136.37 ;
      RECT 24.98 136.37 64.5 136.54 ;
      RECT 23.585 116.16 24.635 135.93 ;
      RECT 21.465 139.525 21.995 157.695 ;
      RECT 21.485 157.695 21.995 159.035 ;
      RECT 21.485 139.325 21.995 139.525 ;
      RECT 23.445 139.16 24.635 158.87 ;
      RECT 30.665 139.525 31.195 157.695 ;
      RECT 30.685 157.695 31.195 159.035 ;
      RECT 30.685 139.325 31.195 139.525 ;
      RECT 26.065 139.525 26.595 157.695 ;
      RECT 26.085 157.695 26.595 159.035 ;
      RECT 26.085 139.325 26.595 139.525 ;
      RECT 26.065 116.525 26.595 134.695 ;
      RECT 26.085 134.695 26.595 136.035 ;
      RECT 26.085 116.325 26.595 116.525 ;
      RECT 30.665 116.525 31.195 134.695 ;
      RECT 30.685 134.695 31.195 136.035 ;
      RECT 30.685 116.325 31.195 116.525 ;
      RECT 28.045 116.16 29.235 135.87 ;
      RECT 28.045 139.16 29.235 158.87 ;
      RECT 35.265 139.525 35.795 157.695 ;
      RECT 35.285 157.695 35.795 159.035 ;
      RECT 35.285 139.325 35.795 139.525 ;
      RECT 35.265 116.525 35.795 134.695 ;
      RECT 35.285 134.695 35.795 136.035 ;
      RECT 35.285 116.325 35.795 116.525 ;
      RECT 37.245 116.16 38.435 135.87 ;
      RECT 32.645 116.16 33.835 135.87 ;
      RECT 37.245 139.16 38.435 158.87 ;
      RECT 32.645 139.16 33.835 158.87 ;
      RECT 44.465 139.525 44.995 157.695 ;
      RECT 44.485 157.695 44.995 159.035 ;
      RECT 44.485 139.325 44.995 139.525 ;
      RECT 39.865 139.525 40.395 157.695 ;
      RECT 39.885 157.695 40.395 159.035 ;
      RECT 39.885 139.325 40.395 139.525 ;
      RECT 39.865 116.525 40.395 134.695 ;
      RECT 39.885 134.695 40.395 136.035 ;
      RECT 39.885 116.325 40.395 116.525 ;
      RECT 44.465 116.525 44.995 134.695 ;
      RECT 44.485 134.695 44.995 136.035 ;
      RECT 44.485 116.325 44.995 116.525 ;
      RECT 41.845 116.16 43.035 135.87 ;
      RECT 41.845 139.16 43.035 158.87 ;
      RECT 49.065 139.525 49.595 157.695 ;
      RECT 49.085 157.695 49.595 159.035 ;
      RECT 49.085 139.325 49.595 139.525 ;
      RECT 49.065 116.525 49.595 134.695 ;
      RECT 49.085 134.695 49.595 136.035 ;
      RECT 49.085 116.325 49.595 116.525 ;
      RECT 51.045 116.16 52.235 135.87 ;
      RECT 46.445 116.16 47.635 135.87 ;
      RECT 51.045 139.16 52.235 158.87 ;
      RECT 46.445 139.16 47.635 158.87 ;
      RECT 58.265 139.525 58.795 157.695 ;
      RECT 58.285 157.695 58.795 159.035 ;
      RECT 58.285 139.325 58.795 139.525 ;
      RECT 53.665 139.525 54.195 157.695 ;
      RECT 53.685 157.695 54.195 159.035 ;
      RECT 27.175 29.77 27.345 36.57 ;
      RECT 26.395 29.78 26.565 36.57 ;
      RECT 31.855 29.775 32.025 36.57 ;
      RECT 31.075 29.78 31.245 36.57 ;
      RECT 30.295 29.77 30.465 36.57 ;
      RECT 29.515 29.78 29.685 36.57 ;
      RECT 28.735 29.775 28.905 36.57 ;
      RECT 27.955 29.78 28.125 36.57 ;
      RECT 28.045 70.16 29.235 89.87 ;
      RECT 28.045 47.16 29.235 66.87 ;
      RECT 35.265 47.525 35.795 65.695 ;
      RECT 35.285 65.695 35.795 67.035 ;
      RECT 35.285 47.325 35.795 47.525 ;
      RECT 35.265 70.525 35.795 88.695 ;
      RECT 35.285 88.695 35.795 90.035 ;
      RECT 35.285 70.325 35.795 70.525 ;
      RECT 38.875 29.78 39.045 36.57 ;
      RECT 38.095 29.775 38.265 36.57 ;
      RECT 37.315 29.78 37.485 36.57 ;
      RECT 36.535 29.77 36.705 36.57 ;
      RECT 35.755 29.78 35.925 36.57 ;
      RECT 34.975 29.775 35.145 36.57 ;
      RECT 34.195 29.78 34.365 36.57 ;
      RECT 33.415 29.77 33.585 36.57 ;
      RECT 32.635 29.78 32.805 36.57 ;
      RECT 37.245 70.16 38.435 89.87 ;
      RECT 32.645 70.16 33.835 89.87 ;
      RECT 37.245 47.16 38.435 66.87 ;
      RECT 32.645 47.16 33.835 66.87 ;
      RECT 45.115 29.78 45.285 36.57 ;
      RECT 39.865 47.525 40.395 65.695 ;
      RECT 39.885 65.695 40.395 67.035 ;
      RECT 39.885 47.325 40.395 47.525 ;
      RECT 44.465 47.525 44.995 65.695 ;
      RECT 44.485 65.695 44.995 67.035 ;
      RECT 44.485 47.325 44.995 47.525 ;
      RECT 44.465 70.525 44.995 88.695 ;
      RECT 44.485 88.695 44.995 90.035 ;
      RECT 44.485 70.325 44.995 70.525 ;
      RECT 39.865 70.525 40.395 88.695 ;
      RECT 39.885 88.695 40.395 90.035 ;
      RECT 39.885 70.325 40.395 70.525 ;
      RECT 44.335 29.77 44.505 36.57 ;
      RECT 43.555 29.78 43.725 36.57 ;
      RECT 42.775 29.775 42.945 36.57 ;
      RECT 41.995 29.78 42.165 36.57 ;
      RECT 41.215 29.77 41.385 36.57 ;
      RECT 40.435 29.78 40.605 36.57 ;
      RECT 39.655 29.77 39.825 36.57 ;
      RECT 41.845 70.16 43.035 89.87 ;
      RECT 41.845 47.16 43.035 66.87 ;
      RECT 49.065 47.525 49.595 65.695 ;
      RECT 49.085 65.695 49.595 67.035 ;
      RECT 49.085 47.325 49.595 47.525 ;
      RECT 49.065 70.525 49.595 88.695 ;
      RECT 49.085 88.695 49.595 90.035 ;
      RECT 49.085 70.325 49.595 70.525 ;
      RECT 51.045 70.16 52.235 89.87 ;
      RECT 46.445 70.16 47.635 89.87 ;
      RECT 51.045 47.16 52.235 66.87 ;
      RECT 46.445 47.16 47.635 66.87 ;
      RECT 54.69 36.19 54.865 39.29 ;
      RECT 54.69 39.29 54.86 39.35 ;
      RECT 54.69 32.56 54.86 36.19 ;
      RECT 53.665 47.525 54.195 65.695 ;
      RECT 53.685 65.695 54.195 67.035 ;
      RECT 53.685 47.325 54.195 47.525 ;
      RECT 58.265 47.525 58.795 65.695 ;
      RECT 58.285 65.695 58.795 67.035 ;
      RECT 58.285 47.325 58.795 47.525 ;
      RECT 58.265 70.525 58.795 88.695 ;
      RECT 58.285 88.695 58.795 90.035 ;
      RECT 58.285 70.325 58.795 70.525 ;
      RECT 53.665 70.525 54.195 88.695 ;
      RECT 53.685 88.695 54.195 90.035 ;
      RECT 53.685 70.325 54.195 70.525 ;
      RECT 55.645 70.16 56.835 89.87 ;
      RECT 58.585 32.62 58.76 35.77 ;
      RECT 58.59 35.77 58.76 39.35 ;
      RECT 58.59 32.56 58.76 32.62 ;
      RECT 57.81 36.19 57.985 39.29 ;
      RECT 57.81 39.29 57.98 39.35 ;
      RECT 57.81 32.56 57.98 36.19 ;
      RECT 57.025 32.62 57.2 35.77 ;
      RECT 57.03 35.77 57.2 39.35 ;
      RECT 57.03 32.56 57.2 32.62 ;
      RECT 56.25 36.19 56.425 39.29 ;
      RECT 56.25 39.29 56.42 39.35 ;
      RECT 56.25 32.56 56.42 36.19 ;
      RECT 55.465 32.62 55.64 35.77 ;
      RECT 55.47 35.77 55.64 39.35 ;
      RECT 55.47 32.56 55.64 32.62 ;
      RECT 55.645 47.16 56.835 66.87 ;
      RECT 53.96 40.41 67.14 40.58 ;
      RECT 53.96 31.835 67.14 32.005 ;
      RECT 53.96 32.005 54.13 40.41 ;
      RECT 66.935 36.275 67.14 40.41 ;
      RECT 66.97 36.065 67.14 36.275 ;
      RECT 66.935 32.005 67.14 36.065 ;
      RECT 64.845 70.16 65.875 89.93 ;
      RECT 64.845 47.16 65.875 66.93 ;
      RECT 62.865 47.525 63.395 65.695 ;
      RECT 62.885 65.695 63.395 67.035 ;
      RECT 62.885 47.325 63.395 47.525 ;
      RECT 62.865 70.525 63.395 88.695 ;
      RECT 62.885 88.695 63.395 90.035 ;
      RECT 62.885 70.325 63.395 70.525 ;
      RECT 60.245 70.16 61.435 89.87 ;
      RECT 65.61 36.19 65.785 39.29 ;
      RECT 65.61 39.29 65.78 39.35 ;
      RECT 65.61 32.56 65.78 36.19 ;
      RECT 64.825 32.62 65 35.77 ;
      RECT 64.83 35.77 65 39.35 ;
      RECT 64.83 32.56 65 32.62 ;
      RECT 64.05 36.19 64.225 39.29 ;
      RECT 64.05 39.29 64.22 39.35 ;
      RECT 64.05 32.56 64.22 36.19 ;
      RECT 63.265 32.62 63.44 35.77 ;
      RECT 63.27 35.77 63.44 39.35 ;
      RECT 63.27 32.56 63.44 32.62 ;
      RECT 62.49 36.19 62.665 39.29 ;
      RECT 62.49 39.29 62.66 39.35 ;
      RECT 62.49 32.56 62.66 36.19 ;
      RECT 61.705 32.62 61.88 35.77 ;
      RECT 61.71 35.77 61.88 39.35 ;
      RECT 61.71 32.56 61.88 32.62 ;
      RECT 60.93 36.19 61.105 39.29 ;
      RECT 39.83 13.99 40 14.725 ;
      RECT 39.83 9.975 40 11.04 ;
      RECT 39.795 4.82 40.025 7.77 ;
      RECT 39.83 7.77 40 8.505 ;
      RECT 39.83 3.755 40 4.82 ;
      RECT 39.795 17.26 40.025 20.21 ;
      RECT 39.83 20.21 40 20.945 ;
      RECT 39.83 16.195 40 17.26 ;
      RECT 49.555 11.04 49.785 13.99 ;
      RECT 49.59 13.99 49.76 14.725 ;
      RECT 49.59 9.975 49.76 11.04 ;
      RECT 48.09 11.04 48.32 13.99 ;
      RECT 48.11 13.99 48.28 14.725 ;
      RECT 48.11 9.975 48.28 11.04 ;
      RECT 49.555 4.82 49.785 7.77 ;
      RECT 49.59 7.77 49.76 8.505 ;
      RECT 49.59 3.755 49.76 4.82 ;
      RECT 48.09 4.82 48.32 7.77 ;
      RECT 48.11 7.77 48.28 8.505 ;
      RECT 48.11 3.755 48.28 4.82 ;
      RECT 49.555 17.26 49.785 20.21 ;
      RECT 49.59 20.21 49.76 20.945 ;
      RECT 49.59 16.195 49.76 17.26 ;
      RECT 48.09 17.26 48.32 20.21 ;
      RECT 48.11 20.21 48.28 20.945 ;
      RECT 48.11 16.195 48.28 17.26 ;
      RECT 59.315 11.04 59.545 13.99 ;
      RECT 59.35 13.99 59.52 14.725 ;
      RECT 59.35 9.975 59.52 11.04 ;
      RECT 57.85 11.04 58.08 13.99 ;
      RECT 57.87 13.99 58.04 14.725 ;
      RECT 57.87 9.975 58.04 11.04 ;
      RECT 59.315 4.82 59.545 7.77 ;
      RECT 59.35 7.77 59.52 8.505 ;
      RECT 59.35 3.755 59.52 4.82 ;
      RECT 57.85 4.82 58.08 7.77 ;
      RECT 57.87 7.77 58.04 8.505 ;
      RECT 57.87 3.755 58.04 4.82 ;
      RECT 57.555 23.48 57.785 26.43 ;
      RECT 57.59 26.43 57.76 27.165 ;
      RECT 57.59 22.415 57.76 23.48 ;
      RECT 59.315 17.26 59.545 20.21 ;
      RECT 59.35 20.21 59.52 20.945 ;
      RECT 59.35 16.195 59.52 17.26 ;
      RECT 57.85 17.26 58.08 20.21 ;
      RECT 57.87 20.21 58.04 20.945 ;
      RECT 57.87 16.195 58.04 17.26 ;
      RECT 57.815 21.735 61.815 21.965 ;
      RECT 61.85 23.48 62.08 26.43 ;
      RECT 61.87 26.43 62.04 27.165 ;
      RECT 61.87 22.415 62.04 23.48 ;
      RECT 63.315 23.48 63.545 26.43 ;
      RECT 63.35 26.43 63.52 27.165 ;
      RECT 63.35 22.415 63.52 23.48 ;
      RECT 63.575 21.735 67.575 21.965 ;
      RECT 67.61 11.04 67.84 13.99 ;
      RECT 67.63 13.99 67.8 14.725 ;
      RECT 67.63 9.975 67.8 11.04 ;
      RECT 67.61 4.82 67.84 7.77 ;
      RECT 67.63 7.77 67.8 8.505 ;
      RECT 67.63 3.755 67.8 4.82 ;
      RECT 67.61 23.48 67.84 26.43 ;
      RECT 67.63 26.43 67.8 27.165 ;
      RECT 67.63 22.415 67.8 23.48 ;
      RECT 67.61 17.26 67.84 20.21 ;
      RECT 67.63 20.21 67.8 20.945 ;
      RECT 67.63 16.195 67.8 17.26 ;
      RECT 1.07 43.27 1.4 43.44 ;
      RECT 1.145 43.44 1.315 43.81 ;
      RECT 4.735 37.425 45.955 37.595 ;
      RECT 4.735 29.43 4.905 37.425 ;
      RECT 45.755 29.43 45.955 37.425 ;
      RECT 4.735 29.23 45.955 29.43 ;
      RECT 8.05 43.27 8.69 43.44 ;
      RECT 6.115 29.78 6.285 36.57 ;
      RECT 12.355 29.78 12.525 36.57 ;
      RECT 11.575 29.77 11.745 36.57 ;
      RECT 10.795 29.78 10.965 36.57 ;
      RECT 10.015 29.775 10.185 36.57 ;
      RECT 9.235 29.78 9.405 36.57 ;
      RECT 8.455 29.77 8.625 36.57 ;
      RECT 7.675 29.78 7.845 36.57 ;
      RECT 6.895 29.775 7.065 36.57 ;
      RECT 14.385 47.16 15.435 66.93 ;
      RECT 16.865 47.525 17.395 65.695 ;
      RECT 16.885 65.695 17.395 67.035 ;
      RECT 16.885 47.325 17.395 47.525 ;
      RECT 18.595 29.78 18.765 36.57 ;
      RECT 17.815 29.77 17.985 36.57 ;
      RECT 17.035 29.78 17.205 36.57 ;
      RECT 16.255 29.77 16.425 36.57 ;
      RECT 15.475 29.78 15.645 36.57 ;
      RECT 14.695 29.77 14.865 36.57 ;
      RECT 13.915 29.78 14.085 36.57 ;
      RECT 13.135 29.775 13.305 36.57 ;
      RECT 18.845 47.16 20.035 66.87 ;
      RECT 13.085 46.99 13.255 67.965 ;
      RECT 13.09 46.74 64.5 46.815 ;
      RECT 13.085 46.815 64.5 46.99 ;
      RECT 15.705 67.34 64.5 68.995 ;
      RECT 23.51 68.995 64.5 69.99 ;
      RECT 23.585 70.16 24.635 89.93 ;
      RECT 21.465 47.525 21.995 65.695 ;
      RECT 21.485 65.695 21.995 67.035 ;
      RECT 21.485 47.325 21.995 47.525 ;
      RECT 25.615 29.775 25.785 36.57 ;
      RECT 24.835 29.78 25.005 36.57 ;
      RECT 24.055 29.77 24.225 36.57 ;
      RECT 23.275 29.78 23.445 36.57 ;
      RECT 22.495 29.775 22.665 36.57 ;
      RECT 21.715 29.78 21.885 36.57 ;
      RECT 20.935 29.77 21.105 36.57 ;
      RECT 20.155 29.78 20.325 36.57 ;
      RECT 19.375 29.775 19.545 36.57 ;
      RECT 23.445 47.16 24.635 66.87 ;
      RECT 26.065 47.525 26.595 65.695 ;
      RECT 26.085 65.695 26.595 67.035 ;
      RECT 26.085 47.325 26.595 47.525 ;
      RECT 30.665 47.525 31.195 65.695 ;
      RECT 30.685 65.695 31.195 67.035 ;
      RECT 30.685 47.325 31.195 47.525 ;
      RECT 30.665 70.525 31.195 88.695 ;
      RECT 30.685 88.695 31.195 90.035 ;
      RECT 30.685 70.325 31.195 70.525 ;
      RECT 26.065 70.525 26.595 88.695 ;
      RECT 26.085 88.695 26.595 90.035 ;
      RECT 26.085 70.325 26.595 70.525 ;
      RECT 69.78 21.235 70.63 22.52 ;
      RECT 69.765 16.165 70.63 21.235 ;
      RECT 69.78 14.915 70.63 16.165 ;
      RECT 67.975 31.06 68.865 40.48 ;
      RECT 67.975 41.315 68.865 41.455 ;
      RECT 68 40.48 68.83 41.315 ;
      RECT 52.32 31.06 53.21 41.455 ;
      RECT 54.16 28.345 70.63 29.3 ;
      RECT 52.32 41.455 68.865 42.495 ;
      RECT 52.32 29.3 68.865 31.06 ;
      RECT 14.515 17.26 14.745 20.21 ;
      RECT 14.55 20.21 14.72 20.945 ;
      RECT 14.55 16.195 14.72 17.26 ;
      RECT 18.81 17.26 19.04 20.21 ;
      RECT 18.83 20.21 19 20.945 ;
      RECT 18.83 16.195 19 17.26 ;
      RECT 14.515 11.04 14.745 13.99 ;
      RECT 14.55 13.99 14.72 14.725 ;
      RECT 14.55 9.975 14.72 11.04 ;
      RECT 18.81 11.04 19.04 13.99 ;
      RECT 18.83 13.99 19 14.725 ;
      RECT 18.83 9.975 19 11.04 ;
      RECT 14.515 4.82 14.745 7.77 ;
      RECT 14.55 7.77 14.72 8.505 ;
      RECT 14.55 3.755 14.72 4.82 ;
      RECT 18.81 4.82 19.04 7.77 ;
      RECT 18.83 7.77 19 8.505 ;
      RECT 18.83 3.755 19 4.82 ;
      RECT 56.82 27.485 68.57 27.715 ;
      RECT 56.82 23.48 57.05 27.485 ;
      RECT 62.58 23.48 62.81 27.485 ;
      RECT 68.34 23.48 68.57 27.485 ;
      RECT 56.85 21.495 57.02 23.48 ;
      RECT 62.61 21.495 62.78 23.48 ;
      RECT 68.37 21.495 68.54 23.48 ;
      RECT 13.78 21.265 68.57 21.495 ;
      RECT 48.82 17.26 49.05 21.265 ;
      RECT 58.58 17.26 58.81 21.265 ;
      RECT 68.34 17.26 68.57 21.265 ;
      RECT 13.78 17.26 14.01 21.265 ;
      RECT 19.54 17.26 19.77 21.265 ;
      RECT 29.3 17.26 29.53 21.265 ;
      RECT 39.06 17.26 39.29 21.265 ;
      RECT 48.85 15.275 49.02 17.26 ;
      RECT 58.61 15.275 58.78 17.26 ;
      RECT 68.37 15.275 68.54 17.26 ;
      RECT 13.81 15.275 13.98 17.26 ;
      RECT 19.57 15.275 19.74 17.26 ;
      RECT 29.33 15.275 29.5 17.26 ;
      RECT 39.09 15.275 39.26 17.26 ;
      RECT 13.78 15.045 68.57 15.275 ;
      RECT 48.82 11.04 49.05 15.045 ;
      RECT 58.58 11.04 58.81 15.045 ;
      RECT 68.34 11.04 68.57 15.045 ;
      RECT 13.78 11.04 14.01 15.045 ;
      RECT 19.54 11.04 19.77 15.045 ;
      RECT 29.3 11.04 29.53 15.045 ;
      RECT 39.06 11.04 39.29 15.045 ;
      RECT 48.85 9.055 49.02 11.04 ;
      RECT 58.61 9.055 58.78 11.04 ;
      RECT 68.37 9.055 68.54 11.04 ;
      RECT 13.81 9.055 13.98 11.04 ;
      RECT 19.57 9.055 19.74 11.04 ;
      RECT 29.33 9.055 29.5 11.04 ;
      RECT 39.09 9.055 39.26 11.04 ;
      RECT 13.78 8.825 68.57 9.055 ;
      RECT 48.82 4.82 49.05 8.825 ;
      RECT 58.58 4.82 58.81 8.825 ;
      RECT 68.34 4.82 68.57 8.825 ;
      RECT 13.78 4.82 14.01 8.825 ;
      RECT 19.54 4.82 19.77 8.825 ;
      RECT 29.3 4.82 29.53 8.825 ;
      RECT 39.06 4.82 39.29 8.825 ;
      RECT 48.85 2.835 49.02 4.82 ;
      RECT 58.61 2.835 58.78 4.82 ;
      RECT 68.37 2.835 68.54 4.82 ;
      RECT 39.26 2.605 48.85 2.635 ;
      RECT 49.02 2.605 58.61 2.635 ;
      RECT 58.78 2.605 68.37 2.635 ;
      RECT 13.81 2.635 68.54 2.835 ;
      RECT 13.81 2.835 13.98 4.82 ;
      RECT 19.57 2.835 19.74 4.82 ;
      RECT 29.33 2.835 29.5 4.82 ;
      RECT 39.09 2.835 39.26 4.82 ;
      RECT 13.98 2.605 19.57 2.635 ;
      RECT 19.74 2.605 29.33 2.635 ;
      RECT 29.5 2.605 39.09 2.635 ;
      RECT 14.775 15.515 18.775 15.745 ;
      RECT 14.775 9.295 18.775 9.525 ;
      RECT 14.775 3.075 18.775 3.305 ;
      RECT 20.275 17.26 20.505 20.21 ;
      RECT 20.31 20.21 20.48 20.945 ;
      RECT 20.31 16.195 20.48 17.26 ;
      RECT 20.275 11.04 20.505 13.99 ;
      RECT 20.31 13.99 20.48 14.725 ;
      RECT 20.31 9.975 20.48 11.04 ;
      RECT 20.275 4.82 20.505 7.77 ;
      RECT 20.31 7.77 20.48 8.505 ;
      RECT 20.31 3.755 20.48 4.82 ;
      RECT 30.035 17.26 30.265 20.21 ;
      RECT 30.07 20.21 30.24 20.945 ;
      RECT 30.07 16.195 30.24 17.26 ;
      RECT 28.57 17.26 28.8 20.21 ;
      RECT 28.59 20.21 28.76 20.945 ;
      RECT 28.59 16.195 28.76 17.26 ;
      RECT 30.035 11.04 30.265 13.99 ;
      RECT 30.07 13.99 30.24 14.725 ;
      RECT 30.07 9.975 30.24 11.04 ;
      RECT 28.57 11.04 28.8 13.99 ;
      RECT 28.59 13.99 28.76 14.725 ;
      RECT 28.59 9.975 28.76 11.04 ;
      RECT 30.035 4.82 30.265 7.77 ;
      RECT 30.07 7.77 30.24 8.505 ;
      RECT 30.07 3.755 30.24 4.82 ;
      RECT 28.57 4.82 28.8 7.77 ;
      RECT 28.59 7.77 28.76 8.505 ;
      RECT 28.59 3.755 28.76 4.82 ;
      RECT 38.33 17.26 38.56 20.21 ;
      RECT 38.35 20.21 38.52 20.945 ;
      RECT 38.35 16.195 38.52 17.26 ;
      RECT 38.33 11.04 38.56 13.99 ;
      RECT 38.35 13.99 38.52 14.725 ;
      RECT 38.35 9.975 38.52 11.04 ;
      RECT 38.33 4.82 38.56 7.77 ;
      RECT 38.35 7.77 38.52 8.505 ;
      RECT 38.35 3.755 38.52 4.82 ;
      RECT 39.795 11.04 40.025 13.99 ;
      RECT 67.265 46.35 68.155 101.315 ;
      RECT 67.265 165.99 68.155 196.835 ;
      RECT 11.105 45.46 68.155 46.35 ;
      RECT 11.1 196.835 68.155 197.725 ;
      RECT 11.1 171.025 11.99 196.835 ;
      RECT 11.125 135.315 22.66 136.165 ;
      RECT 11.105 69.975 22.68 70.865 ;
      RECT 21.79 70.865 22.68 97.45 ;
      RECT 67.29 101.71 68.155 165.59 ;
      RECT 67.29 101.315 68.14 101.71 ;
      RECT 67.29 165.59 68.14 165.99 ;
      RECT 11.125 170.515 11.975 171.025 ;
      RECT 10.77 162.655 11.975 170.515 ;
      RECT 11.105 46.35 11.995 69.975 ;
      RECT 21.81 97.45 22.66 135.315 ;
      RECT 11.125 158.915 11.975 162.655 ;
      RECT 11.125 136.165 12.1 158.915 ;
      RECT 68.875 44.755 70.125 45.995 ;
      RECT 9.135 43.505 70.125 44.755 ;
      RECT 9.15 198.445 70.125 199.695 ;
      RECT 9.15 170.97 10.4 198.445 ;
      RECT 9.17 133.35 20.99 134.54 ;
      RECT 9.135 71.57 21.085 72.82 ;
      RECT 68.905 45.995 70.095 46.185 ;
      RECT 68.875 46.185 70.125 198.445 ;
      RECT 9.2 133.205 14.19 133.35 ;
      RECT 9.135 44.755 10.385 71.57 ;
      RECT 19.8 72.82 21.085 96.895 ;
      RECT 19.565 97.5 20.99 133.145 ;
      RECT 19.8 96.895 20.99 97.5 ;
      RECT 9.17 170.72 10.36 170.97 ;
      RECT 9.17 134.54 10.36 162.655 ;
      RECT 17.835 133.145 20.99 133.35 ;
      RECT 8.51 162.655 10.36 170.72 ;
      RECT 47.31 29.525 48.2 38.695 ;
      RECT 47.31 28.03 48.2 29.215 ;
      RECT 3.13 39.565 48.2 39.585 ;
      RECT 3.13 27.14 48.2 27.16 ;
      RECT 47.33 29.215 48.18 29.525 ;
      RECT 3.1 28.03 4.02 38.695 ;
      RECT 3.1 27.16 48.2 28.03 ;
      RECT 3.1 38.695 48.2 39.565 ;
      RECT 11.65 1 70.65 1.89 ;
      RECT 11.65 22.35 55.05 23.24 ;
      RECT 69.76 1.89 70.65 2.77 ;
      RECT 54.16 23.24 55.05 28.345 ;
      RECT 69.74 22.52 70.63 28.345 ;
      RECT 11.65 1.89 12.54 22.23 ;
      RECT 11.65 22.23 55.03 22.35 ;
      RECT 69.765 3.845 70.63 8.915 ;
      RECT 69.78 2.77 70.63 3.845 ;
      RECT 69.765 9.845 70.63 14.915 ;
      RECT 69.78 8.915 70.63 9.845 ;
    LAYER met3 ;
      RECT 51.44 98.135 75 99.55 ;
      RECT 49.29 0 75 95.985 ;
      RECT 49.29 95.985 75 98.135 ;
      RECT 61.89 175.06 75 190.44 ;
      RECT 59.685 172.855 75 175.06 ;
      RECT 51.44 99.55 75 107.795 ;
      RECT 49.255 110.605 52.885 168.97 ;
      RECT 49.255 168.97 49.375 172.48 ;
      RECT 49.255 107.985 52.885 110.605 ;
      RECT 59.685 107.795 75 172.855 ;
      RECT 43.24 100.45 44.95 101.97 ;
      RECT 43.295 100.395 44.95 100.45 ;
      RECT 43.785 99.905 44.95 100.395 ;
      RECT 43.24 101.97 44.95 102.67 ;
      RECT 49.255 172.48 49.375 190.42 ;
      RECT 43.94 102.67 50.265 107.985 ;
      RECT 37.22 190.42 49.375 190.44 ;
      RECT 0 195.475 75 200 ;
      RECT 37.22 190.44 75 195.475 ;
      RECT 37.22 175.185 37.565 190.42 ;
      RECT 32.33 105.82 42.455 110.785 ;
      RECT 32.33 110.785 42.455 170.295 ;
      RECT 32.33 170.295 37.565 175.185 ;
      RECT 32.33 105.025 37.49 105.82 ;
      RECT 37.295 100.06 37.49 105.025 ;
      RECT 29.925 93.265 31.545 96.21 ;
      RECT 29.925 96.21 30.935 96.82 ;
      RECT 30.4 92.79 31.545 93.265 ;
      RECT 37.295 0 37.49 100.06 ;
      RECT 0 175.73 12.225 195.475 ;
      RECT 0 172.855 12.225 175.73 ;
      RECT 0 102.035 15.1 172.855 ;
      RECT 0 93.79 15.1 102.035 ;
      RECT 0 92.375 23.345 93.79 ;
      RECT 0 0 25.495 90.225 ;
      RECT 0 90.225 23.345 92.375 ;
      RECT 25.41 172.475 25.53 195.475 ;
      RECT 21.9 168.965 25.53 172.475 ;
      RECT 21.9 104.845 25.53 168.965 ;
      RECT 24.52 102.225 25.53 104.845 ;
      RECT 58.49 106.45 75 106.6 ;
      RECT 58.64 106.6 75 106.75 ;
      RECT 58.79 106.75 75 106.9 ;
      RECT 58.94 106.9 75 107.05 ;
      RECT 59.09 107.05 75 107.2 ;
      RECT 59.24 107.2 75 107.35 ;
      RECT 59.39 107.35 75 107.5 ;
      RECT 59.54 107.5 75 107.65 ;
      RECT 59.685 107.65 75 107.795 ;
      RECT 32.33 110.17 41.84 110.32 ;
      RECT 32.33 110.02 41.69 110.17 ;
      RECT 32.33 109.87 41.54 110.02 ;
      RECT 32.33 109.72 41.39 109.87 ;
      RECT 32.33 109.57 41.24 109.72 ;
      RECT 32.33 109.42 41.09 109.57 ;
      RECT 32.33 109.27 40.94 109.42 ;
      RECT 32.33 109.12 40.79 109.27 ;
      RECT 32.33 108.97 40.64 109.12 ;
      RECT 32.33 108.82 40.49 108.97 ;
      RECT 32.33 108.67 40.34 108.82 ;
      RECT 32.33 108.52 40.19 108.67 ;
      RECT 32.33 108.37 40.04 108.52 ;
      RECT 32.33 108.22 39.89 108.37 ;
      RECT 32.33 108.07 39.74 108.22 ;
      RECT 32.33 107.92 39.59 108.07 ;
      RECT 32.33 107.77 39.44 107.92 ;
      RECT 32.33 107.62 39.29 107.77 ;
      RECT 32.33 107.47 39.14 107.62 ;
      RECT 32.33 107.32 38.99 107.47 ;
      RECT 32.33 107.17 38.84 107.32 ;
      RECT 32.33 107.02 38.69 107.17 ;
      RECT 32.33 106.87 38.54 107.02 ;
      RECT 32.33 106.72 38.39 106.87 ;
      RECT 32.33 106.57 38.24 106.72 ;
      RECT 32.33 106.42 38.09 106.57 ;
      RECT 32.33 106.27 37.94 106.42 ;
      RECT 32.33 106.12 37.79 106.27 ;
      RECT 32.33 105.97 37.64 106.12 ;
      RECT 32.33 105.82 37.49 105.97 ;
      RECT 32.39 104.965 37.49 105.025 ;
      RECT 32.54 104.815 37.49 104.965 ;
      RECT 32.69 104.665 37.49 104.815 ;
      RECT 32.84 104.515 37.49 104.665 ;
      RECT 32.99 104.365 37.49 104.515 ;
      RECT 33.14 104.215 37.49 104.365 ;
      RECT 33.29 104.065 37.49 104.215 ;
      RECT 33.44 103.915 37.49 104.065 ;
      RECT 33.59 103.765 37.49 103.915 ;
      RECT 33.74 103.615 37.49 103.765 ;
      RECT 33.89 103.465 37.49 103.615 ;
      RECT 34.04 103.315 37.49 103.465 ;
      RECT 34.19 103.165 37.49 103.315 ;
      RECT 34.34 103.015 37.49 103.165 ;
      RECT 34.49 102.865 37.49 103.015 ;
      RECT 34.64 102.715 37.49 102.865 ;
      RECT 34.79 102.565 37.49 102.715 ;
      RECT 34.94 102.415 37.49 102.565 ;
      RECT 35.09 102.265 37.49 102.415 ;
      RECT 35.24 102.115 37.49 102.265 ;
      RECT 35.39 101.965 37.49 102.115 ;
      RECT 35.54 101.815 37.49 101.965 ;
      RECT 35.69 101.665 37.49 101.815 ;
      RECT 35.84 101.515 37.49 101.665 ;
      RECT 35.99 101.365 37.49 101.515 ;
      RECT 36.14 101.215 37.49 101.365 ;
      RECT 36.29 101.065 37.49 101.215 ;
      RECT 36.44 100.915 37.49 101.065 ;
      RECT 36.59 100.765 37.49 100.915 ;
      RECT 36.74 100.615 37.49 100.765 ;
      RECT 36.89 100.465 37.49 100.615 ;
      RECT 37.04 100.315 37.49 100.465 ;
      RECT 37.19 100.165 37.49 100.315 ;
      RECT 37.34 100.015 37.49 100.165 ;
      RECT 49.44 95.985 75 96.135 ;
      RECT 49.59 96.135 75 96.285 ;
      RECT 49.74 96.285 75 96.435 ;
      RECT 49.89 96.435 75 96.585 ;
      RECT 50.04 96.585 75 96.735 ;
      RECT 50.19 96.735 75 96.885 ;
      RECT 50.34 96.885 75 97.035 ;
      RECT 50.49 97.035 75 97.185 ;
      RECT 50.64 97.185 75 97.335 ;
      RECT 50.79 97.335 75 97.485 ;
      RECT 50.94 97.485 75 97.635 ;
      RECT 51.09 97.635 75 97.785 ;
      RECT 51.24 97.785 75 97.935 ;
      RECT 51.39 97.935 75 98.085 ;
      RECT 51.44 98.085 75 98.135 ;
      RECT 51.59 99.55 75 99.7 ;
      RECT 51.74 99.7 75 99.85 ;
      RECT 51.89 99.85 75 100 ;
      RECT 52.04 100 75 100.15 ;
      RECT 52.19 100.15 75 100.3 ;
      RECT 52.34 100.3 75 100.45 ;
      RECT 52.49 100.45 75 100.6 ;
      RECT 52.64 100.6 75 100.75 ;
      RECT 52.79 100.75 75 100.9 ;
      RECT 52.94 100.9 75 101.05 ;
      RECT 53.09 101.05 75 101.2 ;
      RECT 53.24 101.2 75 101.35 ;
      RECT 53.39 101.35 75 101.5 ;
      RECT 53.54 101.5 75 101.65 ;
      RECT 53.69 101.65 75 101.8 ;
      RECT 53.84 101.8 75 101.95 ;
      RECT 53.99 101.95 75 102.1 ;
      RECT 54.14 102.1 75 102.25 ;
      RECT 54.29 102.25 75 102.4 ;
      RECT 54.44 102.4 75 102.55 ;
      RECT 54.59 102.55 75 102.7 ;
      RECT 54.74 102.7 75 102.85 ;
      RECT 54.89 102.85 75 103 ;
      RECT 55.04 103 75 103.15 ;
      RECT 55.19 103.15 75 103.3 ;
      RECT 55.34 103.3 75 103.45 ;
      RECT 55.49 103.45 75 103.6 ;
      RECT 55.64 103.6 75 103.75 ;
      RECT 55.79 103.75 75 103.9 ;
      RECT 55.94 103.9 75 104.05 ;
      RECT 56.09 104.05 75 104.2 ;
      RECT 56.24 104.2 75 104.35 ;
      RECT 56.39 104.35 75 104.5 ;
      RECT 56.54 104.5 75 104.65 ;
      RECT 56.69 104.65 75 104.8 ;
      RECT 56.84 104.8 75 104.95 ;
      RECT 56.99 104.95 75 105.1 ;
      RECT 57.14 105.1 75 105.25 ;
      RECT 57.29 105.25 75 105.4 ;
      RECT 57.44 105.4 75 105.55 ;
      RECT 57.59 105.55 75 105.7 ;
      RECT 57.74 105.7 75 105.85 ;
      RECT 57.89 105.85 75.105 ;
      RECT 58.04 106 75 106.15 ;
      RECT 58.19 106.15 75 106.3 ;
      RECT 58.34 106.3 75 106.45 ;
      RECT 0 173.155 14.65 173.305 ;
      RECT 0 173.305 14.5 173.455 ;
      RECT 0 173.455 14.35 173.605 ;
      RECT 0 173.605 14.2 173.755 ;
      RECT 0 173.755 14.05 173.905 ;
      RECT 0 173.905 13.9 174.055 ;
      RECT 0 174.055 13.75 174.205 ;
      RECT 0 174.205 13.6 174.355 ;
      RECT 0 174.355 13.45 174.505 ;
      RECT 0 174.505 13.3 174.655 ;
      RECT 0 174.655 13.15 174.805 ;
      RECT 0 174.805 13.0 174.955 ;
      RECT 0 174.955 12.85 175.105 ;
      RECT 0 175.105 12.7 175.255 ;
      RECT 0 175.255 12.55 175.405 ;
      RECT 0 175.405 12.4 175.555 ;
      RECT 0 175.555 12.25 175.705 ;
      RECT 0 175.705 12.225 175.73 ;
      RECT 0 93.79 23.195 93.94 ;
      RECT 0 93.94 23.045 94.09 ;
      RECT 0 94.09 22.895 94.24 ;
      RECT 0 94.24 22.745 94.39 ;
      RECT 0 94.39 22.595 94.54 ;
      RECT 0 94.54 22.445 94.69 ;
      RECT 0 94.69 22.295 94.84 ;
      RECT 0 94.84 22.145 94.99 ;
      RECT 0 94.99 21.995 95.14 ;
      RECT 0 95.14 21.845 95.29 ;
      RECT 0 95.29 21.695 95.44 ;
      RECT 0 95.44 21.545 95.59 ;
      RECT 0 95.59 21.395 95.74 ;
      RECT 0 95.74 21.245 95.89 ;
      RECT 0 95.89 21.095 96.04 ;
      RECT 0 96.04 20.945 96.19 ;
      RECT 0 96.19 20.795 96.34 ;
      RECT 0 96.34 20.645 96.49 ;
      RECT 0 96.49 20.495 96.64 ;
      RECT 0 96.64 20.345 96.79 ;
      RECT 0 96.79 20.195 96.94 ;
      RECT 0 96.94 20.045 97.09 ;
      RECT 0 97.09 19.895 97.24 ;
      RECT 0 97.24 19.745 97.39 ;
      RECT 0 97.39 19.595 97.54 ;
      RECT 0 97.54 19.445 97.69 ;
      RECT 0 97.69 19.295 97.84 ;
      RECT 0 97.84 19.145 97.99 ;
      RECT 0 97.99 18.995 98.14 ;
      RECT 0 98.14 18.845 98.29 ;
      RECT 0 98.29 18.695 98.44 ;
      RECT 0 98.44 18.545 98.59 ;
      RECT 0 98.59 18.395 98.74 ;
      RECT 0 98.74 18.245 98.89 ;
      RECT 0 98.89 18.095 99.04 ;
      RECT 0 99.04 17.945 99.19 ;
      RECT 0 99.19 17.795 99.34 ;
      RECT 0 99.34 17.645 99.49 ;
      RECT 0 99.49 17.495 99.64 ;
      RECT 0 99.64 17.345 99.79 ;
      RECT 0 99.79 17.195 99.94 ;
      RECT 0 99.94 17.045 100.09 ;
      RECT 0 100.09 16.895 100.24 ;
      RECT 0 100.24 16.745 100.39 ;
      RECT 0 100.39 16.595 100.54 ;
      RECT 0 100.54 16.445 100.69 ;
      RECT 0 100.69 16.295 100.84 ;
      RECT 0 100.84 16.145 100.99 ;
      RECT 0 100.99 15.995 101.14 ;
      RECT 0 101.14 15.845 101.29 ;
      RECT 0 101.29 15.695 101.44 ;
      RECT 0 101.44 15.545 101.59 ;
      RECT 0 101.59 15.395 101.74 ;
      RECT 0 101.74 15.245 101.89 ;
      RECT 0 101.89 15.1 102.035 ;
      RECT 0 90.225 25.345 90.375 ;
      RECT 0 90.375 25.195 90.525 ;
      RECT 0 90.525 25.045 90.675 ;
      RECT 0 90.675 24.895 90.825 ;
      RECT 0 90.825 24.745 90.975 ;
      RECT 0 90.975 24.595 91.125 ;
      RECT 0 91.125 24.445 91.275 ;
      RECT 0 91.275 24.295 91.425 ;
      RECT 0 91.425 24.145 91.575 ;
      RECT 0 91.575 23.995 91.725 ;
      RECT 0 91.725 23.845 91.875 ;
      RECT 0 91.875 23.695 92.025 ;
      RECT 0 92.025 23.545 92.175 ;
      RECT 0 92.175 23.395 92.325 ;
      RECT 0 92.325 23.345 92.375 ;
      RECT 37.39 175.245 37.395 175.355 ;
      RECT 37.28 175.095 37.505 175.245 ;
      RECT 37.13 174.945 37.655 175.095 ;
      RECT 36.98 174.795 37.805 174.945 ;
      RECT 36.83 174.645 37.955 174.795 ;
      RECT 36.68 174.495 38.105 174.645 ;
      RECT 36.53 174.345 38.255 174.495 ;
      RECT 36.38 174.195 38.405 174.345 ;
      RECT 36.23 174.045 38.555 174.195 ;
      RECT 36.08 173.895 38.705 174.045 ;
      RECT 35.93 173.745 38.855 173.895 ;
      RECT 35.78 173.595 39.005 173.745 ;
      RECT 35.63 173.445 39.155 173.595 ;
      RECT 35.48 173.295 39.305 173.445 ;
      RECT 35.33 173.145 39.455 173.295 ;
      RECT 35.18 172.995 39.605 173.145 ;
      RECT 35.03 172.845 39.755 172.995 ;
      RECT 34.88 172.695 39.905 172.845 ;
      RECT 34.73 172.545 40.055 172.695 ;
      RECT 34.58 172.395 40.205 172.545 ;
      RECT 34.43 172.245 40.355 172.395 ;
      RECT 34.28 172.095 40.505 172.245 ;
      RECT 34.13 171.945 40.655 172.095 ;
      RECT 33.98 171.795 40.805 171.945 ;
      RECT 33.83 171.645 40.955 171.795 ;
      RECT 33.68 171.495 41.105 171.645 ;
      RECT 33.53 171.345 41.255 171.495 ;
      RECT 33.38 171.195 41.405 171.345 ;
      RECT 33.23 171.045 41.555 171.195 ;
      RECT 33.08 170.895 41.705 171.045 ;
      RECT 32.93 170.745 41.855 170.895 ;
      RECT 32.78 170.595 42.005 170.745 ;
      RECT 32.63 170.445 42.155 170.595 ;
      RECT 32.48 170.295 42.305 170.445 ;
      RECT 32.33 110.77 42.44 110.785 ;
      RECT 32.33 110.62 42.29 110.77 ;
      RECT 32.33 110.47 42.14 110.62 ;
      RECT 32.33 110.32 41.99 110.47 ;
      RECT 37.28 175.095 37.505 175.245 ;
      RECT 37.13 174.945 37.655 175.095 ;
      RECT 36.98 174.795 37.805 174.945 ;
      RECT 36.83 174.645 37.955 174.795 ;
      RECT 36.68 174.495 38.105 174.645 ;
      RECT 36.53 174.345 38.255 174.495 ;
      RECT 36.38 174.195 38.405 174.345 ;
      RECT 36.23 174.045 38.555 174.195 ;
      RECT 36.08 173.895 38.705 174.045 ;
      RECT 35.93 173.745 38.855 173.895 ;
      RECT 35.78 173.595 39.005 173.745 ;
      RECT 35.63 173.445 39.155 173.595 ;
      RECT 35.48 173.295 39.305 173.445 ;
      RECT 35.33 173.145 39.455 173.295 ;
      RECT 35.18 172.995 39.605 173.145 ;
      RECT 35.03 172.845 39.755 172.995 ;
      RECT 34.88 172.695 39.905 172.845 ;
      RECT 34.73 172.545 40.055 172.695 ;
      RECT 34.58 172.395 40.205 172.545 ;
      RECT 34.43 172.245 40.355 172.395 ;
      RECT 34.28 172.095 40.505 172.245 ;
      RECT 34.13 171.945 40.655 172.095 ;
      RECT 33.98 171.795 40.805 171.945 ;
      RECT 33.83 171.645 40.955 171.795 ;
      RECT 33.68 171.495 41.105 171.645 ;
      RECT 33.53 171.345 41.255 171.495 ;
      RECT 33.38 171.195 41.405 171.345 ;
      RECT 33.23 171.045 41.555 171.195 ;
      RECT 33.08 170.895 41.705 171.045 ;
      RECT 32.93 170.745 41.855 170.895 ;
      RECT 32.78 170.595 42.005 170.745 ;
      RECT 32.63 170.445 42.155 170.595 ;
      RECT 32.48 170.295 42.305 170.445 ;
      RECT 32.33 110.77 42.44 110.785 ;
      RECT 32.33 110.62 42.29 110.77 ;
      RECT 32.33 110.47 42.14 110.62 ;
      RECT 32.33 110.32 41.99 110.47 ;
      RECT 32.33 110.17 41.84 110.32 ;
      RECT 32.33 110.02 41.69 110.17 ;
      RECT 32.33 109.87 41.54 110.02 ;
      RECT 32.33 109.72 41.39 109.87 ;
      RECT 32.33 109.57 41.24 109.72 ;
      RECT 32.33 109.42 41.09 109.57 ;
      RECT 32.33 109.27 40.94 109.42 ;
      RECT 32.33 109.12 40.79 109.27 ;
      RECT 32.33 108.97 40.64 109.12 ;
      RECT 32.33 108.82 40.49 108.97 ;
      RECT 32.33 108.67 40.34 108.82 ;
      RECT 32.33 108.52 40.19 108.67 ;
      RECT 32.33 108.37 40.04 108.52 ;
      RECT 32.33 108.22 39.89 108.37 ;
      RECT 32.33 108.07 39.74 108.22 ;
      RECT 32.33 107.92 39.59 108.07 ;
      RECT 32.33 107.77 39.44 107.92 ;
      RECT 32.33 107.62 39.29 107.77 ;
      RECT 32.33 107.47 39.14 107.62 ;
      RECT 32.33 107.32 38.99 107.47 ;
      RECT 32.33 107.17 38.84 107.32 ;
      RECT 32.33 107.02 38.69 107.17 ;
      RECT 32.33 106.87 38.54 107.02 ;
      RECT 32.33 106.72 38.39 106.87 ;
      RECT 32.33 106.57 38.24 106.72 ;
      RECT 32.33 106.42 38.09 106.57 ;
      RECT 32.33 106.27 37.94 106.42 ;
      RECT 32.33 106.12 37.79 106.27 ;
      RECT 32.33 105.97 37.64 106.12 ;
      RECT 32.33 105.82 37.49 105.97 ;
      RECT 32.39 104.965 37.49 105.025 ;
      RECT 32.54 104.815 37.49 104.965 ;
      RECT 32.69 104.665 37.49 104.815 ;
      RECT 32.84 104.515 37.49 104.665 ;
      RECT 32.99 104.365 37.49 104.515 ;
      RECT 33.14 104.215 37.49 104.365 ;
      RECT 33.29 104.065 37.49 104.215 ;
      RECT 33.44 103.915 37.49 104.065 ;
      RECT 33.59 103.765 37.49 103.915 ;
      RECT 33.74 103.615 37.49 103.765 ;
      RECT 33.89 103.465 37.49 103.615 ;
      RECT 34.04 103.315 37.49 103.465 ;
      RECT 34.19 103.165 37.49 103.315 ;
      RECT 34.34 103.015 37.49 103.165 ;
      RECT 34.49 102.865 37.49 103.015 ;
      RECT 34.64 102.715 37.49 102.865 ;
      RECT 34.79 102.565 37.49 102.715 ;
      RECT 34.94 102.415 37.49 102.565 ;
      RECT 35.09 102.265 37.49 102.415 ;
      RECT 35.24 102.115 37.49 102.265 ;
      RECT 35.39 101.965 37.49 102.115 ;
      RECT 35.54 101.815 37.49 101.965 ;
      RECT 35.69 101.665 37.49 101.815 ;
      RECT 35.84 101.515 37.49 101.665 ;
      RECT 35.99 101.365 37.49 101.515 ;
      RECT 36.14 101.215 37.49 101.365 ;
      RECT 36.29 101.065 37.49 101.215 ;
      RECT 36.44 100.915 37.49 101.065 ;
      RECT 36.59 100.765 37.49 100.915 ;
      RECT 36.74 100.615 37.49 100.765 ;
      RECT 36.89 100.465 37.49 100.615 ;
      RECT 37.04 100.315 37.49 100.465 ;
      RECT 37.19 100.165 37.49 100.315 ;
      RECT 37.34 100.015 37.49 100.165 ;
      RECT 37.22 175.27 37.305 175.355 ;
      RECT 37.48 175.27 37.565 175.355 ;
      RECT 59.835 172.855 75 173.005 ;
      RECT 59.985 173.005 75 173.155 ;
      RECT 60.135 173.155 75 173.305 ;
      RECT 60.285 173.305 75 173.455 ;
      RECT 60.435 173.455 75 173.605 ;
      RECT 60.585 173.605 75 173.755 ;
      RECT 60.735 173.755 75 173.905 ;
      RECT 60.885 173.905 75 174.055 ;
      RECT 61.035 174.055 75 174.205 ;
      RECT 61.185 174.205 75 174.355 ;
      RECT 61.335 174.355 75 174.505 ;
      RECT 61.485 174.505 75 174.655 ;
      RECT 61.635 174.655 75 174.805 ;
      RECT 61.785 174.805 75 174.955 ;
      RECT 61.89 174.955 75 175.06 ;
      RECT 0 172.855 14.95 173.005 ;
      RECT 0 173.005 14.8 173.155 ;
      RECT 53.69 101.65 75 101.8 ;
      RECT 53.84 101.8 75 101.95 ;
      RECT 53.99 101.95 75 102.1 ;
      RECT 54.14 102.1 75 102.25 ;
      RECT 54.29 102.25 75 102.4 ;
      RECT 54.44 102.4 75 102.55 ;
      RECT 54.59 102.55 75 102.7 ;
      RECT 54.74 102.7 75 102.85 ;
      RECT 54.89 102.85 75 103 ;
      RECT 55.04 103 75 103.15 ;
      RECT 55.19 103.15 75 103.3 ;
      RECT 55.34 103.3 75 103.45 ;
      RECT 55.49 103.45 75 103.6 ;
      RECT 55.64 103.6 75 103.75 ;
      RECT 55.79 103.75 75 103.9 ;
      RECT 55.94 103.9 75 104.05 ;
      RECT 56.09 104.05 75 104.2 ;
      RECT 56.24 104.2 75 104.35 ;
      RECT 56.39 104.35 75 104.5 ;
      RECT 56.54 104.5 75 104.65 ;
      RECT 56.69 104.65 75 104.8 ;
      RECT 56.84 104.8 75 104.95 ;
      RECT 56.99 104.95 75 105.1 ;
      RECT 57.14 105.1 75 105.25 ;
      RECT 57.29 105.25 75 105.4 ;
      RECT 57.44 105.4 75 105.55 ;
      RECT 57.59 105.55 75 105.7 ;
      RECT 57.74 105.7 75 105.85 ;
      RECT 57.89 105.85 75.105 ;
      RECT 58.04 106 75 106.15 ;
      RECT 58.19 106.15 75 106.3 ;
      RECT 58.34 106.3 75 106.45 ;
      RECT 58.49 106.45 75 106.6 ;
      RECT 58.64 106.6 75 106.75 ;
      RECT 58.79 106.75 75 106.9 ;
      RECT 58.94 106.9 75 107.05 ;
      RECT 59.09 107.05 75 107.2 ;
      RECT 59.24 107.2 75 107.35 ;
      RECT 59.39 107.35 75 107.5 ;
      RECT 59.54 107.5 75 107.65 ;
      RECT 59.685 107.65 75 107.795 ;
      RECT 49.44 95.985 75 96.135 ;
      RECT 49.59 96.135 75 96.285 ;
      RECT 49.74 96.285 75 96.435 ;
      RECT 49.89 96.435 75 96.585 ;
      RECT 50.04 96.585 75 96.735 ;
      RECT 50.19 96.735 75 96.885 ;
      RECT 50.34 96.885 75 97.035 ;
      RECT 50.49 97.035 75 97.185 ;
      RECT 50.64 97.185 75 97.335 ;
      RECT 50.79 97.335 75 97.485 ;
      RECT 50.94 97.485 75 97.635 ;
      RECT 51.09 97.635 75 97.785 ;
      RECT 51.24 97.785 75 97.935 ;
      RECT 51.39 97.935 75 98.085 ;
      RECT 51.44 98.085 75 98.135 ;
      RECT 0 93.79 23.195 93.94 ;
      RECT 0 93.94 23.045 94.09 ;
      RECT 0 94.09 22.895 94.24 ;
      RECT 0 94.24 22.745 94.39 ;
      RECT 0 94.39 22.595 94.54 ;
      RECT 0 94.54 22.445 94.69 ;
      RECT 0 94.69 22.295 94.84 ;
      RECT 0 94.84 22.145 94.99 ;
      RECT 0 94.99 21.995 95.14 ;
      RECT 0 95.14 21.845 95.29 ;
      RECT 0 95.29 21.695 95.44 ;
      RECT 0 95.44 21.545 95.59 ;
      RECT 0 95.59 21.395 95.74 ;
      RECT 0 95.74 21.245 95.89 ;
      RECT 0 95.89 21.095 96.04 ;
      RECT 0 96.04 20.945 96.19 ;
      RECT 0 96.19 20.795 96.34 ;
      RECT 0 96.34 20.645 96.49 ;
      RECT 0 96.49 20.495 96.64 ;
      RECT 0 96.64 20.345 96.79 ;
      RECT 0 96.79 20.195 96.94 ;
      RECT 0 96.94 20.045 97.09 ;
      RECT 0 97.09 19.895 97.24 ;
      RECT 0 97.24 19.745 97.39 ;
      RECT 0 97.39 19.595 97.54 ;
      RECT 0 97.54 19.445 97.69 ;
      RECT 0 97.69 19.295 97.84 ;
      RECT 0 97.84 19.145 97.99 ;
      RECT 0 97.99 18.995 98.14 ;
      RECT 0 98.14 18.845 98.29 ;
      RECT 0 98.29 18.695 98.44 ;
      RECT 0 98.44 18.545 98.59 ;
      RECT 0 98.59 18.395 98.74 ;
      RECT 0 98.74 18.245 98.89 ;
      RECT 0 98.89 18.095 99.04 ;
      RECT 0 99.04 17.945 99.19 ;
      RECT 0 99.19 17.795 99.34 ;
      RECT 0 99.34 17.645 99.49 ;
      RECT 0 99.49 17.495 99.64 ;
      RECT 0 99.64 17.345 99.79 ;
      RECT 0 99.79 17.195 99.94 ;
      RECT 0 99.94 17.045 100.09 ;
      RECT 0 100.09 16.895 100.24 ;
      RECT 0 100.24 16.745 100.39 ;
      RECT 0 100.39 16.595 100.54 ;
      RECT 0 100.54 16.445 100.69 ;
      RECT 0 100.69 16.295 100.84 ;
      RECT 0 100.84 16.145 100.99 ;
      RECT 0 100.99 15.995 101.14 ;
      RECT 0 101.14 15.845 101.29 ;
      RECT 0 101.29 15.695 101.44 ;
      RECT 0 101.44 15.545 101.59 ;
      RECT 0 101.59 15.395 101.74 ;
      RECT 0 101.74 15.245 101.89 ;
      RECT 0 101.89 15.1 102.035 ;
      RECT 0 90.225 25.345 90.375 ;
      RECT 0 90.375 25.195 90.525 ;
      RECT 0 90.525 25.045 90.675 ;
      RECT 0 90.675 24.895 90.825 ;
      RECT 0 90.825 24.745 90.975 ;
      RECT 0 90.975 24.595 91.125 ;
      RECT 0 91.125 24.445 91.275 ;
      RECT 0 91.275 24.295 91.425 ;
      RECT 0 91.425 24.145 91.575 ;
      RECT 0 91.575 23.995 91.725 ;
      RECT 0 91.725 23.845 91.875 ;
      RECT 0 91.875 23.695 92.025 ;
      RECT 0 92.025 23.545 92.175 ;
      RECT 0 92.175 23.395 92.325 ;
      RECT 0 92.325 23.345 92.375 ;
      RECT 37.39 175.245 37.395 175.355 ;
      RECT 44.39 102.97 45.25 103.12 ;
      RECT 44.54 103.12 45.4 103.27 ;
      RECT 44.69 103.27 45.55 103.42 ;
      RECT 44.84 103.42 45.7 103.57 ;
      RECT 44.99 103.57 45.85 103.72 ;
      RECT 45.14 103.72 46.0 103.87 ;
      RECT 45.29 103.87 46.15 104.02 ;
      RECT 45.44 104.02 46.3 104.17 ;
      RECT 45.59 104.17 46.45 104.32 ;
      RECT 45.74 104.32 46.6 104.47 ;
      RECT 45.89 104.47 46.75 104.62 ;
      RECT 46.04 104.62 46.9 104.77 ;
      RECT 46.19 104.77 47.05 104.92 ;
      RECT 46.34 104.92 47.2 105.07 ;
      RECT 46.49 105.07 47.35 105.22 ;
      RECT 46.64 105.22 47.5 105.37 ;
      RECT 46.79 105.37 47.65 105.52 ;
      RECT 46.94 105.52 47.8 105.67 ;
      RECT 47.09 105.67 47.95 105.82 ;
      RECT 47.24 105.82 48.1 105.97 ;
      RECT 47.39 105.97 48.25 106.12 ;
      RECT 47.54 106.12 48.4 106.27 ;
      RECT 47.69 106.27 48.55 106.42 ;
      RECT 47.84 106.42 48.7 106.57 ;
      RECT 47.99 106.57 48.85 106.72 ;
      RECT 48.14 106.72 49.0 106.87 ;
      RECT 48.29 106.87 49.15 107.02 ;
      RECT 48.44 107.02 49.3 107.17 ;
      RECT 48.59 107.17 49.45 107.32 ;
      RECT 48.74 107.32 49.6 107.47 ;
      RECT 48.89 107.47 49.75 107.62 ;
      RECT 49.04 107.62 49.9 107.77 ;
      RECT 49.19 107.77 50.05 107.92 ;
      RECT 49.255 107.92 50.2 107.985 ;
      RECT 49.255 168.97 52.735 169.12 ;
      RECT 49.255 169.12 52.585 169.27 ;
      RECT 49.255 169.27 52.435 169.42 ;
      RECT 49.255 169.42 52.285 169.57 ;
      RECT 49.255 169.57 52.135 169.72 ;
      RECT 49.255 169.72 51.985 169.87 ;
      RECT 49.255 169.87 51.835 170.02 ;
      RECT 49.255 170.02 51.685 170.17 ;
      RECT 49.255 170.17 51.535 170.32 ;
      RECT 49.255 170.32 51.385 170.47 ;
      RECT 49.255 170.47 51.235 170.62 ;
      RECT 49.255 170.62 51.085 170.77 ;
      RECT 49.255 170.77 50.935 170.92 ;
      RECT 49.255 170.92 50.785 171.07 ;
      RECT 49.255 171.07 50.635 171.22 ;
      RECT 49.255 171.22 50.485 171.37 ;
      RECT 49.255 171.37 50.335 171.52 ;
      RECT 49.255 171.52 50.185 171.67 ;
      RECT 49.255 171.67 50.035 171.82 ;
      RECT 49.255 171.82 49.885 171.97 ;
      RECT 49.255 171.97 49.735 172.12 ;
      RECT 49.255 172.12 49.585 172.27 ;
      RECT 49.255 172.27 49.435 172.42 ;
      RECT 49.255 172.42 49.285 172.57 ;
      RECT 49.255 107.985 50.265 108.135 ;
      RECT 49.255 108.135 50.415 108.285 ;
      RECT 49.255 108.285 50.565 108.435 ;
      RECT 49.255 108.435 50.715 108.585 ;
      RECT 49.255 108.585 50.865 108.735 ;
      RECT 49.255 108.735 51.015 108.885 ;
      RECT 49.255 108.885 51.165 109.035 ;
      RECT 49.255 109.035 51.315 109.185 ;
      RECT 49.255 109.185 51.465 109.335 ;
      RECT 49.255 109.335 51.615 109.485 ;
      RECT 49.255 109.485 51.765 109.635 ;
      RECT 49.255 109.635 51.915 109.785 ;
      RECT 49.255 109.785 52.065 109.935 ;
      RECT 49.255 109.935 52.215 110.085 ;
      RECT 49.255 110.085 52.365 110.235 ;
      RECT 49.255 110.235 52.515 110.385 ;
      RECT 49.255 110.385 52.665 110.535 ;
      RECT 49.255 110.535 52.815 110.605 ;
      RECT 0 172.855 14.95 173.005 ;
      RECT 0 173.005 14.8 173.155 ;
      RECT 0 173.155 14.65 173.305 ;
      RECT 0 173.305 14.5 173.455 ;
      RECT 0 173.455 14.35 173.605 ;
      RECT 0 173.605 14.2 173.755 ;
      RECT 0 173.755 14.05 173.905 ;
      RECT 0 173.905 13.9 174.055 ;
      RECT 0 174.055 13.75 174.205 ;
      RECT 0 174.205 13.6 174.355 ;
      RECT 0 174.355 13.45 174.505 ;
      RECT 0 174.505 13.3 174.655 ;
      RECT 0 174.655 13.15 174.805 ;
      RECT 0 174.805 13.0 174.955 ;
      RECT 0 174.955 12.85 175.105 ;
      RECT 0 175.105 12.7 175.255 ;
      RECT 0 175.255 12.55 175.405 ;
      RECT 0 175.405 12.4 175.555 ;
      RECT 0 175.555 12.25 175.705 ;
      RECT 0 175.705 12.225 175.73 ;
      RECT 59.835 172.855 75 173.005 ;
      RECT 59.985 173.005 75 173.155 ;
      RECT 60.135 173.155 75 173.305 ;
      RECT 60.285 173.305 75 173.455 ;
      RECT 60.435 173.455 75 173.605 ;
      RECT 60.585 173.605 75 173.755 ;
      RECT 60.735 173.755 75 173.905 ;
      RECT 60.885 173.905 75 174.055 ;
      RECT 61.035 174.055 75 174.205 ;
      RECT 61.185 174.205 75 174.355 ;
      RECT 61.335 174.355 75 174.505 ;
      RECT 61.485 174.505 75 174.655 ;
      RECT 61.635 174.655 75 174.805 ;
      RECT 61.785 174.805 75 174.955 ;
      RECT 61.89 174.955 75 175.06 ;
      RECT 51.59 99.55 75 99.7 ;
      RECT 51.74 99.7 75 99.85 ;
      RECT 51.89 99.85 75 100 ;
      RECT 52.04 100 75 100.15 ;
      RECT 52.19 100.15 75 100.3 ;
      RECT 52.34 100.3 75 100.45 ;
      RECT 52.49 100.45 75 100.6 ;
      RECT 52.64 100.6 75 100.75 ;
      RECT 52.79 100.75 75 100.9 ;
      RECT 52.94 100.9 75 101.05 ;
      RECT 53.09 101.05 75 101.2 ;
      RECT 53.24 101.2 75 101.35 ;
      RECT 53.39 101.35 75 101.5 ;
      RECT 53.54 101.5 75 101.65 ;
      RECT 29.925 93.265 31.545 96.21 ;
      RECT 43.24 100.45 44.95 101.97 ;
      RECT 21.9 104.845 25.53 168.965 ;
      RECT 37.22 175.355 37.565 190.42 ;
      RECT 49.255 110.605 52.885 168.97 ;
      RECT 37.22 190.42 49.375 190.44 ;
      RECT 0 195.475 75 200 ;
      RECT 0 175.73 12.225 195.475 ;
      RECT 37.22 190.44 75 195.475 ;
      RECT 61.89 175.06 75 190.44 ;
      RECT 59.685 107.795 75 172.855 ;
      RECT 0 102.035 15.1 172.855 ;
      RECT 0 92.375 23.345 93.79 ;
      RECT 0 0 25.495 90.225 ;
      RECT 32.33 110.785 42.455 170.295 ;
      RECT 32.33 105.025 37.49 105.82 ;
      RECT 49.29 0 75 95.985 ;
      RECT 51.44 98.135 75 99.55 ;
      RECT 51.44 0 75 99.55 ;
      RECT 22.05 168.965 25.53 169.115 ;
      RECT 22.2 169.115 25.53 169.265 ;
      RECT 22.35 169.265 25.53 169.415 ;
      RECT 22.5 169.415 25.53 169.565 ;
      RECT 22.65 169.565 25.53 169.715 ;
      RECT 22.8 169.715 25.53 169.865 ;
      RECT 22.95 169.865 25.53 170.015 ;
      RECT 23.1 170.015 25.53 170.165 ;
      RECT 23.25 170.165 25.53 170.315 ;
      RECT 23.4 170.315 25.53 170.465 ;
      RECT 23.55 170.465 25.53 170.615 ;
      RECT 23.7 170.615 25.53 170.765 ;
      RECT 23.85 170.765 25.53 170.915 ;
      RECT 24.0 170.915 25.53 171.065 ;
      RECT 24.15 171.065 25.53 171.215 ;
      RECT 24.3 171.215 25.53 171.365 ;
      RECT 24.45 171.365 25.53 171.515 ;
      RECT 24.6 171.515 25.53 171.665 ;
      RECT 24.75 171.665 25.53 171.815 ;
      RECT 24.9 171.815 25.53 171.965 ;
      RECT 25.05 171.965 25.53 172.115 ;
      RECT 25.2 172.115 25.53 172.265 ;
      RECT 25.35 172.265 25.53 172.415 ;
      RECT 25.5 172.415 25.53 172.565 ;
      RECT 24.52 102.225 25.53 102.375 ;
      RECT 24.37 102.375 25.53 102.525 ;
      RECT 24.22 102.525 25.53 102.675 ;
      RECT 24.07 102.675 25.53 102.825 ;
      RECT 23.92 102.825 25.53 102.975 ;
      RECT 23.77 102.975 25.53 103.125 ;
      RECT 23.62 103.125 25.53 103.275 ;
      RECT 23.47 103.275 25.53 103.425 ;
      RECT 23.32 103.425 25.53 103.575 ;
      RECT 23.17 103.575 25.53 103.725 ;
      RECT 23.02 103.725 25.53 103.875 ;
      RECT 22.87 103.875 25.53 104.025 ;
      RECT 22.72 104.025 25.53 104.175 ;
      RECT 22.57 104.175 25.53 104.325 ;
      RECT 22.42 104.325 25.53 104.475 ;
      RECT 22.27 104.475 25.53 104.625 ;
      RECT 22.12 104.625 25.53 104.775 ;
      RECT 21.97 104.775 25.53 104.845 ;
      RECT 29.925 96.82 30.785 96.97 ;
      RECT 29.775 96.97 30.635 97.12 ;
      RECT 29.625 97.12 30.485 97.27 ;
      RECT 29.475 97.27 30.335 97.42 ;
      RECT 29.325 97.42 30.185 97.57 ;
      RECT 29.175 97.57 30.035 97.72 ;
      RECT 29.025 97.72 29.885 97.87 ;
      RECT 28.875 97.87 29.735 98.02 ;
      RECT 28.725 98.02 29.585 98.17 ;
      RECT 28.575 98.17 29.435 98.32 ;
      RECT 28.425 98.32 29.285 98.47 ;
      RECT 28.275 98.47 29.135 98.62 ;
      RECT 28.125 98.62 28.985 98.77 ;
      RECT 27.975 98.77 28.835 98.92 ;
      RECT 27.825 98.92 28.685 99.07 ;
      RECT 27.675 99.07 28.535 99.22 ;
      RECT 27.525 99.22 28.385 99.37 ;
      RECT 27.375 99.37 28.235 99.52 ;
      RECT 27.225 99.52 28.085 99.67 ;
      RECT 27.075 99.67 27.935 99.82 ;
      RECT 26.925 99.82 27.785 99.97 ;
      RECT 26.775 99.97 27.635 100.12 ;
      RECT 26.625 100.12 27.485 100.27 ;
      RECT 26.475 100.27 27.335 100.42 ;
      RECT 26.325 100.42 27.185 100.57 ;
      RECT 26.175 100.57 27.035 100.72 ;
      RECT 26.025 100.72 26.885 100.87 ;
      RECT 25.875 100.87 26.735 101.02 ;
      RECT 25.725 101.02 26.585 101.17 ;
      RECT 25.575 101.17 26.435 101.32 ;
      RECT 25.425 101.32 26.285 101.47 ;
      RECT 25.275 101.47 26.135 101.62 ;
      RECT 25.125 101.62 25.985 101.77 ;
      RECT 24.975 101.77 25.835 101.92 ;
      RECT 24.825 101.92 25.685 102.07 ;
      RECT 24.675 102.07 25.535 102.22 ;
      RECT 24.525 102.22 25.53 102.225 ;
      RECT 29.925 96.21 31.395 96.36 ;
      RECT 29.925 96.36 31.245 96.51 ;
      RECT 29.925 96.51 31.095 96.66 ;
      RECT 29.925 96.66 30.945 96.81 ;
      RECT 29.925 96.81 30.935 96.82 ;
      RECT 30.4 92.79 31.07 92.94 ;
      RECT 30.25 92.94 31.22 93.09 ;
      RECT 30.1 93.09 31.37 93.24 ;
      RECT 29.95 93.24 31.52 93.265 ;
      RECT 43.39 101.97 44.95 102.12 ;
      RECT 43.54 102.12 44.95 102.27 ;
      RECT 43.69 102.27 44.95 102.42 ;
      RECT 43.84 102.42 44.95 102.57 ;
      RECT 43.94 102.57 44.95 102.67 ;
      RECT 43.295 100.395 44.95 100.425 ;
      RECT 43.265 100.425 44.95 100.45 ;
      RECT 43.785 99.905 44.46 100.055 ;
      RECT 43.635 100.055 44.61 100.205 ;
      RECT 43.485 100.205 44.76 100.355 ;
      RECT 43.335 100.355 44.91 100.395 ;
      RECT 44.09 102.67 44.95 102.82 ;
      RECT 44.24 102.82 45.1 102.97 ;
    LAYER met1 ;
      RECT 0 0 75 200 ;
    LAYER met5 ;
      RECT 0 0 75 200 ;
    LAYER met4 ;
      RECT 0 0 75 200 ;
  END
END sky130_fd_io__top_hvclamp

END LIBRARY
