/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_IO__TOP_GPIO_OVTV2_BLACKBOX_V
`define SKY130_FD_IO__TOP_GPIO_OVTV2_BLACKBOX_V

/**
 * top_gpio_ovtv2: General Purpose I/0.
 *
 * Verilog stub definition (black box without power pins).
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_io__top_gpio_ovtv2 (
           OUT             ,
           OE_N            ,
           HLD_H_N         ,
           ENABLE_H        ,
           ENABLE_INP_H    ,
           ENABLE_VDDA_H   ,
           ENABLE_VDDIO    ,
           ENABLE_VSWITCH_H,
           INP_DIS         ,
           VTRIP_SEL       ,
           HYS_TRIM        ,
           SLOW            ,
           SLEW_CTL        ,
           HLD_OVR         ,
           ANALOG_EN       ,
           ANALOG_SEL      ,
           ANALOG_POL      ,
           DM              ,
           IB_MODE_SEL     ,
           VINREF          ,
           PAD             ,
           PAD_A_NOESD_H   ,
           PAD_A_ESD_0_H   ,
           PAD_A_ESD_1_H   ,
           AMUXBUS_A       ,
           AMUXBUS_B       ,
           IN              ,
           IN_H            ,
           TIE_HI_ESD      ,
           TIE_LO_ESD
       );

input        OUT             ;
input        OE_N            ;
input        HLD_H_N         ;
input        ENABLE_H        ;
input        ENABLE_INP_H    ;
input        ENABLE_VDDA_H   ;
input        ENABLE_VDDIO    ;
input        ENABLE_VSWITCH_H;
input        INP_DIS         ;
input        VTRIP_SEL       ;
input        HYS_TRIM        ;
input        SLOW            ;
input  [1:0] SLEW_CTL        ;
input        HLD_OVR         ;
input        ANALOG_EN       ;
input        ANALOG_SEL      ;
input        ANALOG_POL      ;
input  [2:0] DM              ;
input  [1:0] IB_MODE_SEL     ;
input        VINREF          ;
inout        PAD             ;
inout        PAD_A_NOESD_H   ;
inout        PAD_A_ESD_0_H   ;
inout        PAD_A_ESD_1_H   ;
inout        AMUXBUS_A       ;
inout        AMUXBUS_B       ;
output       IN              ;
output       IN_H            ;
output       TIE_HI_ESD      ;
output       TIE_LO_ESD      ;

// Voltage supply signals
supply1 VDDIO  ;
supply1 VDDIO_Q;
supply1 VDDA   ;
supply1 VCCD   ;
supply1 VSWITCH;
supply1 VCCHIB ;
supply0 VSSA   ;
supply0 VSSD   ;
supply0 VSSIO_Q;
supply0 VSSIO  ;

endmodule

`default_nettype wire
`endif  // SKY130_FD_IO__TOP_GPIO_OVTV2_BLACKBOX_V
