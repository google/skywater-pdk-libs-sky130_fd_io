# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_io__overlay_vssd_hvc
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 1.270000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 8.885000 75.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 1.270000 13.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 2.035000 75.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 1.270000 7.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 14.935000 75.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 0.965000 18.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 1.270000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 19.785000 75.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 70.035000 75.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 1.270000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 1.270000 94.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 19.885000 75.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 1.270000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 64.085000 75.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 1.270000 68.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 1.270000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 1.270000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 36.735000 75.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 47.735000 75.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.645000 75.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.405000 75.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.840000 1.270000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 1.270000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 36.840000 75.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.970000 41.590000 24.395000 46.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000 41.590000 74.290000 46.230000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 24.370000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.415000 41.585000 75.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 1.270000 46.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
    PORT
      LAYER via3 ;
        RECT  1.060000 41.660000  1.260000 41.860000 ;
        RECT  1.060000 42.090000  1.260000 42.290000 ;
        RECT  1.060000 42.520000  1.260000 42.720000 ;
        RECT  1.060000 42.950000  1.260000 43.150000 ;
        RECT  1.060000 43.380000  1.260000 43.580000 ;
        RECT  1.060000 43.810000  1.260000 44.010000 ;
        RECT  1.060000 44.240000  1.260000 44.440000 ;
        RECT  1.060000 44.670000  1.260000 44.870000 ;
        RECT  1.060000 45.100000  1.260000 45.300000 ;
        RECT  1.060000 45.530000  1.260000 45.730000 ;
        RECT  1.060000 45.960000  1.260000 46.160000 ;
        RECT  1.465000 41.660000  1.665000 41.860000 ;
        RECT  1.465000 42.090000  1.665000 42.290000 ;
        RECT  1.465000 42.520000  1.665000 42.720000 ;
        RECT  1.465000 42.950000  1.665000 43.150000 ;
        RECT  1.465000 43.380000  1.665000 43.580000 ;
        RECT  1.465000 43.810000  1.665000 44.010000 ;
        RECT  1.465000 44.240000  1.665000 44.440000 ;
        RECT  1.465000 44.670000  1.665000 44.870000 ;
        RECT  1.465000 45.100000  1.665000 45.300000 ;
        RECT  1.465000 45.530000  1.665000 45.730000 ;
        RECT  1.465000 45.960000  1.665000 46.160000 ;
        RECT  1.870000 41.660000  2.070000 41.860000 ;
        RECT  1.870000 42.090000  2.070000 42.290000 ;
        RECT  1.870000 42.520000  2.070000 42.720000 ;
        RECT  1.870000 42.950000  2.070000 43.150000 ;
        RECT  1.870000 43.380000  2.070000 43.580000 ;
        RECT  1.870000 43.810000  2.070000 44.010000 ;
        RECT  1.870000 44.240000  2.070000 44.440000 ;
        RECT  1.870000 44.670000  2.070000 44.870000 ;
        RECT  1.870000 45.100000  2.070000 45.300000 ;
        RECT  1.870000 45.530000  2.070000 45.730000 ;
        RECT  1.870000 45.960000  2.070000 46.160000 ;
        RECT  2.275000 41.660000  2.475000 41.860000 ;
        RECT  2.275000 42.090000  2.475000 42.290000 ;
        RECT  2.275000 42.520000  2.475000 42.720000 ;
        RECT  2.275000 42.950000  2.475000 43.150000 ;
        RECT  2.275000 43.380000  2.475000 43.580000 ;
        RECT  2.275000 43.810000  2.475000 44.010000 ;
        RECT  2.275000 44.240000  2.475000 44.440000 ;
        RECT  2.275000 44.670000  2.475000 44.870000 ;
        RECT  2.275000 45.100000  2.475000 45.300000 ;
        RECT  2.275000 45.530000  2.475000 45.730000 ;
        RECT  2.275000 45.960000  2.475000 46.160000 ;
        RECT  2.680000 41.660000  2.880000 41.860000 ;
        RECT  2.680000 42.090000  2.880000 42.290000 ;
        RECT  2.680000 42.520000  2.880000 42.720000 ;
        RECT  2.680000 42.950000  2.880000 43.150000 ;
        RECT  2.680000 43.380000  2.880000 43.580000 ;
        RECT  2.680000 43.810000  2.880000 44.010000 ;
        RECT  2.680000 44.240000  2.880000 44.440000 ;
        RECT  2.680000 44.670000  2.880000 44.870000 ;
        RECT  2.680000 45.100000  2.880000 45.300000 ;
        RECT  2.680000 45.530000  2.880000 45.730000 ;
        RECT  2.680000 45.960000  2.880000 46.160000 ;
        RECT  3.085000 41.660000  3.285000 41.860000 ;
        RECT  3.085000 42.090000  3.285000 42.290000 ;
        RECT  3.085000 42.520000  3.285000 42.720000 ;
        RECT  3.085000 42.950000  3.285000 43.150000 ;
        RECT  3.085000 43.380000  3.285000 43.580000 ;
        RECT  3.085000 43.810000  3.285000 44.010000 ;
        RECT  3.085000 44.240000  3.285000 44.440000 ;
        RECT  3.085000 44.670000  3.285000 44.870000 ;
        RECT  3.085000 45.100000  3.285000 45.300000 ;
        RECT  3.085000 45.530000  3.285000 45.730000 ;
        RECT  3.085000 45.960000  3.285000 46.160000 ;
        RECT  3.490000 41.660000  3.690000 41.860000 ;
        RECT  3.490000 42.090000  3.690000 42.290000 ;
        RECT  3.490000 42.520000  3.690000 42.720000 ;
        RECT  3.490000 42.950000  3.690000 43.150000 ;
        RECT  3.490000 43.380000  3.690000 43.580000 ;
        RECT  3.490000 43.810000  3.690000 44.010000 ;
        RECT  3.490000 44.240000  3.690000 44.440000 ;
        RECT  3.490000 44.670000  3.690000 44.870000 ;
        RECT  3.490000 45.100000  3.690000 45.300000 ;
        RECT  3.490000 45.530000  3.690000 45.730000 ;
        RECT  3.490000 45.960000  3.690000 46.160000 ;
        RECT  3.895000 41.660000  4.095000 41.860000 ;
        RECT  3.895000 42.090000  4.095000 42.290000 ;
        RECT  3.895000 42.520000  4.095000 42.720000 ;
        RECT  3.895000 42.950000  4.095000 43.150000 ;
        RECT  3.895000 43.380000  4.095000 43.580000 ;
        RECT  3.895000 43.810000  4.095000 44.010000 ;
        RECT  3.895000 44.240000  4.095000 44.440000 ;
        RECT  3.895000 44.670000  4.095000 44.870000 ;
        RECT  3.895000 45.100000  4.095000 45.300000 ;
        RECT  3.895000 45.530000  4.095000 45.730000 ;
        RECT  3.895000 45.960000  4.095000 46.160000 ;
        RECT  4.300000 41.660000  4.500000 41.860000 ;
        RECT  4.300000 42.090000  4.500000 42.290000 ;
        RECT  4.300000 42.520000  4.500000 42.720000 ;
        RECT  4.300000 42.950000  4.500000 43.150000 ;
        RECT  4.300000 43.380000  4.500000 43.580000 ;
        RECT  4.300000 43.810000  4.500000 44.010000 ;
        RECT  4.300000 44.240000  4.500000 44.440000 ;
        RECT  4.300000 44.670000  4.500000 44.870000 ;
        RECT  4.300000 45.100000  4.500000 45.300000 ;
        RECT  4.300000 45.530000  4.500000 45.730000 ;
        RECT  4.300000 45.960000  4.500000 46.160000 ;
        RECT  4.705000 41.660000  4.905000 41.860000 ;
        RECT  4.705000 42.090000  4.905000 42.290000 ;
        RECT  4.705000 42.520000  4.905000 42.720000 ;
        RECT  4.705000 42.950000  4.905000 43.150000 ;
        RECT  4.705000 43.380000  4.905000 43.580000 ;
        RECT  4.705000 43.810000  4.905000 44.010000 ;
        RECT  4.705000 44.240000  4.905000 44.440000 ;
        RECT  4.705000 44.670000  4.905000 44.870000 ;
        RECT  4.705000 45.100000  4.905000 45.300000 ;
        RECT  4.705000 45.530000  4.905000 45.730000 ;
        RECT  4.705000 45.960000  4.905000 46.160000 ;
        RECT  5.110000 41.660000  5.310000 41.860000 ;
        RECT  5.110000 42.090000  5.310000 42.290000 ;
        RECT  5.110000 42.520000  5.310000 42.720000 ;
        RECT  5.110000 42.950000  5.310000 43.150000 ;
        RECT  5.110000 43.380000  5.310000 43.580000 ;
        RECT  5.110000 43.810000  5.310000 44.010000 ;
        RECT  5.110000 44.240000  5.310000 44.440000 ;
        RECT  5.110000 44.670000  5.310000 44.870000 ;
        RECT  5.110000 45.100000  5.310000 45.300000 ;
        RECT  5.110000 45.530000  5.310000 45.730000 ;
        RECT  5.110000 45.960000  5.310000 46.160000 ;
        RECT  5.515000 41.660000  5.715000 41.860000 ;
        RECT  5.515000 42.090000  5.715000 42.290000 ;
        RECT  5.515000 42.520000  5.715000 42.720000 ;
        RECT  5.515000 42.950000  5.715000 43.150000 ;
        RECT  5.515000 43.380000  5.715000 43.580000 ;
        RECT  5.515000 43.810000  5.715000 44.010000 ;
        RECT  5.515000 44.240000  5.715000 44.440000 ;
        RECT  5.515000 44.670000  5.715000 44.870000 ;
        RECT  5.515000 45.100000  5.715000 45.300000 ;
        RECT  5.515000 45.530000  5.715000 45.730000 ;
        RECT  5.515000 45.960000  5.715000 46.160000 ;
        RECT  5.920000 41.660000  6.120000 41.860000 ;
        RECT  5.920000 42.090000  6.120000 42.290000 ;
        RECT  5.920000 42.520000  6.120000 42.720000 ;
        RECT  5.920000 42.950000  6.120000 43.150000 ;
        RECT  5.920000 43.380000  6.120000 43.580000 ;
        RECT  5.920000 43.810000  6.120000 44.010000 ;
        RECT  5.920000 44.240000  6.120000 44.440000 ;
        RECT  5.920000 44.670000  6.120000 44.870000 ;
        RECT  5.920000 45.100000  6.120000 45.300000 ;
        RECT  5.920000 45.530000  6.120000 45.730000 ;
        RECT  5.920000 45.960000  6.120000 46.160000 ;
        RECT  6.325000 41.660000  6.525000 41.860000 ;
        RECT  6.325000 42.090000  6.525000 42.290000 ;
        RECT  6.325000 42.520000  6.525000 42.720000 ;
        RECT  6.325000 42.950000  6.525000 43.150000 ;
        RECT  6.325000 43.380000  6.525000 43.580000 ;
        RECT  6.325000 43.810000  6.525000 44.010000 ;
        RECT  6.325000 44.240000  6.525000 44.440000 ;
        RECT  6.325000 44.670000  6.525000 44.870000 ;
        RECT  6.325000 45.100000  6.525000 45.300000 ;
        RECT  6.325000 45.530000  6.525000 45.730000 ;
        RECT  6.325000 45.960000  6.525000 46.160000 ;
        RECT  6.730000 41.660000  6.930000 41.860000 ;
        RECT  6.730000 42.090000  6.930000 42.290000 ;
        RECT  6.730000 42.520000  6.930000 42.720000 ;
        RECT  6.730000 42.950000  6.930000 43.150000 ;
        RECT  6.730000 43.380000  6.930000 43.580000 ;
        RECT  6.730000 43.810000  6.930000 44.010000 ;
        RECT  6.730000 44.240000  6.930000 44.440000 ;
        RECT  6.730000 44.670000  6.930000 44.870000 ;
        RECT  6.730000 45.100000  6.930000 45.300000 ;
        RECT  6.730000 45.530000  6.930000 45.730000 ;
        RECT  6.730000 45.960000  6.930000 46.160000 ;
        RECT  7.135000 41.660000  7.335000 41.860000 ;
        RECT  7.135000 42.090000  7.335000 42.290000 ;
        RECT  7.135000 42.520000  7.335000 42.720000 ;
        RECT  7.135000 42.950000  7.335000 43.150000 ;
        RECT  7.135000 43.380000  7.335000 43.580000 ;
        RECT  7.135000 43.810000  7.335000 44.010000 ;
        RECT  7.135000 44.240000  7.335000 44.440000 ;
        RECT  7.135000 44.670000  7.335000 44.870000 ;
        RECT  7.135000 45.100000  7.335000 45.300000 ;
        RECT  7.135000 45.530000  7.335000 45.730000 ;
        RECT  7.135000 45.960000  7.335000 46.160000 ;
        RECT  7.540000 41.660000  7.740000 41.860000 ;
        RECT  7.540000 42.090000  7.740000 42.290000 ;
        RECT  7.540000 42.520000  7.740000 42.720000 ;
        RECT  7.540000 42.950000  7.740000 43.150000 ;
        RECT  7.540000 43.380000  7.740000 43.580000 ;
        RECT  7.540000 43.810000  7.740000 44.010000 ;
        RECT  7.540000 44.240000  7.740000 44.440000 ;
        RECT  7.540000 44.670000  7.740000 44.870000 ;
        RECT  7.540000 45.100000  7.740000 45.300000 ;
        RECT  7.540000 45.530000  7.740000 45.730000 ;
        RECT  7.540000 45.960000  7.740000 46.160000 ;
        RECT  7.945000 41.660000  8.145000 41.860000 ;
        RECT  7.945000 42.090000  8.145000 42.290000 ;
        RECT  7.945000 42.520000  8.145000 42.720000 ;
        RECT  7.945000 42.950000  8.145000 43.150000 ;
        RECT  7.945000 43.380000  8.145000 43.580000 ;
        RECT  7.945000 43.810000  8.145000 44.010000 ;
        RECT  7.945000 44.240000  8.145000 44.440000 ;
        RECT  7.945000 44.670000  8.145000 44.870000 ;
        RECT  7.945000 45.100000  8.145000 45.300000 ;
        RECT  7.945000 45.530000  8.145000 45.730000 ;
        RECT  7.945000 45.960000  8.145000 46.160000 ;
        RECT  8.350000 41.660000  8.550000 41.860000 ;
        RECT  8.350000 42.090000  8.550000 42.290000 ;
        RECT  8.350000 42.520000  8.550000 42.720000 ;
        RECT  8.350000 42.950000  8.550000 43.150000 ;
        RECT  8.350000 43.380000  8.550000 43.580000 ;
        RECT  8.350000 43.810000  8.550000 44.010000 ;
        RECT  8.350000 44.240000  8.550000 44.440000 ;
        RECT  8.350000 44.670000  8.550000 44.870000 ;
        RECT  8.350000 45.100000  8.550000 45.300000 ;
        RECT  8.350000 45.530000  8.550000 45.730000 ;
        RECT  8.350000 45.960000  8.550000 46.160000 ;
        RECT  8.755000 41.660000  8.955000 41.860000 ;
        RECT  8.755000 42.090000  8.955000 42.290000 ;
        RECT  8.755000 42.520000  8.955000 42.720000 ;
        RECT  8.755000 42.950000  8.955000 43.150000 ;
        RECT  8.755000 43.380000  8.955000 43.580000 ;
        RECT  8.755000 43.810000  8.955000 44.010000 ;
        RECT  8.755000 44.240000  8.955000 44.440000 ;
        RECT  8.755000 44.670000  8.955000 44.870000 ;
        RECT  8.755000 45.100000  8.955000 45.300000 ;
        RECT  8.755000 45.530000  8.955000 45.730000 ;
        RECT  8.755000 45.960000  8.955000 46.160000 ;
        RECT  9.160000 41.660000  9.360000 41.860000 ;
        RECT  9.160000 42.090000  9.360000 42.290000 ;
        RECT  9.160000 42.520000  9.360000 42.720000 ;
        RECT  9.160000 42.950000  9.360000 43.150000 ;
        RECT  9.160000 43.380000  9.360000 43.580000 ;
        RECT  9.160000 43.810000  9.360000 44.010000 ;
        RECT  9.160000 44.240000  9.360000 44.440000 ;
        RECT  9.160000 44.670000  9.360000 44.870000 ;
        RECT  9.160000 45.100000  9.360000 45.300000 ;
        RECT  9.160000 45.530000  9.360000 45.730000 ;
        RECT  9.160000 45.960000  9.360000 46.160000 ;
        RECT  9.565000 41.660000  9.765000 41.860000 ;
        RECT  9.565000 42.090000  9.765000 42.290000 ;
        RECT  9.565000 42.520000  9.765000 42.720000 ;
        RECT  9.565000 42.950000  9.765000 43.150000 ;
        RECT  9.565000 43.380000  9.765000 43.580000 ;
        RECT  9.565000 43.810000  9.765000 44.010000 ;
        RECT  9.565000 44.240000  9.765000 44.440000 ;
        RECT  9.565000 44.670000  9.765000 44.870000 ;
        RECT  9.565000 45.100000  9.765000 45.300000 ;
        RECT  9.565000 45.530000  9.765000 45.730000 ;
        RECT  9.565000 45.960000  9.765000 46.160000 ;
        RECT  9.970000 41.660000 10.170000 41.860000 ;
        RECT  9.970000 42.090000 10.170000 42.290000 ;
        RECT  9.970000 42.520000 10.170000 42.720000 ;
        RECT  9.970000 42.950000 10.170000 43.150000 ;
        RECT  9.970000 43.380000 10.170000 43.580000 ;
        RECT  9.970000 43.810000 10.170000 44.010000 ;
        RECT  9.970000 44.240000 10.170000 44.440000 ;
        RECT  9.970000 44.670000 10.170000 44.870000 ;
        RECT  9.970000 45.100000 10.170000 45.300000 ;
        RECT  9.970000 45.530000 10.170000 45.730000 ;
        RECT  9.970000 45.960000 10.170000 46.160000 ;
        RECT 10.375000 41.660000 10.575000 41.860000 ;
        RECT 10.375000 42.090000 10.575000 42.290000 ;
        RECT 10.375000 42.520000 10.575000 42.720000 ;
        RECT 10.375000 42.950000 10.575000 43.150000 ;
        RECT 10.375000 43.380000 10.575000 43.580000 ;
        RECT 10.375000 43.810000 10.575000 44.010000 ;
        RECT 10.375000 44.240000 10.575000 44.440000 ;
        RECT 10.375000 44.670000 10.575000 44.870000 ;
        RECT 10.375000 45.100000 10.575000 45.300000 ;
        RECT 10.375000 45.530000 10.575000 45.730000 ;
        RECT 10.375000 45.960000 10.575000 46.160000 ;
        RECT 10.780000 41.660000 10.980000 41.860000 ;
        RECT 10.780000 42.090000 10.980000 42.290000 ;
        RECT 10.780000 42.520000 10.980000 42.720000 ;
        RECT 10.780000 42.950000 10.980000 43.150000 ;
        RECT 10.780000 43.380000 10.980000 43.580000 ;
        RECT 10.780000 43.810000 10.980000 44.010000 ;
        RECT 10.780000 44.240000 10.980000 44.440000 ;
        RECT 10.780000 44.670000 10.980000 44.870000 ;
        RECT 10.780000 45.100000 10.980000 45.300000 ;
        RECT 10.780000 45.530000 10.980000 45.730000 ;
        RECT 10.780000 45.960000 10.980000 46.160000 ;
        RECT 11.185000 41.660000 11.385000 41.860000 ;
        RECT 11.185000 42.090000 11.385000 42.290000 ;
        RECT 11.185000 42.520000 11.385000 42.720000 ;
        RECT 11.185000 42.950000 11.385000 43.150000 ;
        RECT 11.185000 43.380000 11.385000 43.580000 ;
        RECT 11.185000 43.810000 11.385000 44.010000 ;
        RECT 11.185000 44.240000 11.385000 44.440000 ;
        RECT 11.185000 44.670000 11.385000 44.870000 ;
        RECT 11.185000 45.100000 11.385000 45.300000 ;
        RECT 11.185000 45.530000 11.385000 45.730000 ;
        RECT 11.185000 45.960000 11.385000 46.160000 ;
        RECT 11.590000 41.660000 11.790000 41.860000 ;
        RECT 11.590000 42.090000 11.790000 42.290000 ;
        RECT 11.590000 42.520000 11.790000 42.720000 ;
        RECT 11.590000 42.950000 11.790000 43.150000 ;
        RECT 11.590000 43.380000 11.790000 43.580000 ;
        RECT 11.590000 43.810000 11.790000 44.010000 ;
        RECT 11.590000 44.240000 11.790000 44.440000 ;
        RECT 11.590000 44.670000 11.790000 44.870000 ;
        RECT 11.590000 45.100000 11.790000 45.300000 ;
        RECT 11.590000 45.530000 11.790000 45.730000 ;
        RECT 11.590000 45.960000 11.790000 46.160000 ;
        RECT 11.995000 41.660000 12.195000 41.860000 ;
        RECT 11.995000 42.090000 12.195000 42.290000 ;
        RECT 11.995000 42.520000 12.195000 42.720000 ;
        RECT 11.995000 42.950000 12.195000 43.150000 ;
        RECT 11.995000 43.380000 12.195000 43.580000 ;
        RECT 11.995000 43.810000 12.195000 44.010000 ;
        RECT 11.995000 44.240000 12.195000 44.440000 ;
        RECT 11.995000 44.670000 12.195000 44.870000 ;
        RECT 11.995000 45.100000 12.195000 45.300000 ;
        RECT 11.995000 45.530000 12.195000 45.730000 ;
        RECT 11.995000 45.960000 12.195000 46.160000 ;
        RECT 12.400000 41.660000 12.600000 41.860000 ;
        RECT 12.400000 42.090000 12.600000 42.290000 ;
        RECT 12.400000 42.520000 12.600000 42.720000 ;
        RECT 12.400000 42.950000 12.600000 43.150000 ;
        RECT 12.400000 43.380000 12.600000 43.580000 ;
        RECT 12.400000 43.810000 12.600000 44.010000 ;
        RECT 12.400000 44.240000 12.600000 44.440000 ;
        RECT 12.400000 44.670000 12.600000 44.870000 ;
        RECT 12.400000 45.100000 12.600000 45.300000 ;
        RECT 12.400000 45.530000 12.600000 45.730000 ;
        RECT 12.400000 45.960000 12.600000 46.160000 ;
        RECT 12.805000 41.660000 13.005000 41.860000 ;
        RECT 12.805000 42.090000 13.005000 42.290000 ;
        RECT 12.805000 42.520000 13.005000 42.720000 ;
        RECT 12.805000 42.950000 13.005000 43.150000 ;
        RECT 12.805000 43.380000 13.005000 43.580000 ;
        RECT 12.805000 43.810000 13.005000 44.010000 ;
        RECT 12.805000 44.240000 13.005000 44.440000 ;
        RECT 12.805000 44.670000 13.005000 44.870000 ;
        RECT 12.805000 45.100000 13.005000 45.300000 ;
        RECT 12.805000 45.530000 13.005000 45.730000 ;
        RECT 12.805000 45.960000 13.005000 46.160000 ;
        RECT 13.210000 41.660000 13.410000 41.860000 ;
        RECT 13.210000 42.090000 13.410000 42.290000 ;
        RECT 13.210000 42.520000 13.410000 42.720000 ;
        RECT 13.210000 42.950000 13.410000 43.150000 ;
        RECT 13.210000 43.380000 13.410000 43.580000 ;
        RECT 13.210000 43.810000 13.410000 44.010000 ;
        RECT 13.210000 44.240000 13.410000 44.440000 ;
        RECT 13.210000 44.670000 13.410000 44.870000 ;
        RECT 13.210000 45.100000 13.410000 45.300000 ;
        RECT 13.210000 45.530000 13.410000 45.730000 ;
        RECT 13.210000 45.960000 13.410000 46.160000 ;
        RECT 13.615000 41.660000 13.815000 41.860000 ;
        RECT 13.615000 42.090000 13.815000 42.290000 ;
        RECT 13.615000 42.520000 13.815000 42.720000 ;
        RECT 13.615000 42.950000 13.815000 43.150000 ;
        RECT 13.615000 43.380000 13.815000 43.580000 ;
        RECT 13.615000 43.810000 13.815000 44.010000 ;
        RECT 13.615000 44.240000 13.815000 44.440000 ;
        RECT 13.615000 44.670000 13.815000 44.870000 ;
        RECT 13.615000 45.100000 13.815000 45.300000 ;
        RECT 13.615000 45.530000 13.815000 45.730000 ;
        RECT 13.615000 45.960000 13.815000 46.160000 ;
        RECT 14.020000 41.660000 14.220000 41.860000 ;
        RECT 14.020000 42.090000 14.220000 42.290000 ;
        RECT 14.020000 42.520000 14.220000 42.720000 ;
        RECT 14.020000 42.950000 14.220000 43.150000 ;
        RECT 14.020000 43.380000 14.220000 43.580000 ;
        RECT 14.020000 43.810000 14.220000 44.010000 ;
        RECT 14.020000 44.240000 14.220000 44.440000 ;
        RECT 14.020000 44.670000 14.220000 44.870000 ;
        RECT 14.020000 45.100000 14.220000 45.300000 ;
        RECT 14.020000 45.530000 14.220000 45.730000 ;
        RECT 14.020000 45.960000 14.220000 46.160000 ;
        RECT 14.425000 41.660000 14.625000 41.860000 ;
        RECT 14.425000 42.090000 14.625000 42.290000 ;
        RECT 14.425000 42.520000 14.625000 42.720000 ;
        RECT 14.425000 42.950000 14.625000 43.150000 ;
        RECT 14.425000 43.380000 14.625000 43.580000 ;
        RECT 14.425000 43.810000 14.625000 44.010000 ;
        RECT 14.425000 44.240000 14.625000 44.440000 ;
        RECT 14.425000 44.670000 14.625000 44.870000 ;
        RECT 14.425000 45.100000 14.625000 45.300000 ;
        RECT 14.425000 45.530000 14.625000 45.730000 ;
        RECT 14.425000 45.960000 14.625000 46.160000 ;
        RECT 14.830000 41.660000 15.030000 41.860000 ;
        RECT 14.830000 42.090000 15.030000 42.290000 ;
        RECT 14.830000 42.520000 15.030000 42.720000 ;
        RECT 14.830000 42.950000 15.030000 43.150000 ;
        RECT 14.830000 43.380000 15.030000 43.580000 ;
        RECT 14.830000 43.810000 15.030000 44.010000 ;
        RECT 14.830000 44.240000 15.030000 44.440000 ;
        RECT 14.830000 44.670000 15.030000 44.870000 ;
        RECT 14.830000 45.100000 15.030000 45.300000 ;
        RECT 14.830000 45.530000 15.030000 45.730000 ;
        RECT 14.830000 45.960000 15.030000 46.160000 ;
        RECT 15.235000 41.660000 15.435000 41.860000 ;
        RECT 15.235000 42.090000 15.435000 42.290000 ;
        RECT 15.235000 42.520000 15.435000 42.720000 ;
        RECT 15.235000 42.950000 15.435000 43.150000 ;
        RECT 15.235000 43.380000 15.435000 43.580000 ;
        RECT 15.235000 43.810000 15.435000 44.010000 ;
        RECT 15.235000 44.240000 15.435000 44.440000 ;
        RECT 15.235000 44.670000 15.435000 44.870000 ;
        RECT 15.235000 45.100000 15.435000 45.300000 ;
        RECT 15.235000 45.530000 15.435000 45.730000 ;
        RECT 15.235000 45.960000 15.435000 46.160000 ;
        RECT 15.640000 41.660000 15.840000 41.860000 ;
        RECT 15.640000 42.090000 15.840000 42.290000 ;
        RECT 15.640000 42.520000 15.840000 42.720000 ;
        RECT 15.640000 42.950000 15.840000 43.150000 ;
        RECT 15.640000 43.380000 15.840000 43.580000 ;
        RECT 15.640000 43.810000 15.840000 44.010000 ;
        RECT 15.640000 44.240000 15.840000 44.440000 ;
        RECT 15.640000 44.670000 15.840000 44.870000 ;
        RECT 15.640000 45.100000 15.840000 45.300000 ;
        RECT 15.640000 45.530000 15.840000 45.730000 ;
        RECT 15.640000 45.960000 15.840000 46.160000 ;
        RECT 16.045000 41.660000 16.245000 41.860000 ;
        RECT 16.045000 42.090000 16.245000 42.290000 ;
        RECT 16.045000 42.520000 16.245000 42.720000 ;
        RECT 16.045000 42.950000 16.245000 43.150000 ;
        RECT 16.045000 43.380000 16.245000 43.580000 ;
        RECT 16.045000 43.810000 16.245000 44.010000 ;
        RECT 16.045000 44.240000 16.245000 44.440000 ;
        RECT 16.045000 44.670000 16.245000 44.870000 ;
        RECT 16.045000 45.100000 16.245000 45.300000 ;
        RECT 16.045000 45.530000 16.245000 45.730000 ;
        RECT 16.045000 45.960000 16.245000 46.160000 ;
        RECT 16.450000 41.660000 16.650000 41.860000 ;
        RECT 16.450000 42.090000 16.650000 42.290000 ;
        RECT 16.450000 42.520000 16.650000 42.720000 ;
        RECT 16.450000 42.950000 16.650000 43.150000 ;
        RECT 16.450000 43.380000 16.650000 43.580000 ;
        RECT 16.450000 43.810000 16.650000 44.010000 ;
        RECT 16.450000 44.240000 16.650000 44.440000 ;
        RECT 16.450000 44.670000 16.650000 44.870000 ;
        RECT 16.450000 45.100000 16.650000 45.300000 ;
        RECT 16.450000 45.530000 16.650000 45.730000 ;
        RECT 16.450000 45.960000 16.650000 46.160000 ;
        RECT 16.855000 41.660000 17.055000 41.860000 ;
        RECT 16.855000 42.090000 17.055000 42.290000 ;
        RECT 16.855000 42.520000 17.055000 42.720000 ;
        RECT 16.855000 42.950000 17.055000 43.150000 ;
        RECT 16.855000 43.380000 17.055000 43.580000 ;
        RECT 16.855000 43.810000 17.055000 44.010000 ;
        RECT 16.855000 44.240000 17.055000 44.440000 ;
        RECT 16.855000 44.670000 17.055000 44.870000 ;
        RECT 16.855000 45.100000 17.055000 45.300000 ;
        RECT 16.855000 45.530000 17.055000 45.730000 ;
        RECT 16.855000 45.960000 17.055000 46.160000 ;
        RECT 17.260000 41.660000 17.460000 41.860000 ;
        RECT 17.260000 42.090000 17.460000 42.290000 ;
        RECT 17.260000 42.520000 17.460000 42.720000 ;
        RECT 17.260000 42.950000 17.460000 43.150000 ;
        RECT 17.260000 43.380000 17.460000 43.580000 ;
        RECT 17.260000 43.810000 17.460000 44.010000 ;
        RECT 17.260000 44.240000 17.460000 44.440000 ;
        RECT 17.260000 44.670000 17.460000 44.870000 ;
        RECT 17.260000 45.100000 17.460000 45.300000 ;
        RECT 17.260000 45.530000 17.460000 45.730000 ;
        RECT 17.260000 45.960000 17.460000 46.160000 ;
        RECT 17.665000 41.660000 17.865000 41.860000 ;
        RECT 17.665000 42.090000 17.865000 42.290000 ;
        RECT 17.665000 42.520000 17.865000 42.720000 ;
        RECT 17.665000 42.950000 17.865000 43.150000 ;
        RECT 17.665000 43.380000 17.865000 43.580000 ;
        RECT 17.665000 43.810000 17.865000 44.010000 ;
        RECT 17.665000 44.240000 17.865000 44.440000 ;
        RECT 17.665000 44.670000 17.865000 44.870000 ;
        RECT 17.665000 45.100000 17.865000 45.300000 ;
        RECT 17.665000 45.530000 17.865000 45.730000 ;
        RECT 17.665000 45.960000 17.865000 46.160000 ;
        RECT 18.070000 41.660000 18.270000 41.860000 ;
        RECT 18.070000 42.090000 18.270000 42.290000 ;
        RECT 18.070000 42.520000 18.270000 42.720000 ;
        RECT 18.070000 42.950000 18.270000 43.150000 ;
        RECT 18.070000 43.380000 18.270000 43.580000 ;
        RECT 18.070000 43.810000 18.270000 44.010000 ;
        RECT 18.070000 44.240000 18.270000 44.440000 ;
        RECT 18.070000 44.670000 18.270000 44.870000 ;
        RECT 18.070000 45.100000 18.270000 45.300000 ;
        RECT 18.070000 45.530000 18.270000 45.730000 ;
        RECT 18.070000 45.960000 18.270000 46.160000 ;
        RECT 18.475000 41.660000 18.675000 41.860000 ;
        RECT 18.475000 42.090000 18.675000 42.290000 ;
        RECT 18.475000 42.520000 18.675000 42.720000 ;
        RECT 18.475000 42.950000 18.675000 43.150000 ;
        RECT 18.475000 43.380000 18.675000 43.580000 ;
        RECT 18.475000 43.810000 18.675000 44.010000 ;
        RECT 18.475000 44.240000 18.675000 44.440000 ;
        RECT 18.475000 44.670000 18.675000 44.870000 ;
        RECT 18.475000 45.100000 18.675000 45.300000 ;
        RECT 18.475000 45.530000 18.675000 45.730000 ;
        RECT 18.475000 45.960000 18.675000 46.160000 ;
        RECT 18.880000 41.660000 19.080000 41.860000 ;
        RECT 18.880000 42.090000 19.080000 42.290000 ;
        RECT 18.880000 42.520000 19.080000 42.720000 ;
        RECT 18.880000 42.950000 19.080000 43.150000 ;
        RECT 18.880000 43.380000 19.080000 43.580000 ;
        RECT 18.880000 43.810000 19.080000 44.010000 ;
        RECT 18.880000 44.240000 19.080000 44.440000 ;
        RECT 18.880000 44.670000 19.080000 44.870000 ;
        RECT 18.880000 45.100000 19.080000 45.300000 ;
        RECT 18.880000 45.530000 19.080000 45.730000 ;
        RECT 18.880000 45.960000 19.080000 46.160000 ;
        RECT 19.285000 41.660000 19.485000 41.860000 ;
        RECT 19.285000 42.090000 19.485000 42.290000 ;
        RECT 19.285000 42.520000 19.485000 42.720000 ;
        RECT 19.285000 42.950000 19.485000 43.150000 ;
        RECT 19.285000 43.380000 19.485000 43.580000 ;
        RECT 19.285000 43.810000 19.485000 44.010000 ;
        RECT 19.285000 44.240000 19.485000 44.440000 ;
        RECT 19.285000 44.670000 19.485000 44.870000 ;
        RECT 19.285000 45.100000 19.485000 45.300000 ;
        RECT 19.285000 45.530000 19.485000 45.730000 ;
        RECT 19.285000 45.960000 19.485000 46.160000 ;
        RECT 19.690000 41.660000 19.890000 41.860000 ;
        RECT 19.690000 42.090000 19.890000 42.290000 ;
        RECT 19.690000 42.520000 19.890000 42.720000 ;
        RECT 19.690000 42.950000 19.890000 43.150000 ;
        RECT 19.690000 43.380000 19.890000 43.580000 ;
        RECT 19.690000 43.810000 19.890000 44.010000 ;
        RECT 19.690000 44.240000 19.890000 44.440000 ;
        RECT 19.690000 44.670000 19.890000 44.870000 ;
        RECT 19.690000 45.100000 19.890000 45.300000 ;
        RECT 19.690000 45.530000 19.890000 45.730000 ;
        RECT 19.690000 45.960000 19.890000 46.160000 ;
        RECT 20.095000 41.660000 20.295000 41.860000 ;
        RECT 20.095000 42.090000 20.295000 42.290000 ;
        RECT 20.095000 42.520000 20.295000 42.720000 ;
        RECT 20.095000 42.950000 20.295000 43.150000 ;
        RECT 20.095000 43.380000 20.295000 43.580000 ;
        RECT 20.095000 43.810000 20.295000 44.010000 ;
        RECT 20.095000 44.240000 20.295000 44.440000 ;
        RECT 20.095000 44.670000 20.295000 44.870000 ;
        RECT 20.095000 45.100000 20.295000 45.300000 ;
        RECT 20.095000 45.530000 20.295000 45.730000 ;
        RECT 20.095000 45.960000 20.295000 46.160000 ;
        RECT 20.500000 41.660000 20.700000 41.860000 ;
        RECT 20.500000 42.090000 20.700000 42.290000 ;
        RECT 20.500000 42.520000 20.700000 42.720000 ;
        RECT 20.500000 42.950000 20.700000 43.150000 ;
        RECT 20.500000 43.380000 20.700000 43.580000 ;
        RECT 20.500000 43.810000 20.700000 44.010000 ;
        RECT 20.500000 44.240000 20.700000 44.440000 ;
        RECT 20.500000 44.670000 20.700000 44.870000 ;
        RECT 20.500000 45.100000 20.700000 45.300000 ;
        RECT 20.500000 45.530000 20.700000 45.730000 ;
        RECT 20.500000 45.960000 20.700000 46.160000 ;
        RECT 20.905000 41.660000 21.105000 41.860000 ;
        RECT 20.905000 42.090000 21.105000 42.290000 ;
        RECT 20.905000 42.520000 21.105000 42.720000 ;
        RECT 20.905000 42.950000 21.105000 43.150000 ;
        RECT 20.905000 43.380000 21.105000 43.580000 ;
        RECT 20.905000 43.810000 21.105000 44.010000 ;
        RECT 20.905000 44.240000 21.105000 44.440000 ;
        RECT 20.905000 44.670000 21.105000 44.870000 ;
        RECT 20.905000 45.100000 21.105000 45.300000 ;
        RECT 20.905000 45.530000 21.105000 45.730000 ;
        RECT 20.905000 45.960000 21.105000 46.160000 ;
        RECT 21.305000 41.660000 21.505000 41.860000 ;
        RECT 21.305000 42.090000 21.505000 42.290000 ;
        RECT 21.305000 42.520000 21.505000 42.720000 ;
        RECT 21.305000 42.950000 21.505000 43.150000 ;
        RECT 21.305000 43.380000 21.505000 43.580000 ;
        RECT 21.305000 43.810000 21.505000 44.010000 ;
        RECT 21.305000 44.240000 21.505000 44.440000 ;
        RECT 21.305000 44.670000 21.505000 44.870000 ;
        RECT 21.305000 45.100000 21.505000 45.300000 ;
        RECT 21.305000 45.530000 21.505000 45.730000 ;
        RECT 21.305000 45.960000 21.505000 46.160000 ;
        RECT 21.705000 41.660000 21.905000 41.860000 ;
        RECT 21.705000 42.090000 21.905000 42.290000 ;
        RECT 21.705000 42.520000 21.905000 42.720000 ;
        RECT 21.705000 42.950000 21.905000 43.150000 ;
        RECT 21.705000 43.380000 21.905000 43.580000 ;
        RECT 21.705000 43.810000 21.905000 44.010000 ;
        RECT 21.705000 44.240000 21.905000 44.440000 ;
        RECT 21.705000 44.670000 21.905000 44.870000 ;
        RECT 21.705000 45.100000 21.905000 45.300000 ;
        RECT 21.705000 45.530000 21.905000 45.730000 ;
        RECT 21.705000 45.960000 21.905000 46.160000 ;
        RECT 22.105000 41.660000 22.305000 41.860000 ;
        RECT 22.105000 42.090000 22.305000 42.290000 ;
        RECT 22.105000 42.520000 22.305000 42.720000 ;
        RECT 22.105000 42.950000 22.305000 43.150000 ;
        RECT 22.105000 43.380000 22.305000 43.580000 ;
        RECT 22.105000 43.810000 22.305000 44.010000 ;
        RECT 22.105000 44.240000 22.305000 44.440000 ;
        RECT 22.105000 44.670000 22.305000 44.870000 ;
        RECT 22.105000 45.100000 22.305000 45.300000 ;
        RECT 22.105000 45.530000 22.305000 45.730000 ;
        RECT 22.105000 45.960000 22.305000 46.160000 ;
        RECT 22.505000 41.660000 22.705000 41.860000 ;
        RECT 22.505000 42.090000 22.705000 42.290000 ;
        RECT 22.505000 42.520000 22.705000 42.720000 ;
        RECT 22.505000 42.950000 22.705000 43.150000 ;
        RECT 22.505000 43.380000 22.705000 43.580000 ;
        RECT 22.505000 43.810000 22.705000 44.010000 ;
        RECT 22.505000 44.240000 22.705000 44.440000 ;
        RECT 22.505000 44.670000 22.705000 44.870000 ;
        RECT 22.505000 45.100000 22.705000 45.300000 ;
        RECT 22.505000 45.530000 22.705000 45.730000 ;
        RECT 22.505000 45.960000 22.705000 46.160000 ;
        RECT 22.905000 41.660000 23.105000 41.860000 ;
        RECT 22.905000 42.090000 23.105000 42.290000 ;
        RECT 22.905000 42.520000 23.105000 42.720000 ;
        RECT 22.905000 42.950000 23.105000 43.150000 ;
        RECT 22.905000 43.380000 23.105000 43.580000 ;
        RECT 22.905000 43.810000 23.105000 44.010000 ;
        RECT 22.905000 44.240000 23.105000 44.440000 ;
        RECT 22.905000 44.670000 23.105000 44.870000 ;
        RECT 22.905000 45.100000 23.105000 45.300000 ;
        RECT 22.905000 45.530000 23.105000 45.730000 ;
        RECT 22.905000 45.960000 23.105000 46.160000 ;
        RECT 23.305000 41.660000 23.505000 41.860000 ;
        RECT 23.305000 42.090000 23.505000 42.290000 ;
        RECT 23.305000 42.520000 23.505000 42.720000 ;
        RECT 23.305000 42.950000 23.505000 43.150000 ;
        RECT 23.305000 43.380000 23.505000 43.580000 ;
        RECT 23.305000 43.810000 23.505000 44.010000 ;
        RECT 23.305000 44.240000 23.505000 44.440000 ;
        RECT 23.305000 44.670000 23.505000 44.870000 ;
        RECT 23.305000 45.100000 23.505000 45.300000 ;
        RECT 23.305000 45.530000 23.505000 45.730000 ;
        RECT 23.305000 45.960000 23.505000 46.160000 ;
        RECT 23.705000 41.660000 23.905000 41.860000 ;
        RECT 23.705000 42.090000 23.905000 42.290000 ;
        RECT 23.705000 42.520000 23.905000 42.720000 ;
        RECT 23.705000 42.950000 23.905000 43.150000 ;
        RECT 23.705000 43.380000 23.905000 43.580000 ;
        RECT 23.705000 43.810000 23.905000 44.010000 ;
        RECT 23.705000 44.240000 23.905000 44.440000 ;
        RECT 23.705000 44.670000 23.905000 44.870000 ;
        RECT 23.705000 45.100000 23.905000 45.300000 ;
        RECT 23.705000 45.530000 23.905000 45.730000 ;
        RECT 23.705000 45.960000 23.905000 46.160000 ;
        RECT 24.105000 41.660000 24.305000 41.860000 ;
        RECT 24.105000 42.090000 24.305000 42.290000 ;
        RECT 24.105000 42.520000 24.305000 42.720000 ;
        RECT 24.105000 42.950000 24.305000 43.150000 ;
        RECT 24.105000 43.380000 24.305000 43.580000 ;
        RECT 24.105000 43.810000 24.305000 44.010000 ;
        RECT 24.105000 44.240000 24.305000 44.440000 ;
        RECT 24.105000 44.670000 24.305000 44.870000 ;
        RECT 24.105000 45.100000 24.305000 45.300000 ;
        RECT 24.105000 45.530000 24.305000 45.730000 ;
        RECT 24.105000 45.960000 24.305000 46.160000 ;
        RECT 50.480000 41.660000 50.680000 41.860000 ;
        RECT 50.480000 42.090000 50.680000 42.290000 ;
        RECT 50.480000 42.520000 50.680000 42.720000 ;
        RECT 50.480000 42.950000 50.680000 43.150000 ;
        RECT 50.480000 43.380000 50.680000 43.580000 ;
        RECT 50.480000 43.810000 50.680000 44.010000 ;
        RECT 50.480000 44.240000 50.680000 44.440000 ;
        RECT 50.480000 44.670000 50.680000 44.870000 ;
        RECT 50.480000 45.100000 50.680000 45.300000 ;
        RECT 50.480000 45.530000 50.680000 45.730000 ;
        RECT 50.480000 45.960000 50.680000 46.160000 ;
        RECT 50.890000 41.660000 51.090000 41.860000 ;
        RECT 50.890000 42.090000 51.090000 42.290000 ;
        RECT 50.890000 42.520000 51.090000 42.720000 ;
        RECT 50.890000 42.950000 51.090000 43.150000 ;
        RECT 50.890000 43.380000 51.090000 43.580000 ;
        RECT 50.890000 43.810000 51.090000 44.010000 ;
        RECT 50.890000 44.240000 51.090000 44.440000 ;
        RECT 50.890000 44.670000 51.090000 44.870000 ;
        RECT 50.890000 45.100000 51.090000 45.300000 ;
        RECT 50.890000 45.530000 51.090000 45.730000 ;
        RECT 50.890000 45.960000 51.090000 46.160000 ;
        RECT 51.300000 41.660000 51.500000 41.860000 ;
        RECT 51.300000 42.090000 51.500000 42.290000 ;
        RECT 51.300000 42.520000 51.500000 42.720000 ;
        RECT 51.300000 42.950000 51.500000 43.150000 ;
        RECT 51.300000 43.380000 51.500000 43.580000 ;
        RECT 51.300000 43.810000 51.500000 44.010000 ;
        RECT 51.300000 44.240000 51.500000 44.440000 ;
        RECT 51.300000 44.670000 51.500000 44.870000 ;
        RECT 51.300000 45.100000 51.500000 45.300000 ;
        RECT 51.300000 45.530000 51.500000 45.730000 ;
        RECT 51.300000 45.960000 51.500000 46.160000 ;
        RECT 51.710000 41.660000 51.910000 41.860000 ;
        RECT 51.710000 42.090000 51.910000 42.290000 ;
        RECT 51.710000 42.520000 51.910000 42.720000 ;
        RECT 51.710000 42.950000 51.910000 43.150000 ;
        RECT 51.710000 43.380000 51.910000 43.580000 ;
        RECT 51.710000 43.810000 51.910000 44.010000 ;
        RECT 51.710000 44.240000 51.910000 44.440000 ;
        RECT 51.710000 44.670000 51.910000 44.870000 ;
        RECT 51.710000 45.100000 51.910000 45.300000 ;
        RECT 51.710000 45.530000 51.910000 45.730000 ;
        RECT 51.710000 45.960000 51.910000 46.160000 ;
        RECT 52.120000 41.660000 52.320000 41.860000 ;
        RECT 52.120000 42.090000 52.320000 42.290000 ;
        RECT 52.120000 42.520000 52.320000 42.720000 ;
        RECT 52.120000 42.950000 52.320000 43.150000 ;
        RECT 52.120000 43.380000 52.320000 43.580000 ;
        RECT 52.120000 43.810000 52.320000 44.010000 ;
        RECT 52.120000 44.240000 52.320000 44.440000 ;
        RECT 52.120000 44.670000 52.320000 44.870000 ;
        RECT 52.120000 45.100000 52.320000 45.300000 ;
        RECT 52.120000 45.530000 52.320000 45.730000 ;
        RECT 52.120000 45.960000 52.320000 46.160000 ;
        RECT 52.530000 41.660000 52.730000 41.860000 ;
        RECT 52.530000 42.090000 52.730000 42.290000 ;
        RECT 52.530000 42.520000 52.730000 42.720000 ;
        RECT 52.530000 42.950000 52.730000 43.150000 ;
        RECT 52.530000 43.380000 52.730000 43.580000 ;
        RECT 52.530000 43.810000 52.730000 44.010000 ;
        RECT 52.530000 44.240000 52.730000 44.440000 ;
        RECT 52.530000 44.670000 52.730000 44.870000 ;
        RECT 52.530000 45.100000 52.730000 45.300000 ;
        RECT 52.530000 45.530000 52.730000 45.730000 ;
        RECT 52.530000 45.960000 52.730000 46.160000 ;
        RECT 52.940000 41.660000 53.140000 41.860000 ;
        RECT 52.940000 42.090000 53.140000 42.290000 ;
        RECT 52.940000 42.520000 53.140000 42.720000 ;
        RECT 52.940000 42.950000 53.140000 43.150000 ;
        RECT 52.940000 43.380000 53.140000 43.580000 ;
        RECT 52.940000 43.810000 53.140000 44.010000 ;
        RECT 52.940000 44.240000 53.140000 44.440000 ;
        RECT 52.940000 44.670000 53.140000 44.870000 ;
        RECT 52.940000 45.100000 53.140000 45.300000 ;
        RECT 52.940000 45.530000 53.140000 45.730000 ;
        RECT 52.940000 45.960000 53.140000 46.160000 ;
        RECT 53.345000 41.660000 53.545000 41.860000 ;
        RECT 53.345000 42.090000 53.545000 42.290000 ;
        RECT 53.345000 42.520000 53.545000 42.720000 ;
        RECT 53.345000 42.950000 53.545000 43.150000 ;
        RECT 53.345000 43.380000 53.545000 43.580000 ;
        RECT 53.345000 43.810000 53.545000 44.010000 ;
        RECT 53.345000 44.240000 53.545000 44.440000 ;
        RECT 53.345000 44.670000 53.545000 44.870000 ;
        RECT 53.345000 45.100000 53.545000 45.300000 ;
        RECT 53.345000 45.530000 53.545000 45.730000 ;
        RECT 53.345000 45.960000 53.545000 46.160000 ;
        RECT 53.750000 41.660000 53.950000 41.860000 ;
        RECT 53.750000 42.090000 53.950000 42.290000 ;
        RECT 53.750000 42.520000 53.950000 42.720000 ;
        RECT 53.750000 42.950000 53.950000 43.150000 ;
        RECT 53.750000 43.380000 53.950000 43.580000 ;
        RECT 53.750000 43.810000 53.950000 44.010000 ;
        RECT 53.750000 44.240000 53.950000 44.440000 ;
        RECT 53.750000 44.670000 53.950000 44.870000 ;
        RECT 53.750000 45.100000 53.950000 45.300000 ;
        RECT 53.750000 45.530000 53.950000 45.730000 ;
        RECT 53.750000 45.960000 53.950000 46.160000 ;
        RECT 54.155000 41.660000 54.355000 41.860000 ;
        RECT 54.155000 42.090000 54.355000 42.290000 ;
        RECT 54.155000 42.520000 54.355000 42.720000 ;
        RECT 54.155000 42.950000 54.355000 43.150000 ;
        RECT 54.155000 43.380000 54.355000 43.580000 ;
        RECT 54.155000 43.810000 54.355000 44.010000 ;
        RECT 54.155000 44.240000 54.355000 44.440000 ;
        RECT 54.155000 44.670000 54.355000 44.870000 ;
        RECT 54.155000 45.100000 54.355000 45.300000 ;
        RECT 54.155000 45.530000 54.355000 45.730000 ;
        RECT 54.155000 45.960000 54.355000 46.160000 ;
        RECT 54.560000 41.660000 54.760000 41.860000 ;
        RECT 54.560000 42.090000 54.760000 42.290000 ;
        RECT 54.560000 42.520000 54.760000 42.720000 ;
        RECT 54.560000 42.950000 54.760000 43.150000 ;
        RECT 54.560000 43.380000 54.760000 43.580000 ;
        RECT 54.560000 43.810000 54.760000 44.010000 ;
        RECT 54.560000 44.240000 54.760000 44.440000 ;
        RECT 54.560000 44.670000 54.760000 44.870000 ;
        RECT 54.560000 45.100000 54.760000 45.300000 ;
        RECT 54.560000 45.530000 54.760000 45.730000 ;
        RECT 54.560000 45.960000 54.760000 46.160000 ;
        RECT 54.965000 41.660000 55.165000 41.860000 ;
        RECT 54.965000 42.090000 55.165000 42.290000 ;
        RECT 54.965000 42.520000 55.165000 42.720000 ;
        RECT 54.965000 42.950000 55.165000 43.150000 ;
        RECT 54.965000 43.380000 55.165000 43.580000 ;
        RECT 54.965000 43.810000 55.165000 44.010000 ;
        RECT 54.965000 44.240000 55.165000 44.440000 ;
        RECT 54.965000 44.670000 55.165000 44.870000 ;
        RECT 54.965000 45.100000 55.165000 45.300000 ;
        RECT 54.965000 45.530000 55.165000 45.730000 ;
        RECT 54.965000 45.960000 55.165000 46.160000 ;
        RECT 55.370000 41.660000 55.570000 41.860000 ;
        RECT 55.370000 42.090000 55.570000 42.290000 ;
        RECT 55.370000 42.520000 55.570000 42.720000 ;
        RECT 55.370000 42.950000 55.570000 43.150000 ;
        RECT 55.370000 43.380000 55.570000 43.580000 ;
        RECT 55.370000 43.810000 55.570000 44.010000 ;
        RECT 55.370000 44.240000 55.570000 44.440000 ;
        RECT 55.370000 44.670000 55.570000 44.870000 ;
        RECT 55.370000 45.100000 55.570000 45.300000 ;
        RECT 55.370000 45.530000 55.570000 45.730000 ;
        RECT 55.370000 45.960000 55.570000 46.160000 ;
        RECT 55.775000 41.660000 55.975000 41.860000 ;
        RECT 55.775000 42.090000 55.975000 42.290000 ;
        RECT 55.775000 42.520000 55.975000 42.720000 ;
        RECT 55.775000 42.950000 55.975000 43.150000 ;
        RECT 55.775000 43.380000 55.975000 43.580000 ;
        RECT 55.775000 43.810000 55.975000 44.010000 ;
        RECT 55.775000 44.240000 55.975000 44.440000 ;
        RECT 55.775000 44.670000 55.975000 44.870000 ;
        RECT 55.775000 45.100000 55.975000 45.300000 ;
        RECT 55.775000 45.530000 55.975000 45.730000 ;
        RECT 55.775000 45.960000 55.975000 46.160000 ;
        RECT 56.180000 41.660000 56.380000 41.860000 ;
        RECT 56.180000 42.090000 56.380000 42.290000 ;
        RECT 56.180000 42.520000 56.380000 42.720000 ;
        RECT 56.180000 42.950000 56.380000 43.150000 ;
        RECT 56.180000 43.380000 56.380000 43.580000 ;
        RECT 56.180000 43.810000 56.380000 44.010000 ;
        RECT 56.180000 44.240000 56.380000 44.440000 ;
        RECT 56.180000 44.670000 56.380000 44.870000 ;
        RECT 56.180000 45.100000 56.380000 45.300000 ;
        RECT 56.180000 45.530000 56.380000 45.730000 ;
        RECT 56.180000 45.960000 56.380000 46.160000 ;
        RECT 56.585000 41.660000 56.785000 41.860000 ;
        RECT 56.585000 42.090000 56.785000 42.290000 ;
        RECT 56.585000 42.520000 56.785000 42.720000 ;
        RECT 56.585000 42.950000 56.785000 43.150000 ;
        RECT 56.585000 43.380000 56.785000 43.580000 ;
        RECT 56.585000 43.810000 56.785000 44.010000 ;
        RECT 56.585000 44.240000 56.785000 44.440000 ;
        RECT 56.585000 44.670000 56.785000 44.870000 ;
        RECT 56.585000 45.100000 56.785000 45.300000 ;
        RECT 56.585000 45.530000 56.785000 45.730000 ;
        RECT 56.585000 45.960000 56.785000 46.160000 ;
        RECT 56.990000 41.660000 57.190000 41.860000 ;
        RECT 56.990000 42.090000 57.190000 42.290000 ;
        RECT 56.990000 42.520000 57.190000 42.720000 ;
        RECT 56.990000 42.950000 57.190000 43.150000 ;
        RECT 56.990000 43.380000 57.190000 43.580000 ;
        RECT 56.990000 43.810000 57.190000 44.010000 ;
        RECT 56.990000 44.240000 57.190000 44.440000 ;
        RECT 56.990000 44.670000 57.190000 44.870000 ;
        RECT 56.990000 45.100000 57.190000 45.300000 ;
        RECT 56.990000 45.530000 57.190000 45.730000 ;
        RECT 56.990000 45.960000 57.190000 46.160000 ;
        RECT 57.395000 41.660000 57.595000 41.860000 ;
        RECT 57.395000 42.090000 57.595000 42.290000 ;
        RECT 57.395000 42.520000 57.595000 42.720000 ;
        RECT 57.395000 42.950000 57.595000 43.150000 ;
        RECT 57.395000 43.380000 57.595000 43.580000 ;
        RECT 57.395000 43.810000 57.595000 44.010000 ;
        RECT 57.395000 44.240000 57.595000 44.440000 ;
        RECT 57.395000 44.670000 57.595000 44.870000 ;
        RECT 57.395000 45.100000 57.595000 45.300000 ;
        RECT 57.395000 45.530000 57.595000 45.730000 ;
        RECT 57.395000 45.960000 57.595000 46.160000 ;
        RECT 57.800000 41.660000 58.000000 41.860000 ;
        RECT 57.800000 42.090000 58.000000 42.290000 ;
        RECT 57.800000 42.520000 58.000000 42.720000 ;
        RECT 57.800000 42.950000 58.000000 43.150000 ;
        RECT 57.800000 43.380000 58.000000 43.580000 ;
        RECT 57.800000 43.810000 58.000000 44.010000 ;
        RECT 57.800000 44.240000 58.000000 44.440000 ;
        RECT 57.800000 44.670000 58.000000 44.870000 ;
        RECT 57.800000 45.100000 58.000000 45.300000 ;
        RECT 57.800000 45.530000 58.000000 45.730000 ;
        RECT 57.800000 45.960000 58.000000 46.160000 ;
        RECT 58.205000 41.660000 58.405000 41.860000 ;
        RECT 58.205000 42.090000 58.405000 42.290000 ;
        RECT 58.205000 42.520000 58.405000 42.720000 ;
        RECT 58.205000 42.950000 58.405000 43.150000 ;
        RECT 58.205000 43.380000 58.405000 43.580000 ;
        RECT 58.205000 43.810000 58.405000 44.010000 ;
        RECT 58.205000 44.240000 58.405000 44.440000 ;
        RECT 58.205000 44.670000 58.405000 44.870000 ;
        RECT 58.205000 45.100000 58.405000 45.300000 ;
        RECT 58.205000 45.530000 58.405000 45.730000 ;
        RECT 58.205000 45.960000 58.405000 46.160000 ;
        RECT 58.610000 41.660000 58.810000 41.860000 ;
        RECT 58.610000 42.090000 58.810000 42.290000 ;
        RECT 58.610000 42.520000 58.810000 42.720000 ;
        RECT 58.610000 42.950000 58.810000 43.150000 ;
        RECT 58.610000 43.380000 58.810000 43.580000 ;
        RECT 58.610000 43.810000 58.810000 44.010000 ;
        RECT 58.610000 44.240000 58.810000 44.440000 ;
        RECT 58.610000 44.670000 58.810000 44.870000 ;
        RECT 58.610000 45.100000 58.810000 45.300000 ;
        RECT 58.610000 45.530000 58.810000 45.730000 ;
        RECT 58.610000 45.960000 58.810000 46.160000 ;
        RECT 59.015000 41.660000 59.215000 41.860000 ;
        RECT 59.015000 42.090000 59.215000 42.290000 ;
        RECT 59.015000 42.520000 59.215000 42.720000 ;
        RECT 59.015000 42.950000 59.215000 43.150000 ;
        RECT 59.015000 43.380000 59.215000 43.580000 ;
        RECT 59.015000 43.810000 59.215000 44.010000 ;
        RECT 59.015000 44.240000 59.215000 44.440000 ;
        RECT 59.015000 44.670000 59.215000 44.870000 ;
        RECT 59.015000 45.100000 59.215000 45.300000 ;
        RECT 59.015000 45.530000 59.215000 45.730000 ;
        RECT 59.015000 45.960000 59.215000 46.160000 ;
        RECT 59.420000 41.660000 59.620000 41.860000 ;
        RECT 59.420000 42.090000 59.620000 42.290000 ;
        RECT 59.420000 42.520000 59.620000 42.720000 ;
        RECT 59.420000 42.950000 59.620000 43.150000 ;
        RECT 59.420000 43.380000 59.620000 43.580000 ;
        RECT 59.420000 43.810000 59.620000 44.010000 ;
        RECT 59.420000 44.240000 59.620000 44.440000 ;
        RECT 59.420000 44.670000 59.620000 44.870000 ;
        RECT 59.420000 45.100000 59.620000 45.300000 ;
        RECT 59.420000 45.530000 59.620000 45.730000 ;
        RECT 59.420000 45.960000 59.620000 46.160000 ;
        RECT 59.825000 41.660000 60.025000 41.860000 ;
        RECT 59.825000 42.090000 60.025000 42.290000 ;
        RECT 59.825000 42.520000 60.025000 42.720000 ;
        RECT 59.825000 42.950000 60.025000 43.150000 ;
        RECT 59.825000 43.380000 60.025000 43.580000 ;
        RECT 59.825000 43.810000 60.025000 44.010000 ;
        RECT 59.825000 44.240000 60.025000 44.440000 ;
        RECT 59.825000 44.670000 60.025000 44.870000 ;
        RECT 59.825000 45.100000 60.025000 45.300000 ;
        RECT 59.825000 45.530000 60.025000 45.730000 ;
        RECT 59.825000 45.960000 60.025000 46.160000 ;
        RECT 60.230000 41.660000 60.430000 41.860000 ;
        RECT 60.230000 42.090000 60.430000 42.290000 ;
        RECT 60.230000 42.520000 60.430000 42.720000 ;
        RECT 60.230000 42.950000 60.430000 43.150000 ;
        RECT 60.230000 43.380000 60.430000 43.580000 ;
        RECT 60.230000 43.810000 60.430000 44.010000 ;
        RECT 60.230000 44.240000 60.430000 44.440000 ;
        RECT 60.230000 44.670000 60.430000 44.870000 ;
        RECT 60.230000 45.100000 60.430000 45.300000 ;
        RECT 60.230000 45.530000 60.430000 45.730000 ;
        RECT 60.230000 45.960000 60.430000 46.160000 ;
        RECT 60.635000 41.660000 60.835000 41.860000 ;
        RECT 60.635000 42.090000 60.835000 42.290000 ;
        RECT 60.635000 42.520000 60.835000 42.720000 ;
        RECT 60.635000 42.950000 60.835000 43.150000 ;
        RECT 60.635000 43.380000 60.835000 43.580000 ;
        RECT 60.635000 43.810000 60.835000 44.010000 ;
        RECT 60.635000 44.240000 60.835000 44.440000 ;
        RECT 60.635000 44.670000 60.835000 44.870000 ;
        RECT 60.635000 45.100000 60.835000 45.300000 ;
        RECT 60.635000 45.530000 60.835000 45.730000 ;
        RECT 60.635000 45.960000 60.835000 46.160000 ;
        RECT 61.040000 41.660000 61.240000 41.860000 ;
        RECT 61.040000 42.090000 61.240000 42.290000 ;
        RECT 61.040000 42.520000 61.240000 42.720000 ;
        RECT 61.040000 42.950000 61.240000 43.150000 ;
        RECT 61.040000 43.380000 61.240000 43.580000 ;
        RECT 61.040000 43.810000 61.240000 44.010000 ;
        RECT 61.040000 44.240000 61.240000 44.440000 ;
        RECT 61.040000 44.670000 61.240000 44.870000 ;
        RECT 61.040000 45.100000 61.240000 45.300000 ;
        RECT 61.040000 45.530000 61.240000 45.730000 ;
        RECT 61.040000 45.960000 61.240000 46.160000 ;
        RECT 61.445000 41.660000 61.645000 41.860000 ;
        RECT 61.445000 42.090000 61.645000 42.290000 ;
        RECT 61.445000 42.520000 61.645000 42.720000 ;
        RECT 61.445000 42.950000 61.645000 43.150000 ;
        RECT 61.445000 43.380000 61.645000 43.580000 ;
        RECT 61.445000 43.810000 61.645000 44.010000 ;
        RECT 61.445000 44.240000 61.645000 44.440000 ;
        RECT 61.445000 44.670000 61.645000 44.870000 ;
        RECT 61.445000 45.100000 61.645000 45.300000 ;
        RECT 61.445000 45.530000 61.645000 45.730000 ;
        RECT 61.445000 45.960000 61.645000 46.160000 ;
        RECT 61.850000 41.660000 62.050000 41.860000 ;
        RECT 61.850000 42.090000 62.050000 42.290000 ;
        RECT 61.850000 42.520000 62.050000 42.720000 ;
        RECT 61.850000 42.950000 62.050000 43.150000 ;
        RECT 61.850000 43.380000 62.050000 43.580000 ;
        RECT 61.850000 43.810000 62.050000 44.010000 ;
        RECT 61.850000 44.240000 62.050000 44.440000 ;
        RECT 61.850000 44.670000 62.050000 44.870000 ;
        RECT 61.850000 45.100000 62.050000 45.300000 ;
        RECT 61.850000 45.530000 62.050000 45.730000 ;
        RECT 61.850000 45.960000 62.050000 46.160000 ;
        RECT 62.255000 41.660000 62.455000 41.860000 ;
        RECT 62.255000 42.090000 62.455000 42.290000 ;
        RECT 62.255000 42.520000 62.455000 42.720000 ;
        RECT 62.255000 42.950000 62.455000 43.150000 ;
        RECT 62.255000 43.380000 62.455000 43.580000 ;
        RECT 62.255000 43.810000 62.455000 44.010000 ;
        RECT 62.255000 44.240000 62.455000 44.440000 ;
        RECT 62.255000 44.670000 62.455000 44.870000 ;
        RECT 62.255000 45.100000 62.455000 45.300000 ;
        RECT 62.255000 45.530000 62.455000 45.730000 ;
        RECT 62.255000 45.960000 62.455000 46.160000 ;
        RECT 62.660000 41.660000 62.860000 41.860000 ;
        RECT 62.660000 42.090000 62.860000 42.290000 ;
        RECT 62.660000 42.520000 62.860000 42.720000 ;
        RECT 62.660000 42.950000 62.860000 43.150000 ;
        RECT 62.660000 43.380000 62.860000 43.580000 ;
        RECT 62.660000 43.810000 62.860000 44.010000 ;
        RECT 62.660000 44.240000 62.860000 44.440000 ;
        RECT 62.660000 44.670000 62.860000 44.870000 ;
        RECT 62.660000 45.100000 62.860000 45.300000 ;
        RECT 62.660000 45.530000 62.860000 45.730000 ;
        RECT 62.660000 45.960000 62.860000 46.160000 ;
        RECT 63.065000 41.660000 63.265000 41.860000 ;
        RECT 63.065000 42.090000 63.265000 42.290000 ;
        RECT 63.065000 42.520000 63.265000 42.720000 ;
        RECT 63.065000 42.950000 63.265000 43.150000 ;
        RECT 63.065000 43.380000 63.265000 43.580000 ;
        RECT 63.065000 43.810000 63.265000 44.010000 ;
        RECT 63.065000 44.240000 63.265000 44.440000 ;
        RECT 63.065000 44.670000 63.265000 44.870000 ;
        RECT 63.065000 45.100000 63.265000 45.300000 ;
        RECT 63.065000 45.530000 63.265000 45.730000 ;
        RECT 63.065000 45.960000 63.265000 46.160000 ;
        RECT 63.470000 41.660000 63.670000 41.860000 ;
        RECT 63.470000 42.090000 63.670000 42.290000 ;
        RECT 63.470000 42.520000 63.670000 42.720000 ;
        RECT 63.470000 42.950000 63.670000 43.150000 ;
        RECT 63.470000 43.380000 63.670000 43.580000 ;
        RECT 63.470000 43.810000 63.670000 44.010000 ;
        RECT 63.470000 44.240000 63.670000 44.440000 ;
        RECT 63.470000 44.670000 63.670000 44.870000 ;
        RECT 63.470000 45.100000 63.670000 45.300000 ;
        RECT 63.470000 45.530000 63.670000 45.730000 ;
        RECT 63.470000 45.960000 63.670000 46.160000 ;
        RECT 63.875000 41.660000 64.075000 41.860000 ;
        RECT 63.875000 42.090000 64.075000 42.290000 ;
        RECT 63.875000 42.520000 64.075000 42.720000 ;
        RECT 63.875000 42.950000 64.075000 43.150000 ;
        RECT 63.875000 43.380000 64.075000 43.580000 ;
        RECT 63.875000 43.810000 64.075000 44.010000 ;
        RECT 63.875000 44.240000 64.075000 44.440000 ;
        RECT 63.875000 44.670000 64.075000 44.870000 ;
        RECT 63.875000 45.100000 64.075000 45.300000 ;
        RECT 63.875000 45.530000 64.075000 45.730000 ;
        RECT 63.875000 45.960000 64.075000 46.160000 ;
        RECT 64.280000 41.660000 64.480000 41.860000 ;
        RECT 64.280000 42.090000 64.480000 42.290000 ;
        RECT 64.280000 42.520000 64.480000 42.720000 ;
        RECT 64.280000 42.950000 64.480000 43.150000 ;
        RECT 64.280000 43.380000 64.480000 43.580000 ;
        RECT 64.280000 43.810000 64.480000 44.010000 ;
        RECT 64.280000 44.240000 64.480000 44.440000 ;
        RECT 64.280000 44.670000 64.480000 44.870000 ;
        RECT 64.280000 45.100000 64.480000 45.300000 ;
        RECT 64.280000 45.530000 64.480000 45.730000 ;
        RECT 64.280000 45.960000 64.480000 46.160000 ;
        RECT 64.685000 41.660000 64.885000 41.860000 ;
        RECT 64.685000 42.090000 64.885000 42.290000 ;
        RECT 64.685000 42.520000 64.885000 42.720000 ;
        RECT 64.685000 42.950000 64.885000 43.150000 ;
        RECT 64.685000 43.380000 64.885000 43.580000 ;
        RECT 64.685000 43.810000 64.885000 44.010000 ;
        RECT 64.685000 44.240000 64.885000 44.440000 ;
        RECT 64.685000 44.670000 64.885000 44.870000 ;
        RECT 64.685000 45.100000 64.885000 45.300000 ;
        RECT 64.685000 45.530000 64.885000 45.730000 ;
        RECT 64.685000 45.960000 64.885000 46.160000 ;
        RECT 65.090000 41.660000 65.290000 41.860000 ;
        RECT 65.090000 42.090000 65.290000 42.290000 ;
        RECT 65.090000 42.520000 65.290000 42.720000 ;
        RECT 65.090000 42.950000 65.290000 43.150000 ;
        RECT 65.090000 43.380000 65.290000 43.580000 ;
        RECT 65.090000 43.810000 65.290000 44.010000 ;
        RECT 65.090000 44.240000 65.290000 44.440000 ;
        RECT 65.090000 44.670000 65.290000 44.870000 ;
        RECT 65.090000 45.100000 65.290000 45.300000 ;
        RECT 65.090000 45.530000 65.290000 45.730000 ;
        RECT 65.090000 45.960000 65.290000 46.160000 ;
        RECT 65.495000 41.660000 65.695000 41.860000 ;
        RECT 65.495000 42.090000 65.695000 42.290000 ;
        RECT 65.495000 42.520000 65.695000 42.720000 ;
        RECT 65.495000 42.950000 65.695000 43.150000 ;
        RECT 65.495000 43.380000 65.695000 43.580000 ;
        RECT 65.495000 43.810000 65.695000 44.010000 ;
        RECT 65.495000 44.240000 65.695000 44.440000 ;
        RECT 65.495000 44.670000 65.695000 44.870000 ;
        RECT 65.495000 45.100000 65.695000 45.300000 ;
        RECT 65.495000 45.530000 65.695000 45.730000 ;
        RECT 65.495000 45.960000 65.695000 46.160000 ;
        RECT 65.900000 41.660000 66.100000 41.860000 ;
        RECT 65.900000 42.090000 66.100000 42.290000 ;
        RECT 65.900000 42.520000 66.100000 42.720000 ;
        RECT 65.900000 42.950000 66.100000 43.150000 ;
        RECT 65.900000 43.380000 66.100000 43.580000 ;
        RECT 65.900000 43.810000 66.100000 44.010000 ;
        RECT 65.900000 44.240000 66.100000 44.440000 ;
        RECT 65.900000 44.670000 66.100000 44.870000 ;
        RECT 65.900000 45.100000 66.100000 45.300000 ;
        RECT 65.900000 45.530000 66.100000 45.730000 ;
        RECT 65.900000 45.960000 66.100000 46.160000 ;
        RECT 66.305000 41.660000 66.505000 41.860000 ;
        RECT 66.305000 42.090000 66.505000 42.290000 ;
        RECT 66.305000 42.520000 66.505000 42.720000 ;
        RECT 66.305000 42.950000 66.505000 43.150000 ;
        RECT 66.305000 43.380000 66.505000 43.580000 ;
        RECT 66.305000 43.810000 66.505000 44.010000 ;
        RECT 66.305000 44.240000 66.505000 44.440000 ;
        RECT 66.305000 44.670000 66.505000 44.870000 ;
        RECT 66.305000 45.100000 66.505000 45.300000 ;
        RECT 66.305000 45.530000 66.505000 45.730000 ;
        RECT 66.305000 45.960000 66.505000 46.160000 ;
        RECT 66.710000 41.660000 66.910000 41.860000 ;
        RECT 66.710000 42.090000 66.910000 42.290000 ;
        RECT 66.710000 42.520000 66.910000 42.720000 ;
        RECT 66.710000 42.950000 66.910000 43.150000 ;
        RECT 66.710000 43.380000 66.910000 43.580000 ;
        RECT 66.710000 43.810000 66.910000 44.010000 ;
        RECT 66.710000 44.240000 66.910000 44.440000 ;
        RECT 66.710000 44.670000 66.910000 44.870000 ;
        RECT 66.710000 45.100000 66.910000 45.300000 ;
        RECT 66.710000 45.530000 66.910000 45.730000 ;
        RECT 66.710000 45.960000 66.910000 46.160000 ;
        RECT 67.115000 41.660000 67.315000 41.860000 ;
        RECT 67.115000 42.090000 67.315000 42.290000 ;
        RECT 67.115000 42.520000 67.315000 42.720000 ;
        RECT 67.115000 42.950000 67.315000 43.150000 ;
        RECT 67.115000 43.380000 67.315000 43.580000 ;
        RECT 67.115000 43.810000 67.315000 44.010000 ;
        RECT 67.115000 44.240000 67.315000 44.440000 ;
        RECT 67.115000 44.670000 67.315000 44.870000 ;
        RECT 67.115000 45.100000 67.315000 45.300000 ;
        RECT 67.115000 45.530000 67.315000 45.730000 ;
        RECT 67.115000 45.960000 67.315000 46.160000 ;
        RECT 67.520000 41.660000 67.720000 41.860000 ;
        RECT 67.520000 42.090000 67.720000 42.290000 ;
        RECT 67.520000 42.520000 67.720000 42.720000 ;
        RECT 67.520000 42.950000 67.720000 43.150000 ;
        RECT 67.520000 43.380000 67.720000 43.580000 ;
        RECT 67.520000 43.810000 67.720000 44.010000 ;
        RECT 67.520000 44.240000 67.720000 44.440000 ;
        RECT 67.520000 44.670000 67.720000 44.870000 ;
        RECT 67.520000 45.100000 67.720000 45.300000 ;
        RECT 67.520000 45.530000 67.720000 45.730000 ;
        RECT 67.520000 45.960000 67.720000 46.160000 ;
        RECT 67.925000 41.660000 68.125000 41.860000 ;
        RECT 67.925000 42.090000 68.125000 42.290000 ;
        RECT 67.925000 42.520000 68.125000 42.720000 ;
        RECT 67.925000 42.950000 68.125000 43.150000 ;
        RECT 67.925000 43.380000 68.125000 43.580000 ;
        RECT 67.925000 43.810000 68.125000 44.010000 ;
        RECT 67.925000 44.240000 68.125000 44.440000 ;
        RECT 67.925000 44.670000 68.125000 44.870000 ;
        RECT 67.925000 45.100000 68.125000 45.300000 ;
        RECT 67.925000 45.530000 68.125000 45.730000 ;
        RECT 67.925000 45.960000 68.125000 46.160000 ;
        RECT 68.330000 41.660000 68.530000 41.860000 ;
        RECT 68.330000 42.090000 68.530000 42.290000 ;
        RECT 68.330000 42.520000 68.530000 42.720000 ;
        RECT 68.330000 42.950000 68.530000 43.150000 ;
        RECT 68.330000 43.380000 68.530000 43.580000 ;
        RECT 68.330000 43.810000 68.530000 44.010000 ;
        RECT 68.330000 44.240000 68.530000 44.440000 ;
        RECT 68.330000 44.670000 68.530000 44.870000 ;
        RECT 68.330000 45.100000 68.530000 45.300000 ;
        RECT 68.330000 45.530000 68.530000 45.730000 ;
        RECT 68.330000 45.960000 68.530000 46.160000 ;
        RECT 68.735000 41.660000 68.935000 41.860000 ;
        RECT 68.735000 42.090000 68.935000 42.290000 ;
        RECT 68.735000 42.520000 68.935000 42.720000 ;
        RECT 68.735000 42.950000 68.935000 43.150000 ;
        RECT 68.735000 43.380000 68.935000 43.580000 ;
        RECT 68.735000 43.810000 68.935000 44.010000 ;
        RECT 68.735000 44.240000 68.935000 44.440000 ;
        RECT 68.735000 44.670000 68.935000 44.870000 ;
        RECT 68.735000 45.100000 68.935000 45.300000 ;
        RECT 68.735000 45.530000 68.935000 45.730000 ;
        RECT 68.735000 45.960000 68.935000 46.160000 ;
        RECT 69.140000 41.660000 69.340000 41.860000 ;
        RECT 69.140000 42.090000 69.340000 42.290000 ;
        RECT 69.140000 42.520000 69.340000 42.720000 ;
        RECT 69.140000 42.950000 69.340000 43.150000 ;
        RECT 69.140000 43.380000 69.340000 43.580000 ;
        RECT 69.140000 43.810000 69.340000 44.010000 ;
        RECT 69.140000 44.240000 69.340000 44.440000 ;
        RECT 69.140000 44.670000 69.340000 44.870000 ;
        RECT 69.140000 45.100000 69.340000 45.300000 ;
        RECT 69.140000 45.530000 69.340000 45.730000 ;
        RECT 69.140000 45.960000 69.340000 46.160000 ;
        RECT 69.545000 41.660000 69.745000 41.860000 ;
        RECT 69.545000 42.090000 69.745000 42.290000 ;
        RECT 69.545000 42.520000 69.745000 42.720000 ;
        RECT 69.545000 42.950000 69.745000 43.150000 ;
        RECT 69.545000 43.380000 69.745000 43.580000 ;
        RECT 69.545000 43.810000 69.745000 44.010000 ;
        RECT 69.545000 44.240000 69.745000 44.440000 ;
        RECT 69.545000 44.670000 69.745000 44.870000 ;
        RECT 69.545000 45.100000 69.745000 45.300000 ;
        RECT 69.545000 45.530000 69.745000 45.730000 ;
        RECT 69.545000 45.960000 69.745000 46.160000 ;
        RECT 69.950000 41.660000 70.150000 41.860000 ;
        RECT 69.950000 42.090000 70.150000 42.290000 ;
        RECT 69.950000 42.520000 70.150000 42.720000 ;
        RECT 69.950000 42.950000 70.150000 43.150000 ;
        RECT 69.950000 43.380000 70.150000 43.580000 ;
        RECT 69.950000 43.810000 70.150000 44.010000 ;
        RECT 69.950000 44.240000 70.150000 44.440000 ;
        RECT 69.950000 44.670000 70.150000 44.870000 ;
        RECT 69.950000 45.100000 70.150000 45.300000 ;
        RECT 69.950000 45.530000 70.150000 45.730000 ;
        RECT 69.950000 45.960000 70.150000 46.160000 ;
        RECT 70.355000 41.660000 70.555000 41.860000 ;
        RECT 70.355000 42.090000 70.555000 42.290000 ;
        RECT 70.355000 42.520000 70.555000 42.720000 ;
        RECT 70.355000 42.950000 70.555000 43.150000 ;
        RECT 70.355000 43.380000 70.555000 43.580000 ;
        RECT 70.355000 43.810000 70.555000 44.010000 ;
        RECT 70.355000 44.240000 70.555000 44.440000 ;
        RECT 70.355000 44.670000 70.555000 44.870000 ;
        RECT 70.355000 45.100000 70.555000 45.300000 ;
        RECT 70.355000 45.530000 70.555000 45.730000 ;
        RECT 70.355000 45.960000 70.555000 46.160000 ;
        RECT 70.760000 41.660000 70.960000 41.860000 ;
        RECT 70.760000 42.090000 70.960000 42.290000 ;
        RECT 70.760000 42.520000 70.960000 42.720000 ;
        RECT 70.760000 42.950000 70.960000 43.150000 ;
        RECT 70.760000 43.380000 70.960000 43.580000 ;
        RECT 70.760000 43.810000 70.960000 44.010000 ;
        RECT 70.760000 44.240000 70.960000 44.440000 ;
        RECT 70.760000 44.670000 70.960000 44.870000 ;
        RECT 70.760000 45.100000 70.960000 45.300000 ;
        RECT 70.760000 45.530000 70.960000 45.730000 ;
        RECT 70.760000 45.960000 70.960000 46.160000 ;
        RECT 71.165000 41.660000 71.365000 41.860000 ;
        RECT 71.165000 42.090000 71.365000 42.290000 ;
        RECT 71.165000 42.520000 71.365000 42.720000 ;
        RECT 71.165000 42.950000 71.365000 43.150000 ;
        RECT 71.165000 43.380000 71.365000 43.580000 ;
        RECT 71.165000 43.810000 71.365000 44.010000 ;
        RECT 71.165000 44.240000 71.365000 44.440000 ;
        RECT 71.165000 44.670000 71.365000 44.870000 ;
        RECT 71.165000 45.100000 71.365000 45.300000 ;
        RECT 71.165000 45.530000 71.365000 45.730000 ;
        RECT 71.165000 45.960000 71.365000 46.160000 ;
        RECT 71.570000 41.660000 71.770000 41.860000 ;
        RECT 71.570000 42.090000 71.770000 42.290000 ;
        RECT 71.570000 42.520000 71.770000 42.720000 ;
        RECT 71.570000 42.950000 71.770000 43.150000 ;
        RECT 71.570000 43.380000 71.770000 43.580000 ;
        RECT 71.570000 43.810000 71.770000 44.010000 ;
        RECT 71.570000 44.240000 71.770000 44.440000 ;
        RECT 71.570000 44.670000 71.770000 44.870000 ;
        RECT 71.570000 45.100000 71.770000 45.300000 ;
        RECT 71.570000 45.530000 71.770000 45.730000 ;
        RECT 71.570000 45.960000 71.770000 46.160000 ;
        RECT 71.975000 41.660000 72.175000 41.860000 ;
        RECT 71.975000 42.090000 72.175000 42.290000 ;
        RECT 71.975000 42.520000 72.175000 42.720000 ;
        RECT 71.975000 42.950000 72.175000 43.150000 ;
        RECT 71.975000 43.380000 72.175000 43.580000 ;
        RECT 71.975000 43.810000 72.175000 44.010000 ;
        RECT 71.975000 44.240000 72.175000 44.440000 ;
        RECT 71.975000 44.670000 72.175000 44.870000 ;
        RECT 71.975000 45.100000 72.175000 45.300000 ;
        RECT 71.975000 45.530000 72.175000 45.730000 ;
        RECT 71.975000 45.960000 72.175000 46.160000 ;
        RECT 72.380000 41.660000 72.580000 41.860000 ;
        RECT 72.380000 42.090000 72.580000 42.290000 ;
        RECT 72.380000 42.520000 72.580000 42.720000 ;
        RECT 72.380000 42.950000 72.580000 43.150000 ;
        RECT 72.380000 43.380000 72.580000 43.580000 ;
        RECT 72.380000 43.810000 72.580000 44.010000 ;
        RECT 72.380000 44.240000 72.580000 44.440000 ;
        RECT 72.380000 44.670000 72.580000 44.870000 ;
        RECT 72.380000 45.100000 72.580000 45.300000 ;
        RECT 72.380000 45.530000 72.580000 45.730000 ;
        RECT 72.380000 45.960000 72.580000 46.160000 ;
        RECT 72.785000 41.660000 72.985000 41.860000 ;
        RECT 72.785000 42.090000 72.985000 42.290000 ;
        RECT 72.785000 42.520000 72.985000 42.720000 ;
        RECT 72.785000 42.950000 72.985000 43.150000 ;
        RECT 72.785000 43.380000 72.985000 43.580000 ;
        RECT 72.785000 43.810000 72.985000 44.010000 ;
        RECT 72.785000 44.240000 72.985000 44.440000 ;
        RECT 72.785000 44.670000 72.985000 44.870000 ;
        RECT 72.785000 45.100000 72.985000 45.300000 ;
        RECT 72.785000 45.530000 72.985000 45.730000 ;
        RECT 72.785000 45.960000 72.985000 46.160000 ;
        RECT 73.190000 41.660000 73.390000 41.860000 ;
        RECT 73.190000 42.090000 73.390000 42.290000 ;
        RECT 73.190000 42.520000 73.390000 42.720000 ;
        RECT 73.190000 42.950000 73.390000 43.150000 ;
        RECT 73.190000 43.380000 73.390000 43.580000 ;
        RECT 73.190000 43.810000 73.390000 44.010000 ;
        RECT 73.190000 44.240000 73.390000 44.440000 ;
        RECT 73.190000 44.670000 73.390000 44.870000 ;
        RECT 73.190000 45.100000 73.390000 45.300000 ;
        RECT 73.190000 45.530000 73.390000 45.730000 ;
        RECT 73.190000 45.960000 73.390000 46.160000 ;
        RECT 73.595000 41.660000 73.795000 41.860000 ;
        RECT 73.595000 42.090000 73.795000 42.290000 ;
        RECT 73.595000 42.520000 73.795000 42.720000 ;
        RECT 73.595000 42.950000 73.795000 43.150000 ;
        RECT 73.595000 43.380000 73.795000 43.580000 ;
        RECT 73.595000 43.810000 73.795000 44.010000 ;
        RECT 73.595000 44.240000 73.795000 44.440000 ;
        RECT 73.595000 44.670000 73.795000 44.870000 ;
        RECT 73.595000 45.100000 73.795000 45.300000 ;
        RECT 73.595000 45.530000 73.795000 45.730000 ;
        RECT 73.595000 45.960000 73.795000 46.160000 ;
        RECT 74.000000 41.660000 74.200000 41.860000 ;
        RECT 74.000000 42.090000 74.200000 42.290000 ;
        RECT 74.000000 42.520000 74.200000 42.720000 ;
        RECT 74.000000 42.950000 74.200000 43.150000 ;
        RECT 74.000000 43.380000 74.200000 43.580000 ;
        RECT 74.000000 43.810000 74.200000 44.010000 ;
        RECT 74.000000 44.240000 74.200000 44.440000 ;
        RECT 74.000000 44.670000 74.200000 44.870000 ;
        RECT 74.000000 45.100000 74.200000 45.300000 ;
        RECT 74.000000 45.530000 74.200000 45.730000 ;
        RECT 74.000000 45.960000 74.200000 46.160000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 1.270000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 25.835000 75.000000 30.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 1.270000 30.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 1.270000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 58.235000 75.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 1.270000 62.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 31.885000 75.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 1.270000 35.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met3 ;
      RECT  0.000000  0.000000 75.000000  41.190000 ;
      RECT  0.000000 41.190000  0.570000  46.630000 ;
      RECT  0.000000 46.630000 75.000000 200.000000 ;
      RECT 24.795000 41.190000 49.990000  46.630000 ;
      RECT 74.690000 41.190000 75.000000  46.630000 ;
    LAYER met4 ;
      RECT  0.000000   0.000000  1.670000   1.635000 ;
      RECT  0.000000   7.885000  1.670000   8.485000 ;
      RECT  0.000000  13.935000  1.365000  14.535000 ;
      RECT  0.000000  18.785000  1.365000  19.385000 ;
      RECT  0.000000  24.835000  1.670000  25.435000 ;
      RECT  0.000000  30.885000  1.670000  31.485000 ;
      RECT  0.000000  35.735000  1.670000  36.335000 ;
      RECT  0.000000  40.585000  1.670000  41.185000 ;
      RECT  0.000000  46.635000  1.670000  47.335000 ;
      RECT  0.000000  57.135000  1.670000  57.835000 ;
      RECT  0.000000  63.085000  1.670000  63.685000 ;
      RECT  0.000000  68.935000  1.670000  69.635000 ;
      RECT  0.000000  95.400000 75.000000 175.385000 ;
      RECT  1.365000  13.935000 73.635000  19.385000 ;
      RECT  1.670000   0.000000 73.330000  13.935000 ;
      RECT  1.670000  19.385000 73.330000  41.185000 ;
      RECT  1.670000  46.635000 73.330000  95.400000 ;
      RECT  1.670000 175.385000 73.330000 200.000000 ;
      RECT 24.770000  41.185000 50.015000  46.635000 ;
      RECT 73.330000   0.000000 75.000000   1.635000 ;
      RECT 73.330000   7.885000 75.000000   8.485000 ;
      RECT 73.330000  24.835000 75.000000  25.435000 ;
      RECT 73.330000  30.885000 75.000000  31.485000 ;
      RECT 73.330000  35.735000 75.000000  36.335000 ;
      RECT 73.330000  40.585000 75.000000  41.185000 ;
      RECT 73.330000  46.635000 75.000000  47.335000 ;
      RECT 73.330000  57.135000 75.000000  57.835000 ;
      RECT 73.330000  63.085000 75.000000  63.685000 ;
      RECT 73.330000  68.935000 75.000000  69.635000 ;
      RECT 73.635000  13.935000 75.000000  14.535000 ;
      RECT 73.635000  18.785000 75.000000  19.385000 ;
    LAYER met5 ;
      RECT 0.000000   0.000000 75.000000   1.335000 ;
      RECT 0.000000  95.785000 75.000000 174.985000 ;
      RECT 1.765000  14.235000 73.235000  19.085000 ;
      RECT 2.070000   1.335000 72.930000  14.235000 ;
      RECT 2.070000  19.085000 72.930000  95.785000 ;
      RECT 2.070000 174.985000 72.930000 200.000000 ;
  END
END sky130_fd_io__overlay_vssd_hvc
END LIBRARY
