# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__top_xres4v2
  CLASS BLOCK ;
  FOREIGN sky130_fd_io__top_xres4v2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  75.00000 BY  200.0000 ;
  SYMMETRY R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN DISABLE_PULLUP_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.760000 0.000000 33.020000 0.640000 ;
    END
  END DISABLE_PULLUP_H
  PIN ENABLE_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.285000 0.000000 12.545000 1.470000 ;
    END
  END ENABLE_H
  PIN ENABLE_VDDIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 6.775000 16.895000 7.290000 17.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.775000 17.410000 7.295000 31.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.775000 17.410000 7.400000 17.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.775000 17.515000 7.295000 17.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.775000 17.620000 7.295000 31.295000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.775000 31.400000 7.400000 31.505000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.775000 31.505000 7.150000 31.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.840000 17.345000 7.505000 17.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.925000 31.505000 7.505000 31.655000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.150000 31.880000 7.865000 32.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.290000 16.445000 7.740000 16.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.290000 16.895000 7.870000 17.045000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.295000 17.045000 7.870000 17.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.295000 31.295000 7.880000 31.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.375000 31.955000 7.955000 32.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 16.745000 8.020000 16.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.525000 32.105000 8.105000 32.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.675000 32.255000 8.255000 32.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.740000 15.995000 8.190000 16.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.865000 32.595000 8.450000 33.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.870000 16.585000 8.330000 17.045000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.880000 31.880000 8.595000 32.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.890000 16.295000 8.470000 16.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.125000 32.705000 8.705000 32.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.190000 15.785000 8.400000 15.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.275000 32.855000 8.855000 33.005000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.330000 15.995000 8.920000 16.585000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.400000 0.000000 8.920000 15.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.400000 1.135000 8.920000 15.995000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.450000 33.180000 8.970000 33.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.595000 32.595000 9.180000 33.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.815000 33.395000 22.275000 33.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.970000 33.700000 9.395000 34.125000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.115000 33.695000 22.275000 33.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.180000 33.180000 9.395000 33.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.395000 33.995000 22.275000 34.125000 ;
    END
  END ENABLE_VDDIO
  PIN EN_VDDIO_SIG_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.005000 3.905000 10.350000 4.250000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.045000 4.250000 10.375000 4.580000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.085000 9.250000 10.385000 9.320000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.140000 4.115000 10.440000 4.185000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.165000 9.400000 10.495000 9.730000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.210000 4.045000 10.510000 4.115000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.295000 9.460000 10.595000 9.530000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.335000 9.200000 10.535000 9.400000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.350000 3.575000 10.680000 3.905000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.365000 9.530000 10.665000 9.600000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.375000 3.930000 10.695000 4.250000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.420000 3.835000 10.720000 3.905000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.490000 3.765000 10.790000 3.835000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.495000 9.730000 10.865000 10.100000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.535000 9.400000 10.865000 9.730000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.575000 9.740000 10.875000 9.810000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.645000 9.810000 10.945000 9.880000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.650000 26.610000 10.865000 26.825000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.650000 26.825000 11.125000 27.085000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.650000 27.085000 10.910000 28.005000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.650000 27.085000 11.055000 27.155000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.650000 27.155000 10.985000 27.225000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.650000 27.295000 10.910000 27.300000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.650000 27.300000 10.910000 27.935000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.650000 28.005000 10.980000 28.075000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.650000 28.075000 11.050000 28.145000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.650000 28.150000 11.125000 28.410000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.650000 28.410000 10.865000 28.625000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.655000 26.820000 11.125000 26.825000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.680000 3.435000 10.820000 3.575000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.680000 3.575000 15.025000 3.645000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.695000 3.695000 10.930000 3.930000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.715000 9.880000 11.015000 9.950000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.720000 28.410000 11.125000 28.480000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.725000 26.750000 11.125000 26.820000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.790000 28.480000 11.125000 28.550000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.820000 3.435000 14.885000 3.695000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.865000 10.045000 11.125000 10.100000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.865000 10.100000 11.125000 26.610000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.865000 28.150000 11.125000 31.140000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.865000 28.620000 11.125000 28.625000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.865000 28.625000 11.125000 31.085000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.865000 31.140000 11.180000 31.195000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.865000 31.195000 11.125000 31.455000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.865000 9.730000 11.125000 9.990000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.865000 9.990000 11.125000 27.085000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.910000 27.085000 11.125000 27.300000 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.910000 27.935000 11.125000 28.150000 ;
    END
    PORT
      LAYER met2 ;
        RECT 11.005000 31.265000 11.305000 31.335000 ;
    END
    PORT
      LAYER met2 ;
        RECT 11.125000 31.085000 11.270000 31.230000 ;
    END
    PORT
      LAYER met2 ;
        RECT 11.125000 31.455000 11.260000 31.590000 ;
    END
    PORT
      LAYER met2 ;
        RECT 11.260000 31.480000 11.520000 36.020000 ;
    END
    PORT
      LAYER met2 ;
        RECT 11.260000 31.535000 11.520000 31.590000 ;
    END
    PORT
      LAYER met2 ;
        RECT 11.260000 36.020000 12.150000 36.280000 ;
    END
    PORT
      LAYER met2 ;
        RECT 11.270000 31.230000 11.495000 31.455000 ;
    END
    PORT
      LAYER met2 ;
        RECT 11.495000 31.455000 11.520000 31.480000 ;
    END
    PORT
      LAYER met2 ;
        RECT 14.775000 3.695000 14.875000 3.795000 ;
    END
    PORT
      LAYER met2 ;
        RECT 14.875000 3.795000 15.145000 4.065000 ;
    END
    PORT
      LAYER met2 ;
        RECT 14.885000 3.435000 15.245000 3.795000 ;
    END
    PORT
      LAYER met2 ;
        RECT 14.985000 3.835000 15.285000 3.905000 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.055000 3.905000 15.355000 3.975000 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.145000 4.065000 15.515000 4.435000 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.245000 3.795000 15.515000 4.065000 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.265000 4.115000 15.565000 4.185000 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.335000 4.185000 15.635000 4.255000 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.405000 4.255000 15.705000 4.325000 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.515000 4.065000 15.885000 4.435000 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.515000 4.435000 15.885000 4.805000 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.615000 4.465000 15.915000 4.535000 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.695000 4.545000 28.765000 4.615000 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.765000 4.615000 28.835000 4.685000 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.885000 4.435000 15.995000 4.545000 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.885000 4.755000 28.975000 4.805000 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.060000 4.245000 22.360000 4.545000 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.065000 4.540000 22.940000 4.545000 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.135000 4.470000 22.870000 4.540000 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.205000 4.400000 22.800000 4.470000 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.345000 4.260000 22.660000 4.330000 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.350000 4.255000 22.660000 4.260000 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.360000 0.000000 22.660000 4.245000 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.360000 1.170000 22.660000 4.805000 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.660000 4.260000 22.945000 4.545000 ;
    END
    PORT
      LAYER met2 ;
        RECT 28.655000 4.805000 28.750000 4.900000 ;
    END
    PORT
      LAYER met2 ;
        RECT 28.750000 4.900000 29.080000 5.230000 ;
    END
    PORT
      LAYER met2 ;
        RECT 28.765000 4.545000 29.120000 4.900000 ;
    END
    PORT
      LAYER met2 ;
        RECT 28.865000 4.945000 29.165000 5.015000 ;
    END
    PORT
      LAYER met2 ;
        RECT 28.935000 5.015000 29.235000 5.085000 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.005000 5.085000 29.305000 5.155000 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.080000 5.230000 29.320000 5.470000 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.120000 4.900000 29.450000 5.230000 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.320000 11.030000 29.635000 11.085000 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.320000 11.085000 29.400000 11.165000 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.320000 5.360000 29.580000 11.030000 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.320000 5.415000 29.580000 5.470000 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.320000 5.470000 29.580000 10.975000 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.400000 11.165000 29.770000 11.535000 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.450000 5.230000 29.580000 5.360000 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.530000 11.225000 29.830000 11.295000 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.580000 10.975000 29.770000 11.165000 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.600000 11.295000 29.900000 11.365000 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.770000 11.165000 30.030000 11.425000 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.770000 11.425000 30.030000 15.700000 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.770000 11.480000 30.030000 11.535000 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.770000 11.535000 30.030000 15.645000 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.770000 15.700000 30.085000 15.755000 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.770000 15.755000 29.995000 15.980000 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.840000 15.755000 30.140000 15.825000 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.910000 15.825000 30.210000 15.895000 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.995000 15.980000 30.365000 16.350000 ;
    END
    PORT
      LAYER met2 ;
        RECT 30.030000 15.645000 30.365000 15.980000 ;
    END
    PORT
      LAYER met2 ;
        RECT 30.120000 16.035000 30.420000 16.105000 ;
    END
    PORT
      LAYER met2 ;
        RECT 30.190000 16.105000 30.490000 16.175000 ;
    END
    PORT
      LAYER met2 ;
        RECT 30.365000 15.980000 30.625000 16.240000 ;
    END
    PORT
      LAYER met2 ;
        RECT 30.365000 16.240000 30.625000 16.350000 ;
    END
    PORT
      LAYER met2 ;
        RECT 30.365000 16.350000 30.625000 20.495000 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.735000 4.250000 10.005000 4.520000 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.735000 4.520000 10.050000 4.575000 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.735000 4.520000 9.995000 8.915000 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.735000 4.575000 9.995000 4.630000 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.735000 4.630000 9.995000 8.860000 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.735000 8.915000 10.050000 8.970000 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.735000 8.970000 9.965000 9.200000 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.790000 4.465000 10.105000 4.520000 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.805000 8.970000 10.105000 9.040000 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.860000 4.395000 10.160000 4.465000 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.875000 9.040000 10.175000 9.110000 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.930000 4.325000 10.230000 4.395000 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.965000 9.200000 10.165000 9.400000 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.995000 8.860000 10.335000 9.200000 ;
    END
  END EN_VDDIO_SIG_H
  PIN FILT_IN_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 20.075000 0.000000 21.225000 6.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.075000 3.410000 21.225000 6.820000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.075000 6.820000 21.375000 6.970000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.075000 6.970000 21.525000 7.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.075000 7.120000 21.675000 7.150000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.075000 7.150000 21.060000 8.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.225000 7.150000 21.705000 7.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.375000 7.300000 21.855000 7.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.525000 7.450000 22.005000 7.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.675000 7.600000 22.155000 7.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.825000 7.750000 22.305000 7.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.060000 8.135000 21.340000 8.415000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.225000 6.670000 22.690000 8.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.340000 8.415000 22.905000 9.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.575000 8.500000 23.055000 8.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.725000 8.650000 23.205000 8.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.875000 8.800000 23.355000 8.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 8.950000 23.505000 9.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.175000 9.100000 23.655000 9.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.325000 9.250000 23.805000 9.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.570000 9.495000 24.050000 9.645000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.690000 8.135000 22.970000 8.415000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.720000 9.645000 24.050000 9.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.905000 9.495000 24.050000 9.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.905000 9.980000 24.050000 12.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.970000 8.415000 24.050000 9.495000 ;
    END
  END FILT_IN_H
  PIN INP_SEL_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 24.905000 0.000000 25.135000 9.975000 ;
    END
  END INP_SEL_H
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 6.100000 104.010000 68.800000 166.625000 ;
    END
  END PAD
  PIN PAD_A_ESD_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 17.245000 0.000000 18.910000 3.135000 ;
    END
  END PAD_A_ESD_H
  PIN PULLUP_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.555000 0.000000 15.135000 0.985000 ;
    END
  END PULLUP_H
  PIN TIE_HI_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.505000 0.000000 31.155000 0.330000 ;
    END
  END TIE_HI_ESD
  PIN TIE_LO_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.580000 0.000000 28.230000 0.330000 ;
    END
  END TIE_LO_ESD
  PIN TIE_WEAK_HI_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.860000 70.750000 66.040000 71.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.860000 71.930000 65.990000 72.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.860000 71.930000 66.310000 72.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.860000 72.080000 66.160000 72.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.860000 72.400000 65.990000 94.645000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 71.800000 66.460000 71.930000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.140000 71.650000 66.590000 71.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.290000 71.500000 66.740000 71.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.440000 71.350000 66.890000 71.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590000 71.200000 67.040000 71.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990000 72.210000 66.180000 72.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.040000 69.400000 67.390000 70.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.040000 70.750000 67.490000 70.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180000 71.000000 67.390000 72.210000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.190000 70.600000 67.640000 70.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.340000 70.450000 67.790000 70.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.490000 70.300000 67.940000 70.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640000 70.150000 68.090000 70.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.940000 69.850000 68.390000 70.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.090000 69.700000 68.540000 69.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 68.535000 68.255000 69.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 69.400000 68.840000 69.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 70.035000 68.355000 71.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.540000 69.250000 68.990000 69.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.690000 69.100000 69.140000 69.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990000 68.800000 69.440000 68.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.255000 67.600000 69.190000 68.535000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290000 68.500000 69.740000 68.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.355000 69.085000 69.305000 70.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.440000 68.350000 69.890000 68.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.590000 68.200000 70.040000 68.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.740000 68.050000 70.190000 68.200000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 66.200000 70.590000 67.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190000 67.600000 70.640000 67.750000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.305000 67.800000 70.590000 69.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 67.450000 70.790000 67.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.490000 67.300000 70.940000 67.450000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.640000 67.150000 71.090000 67.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.790000 67.000000 71.240000 67.150000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.940000 66.850000 71.390000 67.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.090000 66.700000 71.540000 66.850000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.240000 66.550000 71.690000 66.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390000 66.400000 71.840000 66.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.590000 64.600000 72.190000 66.200000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.590000 66.200000 72.190000 67.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.840000 65.950000 72.290000 66.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.990000 65.800000 72.440000 65.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.140000 65.650000 72.590000 65.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.290000 65.500000 72.740000 65.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 65.350000 72.890000 65.500000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590000 65.200000 73.040000 65.350000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.740000 65.050000 73.190000 65.200000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.890000 64.900000 73.340000 65.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.190000 0.000000 73.260000 49.320000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.190000 0.725000 73.260000 49.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.190000 49.470000 73.410000 49.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.190000 49.620000 73.560000 49.770000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.190000 49.770000 73.710000 49.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.190000 49.985000 73.925000 64.465000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.190000 64.465000 73.860000 64.530000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.190000 64.465000 73.925000 66.200000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.190000 64.530000 73.795000 64.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.190000 64.595000 73.790000 64.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.260000 49.320000 73.925000 49.985000 ;
    END
  END TIE_WEAK_HI_H
  PIN XRES_H_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.170000 10.145000 28.635000 10.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.170000 10.610000 28.900000 10.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.170000 10.610000 29.050000 10.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.170000 10.910000 28.900000 14.770000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.185000 10.595000 29.200000 10.610000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.335000 10.445000 29.215000 10.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.635000 9.845000 28.935000 10.145000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.900000 10.145000 29.665000 10.910000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.935000 0.000000 29.665000 9.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.935000 4.005000 29.665000 10.145000 ;
    END
  END XRES_H_N
  PIN VCCD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT 0.000000 0.185000 75.000000 199.220000 ;
    LAYER met1 ;
      RECT  0.000000  0.000000 24.625000  10.255000 ;
      RECT  0.000000 10.255000 75.000000 199.210000 ;
      RECT 25.415000  0.000000 75.000000  10.255000 ;
    LAYER met2 ;
      RECT  0.340000  0.000000 12.005000   1.750000 ;
      RECT  0.340000  1.750000 22.080000   3.155000 ;
      RECT  0.340000  3.155000 10.400000   3.295000 ;
      RECT  0.340000  3.295000 10.070000   3.625000 ;
      RECT  0.340000  3.625000  9.725000   3.970000 ;
      RECT  0.340000  3.970000  9.455000   9.480000 ;
      RECT  0.340000  9.480000  9.685000   9.680000 ;
      RECT  0.340000  9.680000  9.885000  10.010000 ;
      RECT  0.340000 10.010000 10.215000  10.380000 ;
      RECT  0.340000 10.380000 10.585000  26.330000 ;
      RECT  0.340000 26.330000 10.370000  28.905000 ;
      RECT  0.340000 28.905000 10.585000  31.735000 ;
      RECT  0.340000 31.735000 10.845000  31.870000 ;
      RECT  0.340000 31.870000 10.980000  36.560000 ;
      RECT  0.340000 36.560000 74.915000 199.210000 ;
      RECT 10.275000  4.860000 15.235000   5.085000 ;
      RECT 10.275000  5.085000 28.375000   5.180000 ;
      RECT 10.275000  5.180000 28.470000   5.510000 ;
      RECT 10.275000  5.510000 28.800000   5.750000 ;
      RECT 10.275000  5.750000 29.040000   8.580000 ;
      RECT 10.615000  8.580000 29.040000   8.920000 ;
      RECT 10.655000  4.530000 14.865000   4.715000 ;
      RECT 10.655000  4.715000 15.235000   4.860000 ;
      RECT 10.815000  8.920000 29.040000   9.120000 ;
      RECT 10.975000  4.210000 14.595000   4.345000 ;
      RECT 10.975000  4.345000 14.865000   4.530000 ;
      RECT 11.145000  9.120000 29.040000   9.450000 ;
      RECT 11.190000 27.580000 74.915000  27.655000 ;
      RECT 11.210000  3.975000 14.495000   4.075000 ;
      RECT 11.210000  4.075000 14.595000   4.210000 ;
      RECT 11.405000  9.450000 29.040000  11.445000 ;
      RECT 11.405000 11.445000 29.120000  11.815000 ;
      RECT 11.405000 11.815000 29.490000  16.260000 ;
      RECT 11.405000 16.260000 29.715000  16.630000 ;
      RECT 11.405000 16.630000 30.085000  20.775000 ;
      RECT 11.405000 20.775000 74.915000  27.580000 ;
      RECT 11.405000 27.655000 74.915000  30.805000 ;
      RECT 11.550000 30.805000 74.915000  30.950000 ;
      RECT 11.775000 30.950000 74.915000  31.175000 ;
      RECT 11.800000 31.175000 74.915000  35.740000 ;
      RECT 12.430000 35.740000 74.915000  36.560000 ;
      RECT 12.825000  0.000000 14.275000   1.265000 ;
      RECT 12.825000  1.265000 22.080000   1.750000 ;
      RECT 15.415000  0.000000 22.080000   1.265000 ;
      RECT 15.525000  3.155000 22.080000   3.515000 ;
      RECT 15.795000  3.515000 22.080000   3.785000 ;
      RECT 16.165000  3.785000 22.080000   3.965000 ;
      RECT 16.165000  3.965000 21.780000   4.155000 ;
      RECT 16.275000  4.155000 21.780000   4.265000 ;
      RECT 22.940000  0.000000 27.300000   0.610000 ;
      RECT 22.940000  0.610000 32.480000   0.920000 ;
      RECT 22.940000  0.920000 74.915000   3.980000 ;
      RECT 23.225000  3.980000 74.915000   4.265000 ;
      RECT 28.510000  0.000000 30.225000   0.610000 ;
      RECT 29.400000  4.265000 74.915000   4.620000 ;
      RECT 29.730000  4.620000 74.915000   4.950000 ;
      RECT 29.860000  4.950000 74.915000  10.695000 ;
      RECT 30.050000 10.695000 74.915000  10.885000 ;
      RECT 30.310000 10.885000 74.915000  15.365000 ;
      RECT 30.645000 15.365000 74.915000  15.700000 ;
      RECT 30.905000 15.700000 74.915000  20.775000 ;
      RECT 31.435000  0.000000 32.480000   0.610000 ;
      RECT 33.300000  0.000000 74.915000   0.920000 ;
    LAYER met3 ;
      RECT  0.965000  0.625000  8.000000  15.385000 ;
      RECT  0.965000 15.385000  7.790000  15.595000 ;
      RECT  0.965000 15.595000  7.340000  16.045000 ;
      RECT  0.965000 16.045000  6.890000  16.495000 ;
      RECT  0.965000 16.495000  6.375000  32.280000 ;
      RECT  0.965000 32.280000  6.750000  32.995000 ;
      RECT  0.965000 32.995000  7.465000  33.580000 ;
      RECT  0.965000 33.580000  8.050000  34.100000 ;
      RECT  0.965000 34.100000  8.570000  34.525000 ;
      RECT  0.965000 34.525000 71.790000  64.200000 ;
      RECT  0.965000 64.200000 70.190000  65.800000 ;
      RECT  0.965000 65.800000 68.790000  67.200000 ;
      RECT  0.965000 67.200000 67.855000  68.135000 ;
      RECT  0.965000 68.135000 66.990000  69.000000 ;
      RECT  0.965000 69.000000 65.640000  70.350000 ;
      RECT  0.965000 70.350000 64.460000  95.045000 ;
      RECT  0.965000 95.045000 74.700000 200.000000 ;
      RECT  7.695000 18.020000 71.790000  30.895000 ;
      RECT  8.270000 17.445000 71.790000  18.020000 ;
      RECT  8.280000 30.895000 71.790000  31.480000 ;
      RECT  8.730000 16.985000 71.790000  17.445000 ;
      RECT  8.995000 31.480000 71.790000  32.195000 ;
      RECT  9.320000  0.625000 16.845000   3.535000 ;
      RECT  9.320000  3.535000 19.675000   8.535000 ;
      RECT  9.320000  8.535000 20.660000   8.815000 ;
      RECT  9.320000  8.815000 20.940000  10.380000 ;
      RECT  9.320000 10.380000 22.505000  12.665000 ;
      RECT  9.320000 12.665000 27.770000  15.170000 ;
      RECT  9.320000 15.170000 71.790000  16.985000 ;
      RECT  9.580000 32.195000 71.790000  32.780000 ;
      RECT  9.795000 32.780000 71.790000  32.995000 ;
      RECT 19.310000  0.625000 19.675000   3.535000 ;
      RECT 21.625000  0.625000 28.535000   6.270000 ;
      RECT 22.675000 32.995000 71.790000  34.525000 ;
      RECT 23.090000  6.270000 28.535000   7.735000 ;
      RECT 23.370000  7.735000 28.535000   8.015000 ;
      RECT 24.450000  8.015000 28.535000   9.445000 ;
      RECT 24.450000  9.445000 28.235000   9.745000 ;
      RECT 24.450000  9.745000 27.770000  12.665000 ;
      RECT 29.300000 11.310000 71.790000  15.170000 ;
      RECT 30.065000  0.625000 71.790000  11.310000 ;
      RECT 66.390000 72.800000 74.700000  95.045000 ;
      RECT 66.580000 72.610000 74.700000  72.800000 ;
      RECT 67.790000 71.400000 74.700000  72.610000 ;
      RECT 68.755000 70.435000 74.700000  71.400000 ;
      RECT 69.705000 69.485000 74.700000  70.435000 ;
      RECT 70.990000 68.200000 74.700000  69.485000 ;
      RECT 72.590000 66.600000 74.700000  68.200000 ;
      RECT 73.660000  0.625000 74.700000  48.920000 ;
      RECT 74.325000 48.920000 74.700000  66.600000 ;
    LAYER met4 ;
      RECT 0.000000  2.035000 75.000000  47.965000 ;
      RECT 0.000000 51.745000 75.000000  52.725000 ;
      RECT 0.000000 56.505000 75.000000 200.000000 ;
    LAYER met5 ;
      RECT  0.000000   2.135000 72.130000  15.035000 ;
      RECT  0.000000  15.035000 72.435000  19.885000 ;
      RECT  0.000000  19.885000 75.000000  24.335000 ;
      RECT  0.000000  24.335000 72.130000  36.835000 ;
      RECT  0.000000  36.835000 75.000000  40.085000 ;
      RECT  0.000000  40.085000 72.130000  96.585000 ;
      RECT  0.000000  96.585000 75.000000 102.410000 ;
      RECT  0.000000 102.410000  4.500000 168.225000 ;
      RECT  0.000000 168.225000 75.000000 200.000000 ;
      RECT 70.400000 102.410000 75.000000 168.225000 ;
  END
END sky130_fd_io__top_xres4v2
END LIBRARY
