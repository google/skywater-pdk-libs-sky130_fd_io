# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__overlay_vddio_lvc
  CLASS PAD ;
  FOREIGN sky130_fd_io__overlay_vddio_lvc ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  75.00000 BY  198.0000 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.630000 17.800000 0.950000 18.120000 ;
      LAYER met4 ;
        RECT 0.630000 17.800000 0.950000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 18.230000 0.950000 18.550000 ;
      LAYER met4 ;
        RECT 0.630000 18.230000 0.950000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 18.660000 0.950000 18.980000 ;
      LAYER met4 ;
        RECT 0.630000 18.660000 0.950000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 19.090000 0.950000 19.410000 ;
      LAYER met4 ;
        RECT 0.630000 19.090000 0.950000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 19.520000 0.950000 19.840000 ;
      LAYER met4 ;
        RECT 0.630000 19.520000 0.950000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 19.950000 0.950000 20.270000 ;
      LAYER met4 ;
        RECT 0.630000 19.950000 0.950000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 20.380000 0.950000 20.700000 ;
      LAYER met4 ;
        RECT 0.630000 20.380000 0.950000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 20.810000 0.950000 21.130000 ;
      LAYER met4 ;
        RECT 0.630000 20.810000 0.950000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 21.240000 0.950000 21.560000 ;
      LAYER met4 ;
        RECT 0.630000 21.240000 0.950000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 21.670000 0.950000 21.990000 ;
      LAYER met4 ;
        RECT 0.630000 21.670000 0.950000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 22.100000 0.950000 22.420000 ;
      LAYER met4 ;
        RECT 0.630000 22.100000 0.950000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 82.795000 0.995000 83.115000 ;
      LAYER met4 ;
        RECT 0.675000 82.795000 0.995000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 83.205000 0.995000 83.525000 ;
      LAYER met4 ;
        RECT 0.675000 83.205000 0.995000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 83.615000 0.995000 83.935000 ;
      LAYER met4 ;
        RECT 0.675000 83.615000 0.995000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 84.025000 0.995000 84.345000 ;
      LAYER met4 ;
        RECT 0.675000 84.025000 0.995000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 84.435000 0.995000 84.755000 ;
      LAYER met4 ;
        RECT 0.675000 84.435000 0.995000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 84.845000 0.995000 85.165000 ;
      LAYER met4 ;
        RECT 0.675000 84.845000 0.995000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 85.255000 0.995000 85.575000 ;
      LAYER met4 ;
        RECT 0.675000 85.255000 0.995000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 85.665000 0.995000 85.985000 ;
      LAYER met4 ;
        RECT 0.675000 85.665000 0.995000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 86.075000 0.995000 86.395000 ;
      LAYER met4 ;
        RECT 0.675000 86.075000 0.995000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 86.485000 0.995000 86.805000 ;
      LAYER met4 ;
        RECT 0.675000 86.485000 0.995000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 86.895000 0.995000 87.215000 ;
      LAYER met4 ;
        RECT 0.675000 86.895000 0.995000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 87.305000 0.995000 87.625000 ;
      LAYER met4 ;
        RECT 0.675000 87.305000 0.995000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 87.715000 0.995000 88.035000 ;
      LAYER met4 ;
        RECT 0.675000 87.715000 0.995000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 88.125000 0.995000 88.445000 ;
      LAYER met4 ;
        RECT 0.675000 88.125000 0.995000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 88.535000 0.995000 88.855000 ;
      LAYER met4 ;
        RECT 0.675000 88.535000 0.995000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 88.945000 0.995000 89.265000 ;
      LAYER met4 ;
        RECT 0.675000 88.945000 0.995000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 89.355000 0.995000 89.675000 ;
      LAYER met4 ;
        RECT 0.675000 89.355000 0.995000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 89.765000 0.995000 90.085000 ;
      LAYER met4 ;
        RECT 0.675000 89.765000 0.995000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 90.175000 0.995000 90.495000 ;
      LAYER met4 ;
        RECT 0.675000 90.175000 0.995000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 90.585000 0.995000 90.905000 ;
      LAYER met4 ;
        RECT 0.675000 90.585000 0.995000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 90.995000 0.995000 91.315000 ;
      LAYER met4 ;
        RECT 0.675000 90.995000 0.995000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 91.405000 0.995000 91.725000 ;
      LAYER met4 ;
        RECT 0.675000 91.405000 0.995000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 91.815000 0.995000 92.135000 ;
      LAYER met4 ;
        RECT 0.675000 91.815000 0.995000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 92.225000 0.995000 92.545000 ;
      LAYER met4 ;
        RECT 0.675000 92.225000 0.995000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675000 92.635000 0.995000 92.955000 ;
      LAYER met4 ;
        RECT 0.675000 92.635000 0.995000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 68.065000 1.105000 68.385000 ;
      LAYER met4 ;
        RECT 0.785000 68.065000 1.105000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 68.475000 1.105000 68.795000 ;
      LAYER met4 ;
        RECT 0.785000 68.475000 1.105000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 68.885000 1.105000 69.205000 ;
      LAYER met4 ;
        RECT 0.785000 68.885000 1.105000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 69.295000 1.105000 69.615000 ;
      LAYER met4 ;
        RECT 0.785000 69.295000 1.105000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 69.705000 1.105000 70.025000 ;
      LAYER met4 ;
        RECT 0.785000 69.705000 1.105000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 70.115000 1.105000 70.435000 ;
      LAYER met4 ;
        RECT 0.785000 70.115000 1.105000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 70.525000 1.105000 70.845000 ;
      LAYER met4 ;
        RECT 0.785000 70.525000 1.105000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 70.935000 1.105000 71.255000 ;
      LAYER met4 ;
        RECT 0.785000 70.935000 1.105000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 71.345000 1.105000 71.665000 ;
      LAYER met4 ;
        RECT 0.785000 71.345000 1.105000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 71.755000 1.105000 72.075000 ;
      LAYER met4 ;
        RECT 0.785000 71.755000 1.105000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 72.165000 1.105000 72.485000 ;
      LAYER met4 ;
        RECT 0.785000 72.165000 1.105000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 72.575000 1.105000 72.895000 ;
      LAYER met4 ;
        RECT 0.785000 72.575000 1.105000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 72.985000 1.105000 73.305000 ;
      LAYER met4 ;
        RECT 0.785000 72.985000 1.105000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 73.390000 1.105000 73.710000 ;
      LAYER met4 ;
        RECT 0.785000 73.390000 1.105000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 73.795000 1.105000 74.115000 ;
      LAYER met4 ;
        RECT 0.785000 73.795000 1.105000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 74.200000 1.105000 74.520000 ;
      LAYER met4 ;
        RECT 0.785000 74.200000 1.105000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 74.605000 1.105000 74.925000 ;
      LAYER met4 ;
        RECT 0.785000 74.605000 1.105000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 75.010000 1.105000 75.330000 ;
      LAYER met4 ;
        RECT 0.785000 75.010000 1.105000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 75.415000 1.105000 75.735000 ;
      LAYER met4 ;
        RECT 0.785000 75.415000 1.105000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 75.820000 1.105000 76.140000 ;
      LAYER met4 ;
        RECT 0.785000 75.820000 1.105000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 76.225000 1.105000 76.545000 ;
      LAYER met4 ;
        RECT 0.785000 76.225000 1.105000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 76.630000 1.105000 76.950000 ;
      LAYER met4 ;
        RECT 0.785000 76.630000 1.105000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 77.035000 1.105000 77.355000 ;
      LAYER met4 ;
        RECT 0.785000 77.035000 1.105000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 77.440000 1.105000 77.760000 ;
      LAYER met4 ;
        RECT 0.785000 77.440000 1.105000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 77.845000 1.105000 78.165000 ;
      LAYER met4 ;
        RECT 0.785000 77.845000 1.105000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 78.250000 1.105000 78.570000 ;
      LAYER met4 ;
        RECT 0.785000 78.250000 1.105000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 78.655000 1.105000 78.975000 ;
      LAYER met4 ;
        RECT 0.785000 78.655000 1.105000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 79.060000 1.105000 79.380000 ;
      LAYER met4 ;
        RECT 0.785000 79.060000 1.105000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 79.465000 1.105000 79.785000 ;
      LAYER met4 ;
        RECT 0.785000 79.465000 1.105000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 79.870000 1.105000 80.190000 ;
      LAYER met4 ;
        RECT 0.785000 79.870000 1.105000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 80.275000 1.105000 80.595000 ;
      LAYER met4 ;
        RECT 0.785000 80.275000 1.105000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 80.680000 1.105000 81.000000 ;
      LAYER met4 ;
        RECT 0.785000 80.680000 1.105000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 81.085000 1.105000 81.405000 ;
      LAYER met4 ;
        RECT 0.785000 81.085000 1.105000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 81.490000 1.105000 81.810000 ;
      LAYER met4 ;
        RECT 0.785000 81.490000 1.105000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 81.895000 1.105000 82.215000 ;
      LAYER met4 ;
        RECT 0.785000 81.895000 1.105000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785000 82.300000 1.105000 82.620000 ;
      LAYER met4 ;
        RECT 0.785000 82.300000 1.105000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035000 17.800000 1.355000 18.120000 ;
      LAYER met4 ;
        RECT 1.035000 17.800000 1.355000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035000 18.230000 1.355000 18.550000 ;
      LAYER met4 ;
        RECT 1.035000 18.230000 1.355000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035000 18.660000 1.355000 18.980000 ;
      LAYER met4 ;
        RECT 1.035000 18.660000 1.355000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035000 19.090000 1.355000 19.410000 ;
      LAYER met4 ;
        RECT 1.035000 19.090000 1.355000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035000 19.520000 1.355000 19.840000 ;
      LAYER met4 ;
        RECT 1.035000 19.520000 1.355000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035000 19.950000 1.355000 20.270000 ;
      LAYER met4 ;
        RECT 1.035000 19.950000 1.355000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035000 20.380000 1.355000 20.700000 ;
      LAYER met4 ;
        RECT 1.035000 20.380000 1.355000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035000 20.810000 1.355000 21.130000 ;
      LAYER met4 ;
        RECT 1.035000 20.810000 1.355000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035000 21.240000 1.355000 21.560000 ;
      LAYER met4 ;
        RECT 1.035000 21.240000 1.355000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035000 21.670000 1.355000 21.990000 ;
      LAYER met4 ;
        RECT 1.035000 21.670000 1.355000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035000 22.100000 1.355000 22.420000 ;
      LAYER met4 ;
        RECT 1.035000 22.100000 1.355000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 82.795000 1.405000 83.115000 ;
      LAYER met4 ;
        RECT 1.085000 82.795000 1.405000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 83.205000 1.405000 83.525000 ;
      LAYER met4 ;
        RECT 1.085000 83.205000 1.405000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 83.615000 1.405000 83.935000 ;
      LAYER met4 ;
        RECT 1.085000 83.615000 1.405000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 84.025000 1.405000 84.345000 ;
      LAYER met4 ;
        RECT 1.085000 84.025000 1.405000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 84.435000 1.405000 84.755000 ;
      LAYER met4 ;
        RECT 1.085000 84.435000 1.405000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 84.845000 1.405000 85.165000 ;
      LAYER met4 ;
        RECT 1.085000 84.845000 1.405000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 85.255000 1.405000 85.575000 ;
      LAYER met4 ;
        RECT 1.085000 85.255000 1.405000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 85.665000 1.405000 85.985000 ;
      LAYER met4 ;
        RECT 1.085000 85.665000 1.405000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 86.075000 1.405000 86.395000 ;
      LAYER met4 ;
        RECT 1.085000 86.075000 1.405000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 86.485000 1.405000 86.805000 ;
      LAYER met4 ;
        RECT 1.085000 86.485000 1.405000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 86.895000 1.405000 87.215000 ;
      LAYER met4 ;
        RECT 1.085000 86.895000 1.405000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 87.305000 1.405000 87.625000 ;
      LAYER met4 ;
        RECT 1.085000 87.305000 1.405000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 87.715000 1.405000 88.035000 ;
      LAYER met4 ;
        RECT 1.085000 87.715000 1.405000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 88.125000 1.405000 88.445000 ;
      LAYER met4 ;
        RECT 1.085000 88.125000 1.405000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 88.535000 1.405000 88.855000 ;
      LAYER met4 ;
        RECT 1.085000 88.535000 1.405000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 88.945000 1.405000 89.265000 ;
      LAYER met4 ;
        RECT 1.085000 88.945000 1.405000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 89.355000 1.405000 89.675000 ;
      LAYER met4 ;
        RECT 1.085000 89.355000 1.405000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 89.765000 1.405000 90.085000 ;
      LAYER met4 ;
        RECT 1.085000 89.765000 1.405000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 90.175000 1.405000 90.495000 ;
      LAYER met4 ;
        RECT 1.085000 90.175000 1.405000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 90.585000 1.405000 90.905000 ;
      LAYER met4 ;
        RECT 1.085000 90.585000 1.405000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 90.995000 1.405000 91.315000 ;
      LAYER met4 ;
        RECT 1.085000 90.995000 1.405000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 91.405000 1.405000 91.725000 ;
      LAYER met4 ;
        RECT 1.085000 91.405000 1.405000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 91.815000 1.405000 92.135000 ;
      LAYER met4 ;
        RECT 1.085000 91.815000 1.405000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 92.225000 1.405000 92.545000 ;
      LAYER met4 ;
        RECT 1.085000 92.225000 1.405000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085000 92.635000 1.405000 92.955000 ;
      LAYER met4 ;
        RECT 1.085000 92.635000 1.405000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 68.065000 1.505000 68.385000 ;
      LAYER met4 ;
        RECT 1.185000 68.065000 1.505000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 68.475000 1.505000 68.795000 ;
      LAYER met4 ;
        RECT 1.185000 68.475000 1.505000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 68.885000 1.505000 69.205000 ;
      LAYER met4 ;
        RECT 1.185000 68.885000 1.505000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 69.295000 1.505000 69.615000 ;
      LAYER met4 ;
        RECT 1.185000 69.295000 1.505000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 69.705000 1.505000 70.025000 ;
      LAYER met4 ;
        RECT 1.185000 69.705000 1.505000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 70.115000 1.505000 70.435000 ;
      LAYER met4 ;
        RECT 1.185000 70.115000 1.505000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 70.525000 1.505000 70.845000 ;
      LAYER met4 ;
        RECT 1.185000 70.525000 1.505000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 70.935000 1.505000 71.255000 ;
      LAYER met4 ;
        RECT 1.185000 70.935000 1.505000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 71.345000 1.505000 71.665000 ;
      LAYER met4 ;
        RECT 1.185000 71.345000 1.505000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 71.755000 1.505000 72.075000 ;
      LAYER met4 ;
        RECT 1.185000 71.755000 1.505000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 72.165000 1.505000 72.485000 ;
      LAYER met4 ;
        RECT 1.185000 72.165000 1.505000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 72.575000 1.505000 72.895000 ;
      LAYER met4 ;
        RECT 1.185000 72.575000 1.505000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 72.985000 1.505000 73.305000 ;
      LAYER met4 ;
        RECT 1.185000 72.985000 1.505000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 73.390000 1.505000 73.710000 ;
      LAYER met4 ;
        RECT 1.185000 73.390000 1.505000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 73.795000 1.505000 74.115000 ;
      LAYER met4 ;
        RECT 1.185000 73.795000 1.505000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 74.200000 1.505000 74.520000 ;
      LAYER met4 ;
        RECT 1.185000 74.200000 1.505000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 74.605000 1.505000 74.925000 ;
      LAYER met4 ;
        RECT 1.185000 74.605000 1.505000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 75.010000 1.505000 75.330000 ;
      LAYER met4 ;
        RECT 1.185000 75.010000 1.505000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 75.415000 1.505000 75.735000 ;
      LAYER met4 ;
        RECT 1.185000 75.415000 1.505000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 75.820000 1.505000 76.140000 ;
      LAYER met4 ;
        RECT 1.185000 75.820000 1.505000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 76.225000 1.505000 76.545000 ;
      LAYER met4 ;
        RECT 1.185000 76.225000 1.505000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 76.630000 1.505000 76.950000 ;
      LAYER met4 ;
        RECT 1.185000 76.630000 1.505000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 77.035000 1.505000 77.355000 ;
      LAYER met4 ;
        RECT 1.185000 77.035000 1.505000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 77.440000 1.505000 77.760000 ;
      LAYER met4 ;
        RECT 1.185000 77.440000 1.505000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 77.845000 1.505000 78.165000 ;
      LAYER met4 ;
        RECT 1.185000 77.845000 1.505000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 78.250000 1.505000 78.570000 ;
      LAYER met4 ;
        RECT 1.185000 78.250000 1.505000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 78.655000 1.505000 78.975000 ;
      LAYER met4 ;
        RECT 1.185000 78.655000 1.505000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 79.060000 1.505000 79.380000 ;
      LAYER met4 ;
        RECT 1.185000 79.060000 1.505000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 79.465000 1.505000 79.785000 ;
      LAYER met4 ;
        RECT 1.185000 79.465000 1.505000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 79.870000 1.505000 80.190000 ;
      LAYER met4 ;
        RECT 1.185000 79.870000 1.505000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 80.275000 1.505000 80.595000 ;
      LAYER met4 ;
        RECT 1.185000 80.275000 1.505000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 80.680000 1.505000 81.000000 ;
      LAYER met4 ;
        RECT 1.185000 80.680000 1.505000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 81.085000 1.505000 81.405000 ;
      LAYER met4 ;
        RECT 1.185000 81.085000 1.505000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 81.490000 1.505000 81.810000 ;
      LAYER met4 ;
        RECT 1.185000 81.490000 1.505000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 81.895000 1.505000 82.215000 ;
      LAYER met4 ;
        RECT 1.185000 81.895000 1.505000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185000 82.300000 1.505000 82.620000 ;
      LAYER met4 ;
        RECT 1.185000 82.300000 1.505000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440000 17.800000 1.760000 18.120000 ;
      LAYER met4 ;
        RECT 1.440000 17.800000 1.760000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440000 18.230000 1.760000 18.550000 ;
      LAYER met4 ;
        RECT 1.440000 18.230000 1.760000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440000 18.660000 1.760000 18.980000 ;
      LAYER met4 ;
        RECT 1.440000 18.660000 1.760000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440000 19.090000 1.760000 19.410000 ;
      LAYER met4 ;
        RECT 1.440000 19.090000 1.760000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440000 19.520000 1.760000 19.840000 ;
      LAYER met4 ;
        RECT 1.440000 19.520000 1.760000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440000 19.950000 1.760000 20.270000 ;
      LAYER met4 ;
        RECT 1.440000 19.950000 1.760000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440000 20.380000 1.760000 20.700000 ;
      LAYER met4 ;
        RECT 1.440000 20.380000 1.760000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440000 20.810000 1.760000 21.130000 ;
      LAYER met4 ;
        RECT 1.440000 20.810000 1.760000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440000 21.240000 1.760000 21.560000 ;
      LAYER met4 ;
        RECT 1.440000 21.240000 1.760000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440000 21.670000 1.760000 21.990000 ;
      LAYER met4 ;
        RECT 1.440000 21.670000 1.760000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440000 22.100000 1.760000 22.420000 ;
      LAYER met4 ;
        RECT 1.440000 22.100000 1.760000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 82.795000 1.815000 83.115000 ;
      LAYER met4 ;
        RECT 1.495000 82.795000 1.815000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 83.205000 1.815000 83.525000 ;
      LAYER met4 ;
        RECT 1.495000 83.205000 1.815000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 83.615000 1.815000 83.935000 ;
      LAYER met4 ;
        RECT 1.495000 83.615000 1.815000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 84.025000 1.815000 84.345000 ;
      LAYER met4 ;
        RECT 1.495000 84.025000 1.815000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 84.435000 1.815000 84.755000 ;
      LAYER met4 ;
        RECT 1.495000 84.435000 1.815000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 84.845000 1.815000 85.165000 ;
      LAYER met4 ;
        RECT 1.495000 84.845000 1.815000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 85.255000 1.815000 85.575000 ;
      LAYER met4 ;
        RECT 1.495000 85.255000 1.815000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 85.665000 1.815000 85.985000 ;
      LAYER met4 ;
        RECT 1.495000 85.665000 1.815000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 86.075000 1.815000 86.395000 ;
      LAYER met4 ;
        RECT 1.495000 86.075000 1.815000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 86.485000 1.815000 86.805000 ;
      LAYER met4 ;
        RECT 1.495000 86.485000 1.815000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 86.895000 1.815000 87.215000 ;
      LAYER met4 ;
        RECT 1.495000 86.895000 1.815000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 87.305000 1.815000 87.625000 ;
      LAYER met4 ;
        RECT 1.495000 87.305000 1.815000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 87.715000 1.815000 88.035000 ;
      LAYER met4 ;
        RECT 1.495000 87.715000 1.815000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 88.125000 1.815000 88.445000 ;
      LAYER met4 ;
        RECT 1.495000 88.125000 1.815000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 88.535000 1.815000 88.855000 ;
      LAYER met4 ;
        RECT 1.495000 88.535000 1.815000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 88.945000 1.815000 89.265000 ;
      LAYER met4 ;
        RECT 1.495000 88.945000 1.815000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 89.355000 1.815000 89.675000 ;
      LAYER met4 ;
        RECT 1.495000 89.355000 1.815000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 89.765000 1.815000 90.085000 ;
      LAYER met4 ;
        RECT 1.495000 89.765000 1.815000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 90.175000 1.815000 90.495000 ;
      LAYER met4 ;
        RECT 1.495000 90.175000 1.815000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 90.585000 1.815000 90.905000 ;
      LAYER met4 ;
        RECT 1.495000 90.585000 1.815000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 90.995000 1.815000 91.315000 ;
      LAYER met4 ;
        RECT 1.495000 90.995000 1.815000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 91.405000 1.815000 91.725000 ;
      LAYER met4 ;
        RECT 1.495000 91.405000 1.815000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 91.815000 1.815000 92.135000 ;
      LAYER met4 ;
        RECT 1.495000 91.815000 1.815000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 92.225000 1.815000 92.545000 ;
      LAYER met4 ;
        RECT 1.495000 92.225000 1.815000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495000 92.635000 1.815000 92.955000 ;
      LAYER met4 ;
        RECT 1.495000 92.635000 1.815000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 68.065000 1.905000 68.385000 ;
      LAYER met4 ;
        RECT 1.585000 68.065000 1.905000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 68.475000 1.905000 68.795000 ;
      LAYER met4 ;
        RECT 1.585000 68.475000 1.905000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 68.885000 1.905000 69.205000 ;
      LAYER met4 ;
        RECT 1.585000 68.885000 1.905000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 69.295000 1.905000 69.615000 ;
      LAYER met4 ;
        RECT 1.585000 69.295000 1.905000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 69.705000 1.905000 70.025000 ;
      LAYER met4 ;
        RECT 1.585000 69.705000 1.905000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 70.115000 1.905000 70.435000 ;
      LAYER met4 ;
        RECT 1.585000 70.115000 1.905000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 70.525000 1.905000 70.845000 ;
      LAYER met4 ;
        RECT 1.585000 70.525000 1.905000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 70.935000 1.905000 71.255000 ;
      LAYER met4 ;
        RECT 1.585000 70.935000 1.905000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 71.345000 1.905000 71.665000 ;
      LAYER met4 ;
        RECT 1.585000 71.345000 1.905000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 71.755000 1.905000 72.075000 ;
      LAYER met4 ;
        RECT 1.585000 71.755000 1.905000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 72.165000 1.905000 72.485000 ;
      LAYER met4 ;
        RECT 1.585000 72.165000 1.905000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 72.575000 1.905000 72.895000 ;
      LAYER met4 ;
        RECT 1.585000 72.575000 1.905000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 72.985000 1.905000 73.305000 ;
      LAYER met4 ;
        RECT 1.585000 72.985000 1.905000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 73.390000 1.905000 73.710000 ;
      LAYER met4 ;
        RECT 1.585000 73.390000 1.905000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 73.795000 1.905000 74.115000 ;
      LAYER met4 ;
        RECT 1.585000 73.795000 1.905000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 74.200000 1.905000 74.520000 ;
      LAYER met4 ;
        RECT 1.585000 74.200000 1.905000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 74.605000 1.905000 74.925000 ;
      LAYER met4 ;
        RECT 1.585000 74.605000 1.905000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 75.010000 1.905000 75.330000 ;
      LAYER met4 ;
        RECT 1.585000 75.010000 1.905000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 75.415000 1.905000 75.735000 ;
      LAYER met4 ;
        RECT 1.585000 75.415000 1.905000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 75.820000 1.905000 76.140000 ;
      LAYER met4 ;
        RECT 1.585000 75.820000 1.905000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 76.225000 1.905000 76.545000 ;
      LAYER met4 ;
        RECT 1.585000 76.225000 1.905000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 76.630000 1.905000 76.950000 ;
      LAYER met4 ;
        RECT 1.585000 76.630000 1.905000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 77.035000 1.905000 77.355000 ;
      LAYER met4 ;
        RECT 1.585000 77.035000 1.905000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 77.440000 1.905000 77.760000 ;
      LAYER met4 ;
        RECT 1.585000 77.440000 1.905000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 77.845000 1.905000 78.165000 ;
      LAYER met4 ;
        RECT 1.585000 77.845000 1.905000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 78.250000 1.905000 78.570000 ;
      LAYER met4 ;
        RECT 1.585000 78.250000 1.905000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 78.655000 1.905000 78.975000 ;
      LAYER met4 ;
        RECT 1.585000 78.655000 1.905000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 79.060000 1.905000 79.380000 ;
      LAYER met4 ;
        RECT 1.585000 79.060000 1.905000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 79.465000 1.905000 79.785000 ;
      LAYER met4 ;
        RECT 1.585000 79.465000 1.905000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 79.870000 1.905000 80.190000 ;
      LAYER met4 ;
        RECT 1.585000 79.870000 1.905000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 80.275000 1.905000 80.595000 ;
      LAYER met4 ;
        RECT 1.585000 80.275000 1.905000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 80.680000 1.905000 81.000000 ;
      LAYER met4 ;
        RECT 1.585000 80.680000 1.905000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 81.085000 1.905000 81.405000 ;
      LAYER met4 ;
        RECT 1.585000 81.085000 1.905000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 81.490000 1.905000 81.810000 ;
      LAYER met4 ;
        RECT 1.585000 81.490000 1.905000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 81.895000 1.905000 82.215000 ;
      LAYER met4 ;
        RECT 1.585000 81.895000 1.905000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585000 82.300000 1.905000 82.620000 ;
      LAYER met4 ;
        RECT 1.585000 82.300000 1.905000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845000 17.800000 2.165000 18.120000 ;
      LAYER met4 ;
        RECT 1.845000 17.800000 2.165000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845000 18.230000 2.165000 18.550000 ;
      LAYER met4 ;
        RECT 1.845000 18.230000 2.165000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845000 18.660000 2.165000 18.980000 ;
      LAYER met4 ;
        RECT 1.845000 18.660000 2.165000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845000 19.090000 2.165000 19.410000 ;
      LAYER met4 ;
        RECT 1.845000 19.090000 2.165000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845000 19.520000 2.165000 19.840000 ;
      LAYER met4 ;
        RECT 1.845000 19.520000 2.165000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845000 19.950000 2.165000 20.270000 ;
      LAYER met4 ;
        RECT 1.845000 19.950000 2.165000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845000 20.380000 2.165000 20.700000 ;
      LAYER met4 ;
        RECT 1.845000 20.380000 2.165000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845000 20.810000 2.165000 21.130000 ;
      LAYER met4 ;
        RECT 1.845000 20.810000 2.165000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845000 21.240000 2.165000 21.560000 ;
      LAYER met4 ;
        RECT 1.845000 21.240000 2.165000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845000 21.670000 2.165000 21.990000 ;
      LAYER met4 ;
        RECT 1.845000 21.670000 2.165000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845000 22.100000 2.165000 22.420000 ;
      LAYER met4 ;
        RECT 1.845000 22.100000 2.165000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 82.795000 2.225000 83.115000 ;
      LAYER met4 ;
        RECT 1.905000 82.795000 2.225000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 83.205000 2.225000 83.525000 ;
      LAYER met4 ;
        RECT 1.905000 83.205000 2.225000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 83.615000 2.225000 83.935000 ;
      LAYER met4 ;
        RECT 1.905000 83.615000 2.225000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 84.025000 2.225000 84.345000 ;
      LAYER met4 ;
        RECT 1.905000 84.025000 2.225000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 84.435000 2.225000 84.755000 ;
      LAYER met4 ;
        RECT 1.905000 84.435000 2.225000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 84.845000 2.225000 85.165000 ;
      LAYER met4 ;
        RECT 1.905000 84.845000 2.225000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 85.255000 2.225000 85.575000 ;
      LAYER met4 ;
        RECT 1.905000 85.255000 2.225000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 85.665000 2.225000 85.985000 ;
      LAYER met4 ;
        RECT 1.905000 85.665000 2.225000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 86.075000 2.225000 86.395000 ;
      LAYER met4 ;
        RECT 1.905000 86.075000 2.225000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 86.485000 2.225000 86.805000 ;
      LAYER met4 ;
        RECT 1.905000 86.485000 2.225000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 86.895000 2.225000 87.215000 ;
      LAYER met4 ;
        RECT 1.905000 86.895000 2.225000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 87.305000 2.225000 87.625000 ;
      LAYER met4 ;
        RECT 1.905000 87.305000 2.225000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 87.715000 2.225000 88.035000 ;
      LAYER met4 ;
        RECT 1.905000 87.715000 2.225000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 88.125000 2.225000 88.445000 ;
      LAYER met4 ;
        RECT 1.905000 88.125000 2.225000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 88.535000 2.225000 88.855000 ;
      LAYER met4 ;
        RECT 1.905000 88.535000 2.225000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 88.945000 2.225000 89.265000 ;
      LAYER met4 ;
        RECT 1.905000 88.945000 2.225000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 89.355000 2.225000 89.675000 ;
      LAYER met4 ;
        RECT 1.905000 89.355000 2.225000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 89.765000 2.225000 90.085000 ;
      LAYER met4 ;
        RECT 1.905000 89.765000 2.225000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 90.175000 2.225000 90.495000 ;
      LAYER met4 ;
        RECT 1.905000 90.175000 2.225000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 90.585000 2.225000 90.905000 ;
      LAYER met4 ;
        RECT 1.905000 90.585000 2.225000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 90.995000 2.225000 91.315000 ;
      LAYER met4 ;
        RECT 1.905000 90.995000 2.225000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 91.405000 2.225000 91.725000 ;
      LAYER met4 ;
        RECT 1.905000 91.405000 2.225000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 91.815000 2.225000 92.135000 ;
      LAYER met4 ;
        RECT 1.905000 91.815000 2.225000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 92.225000 2.225000 92.545000 ;
      LAYER met4 ;
        RECT 1.905000 92.225000 2.225000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905000 92.635000 2.225000 92.955000 ;
      LAYER met4 ;
        RECT 1.905000 92.635000 2.225000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 68.065000 2.305000 68.385000 ;
      LAYER met4 ;
        RECT 1.985000 68.065000 2.305000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 68.475000 2.305000 68.795000 ;
      LAYER met4 ;
        RECT 1.985000 68.475000 2.305000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 68.885000 2.305000 69.205000 ;
      LAYER met4 ;
        RECT 1.985000 68.885000 2.305000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 69.295000 2.305000 69.615000 ;
      LAYER met4 ;
        RECT 1.985000 69.295000 2.305000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 69.705000 2.305000 70.025000 ;
      LAYER met4 ;
        RECT 1.985000 69.705000 2.305000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 70.115000 2.305000 70.435000 ;
      LAYER met4 ;
        RECT 1.985000 70.115000 2.305000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 70.525000 2.305000 70.845000 ;
      LAYER met4 ;
        RECT 1.985000 70.525000 2.305000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 70.935000 2.305000 71.255000 ;
      LAYER met4 ;
        RECT 1.985000 70.935000 2.305000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 71.345000 2.305000 71.665000 ;
      LAYER met4 ;
        RECT 1.985000 71.345000 2.305000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 71.755000 2.305000 72.075000 ;
      LAYER met4 ;
        RECT 1.985000 71.755000 2.305000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 72.165000 2.305000 72.485000 ;
      LAYER met4 ;
        RECT 1.985000 72.165000 2.305000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 72.575000 2.305000 72.895000 ;
      LAYER met4 ;
        RECT 1.985000 72.575000 2.305000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 72.985000 2.305000 73.305000 ;
      LAYER met4 ;
        RECT 1.985000 72.985000 2.305000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 73.390000 2.305000 73.710000 ;
      LAYER met4 ;
        RECT 1.985000 73.390000 2.305000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 73.795000 2.305000 74.115000 ;
      LAYER met4 ;
        RECT 1.985000 73.795000 2.305000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 74.200000 2.305000 74.520000 ;
      LAYER met4 ;
        RECT 1.985000 74.200000 2.305000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 74.605000 2.305000 74.925000 ;
      LAYER met4 ;
        RECT 1.985000 74.605000 2.305000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 75.010000 2.305000 75.330000 ;
      LAYER met4 ;
        RECT 1.985000 75.010000 2.305000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 75.415000 2.305000 75.735000 ;
      LAYER met4 ;
        RECT 1.985000 75.415000 2.305000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 75.820000 2.305000 76.140000 ;
      LAYER met4 ;
        RECT 1.985000 75.820000 2.305000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 76.225000 2.305000 76.545000 ;
      LAYER met4 ;
        RECT 1.985000 76.225000 2.305000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 76.630000 2.305000 76.950000 ;
      LAYER met4 ;
        RECT 1.985000 76.630000 2.305000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 77.035000 2.305000 77.355000 ;
      LAYER met4 ;
        RECT 1.985000 77.035000 2.305000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 77.440000 2.305000 77.760000 ;
      LAYER met4 ;
        RECT 1.985000 77.440000 2.305000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 77.845000 2.305000 78.165000 ;
      LAYER met4 ;
        RECT 1.985000 77.845000 2.305000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 78.250000 2.305000 78.570000 ;
      LAYER met4 ;
        RECT 1.985000 78.250000 2.305000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 78.655000 2.305000 78.975000 ;
      LAYER met4 ;
        RECT 1.985000 78.655000 2.305000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 79.060000 2.305000 79.380000 ;
      LAYER met4 ;
        RECT 1.985000 79.060000 2.305000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 79.465000 2.305000 79.785000 ;
      LAYER met4 ;
        RECT 1.985000 79.465000 2.305000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 79.870000 2.305000 80.190000 ;
      LAYER met4 ;
        RECT 1.985000 79.870000 2.305000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 80.275000 2.305000 80.595000 ;
      LAYER met4 ;
        RECT 1.985000 80.275000 2.305000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 80.680000 2.305000 81.000000 ;
      LAYER met4 ;
        RECT 1.985000 80.680000 2.305000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 81.085000 2.305000 81.405000 ;
      LAYER met4 ;
        RECT 1.985000 81.085000 2.305000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 81.490000 2.305000 81.810000 ;
      LAYER met4 ;
        RECT 1.985000 81.490000 2.305000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 81.895000 2.305000 82.215000 ;
      LAYER met4 ;
        RECT 1.985000 81.895000 2.305000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985000 82.300000 2.305000 82.620000 ;
      LAYER met4 ;
        RECT 1.985000 82.300000 2.305000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 82.795000 10.425000 83.115000 ;
      LAYER met4 ;
        RECT 10.105000 82.795000 10.425000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 83.205000 10.425000 83.525000 ;
      LAYER met4 ;
        RECT 10.105000 83.205000 10.425000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 83.615000 10.425000 83.935000 ;
      LAYER met4 ;
        RECT 10.105000 83.615000 10.425000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 84.025000 10.425000 84.345000 ;
      LAYER met4 ;
        RECT 10.105000 84.025000 10.425000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 84.435000 10.425000 84.755000 ;
      LAYER met4 ;
        RECT 10.105000 84.435000 10.425000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 84.845000 10.425000 85.165000 ;
      LAYER met4 ;
        RECT 10.105000 84.845000 10.425000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 85.255000 10.425000 85.575000 ;
      LAYER met4 ;
        RECT 10.105000 85.255000 10.425000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 85.665000 10.425000 85.985000 ;
      LAYER met4 ;
        RECT 10.105000 85.665000 10.425000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 86.075000 10.425000 86.395000 ;
      LAYER met4 ;
        RECT 10.105000 86.075000 10.425000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 86.485000 10.425000 86.805000 ;
      LAYER met4 ;
        RECT 10.105000 86.485000 10.425000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 86.895000 10.425000 87.215000 ;
      LAYER met4 ;
        RECT 10.105000 86.895000 10.425000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 87.305000 10.425000 87.625000 ;
      LAYER met4 ;
        RECT 10.105000 87.305000 10.425000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 87.715000 10.425000 88.035000 ;
      LAYER met4 ;
        RECT 10.105000 87.715000 10.425000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 88.125000 10.425000 88.445000 ;
      LAYER met4 ;
        RECT 10.105000 88.125000 10.425000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 88.535000 10.425000 88.855000 ;
      LAYER met4 ;
        RECT 10.105000 88.535000 10.425000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 88.945000 10.425000 89.265000 ;
      LAYER met4 ;
        RECT 10.105000 88.945000 10.425000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 89.355000 10.425000 89.675000 ;
      LAYER met4 ;
        RECT 10.105000 89.355000 10.425000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 89.765000 10.425000 90.085000 ;
      LAYER met4 ;
        RECT 10.105000 89.765000 10.425000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 90.175000 10.425000 90.495000 ;
      LAYER met4 ;
        RECT 10.105000 90.175000 10.425000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 90.585000 10.425000 90.905000 ;
      LAYER met4 ;
        RECT 10.105000 90.585000 10.425000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 90.995000 10.425000 91.315000 ;
      LAYER met4 ;
        RECT 10.105000 90.995000 10.425000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 91.405000 10.425000 91.725000 ;
      LAYER met4 ;
        RECT 10.105000 91.405000 10.425000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 91.815000 10.425000 92.135000 ;
      LAYER met4 ;
        RECT 10.105000 91.815000 10.425000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 92.225000 10.425000 92.545000 ;
      LAYER met4 ;
        RECT 10.105000 92.225000 10.425000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105000 92.635000 10.425000 92.955000 ;
      LAYER met4 ;
        RECT 10.105000 92.635000 10.425000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350000 17.800000 10.670000 18.120000 ;
      LAYER met4 ;
        RECT 10.350000 17.800000 10.670000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350000 18.230000 10.670000 18.550000 ;
      LAYER met4 ;
        RECT 10.350000 18.230000 10.670000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350000 18.660000 10.670000 18.980000 ;
      LAYER met4 ;
        RECT 10.350000 18.660000 10.670000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350000 19.090000 10.670000 19.410000 ;
      LAYER met4 ;
        RECT 10.350000 19.090000 10.670000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350000 19.520000 10.670000 19.840000 ;
      LAYER met4 ;
        RECT 10.350000 19.520000 10.670000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350000 19.950000 10.670000 20.270000 ;
      LAYER met4 ;
        RECT 10.350000 19.950000 10.670000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350000 20.380000 10.670000 20.700000 ;
      LAYER met4 ;
        RECT 10.350000 20.380000 10.670000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350000 20.810000 10.670000 21.130000 ;
      LAYER met4 ;
        RECT 10.350000 20.810000 10.670000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350000 21.240000 10.670000 21.560000 ;
      LAYER met4 ;
        RECT 10.350000 21.240000 10.670000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350000 21.670000 10.670000 21.990000 ;
      LAYER met4 ;
        RECT 10.350000 21.670000 10.670000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350000 22.100000 10.670000 22.420000 ;
      LAYER met4 ;
        RECT 10.350000 22.100000 10.670000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 68.065000 10.705000 68.385000 ;
      LAYER met4 ;
        RECT 10.385000 68.065000 10.705000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 68.475000 10.705000 68.795000 ;
      LAYER met4 ;
        RECT 10.385000 68.475000 10.705000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 68.885000 10.705000 69.205000 ;
      LAYER met4 ;
        RECT 10.385000 68.885000 10.705000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 69.295000 10.705000 69.615000 ;
      LAYER met4 ;
        RECT 10.385000 69.295000 10.705000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 69.705000 10.705000 70.025000 ;
      LAYER met4 ;
        RECT 10.385000 69.705000 10.705000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 70.115000 10.705000 70.435000 ;
      LAYER met4 ;
        RECT 10.385000 70.115000 10.705000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 70.525000 10.705000 70.845000 ;
      LAYER met4 ;
        RECT 10.385000 70.525000 10.705000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 70.935000 10.705000 71.255000 ;
      LAYER met4 ;
        RECT 10.385000 70.935000 10.705000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 71.345000 10.705000 71.665000 ;
      LAYER met4 ;
        RECT 10.385000 71.345000 10.705000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 71.755000 10.705000 72.075000 ;
      LAYER met4 ;
        RECT 10.385000 71.755000 10.705000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 72.165000 10.705000 72.485000 ;
      LAYER met4 ;
        RECT 10.385000 72.165000 10.705000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 72.575000 10.705000 72.895000 ;
      LAYER met4 ;
        RECT 10.385000 72.575000 10.705000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 72.985000 10.705000 73.305000 ;
      LAYER met4 ;
        RECT 10.385000 72.985000 10.705000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 73.390000 10.705000 73.710000 ;
      LAYER met4 ;
        RECT 10.385000 73.390000 10.705000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 73.795000 10.705000 74.115000 ;
      LAYER met4 ;
        RECT 10.385000 73.795000 10.705000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 74.200000 10.705000 74.520000 ;
      LAYER met4 ;
        RECT 10.385000 74.200000 10.705000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 74.605000 10.705000 74.925000 ;
      LAYER met4 ;
        RECT 10.385000 74.605000 10.705000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 75.010000 10.705000 75.330000 ;
      LAYER met4 ;
        RECT 10.385000 75.010000 10.705000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 75.415000 10.705000 75.735000 ;
      LAYER met4 ;
        RECT 10.385000 75.415000 10.705000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 75.820000 10.705000 76.140000 ;
      LAYER met4 ;
        RECT 10.385000 75.820000 10.705000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 76.225000 10.705000 76.545000 ;
      LAYER met4 ;
        RECT 10.385000 76.225000 10.705000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 76.630000 10.705000 76.950000 ;
      LAYER met4 ;
        RECT 10.385000 76.630000 10.705000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 77.035000 10.705000 77.355000 ;
      LAYER met4 ;
        RECT 10.385000 77.035000 10.705000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 77.440000 10.705000 77.760000 ;
      LAYER met4 ;
        RECT 10.385000 77.440000 10.705000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 77.845000 10.705000 78.165000 ;
      LAYER met4 ;
        RECT 10.385000 77.845000 10.705000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 78.250000 10.705000 78.570000 ;
      LAYER met4 ;
        RECT 10.385000 78.250000 10.705000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 78.655000 10.705000 78.975000 ;
      LAYER met4 ;
        RECT 10.385000 78.655000 10.705000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 79.060000 10.705000 79.380000 ;
      LAYER met4 ;
        RECT 10.385000 79.060000 10.705000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 79.465000 10.705000 79.785000 ;
      LAYER met4 ;
        RECT 10.385000 79.465000 10.705000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 79.870000 10.705000 80.190000 ;
      LAYER met4 ;
        RECT 10.385000 79.870000 10.705000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 80.275000 10.705000 80.595000 ;
      LAYER met4 ;
        RECT 10.385000 80.275000 10.705000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 80.680000 10.705000 81.000000 ;
      LAYER met4 ;
        RECT 10.385000 80.680000 10.705000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 81.085000 10.705000 81.405000 ;
      LAYER met4 ;
        RECT 10.385000 81.085000 10.705000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 81.490000 10.705000 81.810000 ;
      LAYER met4 ;
        RECT 10.385000 81.490000 10.705000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 81.895000 10.705000 82.215000 ;
      LAYER met4 ;
        RECT 10.385000 81.895000 10.705000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385000 82.300000 10.705000 82.620000 ;
      LAYER met4 ;
        RECT 10.385000 82.300000 10.705000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 82.795000 10.835000 83.115000 ;
      LAYER met4 ;
        RECT 10.515000 82.795000 10.835000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 83.205000 10.835000 83.525000 ;
      LAYER met4 ;
        RECT 10.515000 83.205000 10.835000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 83.615000 10.835000 83.935000 ;
      LAYER met4 ;
        RECT 10.515000 83.615000 10.835000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 84.025000 10.835000 84.345000 ;
      LAYER met4 ;
        RECT 10.515000 84.025000 10.835000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 84.435000 10.835000 84.755000 ;
      LAYER met4 ;
        RECT 10.515000 84.435000 10.835000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 84.845000 10.835000 85.165000 ;
      LAYER met4 ;
        RECT 10.515000 84.845000 10.835000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 85.255000 10.835000 85.575000 ;
      LAYER met4 ;
        RECT 10.515000 85.255000 10.835000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 85.665000 10.835000 85.985000 ;
      LAYER met4 ;
        RECT 10.515000 85.665000 10.835000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 86.075000 10.835000 86.395000 ;
      LAYER met4 ;
        RECT 10.515000 86.075000 10.835000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 86.485000 10.835000 86.805000 ;
      LAYER met4 ;
        RECT 10.515000 86.485000 10.835000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 86.895000 10.835000 87.215000 ;
      LAYER met4 ;
        RECT 10.515000 86.895000 10.835000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 87.305000 10.835000 87.625000 ;
      LAYER met4 ;
        RECT 10.515000 87.305000 10.835000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 87.715000 10.835000 88.035000 ;
      LAYER met4 ;
        RECT 10.515000 87.715000 10.835000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 88.125000 10.835000 88.445000 ;
      LAYER met4 ;
        RECT 10.515000 88.125000 10.835000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 88.535000 10.835000 88.855000 ;
      LAYER met4 ;
        RECT 10.515000 88.535000 10.835000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 88.945000 10.835000 89.265000 ;
      LAYER met4 ;
        RECT 10.515000 88.945000 10.835000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 89.355000 10.835000 89.675000 ;
      LAYER met4 ;
        RECT 10.515000 89.355000 10.835000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 89.765000 10.835000 90.085000 ;
      LAYER met4 ;
        RECT 10.515000 89.765000 10.835000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 90.175000 10.835000 90.495000 ;
      LAYER met4 ;
        RECT 10.515000 90.175000 10.835000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 90.585000 10.835000 90.905000 ;
      LAYER met4 ;
        RECT 10.515000 90.585000 10.835000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 90.995000 10.835000 91.315000 ;
      LAYER met4 ;
        RECT 10.515000 90.995000 10.835000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 91.405000 10.835000 91.725000 ;
      LAYER met4 ;
        RECT 10.515000 91.405000 10.835000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 91.815000 10.835000 92.135000 ;
      LAYER met4 ;
        RECT 10.515000 91.815000 10.835000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 92.225000 10.835000 92.545000 ;
      LAYER met4 ;
        RECT 10.515000 92.225000 10.835000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515000 92.635000 10.835000 92.955000 ;
      LAYER met4 ;
        RECT 10.515000 92.635000 10.835000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755000 17.800000 11.075000 18.120000 ;
      LAYER met4 ;
        RECT 10.755000 17.800000 11.075000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755000 18.230000 11.075000 18.550000 ;
      LAYER met4 ;
        RECT 10.755000 18.230000 11.075000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755000 18.660000 11.075000 18.980000 ;
      LAYER met4 ;
        RECT 10.755000 18.660000 11.075000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755000 19.090000 11.075000 19.410000 ;
      LAYER met4 ;
        RECT 10.755000 19.090000 11.075000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755000 19.520000 11.075000 19.840000 ;
      LAYER met4 ;
        RECT 10.755000 19.520000 11.075000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755000 19.950000 11.075000 20.270000 ;
      LAYER met4 ;
        RECT 10.755000 19.950000 11.075000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755000 20.380000 11.075000 20.700000 ;
      LAYER met4 ;
        RECT 10.755000 20.380000 11.075000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755000 20.810000 11.075000 21.130000 ;
      LAYER met4 ;
        RECT 10.755000 20.810000 11.075000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755000 21.240000 11.075000 21.560000 ;
      LAYER met4 ;
        RECT 10.755000 21.240000 11.075000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755000 21.670000 11.075000 21.990000 ;
      LAYER met4 ;
        RECT 10.755000 21.670000 11.075000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755000 22.100000 11.075000 22.420000 ;
      LAYER met4 ;
        RECT 10.755000 22.100000 11.075000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 68.065000 11.105000 68.385000 ;
      LAYER met4 ;
        RECT 10.785000 68.065000 11.105000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 68.475000 11.105000 68.795000 ;
      LAYER met4 ;
        RECT 10.785000 68.475000 11.105000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 68.885000 11.105000 69.205000 ;
      LAYER met4 ;
        RECT 10.785000 68.885000 11.105000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 69.295000 11.105000 69.615000 ;
      LAYER met4 ;
        RECT 10.785000 69.295000 11.105000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 69.705000 11.105000 70.025000 ;
      LAYER met4 ;
        RECT 10.785000 69.705000 11.105000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 70.115000 11.105000 70.435000 ;
      LAYER met4 ;
        RECT 10.785000 70.115000 11.105000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 70.525000 11.105000 70.845000 ;
      LAYER met4 ;
        RECT 10.785000 70.525000 11.105000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 70.935000 11.105000 71.255000 ;
      LAYER met4 ;
        RECT 10.785000 70.935000 11.105000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 71.345000 11.105000 71.665000 ;
      LAYER met4 ;
        RECT 10.785000 71.345000 11.105000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 71.755000 11.105000 72.075000 ;
      LAYER met4 ;
        RECT 10.785000 71.755000 11.105000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 72.165000 11.105000 72.485000 ;
      LAYER met4 ;
        RECT 10.785000 72.165000 11.105000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 72.575000 11.105000 72.895000 ;
      LAYER met4 ;
        RECT 10.785000 72.575000 11.105000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 72.985000 11.105000 73.305000 ;
      LAYER met4 ;
        RECT 10.785000 72.985000 11.105000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 73.390000 11.105000 73.710000 ;
      LAYER met4 ;
        RECT 10.785000 73.390000 11.105000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 73.795000 11.105000 74.115000 ;
      LAYER met4 ;
        RECT 10.785000 73.795000 11.105000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 74.200000 11.105000 74.520000 ;
      LAYER met4 ;
        RECT 10.785000 74.200000 11.105000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 74.605000 11.105000 74.925000 ;
      LAYER met4 ;
        RECT 10.785000 74.605000 11.105000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 75.010000 11.105000 75.330000 ;
      LAYER met4 ;
        RECT 10.785000 75.010000 11.105000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 75.415000 11.105000 75.735000 ;
      LAYER met4 ;
        RECT 10.785000 75.415000 11.105000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 75.820000 11.105000 76.140000 ;
      LAYER met4 ;
        RECT 10.785000 75.820000 11.105000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 76.225000 11.105000 76.545000 ;
      LAYER met4 ;
        RECT 10.785000 76.225000 11.105000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 76.630000 11.105000 76.950000 ;
      LAYER met4 ;
        RECT 10.785000 76.630000 11.105000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 77.035000 11.105000 77.355000 ;
      LAYER met4 ;
        RECT 10.785000 77.035000 11.105000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 77.440000 11.105000 77.760000 ;
      LAYER met4 ;
        RECT 10.785000 77.440000 11.105000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 77.845000 11.105000 78.165000 ;
      LAYER met4 ;
        RECT 10.785000 77.845000 11.105000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 78.250000 11.105000 78.570000 ;
      LAYER met4 ;
        RECT 10.785000 78.250000 11.105000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 78.655000 11.105000 78.975000 ;
      LAYER met4 ;
        RECT 10.785000 78.655000 11.105000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 79.060000 11.105000 79.380000 ;
      LAYER met4 ;
        RECT 10.785000 79.060000 11.105000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 79.465000 11.105000 79.785000 ;
      LAYER met4 ;
        RECT 10.785000 79.465000 11.105000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 79.870000 11.105000 80.190000 ;
      LAYER met4 ;
        RECT 10.785000 79.870000 11.105000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 80.275000 11.105000 80.595000 ;
      LAYER met4 ;
        RECT 10.785000 80.275000 11.105000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 80.680000 11.105000 81.000000 ;
      LAYER met4 ;
        RECT 10.785000 80.680000 11.105000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 81.085000 11.105000 81.405000 ;
      LAYER met4 ;
        RECT 10.785000 81.085000 11.105000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 81.490000 11.105000 81.810000 ;
      LAYER met4 ;
        RECT 10.785000 81.490000 11.105000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 81.895000 11.105000 82.215000 ;
      LAYER met4 ;
        RECT 10.785000 81.895000 11.105000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 82.300000 11.105000 82.620000 ;
      LAYER met4 ;
        RECT 10.785000 82.300000 11.105000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 82.795000 11.245000 83.115000 ;
      LAYER met4 ;
        RECT 10.925000 82.795000 11.245000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 83.205000 11.245000 83.525000 ;
      LAYER met4 ;
        RECT 10.925000 83.205000 11.245000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 83.615000 11.245000 83.935000 ;
      LAYER met4 ;
        RECT 10.925000 83.615000 11.245000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 84.025000 11.245000 84.345000 ;
      LAYER met4 ;
        RECT 10.925000 84.025000 11.245000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 84.435000 11.245000 84.755000 ;
      LAYER met4 ;
        RECT 10.925000 84.435000 11.245000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 84.845000 11.245000 85.165000 ;
      LAYER met4 ;
        RECT 10.925000 84.845000 11.245000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 85.255000 11.245000 85.575000 ;
      LAYER met4 ;
        RECT 10.925000 85.255000 11.245000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 85.665000 11.245000 85.985000 ;
      LAYER met4 ;
        RECT 10.925000 85.665000 11.245000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 86.075000 11.245000 86.395000 ;
      LAYER met4 ;
        RECT 10.925000 86.075000 11.245000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 86.485000 11.245000 86.805000 ;
      LAYER met4 ;
        RECT 10.925000 86.485000 11.245000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 86.895000 11.245000 87.215000 ;
      LAYER met4 ;
        RECT 10.925000 86.895000 11.245000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 87.305000 11.245000 87.625000 ;
      LAYER met4 ;
        RECT 10.925000 87.305000 11.245000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 87.715000 11.245000 88.035000 ;
      LAYER met4 ;
        RECT 10.925000 87.715000 11.245000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 88.125000 11.245000 88.445000 ;
      LAYER met4 ;
        RECT 10.925000 88.125000 11.245000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 88.535000 11.245000 88.855000 ;
      LAYER met4 ;
        RECT 10.925000 88.535000 11.245000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 88.945000 11.245000 89.265000 ;
      LAYER met4 ;
        RECT 10.925000 88.945000 11.245000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 89.355000 11.245000 89.675000 ;
      LAYER met4 ;
        RECT 10.925000 89.355000 11.245000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 89.765000 11.245000 90.085000 ;
      LAYER met4 ;
        RECT 10.925000 89.765000 11.245000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 90.175000 11.245000 90.495000 ;
      LAYER met4 ;
        RECT 10.925000 90.175000 11.245000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 90.585000 11.245000 90.905000 ;
      LAYER met4 ;
        RECT 10.925000 90.585000 11.245000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 90.995000 11.245000 91.315000 ;
      LAYER met4 ;
        RECT 10.925000 90.995000 11.245000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 91.405000 11.245000 91.725000 ;
      LAYER met4 ;
        RECT 10.925000 91.405000 11.245000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 91.815000 11.245000 92.135000 ;
      LAYER met4 ;
        RECT 10.925000 91.815000 11.245000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 92.225000 11.245000 92.545000 ;
      LAYER met4 ;
        RECT 10.925000 92.225000 11.245000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925000 92.635000 11.245000 92.955000 ;
      LAYER met4 ;
        RECT 10.925000 92.635000 11.245000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160000 17.800000 11.480000 18.120000 ;
      LAYER met4 ;
        RECT 11.160000 17.800000 11.480000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160000 18.230000 11.480000 18.550000 ;
      LAYER met4 ;
        RECT 11.160000 18.230000 11.480000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160000 18.660000 11.480000 18.980000 ;
      LAYER met4 ;
        RECT 11.160000 18.660000 11.480000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160000 19.090000 11.480000 19.410000 ;
      LAYER met4 ;
        RECT 11.160000 19.090000 11.480000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160000 19.520000 11.480000 19.840000 ;
      LAYER met4 ;
        RECT 11.160000 19.520000 11.480000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160000 19.950000 11.480000 20.270000 ;
      LAYER met4 ;
        RECT 11.160000 19.950000 11.480000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160000 20.380000 11.480000 20.700000 ;
      LAYER met4 ;
        RECT 11.160000 20.380000 11.480000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160000 20.810000 11.480000 21.130000 ;
      LAYER met4 ;
        RECT 11.160000 20.810000 11.480000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160000 21.240000 11.480000 21.560000 ;
      LAYER met4 ;
        RECT 11.160000 21.240000 11.480000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160000 21.670000 11.480000 21.990000 ;
      LAYER met4 ;
        RECT 11.160000 21.670000 11.480000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160000 22.100000 11.480000 22.420000 ;
      LAYER met4 ;
        RECT 11.160000 22.100000 11.480000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 68.065000 11.505000 68.385000 ;
      LAYER met4 ;
        RECT 11.185000 68.065000 11.505000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 68.475000 11.505000 68.795000 ;
      LAYER met4 ;
        RECT 11.185000 68.475000 11.505000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 68.885000 11.505000 69.205000 ;
      LAYER met4 ;
        RECT 11.185000 68.885000 11.505000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 69.295000 11.505000 69.615000 ;
      LAYER met4 ;
        RECT 11.185000 69.295000 11.505000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 69.705000 11.505000 70.025000 ;
      LAYER met4 ;
        RECT 11.185000 69.705000 11.505000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 70.115000 11.505000 70.435000 ;
      LAYER met4 ;
        RECT 11.185000 70.115000 11.505000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 70.525000 11.505000 70.845000 ;
      LAYER met4 ;
        RECT 11.185000 70.525000 11.505000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 70.935000 11.505000 71.255000 ;
      LAYER met4 ;
        RECT 11.185000 70.935000 11.505000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 71.345000 11.505000 71.665000 ;
      LAYER met4 ;
        RECT 11.185000 71.345000 11.505000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 71.755000 11.505000 72.075000 ;
      LAYER met4 ;
        RECT 11.185000 71.755000 11.505000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 72.165000 11.505000 72.485000 ;
      LAYER met4 ;
        RECT 11.185000 72.165000 11.505000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 72.575000 11.505000 72.895000 ;
      LAYER met4 ;
        RECT 11.185000 72.575000 11.505000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 72.985000 11.505000 73.305000 ;
      LAYER met4 ;
        RECT 11.185000 72.985000 11.505000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 73.390000 11.505000 73.710000 ;
      LAYER met4 ;
        RECT 11.185000 73.390000 11.505000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 73.795000 11.505000 74.115000 ;
      LAYER met4 ;
        RECT 11.185000 73.795000 11.505000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 74.200000 11.505000 74.520000 ;
      LAYER met4 ;
        RECT 11.185000 74.200000 11.505000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 74.605000 11.505000 74.925000 ;
      LAYER met4 ;
        RECT 11.185000 74.605000 11.505000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 75.010000 11.505000 75.330000 ;
      LAYER met4 ;
        RECT 11.185000 75.010000 11.505000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 75.415000 11.505000 75.735000 ;
      LAYER met4 ;
        RECT 11.185000 75.415000 11.505000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 75.820000 11.505000 76.140000 ;
      LAYER met4 ;
        RECT 11.185000 75.820000 11.505000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 76.225000 11.505000 76.545000 ;
      LAYER met4 ;
        RECT 11.185000 76.225000 11.505000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 76.630000 11.505000 76.950000 ;
      LAYER met4 ;
        RECT 11.185000 76.630000 11.505000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 77.035000 11.505000 77.355000 ;
      LAYER met4 ;
        RECT 11.185000 77.035000 11.505000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 77.440000 11.505000 77.760000 ;
      LAYER met4 ;
        RECT 11.185000 77.440000 11.505000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 77.845000 11.505000 78.165000 ;
      LAYER met4 ;
        RECT 11.185000 77.845000 11.505000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 78.250000 11.505000 78.570000 ;
      LAYER met4 ;
        RECT 11.185000 78.250000 11.505000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 78.655000 11.505000 78.975000 ;
      LAYER met4 ;
        RECT 11.185000 78.655000 11.505000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 79.060000 11.505000 79.380000 ;
      LAYER met4 ;
        RECT 11.185000 79.060000 11.505000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 79.465000 11.505000 79.785000 ;
      LAYER met4 ;
        RECT 11.185000 79.465000 11.505000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 79.870000 11.505000 80.190000 ;
      LAYER met4 ;
        RECT 11.185000 79.870000 11.505000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 80.275000 11.505000 80.595000 ;
      LAYER met4 ;
        RECT 11.185000 80.275000 11.505000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 80.680000 11.505000 81.000000 ;
      LAYER met4 ;
        RECT 11.185000 80.680000 11.505000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 81.085000 11.505000 81.405000 ;
      LAYER met4 ;
        RECT 11.185000 81.085000 11.505000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 81.490000 11.505000 81.810000 ;
      LAYER met4 ;
        RECT 11.185000 81.490000 11.505000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 81.895000 11.505000 82.215000 ;
      LAYER met4 ;
        RECT 11.185000 81.895000 11.505000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185000 82.300000 11.505000 82.620000 ;
      LAYER met4 ;
        RECT 11.185000 82.300000 11.505000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 82.795000 11.655000 83.115000 ;
      LAYER met4 ;
        RECT 11.335000 82.795000 11.655000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 83.205000 11.655000 83.525000 ;
      LAYER met4 ;
        RECT 11.335000 83.205000 11.655000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 83.615000 11.655000 83.935000 ;
      LAYER met4 ;
        RECT 11.335000 83.615000 11.655000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 84.025000 11.655000 84.345000 ;
      LAYER met4 ;
        RECT 11.335000 84.025000 11.655000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 84.435000 11.655000 84.755000 ;
      LAYER met4 ;
        RECT 11.335000 84.435000 11.655000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 84.845000 11.655000 85.165000 ;
      LAYER met4 ;
        RECT 11.335000 84.845000 11.655000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 85.255000 11.655000 85.575000 ;
      LAYER met4 ;
        RECT 11.335000 85.255000 11.655000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 85.665000 11.655000 85.985000 ;
      LAYER met4 ;
        RECT 11.335000 85.665000 11.655000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 86.075000 11.655000 86.395000 ;
      LAYER met4 ;
        RECT 11.335000 86.075000 11.655000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 86.485000 11.655000 86.805000 ;
      LAYER met4 ;
        RECT 11.335000 86.485000 11.655000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 86.895000 11.655000 87.215000 ;
      LAYER met4 ;
        RECT 11.335000 86.895000 11.655000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 87.305000 11.655000 87.625000 ;
      LAYER met4 ;
        RECT 11.335000 87.305000 11.655000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 87.715000 11.655000 88.035000 ;
      LAYER met4 ;
        RECT 11.335000 87.715000 11.655000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 88.125000 11.655000 88.445000 ;
      LAYER met4 ;
        RECT 11.335000 88.125000 11.655000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 88.535000 11.655000 88.855000 ;
      LAYER met4 ;
        RECT 11.335000 88.535000 11.655000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 88.945000 11.655000 89.265000 ;
      LAYER met4 ;
        RECT 11.335000 88.945000 11.655000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 89.355000 11.655000 89.675000 ;
      LAYER met4 ;
        RECT 11.335000 89.355000 11.655000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 89.765000 11.655000 90.085000 ;
      LAYER met4 ;
        RECT 11.335000 89.765000 11.655000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 90.175000 11.655000 90.495000 ;
      LAYER met4 ;
        RECT 11.335000 90.175000 11.655000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 90.585000 11.655000 90.905000 ;
      LAYER met4 ;
        RECT 11.335000 90.585000 11.655000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 90.995000 11.655000 91.315000 ;
      LAYER met4 ;
        RECT 11.335000 90.995000 11.655000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 91.405000 11.655000 91.725000 ;
      LAYER met4 ;
        RECT 11.335000 91.405000 11.655000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 91.815000 11.655000 92.135000 ;
      LAYER met4 ;
        RECT 11.335000 91.815000 11.655000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 92.225000 11.655000 92.545000 ;
      LAYER met4 ;
        RECT 11.335000 92.225000 11.655000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335000 92.635000 11.655000 92.955000 ;
      LAYER met4 ;
        RECT 11.335000 92.635000 11.655000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565000 17.800000 11.885000 18.120000 ;
      LAYER met4 ;
        RECT 11.565000 17.800000 11.885000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565000 18.230000 11.885000 18.550000 ;
      LAYER met4 ;
        RECT 11.565000 18.230000 11.885000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565000 18.660000 11.885000 18.980000 ;
      LAYER met4 ;
        RECT 11.565000 18.660000 11.885000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565000 19.090000 11.885000 19.410000 ;
      LAYER met4 ;
        RECT 11.565000 19.090000 11.885000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565000 19.520000 11.885000 19.840000 ;
      LAYER met4 ;
        RECT 11.565000 19.520000 11.885000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565000 19.950000 11.885000 20.270000 ;
      LAYER met4 ;
        RECT 11.565000 19.950000 11.885000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565000 20.380000 11.885000 20.700000 ;
      LAYER met4 ;
        RECT 11.565000 20.380000 11.885000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565000 20.810000 11.885000 21.130000 ;
      LAYER met4 ;
        RECT 11.565000 20.810000 11.885000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565000 21.240000 11.885000 21.560000 ;
      LAYER met4 ;
        RECT 11.565000 21.240000 11.885000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565000 21.670000 11.885000 21.990000 ;
      LAYER met4 ;
        RECT 11.565000 21.670000 11.885000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565000 22.100000 11.885000 22.420000 ;
      LAYER met4 ;
        RECT 11.565000 22.100000 11.885000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 68.065000 11.905000 68.385000 ;
      LAYER met4 ;
        RECT 11.585000 68.065000 11.905000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 68.475000 11.905000 68.795000 ;
      LAYER met4 ;
        RECT 11.585000 68.475000 11.905000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 68.885000 11.905000 69.205000 ;
      LAYER met4 ;
        RECT 11.585000 68.885000 11.905000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 69.295000 11.905000 69.615000 ;
      LAYER met4 ;
        RECT 11.585000 69.295000 11.905000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 69.705000 11.905000 70.025000 ;
      LAYER met4 ;
        RECT 11.585000 69.705000 11.905000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 70.115000 11.905000 70.435000 ;
      LAYER met4 ;
        RECT 11.585000 70.115000 11.905000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 70.525000 11.905000 70.845000 ;
      LAYER met4 ;
        RECT 11.585000 70.525000 11.905000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 70.935000 11.905000 71.255000 ;
      LAYER met4 ;
        RECT 11.585000 70.935000 11.905000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 71.345000 11.905000 71.665000 ;
      LAYER met4 ;
        RECT 11.585000 71.345000 11.905000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 71.755000 11.905000 72.075000 ;
      LAYER met4 ;
        RECT 11.585000 71.755000 11.905000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 72.165000 11.905000 72.485000 ;
      LAYER met4 ;
        RECT 11.585000 72.165000 11.905000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 72.575000 11.905000 72.895000 ;
      LAYER met4 ;
        RECT 11.585000 72.575000 11.905000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 72.985000 11.905000 73.305000 ;
      LAYER met4 ;
        RECT 11.585000 72.985000 11.905000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 73.390000 11.905000 73.710000 ;
      LAYER met4 ;
        RECT 11.585000 73.390000 11.905000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 73.795000 11.905000 74.115000 ;
      LAYER met4 ;
        RECT 11.585000 73.795000 11.905000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 74.200000 11.905000 74.520000 ;
      LAYER met4 ;
        RECT 11.585000 74.200000 11.905000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 74.605000 11.905000 74.925000 ;
      LAYER met4 ;
        RECT 11.585000 74.605000 11.905000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 75.010000 11.905000 75.330000 ;
      LAYER met4 ;
        RECT 11.585000 75.010000 11.905000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 75.415000 11.905000 75.735000 ;
      LAYER met4 ;
        RECT 11.585000 75.415000 11.905000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 75.820000 11.905000 76.140000 ;
      LAYER met4 ;
        RECT 11.585000 75.820000 11.905000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 76.225000 11.905000 76.545000 ;
      LAYER met4 ;
        RECT 11.585000 76.225000 11.905000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 76.630000 11.905000 76.950000 ;
      LAYER met4 ;
        RECT 11.585000 76.630000 11.905000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 77.035000 11.905000 77.355000 ;
      LAYER met4 ;
        RECT 11.585000 77.035000 11.905000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 77.440000 11.905000 77.760000 ;
      LAYER met4 ;
        RECT 11.585000 77.440000 11.905000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 77.845000 11.905000 78.165000 ;
      LAYER met4 ;
        RECT 11.585000 77.845000 11.905000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 78.250000 11.905000 78.570000 ;
      LAYER met4 ;
        RECT 11.585000 78.250000 11.905000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 78.655000 11.905000 78.975000 ;
      LAYER met4 ;
        RECT 11.585000 78.655000 11.905000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 79.060000 11.905000 79.380000 ;
      LAYER met4 ;
        RECT 11.585000 79.060000 11.905000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 79.465000 11.905000 79.785000 ;
      LAYER met4 ;
        RECT 11.585000 79.465000 11.905000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 79.870000 11.905000 80.190000 ;
      LAYER met4 ;
        RECT 11.585000 79.870000 11.905000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 80.275000 11.905000 80.595000 ;
      LAYER met4 ;
        RECT 11.585000 80.275000 11.905000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 80.680000 11.905000 81.000000 ;
      LAYER met4 ;
        RECT 11.585000 80.680000 11.905000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 81.085000 11.905000 81.405000 ;
      LAYER met4 ;
        RECT 11.585000 81.085000 11.905000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 81.490000 11.905000 81.810000 ;
      LAYER met4 ;
        RECT 11.585000 81.490000 11.905000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 81.895000 11.905000 82.215000 ;
      LAYER met4 ;
        RECT 11.585000 81.895000 11.905000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585000 82.300000 11.905000 82.620000 ;
      LAYER met4 ;
        RECT 11.585000 82.300000 11.905000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 82.795000 12.065000 83.115000 ;
      LAYER met4 ;
        RECT 11.745000 82.795000 12.065000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 83.205000 12.065000 83.525000 ;
      LAYER met4 ;
        RECT 11.745000 83.205000 12.065000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 83.615000 12.065000 83.935000 ;
      LAYER met4 ;
        RECT 11.745000 83.615000 12.065000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 84.025000 12.065000 84.345000 ;
      LAYER met4 ;
        RECT 11.745000 84.025000 12.065000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 84.435000 12.065000 84.755000 ;
      LAYER met4 ;
        RECT 11.745000 84.435000 12.065000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 84.845000 12.065000 85.165000 ;
      LAYER met4 ;
        RECT 11.745000 84.845000 12.065000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 85.255000 12.065000 85.575000 ;
      LAYER met4 ;
        RECT 11.745000 85.255000 12.065000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 85.665000 12.065000 85.985000 ;
      LAYER met4 ;
        RECT 11.745000 85.665000 12.065000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 86.075000 12.065000 86.395000 ;
      LAYER met4 ;
        RECT 11.745000 86.075000 12.065000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 86.485000 12.065000 86.805000 ;
      LAYER met4 ;
        RECT 11.745000 86.485000 12.065000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 86.895000 12.065000 87.215000 ;
      LAYER met4 ;
        RECT 11.745000 86.895000 12.065000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 87.305000 12.065000 87.625000 ;
      LAYER met4 ;
        RECT 11.745000 87.305000 12.065000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 87.715000 12.065000 88.035000 ;
      LAYER met4 ;
        RECT 11.745000 87.715000 12.065000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 88.125000 12.065000 88.445000 ;
      LAYER met4 ;
        RECT 11.745000 88.125000 12.065000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 88.535000 12.065000 88.855000 ;
      LAYER met4 ;
        RECT 11.745000 88.535000 12.065000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 88.945000 12.065000 89.265000 ;
      LAYER met4 ;
        RECT 11.745000 88.945000 12.065000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 89.355000 12.065000 89.675000 ;
      LAYER met4 ;
        RECT 11.745000 89.355000 12.065000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 89.765000 12.065000 90.085000 ;
      LAYER met4 ;
        RECT 11.745000 89.765000 12.065000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 90.175000 12.065000 90.495000 ;
      LAYER met4 ;
        RECT 11.745000 90.175000 12.065000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 90.585000 12.065000 90.905000 ;
      LAYER met4 ;
        RECT 11.745000 90.585000 12.065000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 90.995000 12.065000 91.315000 ;
      LAYER met4 ;
        RECT 11.745000 90.995000 12.065000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 91.405000 12.065000 91.725000 ;
      LAYER met4 ;
        RECT 11.745000 91.405000 12.065000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 91.815000 12.065000 92.135000 ;
      LAYER met4 ;
        RECT 11.745000 91.815000 12.065000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 92.225000 12.065000 92.545000 ;
      LAYER met4 ;
        RECT 11.745000 92.225000 12.065000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745000 92.635000 12.065000 92.955000 ;
      LAYER met4 ;
        RECT 11.745000 92.635000 12.065000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970000 17.800000 12.290000 18.120000 ;
      LAYER met4 ;
        RECT 11.970000 17.800000 12.290000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970000 18.230000 12.290000 18.550000 ;
      LAYER met4 ;
        RECT 11.970000 18.230000 12.290000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970000 18.660000 12.290000 18.980000 ;
      LAYER met4 ;
        RECT 11.970000 18.660000 12.290000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970000 19.090000 12.290000 19.410000 ;
      LAYER met4 ;
        RECT 11.970000 19.090000 12.290000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970000 19.520000 12.290000 19.840000 ;
      LAYER met4 ;
        RECT 11.970000 19.520000 12.290000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970000 19.950000 12.290000 20.270000 ;
      LAYER met4 ;
        RECT 11.970000 19.950000 12.290000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970000 20.380000 12.290000 20.700000 ;
      LAYER met4 ;
        RECT 11.970000 20.380000 12.290000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970000 20.810000 12.290000 21.130000 ;
      LAYER met4 ;
        RECT 11.970000 20.810000 12.290000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970000 21.240000 12.290000 21.560000 ;
      LAYER met4 ;
        RECT 11.970000 21.240000 12.290000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970000 21.670000 12.290000 21.990000 ;
      LAYER met4 ;
        RECT 11.970000 21.670000 12.290000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970000 22.100000 12.290000 22.420000 ;
      LAYER met4 ;
        RECT 11.970000 22.100000 12.290000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 68.065000 12.305000 68.385000 ;
      LAYER met4 ;
        RECT 11.985000 68.065000 12.305000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 68.475000 12.305000 68.795000 ;
      LAYER met4 ;
        RECT 11.985000 68.475000 12.305000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 68.885000 12.305000 69.205000 ;
      LAYER met4 ;
        RECT 11.985000 68.885000 12.305000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 69.295000 12.305000 69.615000 ;
      LAYER met4 ;
        RECT 11.985000 69.295000 12.305000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 69.705000 12.305000 70.025000 ;
      LAYER met4 ;
        RECT 11.985000 69.705000 12.305000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 70.115000 12.305000 70.435000 ;
      LAYER met4 ;
        RECT 11.985000 70.115000 12.305000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 70.525000 12.305000 70.845000 ;
      LAYER met4 ;
        RECT 11.985000 70.525000 12.305000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 70.935000 12.305000 71.255000 ;
      LAYER met4 ;
        RECT 11.985000 70.935000 12.305000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 71.345000 12.305000 71.665000 ;
      LAYER met4 ;
        RECT 11.985000 71.345000 12.305000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 71.755000 12.305000 72.075000 ;
      LAYER met4 ;
        RECT 11.985000 71.755000 12.305000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 72.165000 12.305000 72.485000 ;
      LAYER met4 ;
        RECT 11.985000 72.165000 12.305000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 72.575000 12.305000 72.895000 ;
      LAYER met4 ;
        RECT 11.985000 72.575000 12.305000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 72.985000 12.305000 73.305000 ;
      LAYER met4 ;
        RECT 11.985000 72.985000 12.305000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 73.390000 12.305000 73.710000 ;
      LAYER met4 ;
        RECT 11.985000 73.390000 12.305000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 73.795000 12.305000 74.115000 ;
      LAYER met4 ;
        RECT 11.985000 73.795000 12.305000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 74.200000 12.305000 74.520000 ;
      LAYER met4 ;
        RECT 11.985000 74.200000 12.305000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 74.605000 12.305000 74.925000 ;
      LAYER met4 ;
        RECT 11.985000 74.605000 12.305000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 75.010000 12.305000 75.330000 ;
      LAYER met4 ;
        RECT 11.985000 75.010000 12.305000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 75.415000 12.305000 75.735000 ;
      LAYER met4 ;
        RECT 11.985000 75.415000 12.305000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 75.820000 12.305000 76.140000 ;
      LAYER met4 ;
        RECT 11.985000 75.820000 12.305000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 76.225000 12.305000 76.545000 ;
      LAYER met4 ;
        RECT 11.985000 76.225000 12.305000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 76.630000 12.305000 76.950000 ;
      LAYER met4 ;
        RECT 11.985000 76.630000 12.305000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 77.035000 12.305000 77.355000 ;
      LAYER met4 ;
        RECT 11.985000 77.035000 12.305000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 77.440000 12.305000 77.760000 ;
      LAYER met4 ;
        RECT 11.985000 77.440000 12.305000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 77.845000 12.305000 78.165000 ;
      LAYER met4 ;
        RECT 11.985000 77.845000 12.305000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 78.250000 12.305000 78.570000 ;
      LAYER met4 ;
        RECT 11.985000 78.250000 12.305000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 78.655000 12.305000 78.975000 ;
      LAYER met4 ;
        RECT 11.985000 78.655000 12.305000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 79.060000 12.305000 79.380000 ;
      LAYER met4 ;
        RECT 11.985000 79.060000 12.305000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 79.465000 12.305000 79.785000 ;
      LAYER met4 ;
        RECT 11.985000 79.465000 12.305000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 79.870000 12.305000 80.190000 ;
      LAYER met4 ;
        RECT 11.985000 79.870000 12.305000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 80.275000 12.305000 80.595000 ;
      LAYER met4 ;
        RECT 11.985000 80.275000 12.305000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 80.680000 12.305000 81.000000 ;
      LAYER met4 ;
        RECT 11.985000 80.680000 12.305000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 81.085000 12.305000 81.405000 ;
      LAYER met4 ;
        RECT 11.985000 81.085000 12.305000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 81.490000 12.305000 81.810000 ;
      LAYER met4 ;
        RECT 11.985000 81.490000 12.305000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 81.895000 12.305000 82.215000 ;
      LAYER met4 ;
        RECT 11.985000 81.895000 12.305000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985000 82.300000 12.305000 82.620000 ;
      LAYER met4 ;
        RECT 11.985000 82.300000 12.305000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 82.795000 12.475000 83.115000 ;
      LAYER met4 ;
        RECT 12.155000 82.795000 12.475000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 83.205000 12.475000 83.525000 ;
      LAYER met4 ;
        RECT 12.155000 83.205000 12.475000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 83.615000 12.475000 83.935000 ;
      LAYER met4 ;
        RECT 12.155000 83.615000 12.475000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 84.025000 12.475000 84.345000 ;
      LAYER met4 ;
        RECT 12.155000 84.025000 12.475000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 84.435000 12.475000 84.755000 ;
      LAYER met4 ;
        RECT 12.155000 84.435000 12.475000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 84.845000 12.475000 85.165000 ;
      LAYER met4 ;
        RECT 12.155000 84.845000 12.475000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 85.255000 12.475000 85.575000 ;
      LAYER met4 ;
        RECT 12.155000 85.255000 12.475000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 85.665000 12.475000 85.985000 ;
      LAYER met4 ;
        RECT 12.155000 85.665000 12.475000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 86.075000 12.475000 86.395000 ;
      LAYER met4 ;
        RECT 12.155000 86.075000 12.475000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 86.485000 12.475000 86.805000 ;
      LAYER met4 ;
        RECT 12.155000 86.485000 12.475000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 86.895000 12.475000 87.215000 ;
      LAYER met4 ;
        RECT 12.155000 86.895000 12.475000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 87.305000 12.475000 87.625000 ;
      LAYER met4 ;
        RECT 12.155000 87.305000 12.475000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 87.715000 12.475000 88.035000 ;
      LAYER met4 ;
        RECT 12.155000 87.715000 12.475000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 88.125000 12.475000 88.445000 ;
      LAYER met4 ;
        RECT 12.155000 88.125000 12.475000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 88.535000 12.475000 88.855000 ;
      LAYER met4 ;
        RECT 12.155000 88.535000 12.475000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 88.945000 12.475000 89.265000 ;
      LAYER met4 ;
        RECT 12.155000 88.945000 12.475000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 89.355000 12.475000 89.675000 ;
      LAYER met4 ;
        RECT 12.155000 89.355000 12.475000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 89.765000 12.475000 90.085000 ;
      LAYER met4 ;
        RECT 12.155000 89.765000 12.475000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 90.175000 12.475000 90.495000 ;
      LAYER met4 ;
        RECT 12.155000 90.175000 12.475000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 90.585000 12.475000 90.905000 ;
      LAYER met4 ;
        RECT 12.155000 90.585000 12.475000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 90.995000 12.475000 91.315000 ;
      LAYER met4 ;
        RECT 12.155000 90.995000 12.475000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 91.405000 12.475000 91.725000 ;
      LAYER met4 ;
        RECT 12.155000 91.405000 12.475000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 91.815000 12.475000 92.135000 ;
      LAYER met4 ;
        RECT 12.155000 91.815000 12.475000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 92.225000 12.475000 92.545000 ;
      LAYER met4 ;
        RECT 12.155000 92.225000 12.475000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155000 92.635000 12.475000 92.955000 ;
      LAYER met4 ;
        RECT 12.155000 92.635000 12.475000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375000 17.800000 12.695000 18.120000 ;
      LAYER met4 ;
        RECT 12.375000 17.800000 12.695000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375000 18.230000 12.695000 18.550000 ;
      LAYER met4 ;
        RECT 12.375000 18.230000 12.695000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375000 18.660000 12.695000 18.980000 ;
      LAYER met4 ;
        RECT 12.375000 18.660000 12.695000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375000 19.090000 12.695000 19.410000 ;
      LAYER met4 ;
        RECT 12.375000 19.090000 12.695000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375000 19.520000 12.695000 19.840000 ;
      LAYER met4 ;
        RECT 12.375000 19.520000 12.695000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375000 19.950000 12.695000 20.270000 ;
      LAYER met4 ;
        RECT 12.375000 19.950000 12.695000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375000 20.380000 12.695000 20.700000 ;
      LAYER met4 ;
        RECT 12.375000 20.380000 12.695000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375000 20.810000 12.695000 21.130000 ;
      LAYER met4 ;
        RECT 12.375000 20.810000 12.695000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375000 21.240000 12.695000 21.560000 ;
      LAYER met4 ;
        RECT 12.375000 21.240000 12.695000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375000 21.670000 12.695000 21.990000 ;
      LAYER met4 ;
        RECT 12.375000 21.670000 12.695000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375000 22.100000 12.695000 22.420000 ;
      LAYER met4 ;
        RECT 12.375000 22.100000 12.695000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 68.065000 12.705000 68.385000 ;
      LAYER met4 ;
        RECT 12.385000 68.065000 12.705000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 68.475000 12.705000 68.795000 ;
      LAYER met4 ;
        RECT 12.385000 68.475000 12.705000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 68.885000 12.705000 69.205000 ;
      LAYER met4 ;
        RECT 12.385000 68.885000 12.705000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 69.295000 12.705000 69.615000 ;
      LAYER met4 ;
        RECT 12.385000 69.295000 12.705000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 69.705000 12.705000 70.025000 ;
      LAYER met4 ;
        RECT 12.385000 69.705000 12.705000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 70.115000 12.705000 70.435000 ;
      LAYER met4 ;
        RECT 12.385000 70.115000 12.705000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 70.525000 12.705000 70.845000 ;
      LAYER met4 ;
        RECT 12.385000 70.525000 12.705000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 70.935000 12.705000 71.255000 ;
      LAYER met4 ;
        RECT 12.385000 70.935000 12.705000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 71.345000 12.705000 71.665000 ;
      LAYER met4 ;
        RECT 12.385000 71.345000 12.705000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 71.755000 12.705000 72.075000 ;
      LAYER met4 ;
        RECT 12.385000 71.755000 12.705000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 72.165000 12.705000 72.485000 ;
      LAYER met4 ;
        RECT 12.385000 72.165000 12.705000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 72.575000 12.705000 72.895000 ;
      LAYER met4 ;
        RECT 12.385000 72.575000 12.705000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 72.985000 12.705000 73.305000 ;
      LAYER met4 ;
        RECT 12.385000 72.985000 12.705000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 73.390000 12.705000 73.710000 ;
      LAYER met4 ;
        RECT 12.385000 73.390000 12.705000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 73.795000 12.705000 74.115000 ;
      LAYER met4 ;
        RECT 12.385000 73.795000 12.705000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 74.200000 12.705000 74.520000 ;
      LAYER met4 ;
        RECT 12.385000 74.200000 12.705000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 74.605000 12.705000 74.925000 ;
      LAYER met4 ;
        RECT 12.385000 74.605000 12.705000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 75.010000 12.705000 75.330000 ;
      LAYER met4 ;
        RECT 12.385000 75.010000 12.705000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 75.415000 12.705000 75.735000 ;
      LAYER met4 ;
        RECT 12.385000 75.415000 12.705000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 75.820000 12.705000 76.140000 ;
      LAYER met4 ;
        RECT 12.385000 75.820000 12.705000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 76.225000 12.705000 76.545000 ;
      LAYER met4 ;
        RECT 12.385000 76.225000 12.705000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 76.630000 12.705000 76.950000 ;
      LAYER met4 ;
        RECT 12.385000 76.630000 12.705000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 77.035000 12.705000 77.355000 ;
      LAYER met4 ;
        RECT 12.385000 77.035000 12.705000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 77.440000 12.705000 77.760000 ;
      LAYER met4 ;
        RECT 12.385000 77.440000 12.705000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 77.845000 12.705000 78.165000 ;
      LAYER met4 ;
        RECT 12.385000 77.845000 12.705000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 78.250000 12.705000 78.570000 ;
      LAYER met4 ;
        RECT 12.385000 78.250000 12.705000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 78.655000 12.705000 78.975000 ;
      LAYER met4 ;
        RECT 12.385000 78.655000 12.705000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 79.060000 12.705000 79.380000 ;
      LAYER met4 ;
        RECT 12.385000 79.060000 12.705000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 79.465000 12.705000 79.785000 ;
      LAYER met4 ;
        RECT 12.385000 79.465000 12.705000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 79.870000 12.705000 80.190000 ;
      LAYER met4 ;
        RECT 12.385000 79.870000 12.705000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 80.275000 12.705000 80.595000 ;
      LAYER met4 ;
        RECT 12.385000 80.275000 12.705000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 80.680000 12.705000 81.000000 ;
      LAYER met4 ;
        RECT 12.385000 80.680000 12.705000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 81.085000 12.705000 81.405000 ;
      LAYER met4 ;
        RECT 12.385000 81.085000 12.705000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 81.490000 12.705000 81.810000 ;
      LAYER met4 ;
        RECT 12.385000 81.490000 12.705000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 81.895000 12.705000 82.215000 ;
      LAYER met4 ;
        RECT 12.385000 81.895000 12.705000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385000 82.300000 12.705000 82.620000 ;
      LAYER met4 ;
        RECT 12.385000 82.300000 12.705000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 82.795000 12.885000 83.115000 ;
      LAYER met4 ;
        RECT 12.565000 82.795000 12.885000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 83.205000 12.885000 83.525000 ;
      LAYER met4 ;
        RECT 12.565000 83.205000 12.885000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 83.615000 12.885000 83.935000 ;
      LAYER met4 ;
        RECT 12.565000 83.615000 12.885000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 84.025000 12.885000 84.345000 ;
      LAYER met4 ;
        RECT 12.565000 84.025000 12.885000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 84.435000 12.885000 84.755000 ;
      LAYER met4 ;
        RECT 12.565000 84.435000 12.885000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 84.845000 12.885000 85.165000 ;
      LAYER met4 ;
        RECT 12.565000 84.845000 12.885000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 85.255000 12.885000 85.575000 ;
      LAYER met4 ;
        RECT 12.565000 85.255000 12.885000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 85.665000 12.885000 85.985000 ;
      LAYER met4 ;
        RECT 12.565000 85.665000 12.885000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 86.075000 12.885000 86.395000 ;
      LAYER met4 ;
        RECT 12.565000 86.075000 12.885000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 86.485000 12.885000 86.805000 ;
      LAYER met4 ;
        RECT 12.565000 86.485000 12.885000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 86.895000 12.885000 87.215000 ;
      LAYER met4 ;
        RECT 12.565000 86.895000 12.885000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 87.305000 12.885000 87.625000 ;
      LAYER met4 ;
        RECT 12.565000 87.305000 12.885000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 87.715000 12.885000 88.035000 ;
      LAYER met4 ;
        RECT 12.565000 87.715000 12.885000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 88.125000 12.885000 88.445000 ;
      LAYER met4 ;
        RECT 12.565000 88.125000 12.885000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 88.535000 12.885000 88.855000 ;
      LAYER met4 ;
        RECT 12.565000 88.535000 12.885000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 88.945000 12.885000 89.265000 ;
      LAYER met4 ;
        RECT 12.565000 88.945000 12.885000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 89.355000 12.885000 89.675000 ;
      LAYER met4 ;
        RECT 12.565000 89.355000 12.885000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 89.765000 12.885000 90.085000 ;
      LAYER met4 ;
        RECT 12.565000 89.765000 12.885000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 90.175000 12.885000 90.495000 ;
      LAYER met4 ;
        RECT 12.565000 90.175000 12.885000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 90.585000 12.885000 90.905000 ;
      LAYER met4 ;
        RECT 12.565000 90.585000 12.885000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 90.995000 12.885000 91.315000 ;
      LAYER met4 ;
        RECT 12.565000 90.995000 12.885000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 91.405000 12.885000 91.725000 ;
      LAYER met4 ;
        RECT 12.565000 91.405000 12.885000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 91.815000 12.885000 92.135000 ;
      LAYER met4 ;
        RECT 12.565000 91.815000 12.885000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 92.225000 12.885000 92.545000 ;
      LAYER met4 ;
        RECT 12.565000 92.225000 12.885000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565000 92.635000 12.885000 92.955000 ;
      LAYER met4 ;
        RECT 12.565000 92.635000 12.885000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 17.800000 13.100000 18.120000 ;
      LAYER met4 ;
        RECT 12.780000 17.800000 13.100000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 18.230000 13.100000 18.550000 ;
      LAYER met4 ;
        RECT 12.780000 18.230000 13.100000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 18.660000 13.100000 18.980000 ;
      LAYER met4 ;
        RECT 12.780000 18.660000 13.100000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 19.090000 13.100000 19.410000 ;
      LAYER met4 ;
        RECT 12.780000 19.090000 13.100000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 19.520000 13.100000 19.840000 ;
      LAYER met4 ;
        RECT 12.780000 19.520000 13.100000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 19.950000 13.100000 20.270000 ;
      LAYER met4 ;
        RECT 12.780000 19.950000 13.100000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 20.380000 13.100000 20.700000 ;
      LAYER met4 ;
        RECT 12.780000 20.380000 13.100000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 20.810000 13.100000 21.130000 ;
      LAYER met4 ;
        RECT 12.780000 20.810000 13.100000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 21.240000 13.100000 21.560000 ;
      LAYER met4 ;
        RECT 12.780000 21.240000 13.100000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 21.670000 13.100000 21.990000 ;
      LAYER met4 ;
        RECT 12.780000 21.670000 13.100000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 22.100000 13.100000 22.420000 ;
      LAYER met4 ;
        RECT 12.780000 22.100000 13.100000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 68.065000 13.105000 68.385000 ;
      LAYER met4 ;
        RECT 12.785000 68.065000 13.105000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 68.475000 13.105000 68.795000 ;
      LAYER met4 ;
        RECT 12.785000 68.475000 13.105000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 68.885000 13.105000 69.205000 ;
      LAYER met4 ;
        RECT 12.785000 68.885000 13.105000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 69.295000 13.105000 69.615000 ;
      LAYER met4 ;
        RECT 12.785000 69.295000 13.105000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 69.705000 13.105000 70.025000 ;
      LAYER met4 ;
        RECT 12.785000 69.705000 13.105000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 70.115000 13.105000 70.435000 ;
      LAYER met4 ;
        RECT 12.785000 70.115000 13.105000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 70.525000 13.105000 70.845000 ;
      LAYER met4 ;
        RECT 12.785000 70.525000 13.105000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 70.935000 13.105000 71.255000 ;
      LAYER met4 ;
        RECT 12.785000 70.935000 13.105000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 71.345000 13.105000 71.665000 ;
      LAYER met4 ;
        RECT 12.785000 71.345000 13.105000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 71.755000 13.105000 72.075000 ;
      LAYER met4 ;
        RECT 12.785000 71.755000 13.105000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 72.165000 13.105000 72.485000 ;
      LAYER met4 ;
        RECT 12.785000 72.165000 13.105000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 72.575000 13.105000 72.895000 ;
      LAYER met4 ;
        RECT 12.785000 72.575000 13.105000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 72.985000 13.105000 73.305000 ;
      LAYER met4 ;
        RECT 12.785000 72.985000 13.105000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 73.390000 13.105000 73.710000 ;
      LAYER met4 ;
        RECT 12.785000 73.390000 13.105000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 73.795000 13.105000 74.115000 ;
      LAYER met4 ;
        RECT 12.785000 73.795000 13.105000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 74.200000 13.105000 74.520000 ;
      LAYER met4 ;
        RECT 12.785000 74.200000 13.105000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 74.605000 13.105000 74.925000 ;
      LAYER met4 ;
        RECT 12.785000 74.605000 13.105000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 75.010000 13.105000 75.330000 ;
      LAYER met4 ;
        RECT 12.785000 75.010000 13.105000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 75.415000 13.105000 75.735000 ;
      LAYER met4 ;
        RECT 12.785000 75.415000 13.105000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 75.820000 13.105000 76.140000 ;
      LAYER met4 ;
        RECT 12.785000 75.820000 13.105000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 76.225000 13.105000 76.545000 ;
      LAYER met4 ;
        RECT 12.785000 76.225000 13.105000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 76.630000 13.105000 76.950000 ;
      LAYER met4 ;
        RECT 12.785000 76.630000 13.105000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 77.035000 13.105000 77.355000 ;
      LAYER met4 ;
        RECT 12.785000 77.035000 13.105000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 77.440000 13.105000 77.760000 ;
      LAYER met4 ;
        RECT 12.785000 77.440000 13.105000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 77.845000 13.105000 78.165000 ;
      LAYER met4 ;
        RECT 12.785000 77.845000 13.105000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 78.250000 13.105000 78.570000 ;
      LAYER met4 ;
        RECT 12.785000 78.250000 13.105000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 78.655000 13.105000 78.975000 ;
      LAYER met4 ;
        RECT 12.785000 78.655000 13.105000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 79.060000 13.105000 79.380000 ;
      LAYER met4 ;
        RECT 12.785000 79.060000 13.105000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 79.465000 13.105000 79.785000 ;
      LAYER met4 ;
        RECT 12.785000 79.465000 13.105000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 79.870000 13.105000 80.190000 ;
      LAYER met4 ;
        RECT 12.785000 79.870000 13.105000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 80.275000 13.105000 80.595000 ;
      LAYER met4 ;
        RECT 12.785000 80.275000 13.105000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 80.680000 13.105000 81.000000 ;
      LAYER met4 ;
        RECT 12.785000 80.680000 13.105000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 81.085000 13.105000 81.405000 ;
      LAYER met4 ;
        RECT 12.785000 81.085000 13.105000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 81.490000 13.105000 81.810000 ;
      LAYER met4 ;
        RECT 12.785000 81.490000 13.105000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 81.895000 13.105000 82.215000 ;
      LAYER met4 ;
        RECT 12.785000 81.895000 13.105000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785000 82.300000 13.105000 82.620000 ;
      LAYER met4 ;
        RECT 12.785000 82.300000 13.105000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 82.795000 13.290000 83.115000 ;
      LAYER met4 ;
        RECT 12.970000 82.795000 13.290000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 83.205000 13.290000 83.525000 ;
      LAYER met4 ;
        RECT 12.970000 83.205000 13.290000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 83.615000 13.290000 83.935000 ;
      LAYER met4 ;
        RECT 12.970000 83.615000 13.290000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 84.025000 13.290000 84.345000 ;
      LAYER met4 ;
        RECT 12.970000 84.025000 13.290000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 84.435000 13.290000 84.755000 ;
      LAYER met4 ;
        RECT 12.970000 84.435000 13.290000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 84.845000 13.290000 85.165000 ;
      LAYER met4 ;
        RECT 12.970000 84.845000 13.290000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 85.255000 13.290000 85.575000 ;
      LAYER met4 ;
        RECT 12.970000 85.255000 13.290000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 85.665000 13.290000 85.985000 ;
      LAYER met4 ;
        RECT 12.970000 85.665000 13.290000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 86.075000 13.290000 86.395000 ;
      LAYER met4 ;
        RECT 12.970000 86.075000 13.290000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 86.485000 13.290000 86.805000 ;
      LAYER met4 ;
        RECT 12.970000 86.485000 13.290000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 86.895000 13.290000 87.215000 ;
      LAYER met4 ;
        RECT 12.970000 86.895000 13.290000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 87.305000 13.290000 87.625000 ;
      LAYER met4 ;
        RECT 12.970000 87.305000 13.290000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 87.715000 13.290000 88.035000 ;
      LAYER met4 ;
        RECT 12.970000 87.715000 13.290000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 88.125000 13.290000 88.445000 ;
      LAYER met4 ;
        RECT 12.970000 88.125000 13.290000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 88.535000 13.290000 88.855000 ;
      LAYER met4 ;
        RECT 12.970000 88.535000 13.290000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 88.945000 13.290000 89.265000 ;
      LAYER met4 ;
        RECT 12.970000 88.945000 13.290000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 89.355000 13.290000 89.675000 ;
      LAYER met4 ;
        RECT 12.970000 89.355000 13.290000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 89.765000 13.290000 90.085000 ;
      LAYER met4 ;
        RECT 12.970000 89.765000 13.290000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 90.175000 13.290000 90.495000 ;
      LAYER met4 ;
        RECT 12.970000 90.175000 13.290000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 90.585000 13.290000 90.905000 ;
      LAYER met4 ;
        RECT 12.970000 90.585000 13.290000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 90.995000 13.290000 91.315000 ;
      LAYER met4 ;
        RECT 12.970000 90.995000 13.290000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 91.405000 13.290000 91.725000 ;
      LAYER met4 ;
        RECT 12.970000 91.405000 13.290000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 91.815000 13.290000 92.135000 ;
      LAYER met4 ;
        RECT 12.970000 91.815000 13.290000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 92.225000 13.290000 92.545000 ;
      LAYER met4 ;
        RECT 12.970000 92.225000 13.290000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970000 92.635000 13.290000 92.955000 ;
      LAYER met4 ;
        RECT 12.970000 92.635000 13.290000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 17.800000 13.505000 18.120000 ;
      LAYER met4 ;
        RECT 13.185000 17.800000 13.505000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 18.230000 13.505000 18.550000 ;
      LAYER met4 ;
        RECT 13.185000 18.230000 13.505000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 18.660000 13.505000 18.980000 ;
      LAYER met4 ;
        RECT 13.185000 18.660000 13.505000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 19.090000 13.505000 19.410000 ;
      LAYER met4 ;
        RECT 13.185000 19.090000 13.505000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 19.520000 13.505000 19.840000 ;
      LAYER met4 ;
        RECT 13.185000 19.520000 13.505000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 19.950000 13.505000 20.270000 ;
      LAYER met4 ;
        RECT 13.185000 19.950000 13.505000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 20.380000 13.505000 20.700000 ;
      LAYER met4 ;
        RECT 13.185000 20.380000 13.505000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 20.810000 13.505000 21.130000 ;
      LAYER met4 ;
        RECT 13.185000 20.810000 13.505000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 21.240000 13.505000 21.560000 ;
      LAYER met4 ;
        RECT 13.185000 21.240000 13.505000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 21.670000 13.505000 21.990000 ;
      LAYER met4 ;
        RECT 13.185000 21.670000 13.505000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 22.100000 13.505000 22.420000 ;
      LAYER met4 ;
        RECT 13.185000 22.100000 13.505000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 68.065000 13.505000 68.385000 ;
      LAYER met4 ;
        RECT 13.185000 68.065000 13.505000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 68.475000 13.505000 68.795000 ;
      LAYER met4 ;
        RECT 13.185000 68.475000 13.505000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 68.885000 13.505000 69.205000 ;
      LAYER met4 ;
        RECT 13.185000 68.885000 13.505000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 69.295000 13.505000 69.615000 ;
      LAYER met4 ;
        RECT 13.185000 69.295000 13.505000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 69.705000 13.505000 70.025000 ;
      LAYER met4 ;
        RECT 13.185000 69.705000 13.505000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 70.115000 13.505000 70.435000 ;
      LAYER met4 ;
        RECT 13.185000 70.115000 13.505000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 70.525000 13.505000 70.845000 ;
      LAYER met4 ;
        RECT 13.185000 70.525000 13.505000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 70.935000 13.505000 71.255000 ;
      LAYER met4 ;
        RECT 13.185000 70.935000 13.505000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 71.345000 13.505000 71.665000 ;
      LAYER met4 ;
        RECT 13.185000 71.345000 13.505000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 71.755000 13.505000 72.075000 ;
      LAYER met4 ;
        RECT 13.185000 71.755000 13.505000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 72.165000 13.505000 72.485000 ;
      LAYER met4 ;
        RECT 13.185000 72.165000 13.505000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 72.575000 13.505000 72.895000 ;
      LAYER met4 ;
        RECT 13.185000 72.575000 13.505000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 72.985000 13.505000 73.305000 ;
      LAYER met4 ;
        RECT 13.185000 72.985000 13.505000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 73.390000 13.505000 73.710000 ;
      LAYER met4 ;
        RECT 13.185000 73.390000 13.505000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 73.795000 13.505000 74.115000 ;
      LAYER met4 ;
        RECT 13.185000 73.795000 13.505000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 74.200000 13.505000 74.520000 ;
      LAYER met4 ;
        RECT 13.185000 74.200000 13.505000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 74.605000 13.505000 74.925000 ;
      LAYER met4 ;
        RECT 13.185000 74.605000 13.505000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 75.010000 13.505000 75.330000 ;
      LAYER met4 ;
        RECT 13.185000 75.010000 13.505000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 75.415000 13.505000 75.735000 ;
      LAYER met4 ;
        RECT 13.185000 75.415000 13.505000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 75.820000 13.505000 76.140000 ;
      LAYER met4 ;
        RECT 13.185000 75.820000 13.505000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 76.225000 13.505000 76.545000 ;
      LAYER met4 ;
        RECT 13.185000 76.225000 13.505000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 76.630000 13.505000 76.950000 ;
      LAYER met4 ;
        RECT 13.185000 76.630000 13.505000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 77.035000 13.505000 77.355000 ;
      LAYER met4 ;
        RECT 13.185000 77.035000 13.505000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 77.440000 13.505000 77.760000 ;
      LAYER met4 ;
        RECT 13.185000 77.440000 13.505000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 77.845000 13.505000 78.165000 ;
      LAYER met4 ;
        RECT 13.185000 77.845000 13.505000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 78.250000 13.505000 78.570000 ;
      LAYER met4 ;
        RECT 13.185000 78.250000 13.505000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 78.655000 13.505000 78.975000 ;
      LAYER met4 ;
        RECT 13.185000 78.655000 13.505000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 79.060000 13.505000 79.380000 ;
      LAYER met4 ;
        RECT 13.185000 79.060000 13.505000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 79.465000 13.505000 79.785000 ;
      LAYER met4 ;
        RECT 13.185000 79.465000 13.505000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 79.870000 13.505000 80.190000 ;
      LAYER met4 ;
        RECT 13.185000 79.870000 13.505000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 80.275000 13.505000 80.595000 ;
      LAYER met4 ;
        RECT 13.185000 80.275000 13.505000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 80.680000 13.505000 81.000000 ;
      LAYER met4 ;
        RECT 13.185000 80.680000 13.505000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 81.085000 13.505000 81.405000 ;
      LAYER met4 ;
        RECT 13.185000 81.085000 13.505000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 81.490000 13.505000 81.810000 ;
      LAYER met4 ;
        RECT 13.185000 81.490000 13.505000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 81.895000 13.505000 82.215000 ;
      LAYER met4 ;
        RECT 13.185000 81.895000 13.505000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 82.300000 13.505000 82.620000 ;
      LAYER met4 ;
        RECT 13.185000 82.300000 13.505000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 82.795000 13.695000 83.115000 ;
      LAYER met4 ;
        RECT 13.375000 82.795000 13.695000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 83.205000 13.695000 83.525000 ;
      LAYER met4 ;
        RECT 13.375000 83.205000 13.695000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 83.615000 13.695000 83.935000 ;
      LAYER met4 ;
        RECT 13.375000 83.615000 13.695000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 84.025000 13.695000 84.345000 ;
      LAYER met4 ;
        RECT 13.375000 84.025000 13.695000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 84.435000 13.695000 84.755000 ;
      LAYER met4 ;
        RECT 13.375000 84.435000 13.695000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 84.845000 13.695000 85.165000 ;
      LAYER met4 ;
        RECT 13.375000 84.845000 13.695000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 85.255000 13.695000 85.575000 ;
      LAYER met4 ;
        RECT 13.375000 85.255000 13.695000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 85.665000 13.695000 85.985000 ;
      LAYER met4 ;
        RECT 13.375000 85.665000 13.695000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 86.075000 13.695000 86.395000 ;
      LAYER met4 ;
        RECT 13.375000 86.075000 13.695000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 86.485000 13.695000 86.805000 ;
      LAYER met4 ;
        RECT 13.375000 86.485000 13.695000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 86.895000 13.695000 87.215000 ;
      LAYER met4 ;
        RECT 13.375000 86.895000 13.695000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 87.305000 13.695000 87.625000 ;
      LAYER met4 ;
        RECT 13.375000 87.305000 13.695000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 87.715000 13.695000 88.035000 ;
      LAYER met4 ;
        RECT 13.375000 87.715000 13.695000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 88.125000 13.695000 88.445000 ;
      LAYER met4 ;
        RECT 13.375000 88.125000 13.695000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 88.535000 13.695000 88.855000 ;
      LAYER met4 ;
        RECT 13.375000 88.535000 13.695000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 88.945000 13.695000 89.265000 ;
      LAYER met4 ;
        RECT 13.375000 88.945000 13.695000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 89.355000 13.695000 89.675000 ;
      LAYER met4 ;
        RECT 13.375000 89.355000 13.695000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 89.765000 13.695000 90.085000 ;
      LAYER met4 ;
        RECT 13.375000 89.765000 13.695000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 90.175000 13.695000 90.495000 ;
      LAYER met4 ;
        RECT 13.375000 90.175000 13.695000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 90.585000 13.695000 90.905000 ;
      LAYER met4 ;
        RECT 13.375000 90.585000 13.695000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 90.995000 13.695000 91.315000 ;
      LAYER met4 ;
        RECT 13.375000 90.995000 13.695000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 91.405000 13.695000 91.725000 ;
      LAYER met4 ;
        RECT 13.375000 91.405000 13.695000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 91.815000 13.695000 92.135000 ;
      LAYER met4 ;
        RECT 13.375000 91.815000 13.695000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 92.225000 13.695000 92.545000 ;
      LAYER met4 ;
        RECT 13.375000 92.225000 13.695000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375000 92.635000 13.695000 92.955000 ;
      LAYER met4 ;
        RECT 13.375000 92.635000 13.695000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 68.065000 13.905000 68.385000 ;
      LAYER met4 ;
        RECT 13.585000 68.065000 13.905000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 68.475000 13.905000 68.795000 ;
      LAYER met4 ;
        RECT 13.585000 68.475000 13.905000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 68.885000 13.905000 69.205000 ;
      LAYER met4 ;
        RECT 13.585000 68.885000 13.905000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 69.295000 13.905000 69.615000 ;
      LAYER met4 ;
        RECT 13.585000 69.295000 13.905000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 69.705000 13.905000 70.025000 ;
      LAYER met4 ;
        RECT 13.585000 69.705000 13.905000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 70.115000 13.905000 70.435000 ;
      LAYER met4 ;
        RECT 13.585000 70.115000 13.905000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 70.525000 13.905000 70.845000 ;
      LAYER met4 ;
        RECT 13.585000 70.525000 13.905000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 70.935000 13.905000 71.255000 ;
      LAYER met4 ;
        RECT 13.585000 70.935000 13.905000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 71.345000 13.905000 71.665000 ;
      LAYER met4 ;
        RECT 13.585000 71.345000 13.905000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 71.755000 13.905000 72.075000 ;
      LAYER met4 ;
        RECT 13.585000 71.755000 13.905000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 72.165000 13.905000 72.485000 ;
      LAYER met4 ;
        RECT 13.585000 72.165000 13.905000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 72.575000 13.905000 72.895000 ;
      LAYER met4 ;
        RECT 13.585000 72.575000 13.905000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 72.985000 13.905000 73.305000 ;
      LAYER met4 ;
        RECT 13.585000 72.985000 13.905000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 73.390000 13.905000 73.710000 ;
      LAYER met4 ;
        RECT 13.585000 73.390000 13.905000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 73.795000 13.905000 74.115000 ;
      LAYER met4 ;
        RECT 13.585000 73.795000 13.905000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 74.200000 13.905000 74.520000 ;
      LAYER met4 ;
        RECT 13.585000 74.200000 13.905000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 74.605000 13.905000 74.925000 ;
      LAYER met4 ;
        RECT 13.585000 74.605000 13.905000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 75.010000 13.905000 75.330000 ;
      LAYER met4 ;
        RECT 13.585000 75.010000 13.905000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 75.415000 13.905000 75.735000 ;
      LAYER met4 ;
        RECT 13.585000 75.415000 13.905000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 75.820000 13.905000 76.140000 ;
      LAYER met4 ;
        RECT 13.585000 75.820000 13.905000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 76.225000 13.905000 76.545000 ;
      LAYER met4 ;
        RECT 13.585000 76.225000 13.905000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 76.630000 13.905000 76.950000 ;
      LAYER met4 ;
        RECT 13.585000 76.630000 13.905000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 77.035000 13.905000 77.355000 ;
      LAYER met4 ;
        RECT 13.585000 77.035000 13.905000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 77.440000 13.905000 77.760000 ;
      LAYER met4 ;
        RECT 13.585000 77.440000 13.905000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 77.845000 13.905000 78.165000 ;
      LAYER met4 ;
        RECT 13.585000 77.845000 13.905000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 78.250000 13.905000 78.570000 ;
      LAYER met4 ;
        RECT 13.585000 78.250000 13.905000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 78.655000 13.905000 78.975000 ;
      LAYER met4 ;
        RECT 13.585000 78.655000 13.905000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 79.060000 13.905000 79.380000 ;
      LAYER met4 ;
        RECT 13.585000 79.060000 13.905000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 79.465000 13.905000 79.785000 ;
      LAYER met4 ;
        RECT 13.585000 79.465000 13.905000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 79.870000 13.905000 80.190000 ;
      LAYER met4 ;
        RECT 13.585000 79.870000 13.905000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 80.275000 13.905000 80.595000 ;
      LAYER met4 ;
        RECT 13.585000 80.275000 13.905000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 80.680000 13.905000 81.000000 ;
      LAYER met4 ;
        RECT 13.585000 80.680000 13.905000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 81.085000 13.905000 81.405000 ;
      LAYER met4 ;
        RECT 13.585000 81.085000 13.905000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 81.490000 13.905000 81.810000 ;
      LAYER met4 ;
        RECT 13.585000 81.490000 13.905000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 81.895000 13.905000 82.215000 ;
      LAYER met4 ;
        RECT 13.585000 81.895000 13.905000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585000 82.300000 13.905000 82.620000 ;
      LAYER met4 ;
        RECT 13.585000 82.300000 13.905000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590000 17.800000 13.910000 18.120000 ;
      LAYER met4 ;
        RECT 13.590000 17.800000 13.910000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590000 18.230000 13.910000 18.550000 ;
      LAYER met4 ;
        RECT 13.590000 18.230000 13.910000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590000 18.660000 13.910000 18.980000 ;
      LAYER met4 ;
        RECT 13.590000 18.660000 13.910000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590000 19.090000 13.910000 19.410000 ;
      LAYER met4 ;
        RECT 13.590000 19.090000 13.910000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590000 19.520000 13.910000 19.840000 ;
      LAYER met4 ;
        RECT 13.590000 19.520000 13.910000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590000 19.950000 13.910000 20.270000 ;
      LAYER met4 ;
        RECT 13.590000 19.950000 13.910000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590000 20.380000 13.910000 20.700000 ;
      LAYER met4 ;
        RECT 13.590000 20.380000 13.910000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590000 20.810000 13.910000 21.130000 ;
      LAYER met4 ;
        RECT 13.590000 20.810000 13.910000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590000 21.240000 13.910000 21.560000 ;
      LAYER met4 ;
        RECT 13.590000 21.240000 13.910000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590000 21.670000 13.910000 21.990000 ;
      LAYER met4 ;
        RECT 13.590000 21.670000 13.910000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590000 22.100000 13.910000 22.420000 ;
      LAYER met4 ;
        RECT 13.590000 22.100000 13.910000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 82.795000 14.100000 83.115000 ;
      LAYER met4 ;
        RECT 13.780000 82.795000 14.100000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 83.205000 14.100000 83.525000 ;
      LAYER met4 ;
        RECT 13.780000 83.205000 14.100000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 83.615000 14.100000 83.935000 ;
      LAYER met4 ;
        RECT 13.780000 83.615000 14.100000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 84.025000 14.100000 84.345000 ;
      LAYER met4 ;
        RECT 13.780000 84.025000 14.100000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 84.435000 14.100000 84.755000 ;
      LAYER met4 ;
        RECT 13.780000 84.435000 14.100000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 84.845000 14.100000 85.165000 ;
      LAYER met4 ;
        RECT 13.780000 84.845000 14.100000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 85.255000 14.100000 85.575000 ;
      LAYER met4 ;
        RECT 13.780000 85.255000 14.100000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 85.665000 14.100000 85.985000 ;
      LAYER met4 ;
        RECT 13.780000 85.665000 14.100000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 86.075000 14.100000 86.395000 ;
      LAYER met4 ;
        RECT 13.780000 86.075000 14.100000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 86.485000 14.100000 86.805000 ;
      LAYER met4 ;
        RECT 13.780000 86.485000 14.100000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 86.895000 14.100000 87.215000 ;
      LAYER met4 ;
        RECT 13.780000 86.895000 14.100000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 87.305000 14.100000 87.625000 ;
      LAYER met4 ;
        RECT 13.780000 87.305000 14.100000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 87.715000 14.100000 88.035000 ;
      LAYER met4 ;
        RECT 13.780000 87.715000 14.100000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 88.125000 14.100000 88.445000 ;
      LAYER met4 ;
        RECT 13.780000 88.125000 14.100000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 88.535000 14.100000 88.855000 ;
      LAYER met4 ;
        RECT 13.780000 88.535000 14.100000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 88.945000 14.100000 89.265000 ;
      LAYER met4 ;
        RECT 13.780000 88.945000 14.100000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 89.355000 14.100000 89.675000 ;
      LAYER met4 ;
        RECT 13.780000 89.355000 14.100000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 89.765000 14.100000 90.085000 ;
      LAYER met4 ;
        RECT 13.780000 89.765000 14.100000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 90.175000 14.100000 90.495000 ;
      LAYER met4 ;
        RECT 13.780000 90.175000 14.100000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 90.585000 14.100000 90.905000 ;
      LAYER met4 ;
        RECT 13.780000 90.585000 14.100000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 90.995000 14.100000 91.315000 ;
      LAYER met4 ;
        RECT 13.780000 90.995000 14.100000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 91.405000 14.100000 91.725000 ;
      LAYER met4 ;
        RECT 13.780000 91.405000 14.100000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 91.815000 14.100000 92.135000 ;
      LAYER met4 ;
        RECT 13.780000 91.815000 14.100000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 92.225000 14.100000 92.545000 ;
      LAYER met4 ;
        RECT 13.780000 92.225000 14.100000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780000 92.635000 14.100000 92.955000 ;
      LAYER met4 ;
        RECT 13.780000 92.635000 14.100000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 68.065000 14.305000 68.385000 ;
      LAYER met4 ;
        RECT 13.985000 68.065000 14.305000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 68.475000 14.305000 68.795000 ;
      LAYER met4 ;
        RECT 13.985000 68.475000 14.305000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 68.885000 14.305000 69.205000 ;
      LAYER met4 ;
        RECT 13.985000 68.885000 14.305000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 69.295000 14.305000 69.615000 ;
      LAYER met4 ;
        RECT 13.985000 69.295000 14.305000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 69.705000 14.305000 70.025000 ;
      LAYER met4 ;
        RECT 13.985000 69.705000 14.305000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 70.115000 14.305000 70.435000 ;
      LAYER met4 ;
        RECT 13.985000 70.115000 14.305000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 70.525000 14.305000 70.845000 ;
      LAYER met4 ;
        RECT 13.985000 70.525000 14.305000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 70.935000 14.305000 71.255000 ;
      LAYER met4 ;
        RECT 13.985000 70.935000 14.305000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 71.345000 14.305000 71.665000 ;
      LAYER met4 ;
        RECT 13.985000 71.345000 14.305000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 71.755000 14.305000 72.075000 ;
      LAYER met4 ;
        RECT 13.985000 71.755000 14.305000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 72.165000 14.305000 72.485000 ;
      LAYER met4 ;
        RECT 13.985000 72.165000 14.305000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 72.575000 14.305000 72.895000 ;
      LAYER met4 ;
        RECT 13.985000 72.575000 14.305000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 72.985000 14.305000 73.305000 ;
      LAYER met4 ;
        RECT 13.985000 72.985000 14.305000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 73.390000 14.305000 73.710000 ;
      LAYER met4 ;
        RECT 13.985000 73.390000 14.305000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 73.795000 14.305000 74.115000 ;
      LAYER met4 ;
        RECT 13.985000 73.795000 14.305000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 74.200000 14.305000 74.520000 ;
      LAYER met4 ;
        RECT 13.985000 74.200000 14.305000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 74.605000 14.305000 74.925000 ;
      LAYER met4 ;
        RECT 13.985000 74.605000 14.305000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 75.010000 14.305000 75.330000 ;
      LAYER met4 ;
        RECT 13.985000 75.010000 14.305000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 75.415000 14.305000 75.735000 ;
      LAYER met4 ;
        RECT 13.985000 75.415000 14.305000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 75.820000 14.305000 76.140000 ;
      LAYER met4 ;
        RECT 13.985000 75.820000 14.305000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 76.225000 14.305000 76.545000 ;
      LAYER met4 ;
        RECT 13.985000 76.225000 14.305000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 76.630000 14.305000 76.950000 ;
      LAYER met4 ;
        RECT 13.985000 76.630000 14.305000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 77.035000 14.305000 77.355000 ;
      LAYER met4 ;
        RECT 13.985000 77.035000 14.305000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 77.440000 14.305000 77.760000 ;
      LAYER met4 ;
        RECT 13.985000 77.440000 14.305000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 77.845000 14.305000 78.165000 ;
      LAYER met4 ;
        RECT 13.985000 77.845000 14.305000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 78.250000 14.305000 78.570000 ;
      LAYER met4 ;
        RECT 13.985000 78.250000 14.305000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 78.655000 14.305000 78.975000 ;
      LAYER met4 ;
        RECT 13.985000 78.655000 14.305000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 79.060000 14.305000 79.380000 ;
      LAYER met4 ;
        RECT 13.985000 79.060000 14.305000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 79.465000 14.305000 79.785000 ;
      LAYER met4 ;
        RECT 13.985000 79.465000 14.305000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 79.870000 14.305000 80.190000 ;
      LAYER met4 ;
        RECT 13.985000 79.870000 14.305000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 80.275000 14.305000 80.595000 ;
      LAYER met4 ;
        RECT 13.985000 80.275000 14.305000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 80.680000 14.305000 81.000000 ;
      LAYER met4 ;
        RECT 13.985000 80.680000 14.305000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 81.085000 14.305000 81.405000 ;
      LAYER met4 ;
        RECT 13.985000 81.085000 14.305000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 81.490000 14.305000 81.810000 ;
      LAYER met4 ;
        RECT 13.985000 81.490000 14.305000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 81.895000 14.305000 82.215000 ;
      LAYER met4 ;
        RECT 13.985000 81.895000 14.305000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985000 82.300000 14.305000 82.620000 ;
      LAYER met4 ;
        RECT 13.985000 82.300000 14.305000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995000 17.800000 14.315000 18.120000 ;
      LAYER met4 ;
        RECT 13.995000 17.800000 14.315000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995000 18.230000 14.315000 18.550000 ;
      LAYER met4 ;
        RECT 13.995000 18.230000 14.315000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995000 18.660000 14.315000 18.980000 ;
      LAYER met4 ;
        RECT 13.995000 18.660000 14.315000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995000 19.090000 14.315000 19.410000 ;
      LAYER met4 ;
        RECT 13.995000 19.090000 14.315000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995000 19.520000 14.315000 19.840000 ;
      LAYER met4 ;
        RECT 13.995000 19.520000 14.315000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995000 19.950000 14.315000 20.270000 ;
      LAYER met4 ;
        RECT 13.995000 19.950000 14.315000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995000 20.380000 14.315000 20.700000 ;
      LAYER met4 ;
        RECT 13.995000 20.380000 14.315000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995000 20.810000 14.315000 21.130000 ;
      LAYER met4 ;
        RECT 13.995000 20.810000 14.315000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995000 21.240000 14.315000 21.560000 ;
      LAYER met4 ;
        RECT 13.995000 21.240000 14.315000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995000 21.670000 14.315000 21.990000 ;
      LAYER met4 ;
        RECT 13.995000 21.670000 14.315000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995000 22.100000 14.315000 22.420000 ;
      LAYER met4 ;
        RECT 13.995000 22.100000 14.315000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.260000 90.955000 14.580000 91.275000 ;
      LAYER met4 ;
        RECT 14.260000 90.955000 14.580000 91.275000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.260000 91.385000 14.580000 91.705000 ;
      LAYER met4 ;
        RECT 14.260000 91.385000 14.580000 91.705000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.280000 88.350000 14.600000 88.670000 ;
      LAYER met4 ;
        RECT 14.280000 88.350000 14.600000 88.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.280000 88.775000 14.600000 89.095000 ;
      LAYER met4 ;
        RECT 14.280000 88.775000 14.600000 89.095000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.280000 89.205000 14.600000 89.525000 ;
      LAYER met4 ;
        RECT 14.280000 89.205000 14.600000 89.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.280000 89.635000 14.600000 89.955000 ;
      LAYER met4 ;
        RECT 14.280000 89.635000 14.600000 89.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.280000 90.065000 14.600000 90.385000 ;
      LAYER met4 ;
        RECT 14.280000 90.065000 14.600000 90.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.280000 90.495000 14.600000 90.815000 ;
      LAYER met4 ;
        RECT 14.280000 90.495000 14.600000 90.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 68.065000 14.705000 68.385000 ;
      LAYER met4 ;
        RECT 14.385000 68.065000 14.705000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 68.475000 14.705000 68.795000 ;
      LAYER met4 ;
        RECT 14.385000 68.475000 14.705000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 68.885000 14.705000 69.205000 ;
      LAYER met4 ;
        RECT 14.385000 68.885000 14.705000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 69.295000 14.705000 69.615000 ;
      LAYER met4 ;
        RECT 14.385000 69.295000 14.705000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 69.705000 14.705000 70.025000 ;
      LAYER met4 ;
        RECT 14.385000 69.705000 14.705000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 70.115000 14.705000 70.435000 ;
      LAYER met4 ;
        RECT 14.385000 70.115000 14.705000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 70.525000 14.705000 70.845000 ;
      LAYER met4 ;
        RECT 14.385000 70.525000 14.705000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 70.935000 14.705000 71.255000 ;
      LAYER met4 ;
        RECT 14.385000 70.935000 14.705000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 71.345000 14.705000 71.665000 ;
      LAYER met4 ;
        RECT 14.385000 71.345000 14.705000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 71.755000 14.705000 72.075000 ;
      LAYER met4 ;
        RECT 14.385000 71.755000 14.705000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 72.165000 14.705000 72.485000 ;
      LAYER met4 ;
        RECT 14.385000 72.165000 14.705000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 72.575000 14.705000 72.895000 ;
      LAYER met4 ;
        RECT 14.385000 72.575000 14.705000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 72.985000 14.705000 73.305000 ;
      LAYER met4 ;
        RECT 14.385000 72.985000 14.705000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 73.390000 14.705000 73.710000 ;
      LAYER met4 ;
        RECT 14.385000 73.390000 14.705000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 73.795000 14.705000 74.115000 ;
      LAYER met4 ;
        RECT 14.385000 73.795000 14.705000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 74.200000 14.705000 74.520000 ;
      LAYER met4 ;
        RECT 14.385000 74.200000 14.705000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 74.605000 14.705000 74.925000 ;
      LAYER met4 ;
        RECT 14.385000 74.605000 14.705000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 75.010000 14.705000 75.330000 ;
      LAYER met4 ;
        RECT 14.385000 75.010000 14.705000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 75.415000 14.705000 75.735000 ;
      LAYER met4 ;
        RECT 14.385000 75.415000 14.705000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 75.820000 14.705000 76.140000 ;
      LAYER met4 ;
        RECT 14.385000 75.820000 14.705000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 76.225000 14.705000 76.545000 ;
      LAYER met4 ;
        RECT 14.385000 76.225000 14.705000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 76.630000 14.705000 76.950000 ;
      LAYER met4 ;
        RECT 14.385000 76.630000 14.705000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 77.035000 14.705000 77.355000 ;
      LAYER met4 ;
        RECT 14.385000 77.035000 14.705000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 77.440000 14.705000 77.760000 ;
      LAYER met4 ;
        RECT 14.385000 77.440000 14.705000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 77.845000 14.705000 78.165000 ;
      LAYER met4 ;
        RECT 14.385000 77.845000 14.705000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 78.250000 14.705000 78.570000 ;
      LAYER met4 ;
        RECT 14.385000 78.250000 14.705000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 78.655000 14.705000 78.975000 ;
      LAYER met4 ;
        RECT 14.385000 78.655000 14.705000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 79.060000 14.705000 79.380000 ;
      LAYER met4 ;
        RECT 14.385000 79.060000 14.705000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 79.465000 14.705000 79.785000 ;
      LAYER met4 ;
        RECT 14.385000 79.465000 14.705000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 79.870000 14.705000 80.190000 ;
      LAYER met4 ;
        RECT 14.385000 79.870000 14.705000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 80.275000 14.705000 80.595000 ;
      LAYER met4 ;
        RECT 14.385000 80.275000 14.705000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 80.680000 14.705000 81.000000 ;
      LAYER met4 ;
        RECT 14.385000 80.680000 14.705000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 81.085000 14.705000 81.405000 ;
      LAYER met4 ;
        RECT 14.385000 81.085000 14.705000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 81.490000 14.705000 81.810000 ;
      LAYER met4 ;
        RECT 14.385000 81.490000 14.705000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 81.895000 14.705000 82.215000 ;
      LAYER met4 ;
        RECT 14.385000 81.895000 14.705000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385000 82.300000 14.705000 82.620000 ;
      LAYER met4 ;
        RECT 14.385000 82.300000 14.705000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400000 17.800000 14.720000 18.120000 ;
      LAYER met4 ;
        RECT 14.400000 17.800000 14.720000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400000 18.230000 14.720000 18.550000 ;
      LAYER met4 ;
        RECT 14.400000 18.230000 14.720000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400000 18.660000 14.720000 18.980000 ;
      LAYER met4 ;
        RECT 14.400000 18.660000 14.720000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400000 19.090000 14.720000 19.410000 ;
      LAYER met4 ;
        RECT 14.400000 19.090000 14.720000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400000 19.520000 14.720000 19.840000 ;
      LAYER met4 ;
        RECT 14.400000 19.520000 14.720000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400000 19.950000 14.720000 20.270000 ;
      LAYER met4 ;
        RECT 14.400000 19.950000 14.720000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400000 20.380000 14.720000 20.700000 ;
      LAYER met4 ;
        RECT 14.400000 20.380000 14.720000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400000 20.810000 14.720000 21.130000 ;
      LAYER met4 ;
        RECT 14.400000 20.810000 14.720000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400000 21.240000 14.720000 21.560000 ;
      LAYER met4 ;
        RECT 14.400000 21.240000 14.720000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400000 21.670000 14.720000 21.990000 ;
      LAYER met4 ;
        RECT 14.400000 21.670000 14.720000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400000 22.100000 14.720000 22.420000 ;
      LAYER met4 ;
        RECT 14.400000 22.100000 14.720000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405000 82.995000 14.725000 83.315000 ;
      LAYER met4 ;
        RECT 14.405000 82.995000 14.725000 83.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405000 83.395000 14.725000 83.715000 ;
      LAYER met4 ;
        RECT 14.405000 83.395000 14.725000 83.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405000 83.795000 14.725000 84.115000 ;
      LAYER met4 ;
        RECT 14.405000 83.795000 14.725000 84.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405000 84.195000 14.725000 84.515000 ;
      LAYER met4 ;
        RECT 14.405000 84.195000 14.725000 84.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405000 84.595000 14.725000 84.915000 ;
      LAYER met4 ;
        RECT 14.405000 84.595000 14.725000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405000 84.995000 14.725000 85.315000 ;
      LAYER met4 ;
        RECT 14.405000 84.995000 14.725000 85.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405000 85.395000 14.725000 85.715000 ;
      LAYER met4 ;
        RECT 14.405000 85.395000 14.725000 85.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405000 85.795000 14.725000 86.115000 ;
      LAYER met4 ;
        RECT 14.405000 85.795000 14.725000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405000 86.195000 14.725000 86.515000 ;
      LAYER met4 ;
        RECT 14.405000 86.195000 14.725000 86.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405000 86.600000 14.725000 86.920000 ;
      LAYER met4 ;
        RECT 14.405000 86.600000 14.725000 86.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405000 87.005000 14.725000 87.325000 ;
      LAYER met4 ;
        RECT 14.405000 87.005000 14.725000 87.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405000 87.410000 14.725000 87.730000 ;
      LAYER met4 ;
        RECT 14.405000 87.410000 14.725000 87.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405000 87.815000 14.725000 88.135000 ;
      LAYER met4 ;
        RECT 14.405000 87.815000 14.725000 88.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.690000 88.350000 15.010000 88.670000 ;
      LAYER met4 ;
        RECT 14.690000 88.350000 15.010000 88.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.690000 88.775000 15.010000 89.095000 ;
      LAYER met4 ;
        RECT 14.690000 88.775000 15.010000 89.095000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.690000 89.205000 15.010000 89.525000 ;
      LAYER met4 ;
        RECT 14.690000 89.205000 15.010000 89.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.690000 89.635000 15.010000 89.955000 ;
      LAYER met4 ;
        RECT 14.690000 89.635000 15.010000 89.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.690000 90.065000 15.010000 90.385000 ;
      LAYER met4 ;
        RECT 14.690000 90.065000 15.010000 90.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.690000 90.495000 15.010000 90.815000 ;
      LAYER met4 ;
        RECT 14.690000 90.495000 15.010000 90.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 68.065000 15.105000 68.385000 ;
      LAYER met4 ;
        RECT 14.785000 68.065000 15.105000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 68.475000 15.105000 68.795000 ;
      LAYER met4 ;
        RECT 14.785000 68.475000 15.105000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 68.885000 15.105000 69.205000 ;
      LAYER met4 ;
        RECT 14.785000 68.885000 15.105000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 69.295000 15.105000 69.615000 ;
      LAYER met4 ;
        RECT 14.785000 69.295000 15.105000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 69.705000 15.105000 70.025000 ;
      LAYER met4 ;
        RECT 14.785000 69.705000 15.105000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 70.115000 15.105000 70.435000 ;
      LAYER met4 ;
        RECT 14.785000 70.115000 15.105000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 70.525000 15.105000 70.845000 ;
      LAYER met4 ;
        RECT 14.785000 70.525000 15.105000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 70.935000 15.105000 71.255000 ;
      LAYER met4 ;
        RECT 14.785000 70.935000 15.105000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 71.345000 15.105000 71.665000 ;
      LAYER met4 ;
        RECT 14.785000 71.345000 15.105000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 71.755000 15.105000 72.075000 ;
      LAYER met4 ;
        RECT 14.785000 71.755000 15.105000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 72.165000 15.105000 72.485000 ;
      LAYER met4 ;
        RECT 14.785000 72.165000 15.105000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 72.575000 15.105000 72.895000 ;
      LAYER met4 ;
        RECT 14.785000 72.575000 15.105000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 72.985000 15.105000 73.305000 ;
      LAYER met4 ;
        RECT 14.785000 72.985000 15.105000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 73.390000 15.105000 73.710000 ;
      LAYER met4 ;
        RECT 14.785000 73.390000 15.105000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 73.795000 15.105000 74.115000 ;
      LAYER met4 ;
        RECT 14.785000 73.795000 15.105000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 74.200000 15.105000 74.520000 ;
      LAYER met4 ;
        RECT 14.785000 74.200000 15.105000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 74.605000 15.105000 74.925000 ;
      LAYER met4 ;
        RECT 14.785000 74.605000 15.105000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 75.010000 15.105000 75.330000 ;
      LAYER met4 ;
        RECT 14.785000 75.010000 15.105000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 75.415000 15.105000 75.735000 ;
      LAYER met4 ;
        RECT 14.785000 75.415000 15.105000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 75.820000 15.105000 76.140000 ;
      LAYER met4 ;
        RECT 14.785000 75.820000 15.105000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 76.225000 15.105000 76.545000 ;
      LAYER met4 ;
        RECT 14.785000 76.225000 15.105000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 76.630000 15.105000 76.950000 ;
      LAYER met4 ;
        RECT 14.785000 76.630000 15.105000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 77.035000 15.105000 77.355000 ;
      LAYER met4 ;
        RECT 14.785000 77.035000 15.105000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 77.440000 15.105000 77.760000 ;
      LAYER met4 ;
        RECT 14.785000 77.440000 15.105000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 77.845000 15.105000 78.165000 ;
      LAYER met4 ;
        RECT 14.785000 77.845000 15.105000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 78.250000 15.105000 78.570000 ;
      LAYER met4 ;
        RECT 14.785000 78.250000 15.105000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 78.655000 15.105000 78.975000 ;
      LAYER met4 ;
        RECT 14.785000 78.655000 15.105000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 79.060000 15.105000 79.380000 ;
      LAYER met4 ;
        RECT 14.785000 79.060000 15.105000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 79.465000 15.105000 79.785000 ;
      LAYER met4 ;
        RECT 14.785000 79.465000 15.105000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 79.870000 15.105000 80.190000 ;
      LAYER met4 ;
        RECT 14.785000 79.870000 15.105000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 80.275000 15.105000 80.595000 ;
      LAYER met4 ;
        RECT 14.785000 80.275000 15.105000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 80.680000 15.105000 81.000000 ;
      LAYER met4 ;
        RECT 14.785000 80.680000 15.105000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 81.085000 15.105000 81.405000 ;
      LAYER met4 ;
        RECT 14.785000 81.085000 15.105000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 81.490000 15.105000 81.810000 ;
      LAYER met4 ;
        RECT 14.785000 81.490000 15.105000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 81.895000 15.105000 82.215000 ;
      LAYER met4 ;
        RECT 14.785000 81.895000 15.105000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785000 82.300000 15.105000 82.620000 ;
      LAYER met4 ;
        RECT 14.785000 82.300000 15.105000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805000 17.800000 15.125000 18.120000 ;
      LAYER met4 ;
        RECT 14.805000 17.800000 15.125000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805000 18.230000 15.125000 18.550000 ;
      LAYER met4 ;
        RECT 14.805000 18.230000 15.125000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805000 18.660000 15.125000 18.980000 ;
      LAYER met4 ;
        RECT 14.805000 18.660000 15.125000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805000 19.090000 15.125000 19.410000 ;
      LAYER met4 ;
        RECT 14.805000 19.090000 15.125000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805000 19.520000 15.125000 19.840000 ;
      LAYER met4 ;
        RECT 14.805000 19.520000 15.125000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805000 19.950000 15.125000 20.270000 ;
      LAYER met4 ;
        RECT 14.805000 19.950000 15.125000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805000 20.380000 15.125000 20.700000 ;
      LAYER met4 ;
        RECT 14.805000 20.380000 15.125000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805000 20.810000 15.125000 21.130000 ;
      LAYER met4 ;
        RECT 14.805000 20.810000 15.125000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805000 21.240000 15.125000 21.560000 ;
      LAYER met4 ;
        RECT 14.805000 21.240000 15.125000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805000 21.670000 15.125000 21.990000 ;
      LAYER met4 ;
        RECT 14.805000 21.670000 15.125000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805000 22.100000 15.125000 22.420000 ;
      LAYER met4 ;
        RECT 14.805000 22.100000 15.125000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815000 82.995000 15.135000 83.315000 ;
      LAYER met4 ;
        RECT 14.815000 82.995000 15.135000 83.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815000 83.395000 15.135000 83.715000 ;
      LAYER met4 ;
        RECT 14.815000 83.395000 15.135000 83.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815000 83.795000 15.135000 84.115000 ;
      LAYER met4 ;
        RECT 14.815000 83.795000 15.135000 84.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815000 84.195000 15.135000 84.515000 ;
      LAYER met4 ;
        RECT 14.815000 84.195000 15.135000 84.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815000 84.595000 15.135000 84.915000 ;
      LAYER met4 ;
        RECT 14.815000 84.595000 15.135000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815000 84.995000 15.135000 85.315000 ;
      LAYER met4 ;
        RECT 14.815000 84.995000 15.135000 85.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815000 85.395000 15.135000 85.715000 ;
      LAYER met4 ;
        RECT 14.815000 85.395000 15.135000 85.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815000 85.795000 15.135000 86.115000 ;
      LAYER met4 ;
        RECT 14.815000 85.795000 15.135000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815000 86.195000 15.135000 86.515000 ;
      LAYER met4 ;
        RECT 14.815000 86.195000 15.135000 86.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815000 86.600000 15.135000 86.920000 ;
      LAYER met4 ;
        RECT 14.815000 86.600000 15.135000 86.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815000 87.005000 15.135000 87.325000 ;
      LAYER met4 ;
        RECT 14.815000 87.005000 15.135000 87.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815000 87.410000 15.135000 87.730000 ;
      LAYER met4 ;
        RECT 14.815000 87.410000 15.135000 87.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815000 87.815000 15.135000 88.135000 ;
      LAYER met4 ;
        RECT 14.815000 87.815000 15.135000 88.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.040000 90.955000 15.360000 91.275000 ;
      LAYER met4 ;
        RECT 15.040000 90.955000 15.360000 91.275000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.040000 91.385000 15.360000 91.705000 ;
      LAYER met4 ;
        RECT 15.040000 91.385000 15.360000 91.705000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.100000 88.350000 15.420000 88.670000 ;
      LAYER met4 ;
        RECT 15.100000 88.350000 15.420000 88.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.100000 88.775000 15.420000 89.095000 ;
      LAYER met4 ;
        RECT 15.100000 88.775000 15.420000 89.095000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.100000 89.205000 15.420000 89.525000 ;
      LAYER met4 ;
        RECT 15.100000 89.205000 15.420000 89.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.100000 89.635000 15.420000 89.955000 ;
      LAYER met4 ;
        RECT 15.100000 89.635000 15.420000 89.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.100000 90.065000 15.420000 90.385000 ;
      LAYER met4 ;
        RECT 15.100000 90.065000 15.420000 90.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.100000 90.495000 15.420000 90.815000 ;
      LAYER met4 ;
        RECT 15.100000 90.495000 15.420000 90.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 68.065000 15.505000 68.385000 ;
      LAYER met4 ;
        RECT 15.185000 68.065000 15.505000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 68.475000 15.505000 68.795000 ;
      LAYER met4 ;
        RECT 15.185000 68.475000 15.505000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 68.885000 15.505000 69.205000 ;
      LAYER met4 ;
        RECT 15.185000 68.885000 15.505000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 69.295000 15.505000 69.615000 ;
      LAYER met4 ;
        RECT 15.185000 69.295000 15.505000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 69.705000 15.505000 70.025000 ;
      LAYER met4 ;
        RECT 15.185000 69.705000 15.505000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 70.115000 15.505000 70.435000 ;
      LAYER met4 ;
        RECT 15.185000 70.115000 15.505000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 70.525000 15.505000 70.845000 ;
      LAYER met4 ;
        RECT 15.185000 70.525000 15.505000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 70.935000 15.505000 71.255000 ;
      LAYER met4 ;
        RECT 15.185000 70.935000 15.505000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 71.345000 15.505000 71.665000 ;
      LAYER met4 ;
        RECT 15.185000 71.345000 15.505000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 71.755000 15.505000 72.075000 ;
      LAYER met4 ;
        RECT 15.185000 71.755000 15.505000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 72.165000 15.505000 72.485000 ;
      LAYER met4 ;
        RECT 15.185000 72.165000 15.505000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 72.575000 15.505000 72.895000 ;
      LAYER met4 ;
        RECT 15.185000 72.575000 15.505000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 72.985000 15.505000 73.305000 ;
      LAYER met4 ;
        RECT 15.185000 72.985000 15.505000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 73.390000 15.505000 73.710000 ;
      LAYER met4 ;
        RECT 15.185000 73.390000 15.505000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 73.795000 15.505000 74.115000 ;
      LAYER met4 ;
        RECT 15.185000 73.795000 15.505000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 74.200000 15.505000 74.520000 ;
      LAYER met4 ;
        RECT 15.185000 74.200000 15.505000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 74.605000 15.505000 74.925000 ;
      LAYER met4 ;
        RECT 15.185000 74.605000 15.505000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 75.010000 15.505000 75.330000 ;
      LAYER met4 ;
        RECT 15.185000 75.010000 15.505000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 75.415000 15.505000 75.735000 ;
      LAYER met4 ;
        RECT 15.185000 75.415000 15.505000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 75.820000 15.505000 76.140000 ;
      LAYER met4 ;
        RECT 15.185000 75.820000 15.505000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 76.225000 15.505000 76.545000 ;
      LAYER met4 ;
        RECT 15.185000 76.225000 15.505000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 76.630000 15.505000 76.950000 ;
      LAYER met4 ;
        RECT 15.185000 76.630000 15.505000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 77.035000 15.505000 77.355000 ;
      LAYER met4 ;
        RECT 15.185000 77.035000 15.505000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 77.440000 15.505000 77.760000 ;
      LAYER met4 ;
        RECT 15.185000 77.440000 15.505000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 77.845000 15.505000 78.165000 ;
      LAYER met4 ;
        RECT 15.185000 77.845000 15.505000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 78.250000 15.505000 78.570000 ;
      LAYER met4 ;
        RECT 15.185000 78.250000 15.505000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 78.655000 15.505000 78.975000 ;
      LAYER met4 ;
        RECT 15.185000 78.655000 15.505000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 79.060000 15.505000 79.380000 ;
      LAYER met4 ;
        RECT 15.185000 79.060000 15.505000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 79.465000 15.505000 79.785000 ;
      LAYER met4 ;
        RECT 15.185000 79.465000 15.505000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 79.870000 15.505000 80.190000 ;
      LAYER met4 ;
        RECT 15.185000 79.870000 15.505000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 80.275000 15.505000 80.595000 ;
      LAYER met4 ;
        RECT 15.185000 80.275000 15.505000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 80.680000 15.505000 81.000000 ;
      LAYER met4 ;
        RECT 15.185000 80.680000 15.505000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 81.085000 15.505000 81.405000 ;
      LAYER met4 ;
        RECT 15.185000 81.085000 15.505000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 81.490000 15.505000 81.810000 ;
      LAYER met4 ;
        RECT 15.185000 81.490000 15.505000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 81.895000 15.505000 82.215000 ;
      LAYER met4 ;
        RECT 15.185000 81.895000 15.505000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185000 82.300000 15.505000 82.620000 ;
      LAYER met4 ;
        RECT 15.185000 82.300000 15.505000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210000 17.800000 15.530000 18.120000 ;
      LAYER met4 ;
        RECT 15.210000 17.800000 15.530000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210000 18.230000 15.530000 18.550000 ;
      LAYER met4 ;
        RECT 15.210000 18.230000 15.530000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210000 18.660000 15.530000 18.980000 ;
      LAYER met4 ;
        RECT 15.210000 18.660000 15.530000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210000 19.090000 15.530000 19.410000 ;
      LAYER met4 ;
        RECT 15.210000 19.090000 15.530000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210000 19.520000 15.530000 19.840000 ;
      LAYER met4 ;
        RECT 15.210000 19.520000 15.530000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210000 19.950000 15.530000 20.270000 ;
      LAYER met4 ;
        RECT 15.210000 19.950000 15.530000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210000 20.380000 15.530000 20.700000 ;
      LAYER met4 ;
        RECT 15.210000 20.380000 15.530000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210000 20.810000 15.530000 21.130000 ;
      LAYER met4 ;
        RECT 15.210000 20.810000 15.530000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210000 21.240000 15.530000 21.560000 ;
      LAYER met4 ;
        RECT 15.210000 21.240000 15.530000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210000 21.670000 15.530000 21.990000 ;
      LAYER met4 ;
        RECT 15.210000 21.670000 15.530000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210000 22.100000 15.530000 22.420000 ;
      LAYER met4 ;
        RECT 15.210000 22.100000 15.530000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225000 82.995000 15.545000 83.315000 ;
      LAYER met4 ;
        RECT 15.225000 82.995000 15.545000 83.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225000 83.395000 15.545000 83.715000 ;
      LAYER met4 ;
        RECT 15.225000 83.395000 15.545000 83.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225000 83.795000 15.545000 84.115000 ;
      LAYER met4 ;
        RECT 15.225000 83.795000 15.545000 84.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225000 84.195000 15.545000 84.515000 ;
      LAYER met4 ;
        RECT 15.225000 84.195000 15.545000 84.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225000 84.595000 15.545000 84.915000 ;
      LAYER met4 ;
        RECT 15.225000 84.595000 15.545000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225000 84.995000 15.545000 85.315000 ;
      LAYER met4 ;
        RECT 15.225000 84.995000 15.545000 85.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225000 85.395000 15.545000 85.715000 ;
      LAYER met4 ;
        RECT 15.225000 85.395000 15.545000 85.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225000 85.795000 15.545000 86.115000 ;
      LAYER met4 ;
        RECT 15.225000 85.795000 15.545000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225000 86.195000 15.545000 86.515000 ;
      LAYER met4 ;
        RECT 15.225000 86.195000 15.545000 86.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225000 86.600000 15.545000 86.920000 ;
      LAYER met4 ;
        RECT 15.225000 86.600000 15.545000 86.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225000 87.005000 15.545000 87.325000 ;
      LAYER met4 ;
        RECT 15.225000 87.005000 15.545000 87.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225000 87.410000 15.545000 87.730000 ;
      LAYER met4 ;
        RECT 15.225000 87.410000 15.545000 87.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225000 87.815000 15.545000 88.135000 ;
      LAYER met4 ;
        RECT 15.225000 87.815000 15.545000 88.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.510000 88.350000 15.830000 88.670000 ;
      LAYER met4 ;
        RECT 15.510000 88.350000 15.830000 88.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.510000 88.775000 15.830000 89.095000 ;
      LAYER met4 ;
        RECT 15.510000 88.775000 15.830000 89.095000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.510000 89.205000 15.830000 89.525000 ;
      LAYER met4 ;
        RECT 15.510000 89.205000 15.830000 89.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.510000 89.635000 15.830000 89.955000 ;
      LAYER met4 ;
        RECT 15.510000 89.635000 15.830000 89.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.510000 90.065000 15.830000 90.385000 ;
      LAYER met4 ;
        RECT 15.510000 90.065000 15.830000 90.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.510000 90.495000 15.830000 90.815000 ;
      LAYER met4 ;
        RECT 15.510000 90.495000 15.830000 90.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 68.065000 15.905000 68.385000 ;
      LAYER met4 ;
        RECT 15.585000 68.065000 15.905000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 68.475000 15.905000 68.795000 ;
      LAYER met4 ;
        RECT 15.585000 68.475000 15.905000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 68.885000 15.905000 69.205000 ;
      LAYER met4 ;
        RECT 15.585000 68.885000 15.905000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 69.295000 15.905000 69.615000 ;
      LAYER met4 ;
        RECT 15.585000 69.295000 15.905000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 69.705000 15.905000 70.025000 ;
      LAYER met4 ;
        RECT 15.585000 69.705000 15.905000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 70.115000 15.905000 70.435000 ;
      LAYER met4 ;
        RECT 15.585000 70.115000 15.905000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 70.525000 15.905000 70.845000 ;
      LAYER met4 ;
        RECT 15.585000 70.525000 15.905000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 70.935000 15.905000 71.255000 ;
      LAYER met4 ;
        RECT 15.585000 70.935000 15.905000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 71.345000 15.905000 71.665000 ;
      LAYER met4 ;
        RECT 15.585000 71.345000 15.905000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 71.755000 15.905000 72.075000 ;
      LAYER met4 ;
        RECT 15.585000 71.755000 15.905000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 72.165000 15.905000 72.485000 ;
      LAYER met4 ;
        RECT 15.585000 72.165000 15.905000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 72.575000 15.905000 72.895000 ;
      LAYER met4 ;
        RECT 15.585000 72.575000 15.905000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 72.985000 15.905000 73.305000 ;
      LAYER met4 ;
        RECT 15.585000 72.985000 15.905000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 73.390000 15.905000 73.710000 ;
      LAYER met4 ;
        RECT 15.585000 73.390000 15.905000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 73.795000 15.905000 74.115000 ;
      LAYER met4 ;
        RECT 15.585000 73.795000 15.905000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 74.200000 15.905000 74.520000 ;
      LAYER met4 ;
        RECT 15.585000 74.200000 15.905000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 74.605000 15.905000 74.925000 ;
      LAYER met4 ;
        RECT 15.585000 74.605000 15.905000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 75.010000 15.905000 75.330000 ;
      LAYER met4 ;
        RECT 15.585000 75.010000 15.905000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 75.415000 15.905000 75.735000 ;
      LAYER met4 ;
        RECT 15.585000 75.415000 15.905000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 75.820000 15.905000 76.140000 ;
      LAYER met4 ;
        RECT 15.585000 75.820000 15.905000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 76.225000 15.905000 76.545000 ;
      LAYER met4 ;
        RECT 15.585000 76.225000 15.905000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 76.630000 15.905000 76.950000 ;
      LAYER met4 ;
        RECT 15.585000 76.630000 15.905000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 77.035000 15.905000 77.355000 ;
      LAYER met4 ;
        RECT 15.585000 77.035000 15.905000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 77.440000 15.905000 77.760000 ;
      LAYER met4 ;
        RECT 15.585000 77.440000 15.905000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 77.845000 15.905000 78.165000 ;
      LAYER met4 ;
        RECT 15.585000 77.845000 15.905000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 78.250000 15.905000 78.570000 ;
      LAYER met4 ;
        RECT 15.585000 78.250000 15.905000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 78.655000 15.905000 78.975000 ;
      LAYER met4 ;
        RECT 15.585000 78.655000 15.905000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 79.060000 15.905000 79.380000 ;
      LAYER met4 ;
        RECT 15.585000 79.060000 15.905000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 79.465000 15.905000 79.785000 ;
      LAYER met4 ;
        RECT 15.585000 79.465000 15.905000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 79.870000 15.905000 80.190000 ;
      LAYER met4 ;
        RECT 15.585000 79.870000 15.905000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 80.275000 15.905000 80.595000 ;
      LAYER met4 ;
        RECT 15.585000 80.275000 15.905000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 80.680000 15.905000 81.000000 ;
      LAYER met4 ;
        RECT 15.585000 80.680000 15.905000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 81.085000 15.905000 81.405000 ;
      LAYER met4 ;
        RECT 15.585000 81.085000 15.905000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 81.490000 15.905000 81.810000 ;
      LAYER met4 ;
        RECT 15.585000 81.490000 15.905000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 81.895000 15.905000 82.215000 ;
      LAYER met4 ;
        RECT 15.585000 81.895000 15.905000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585000 82.300000 15.905000 82.620000 ;
      LAYER met4 ;
        RECT 15.585000 82.300000 15.905000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615000 17.800000 15.935000 18.120000 ;
      LAYER met4 ;
        RECT 15.615000 17.800000 15.935000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615000 18.230000 15.935000 18.550000 ;
      LAYER met4 ;
        RECT 15.615000 18.230000 15.935000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615000 18.660000 15.935000 18.980000 ;
      LAYER met4 ;
        RECT 15.615000 18.660000 15.935000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615000 19.090000 15.935000 19.410000 ;
      LAYER met4 ;
        RECT 15.615000 19.090000 15.935000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615000 19.520000 15.935000 19.840000 ;
      LAYER met4 ;
        RECT 15.615000 19.520000 15.935000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615000 19.950000 15.935000 20.270000 ;
      LAYER met4 ;
        RECT 15.615000 19.950000 15.935000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615000 20.380000 15.935000 20.700000 ;
      LAYER met4 ;
        RECT 15.615000 20.380000 15.935000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615000 20.810000 15.935000 21.130000 ;
      LAYER met4 ;
        RECT 15.615000 20.810000 15.935000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615000 21.240000 15.935000 21.560000 ;
      LAYER met4 ;
        RECT 15.615000 21.240000 15.935000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615000 21.670000 15.935000 21.990000 ;
      LAYER met4 ;
        RECT 15.615000 21.670000 15.935000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615000 22.100000 15.935000 22.420000 ;
      LAYER met4 ;
        RECT 15.615000 22.100000 15.935000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635000 82.995000 15.955000 83.315000 ;
      LAYER met4 ;
        RECT 15.635000 82.995000 15.955000 83.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635000 83.395000 15.955000 83.715000 ;
      LAYER met4 ;
        RECT 15.635000 83.395000 15.955000 83.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635000 83.795000 15.955000 84.115000 ;
      LAYER met4 ;
        RECT 15.635000 83.795000 15.955000 84.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635000 84.195000 15.955000 84.515000 ;
      LAYER met4 ;
        RECT 15.635000 84.195000 15.955000 84.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635000 84.595000 15.955000 84.915000 ;
      LAYER met4 ;
        RECT 15.635000 84.595000 15.955000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635000 84.995000 15.955000 85.315000 ;
      LAYER met4 ;
        RECT 15.635000 84.995000 15.955000 85.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635000 85.395000 15.955000 85.715000 ;
      LAYER met4 ;
        RECT 15.635000 85.395000 15.955000 85.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635000 85.795000 15.955000 86.115000 ;
      LAYER met4 ;
        RECT 15.635000 85.795000 15.955000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635000 86.195000 15.955000 86.515000 ;
      LAYER met4 ;
        RECT 15.635000 86.195000 15.955000 86.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635000 86.600000 15.955000 86.920000 ;
      LAYER met4 ;
        RECT 15.635000 86.600000 15.955000 86.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635000 87.005000 15.955000 87.325000 ;
      LAYER met4 ;
        RECT 15.635000 87.005000 15.955000 87.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635000 87.410000 15.955000 87.730000 ;
      LAYER met4 ;
        RECT 15.635000 87.410000 15.955000 87.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635000 87.815000 15.955000 88.135000 ;
      LAYER met4 ;
        RECT 15.635000 87.815000 15.955000 88.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.920000 88.350000 16.240000 88.670000 ;
      LAYER met4 ;
        RECT 15.920000 88.350000 16.240000 88.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.920000 88.775000 16.240000 89.095000 ;
      LAYER met4 ;
        RECT 15.920000 88.775000 16.240000 89.095000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.920000 89.205000 16.240000 89.525000 ;
      LAYER met4 ;
        RECT 15.920000 89.205000 16.240000 89.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.920000 89.635000 16.240000 89.955000 ;
      LAYER met4 ;
        RECT 15.920000 89.635000 16.240000 89.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.920000 90.065000 16.240000 90.385000 ;
      LAYER met4 ;
        RECT 15.920000 90.065000 16.240000 90.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.920000 90.495000 16.240000 90.815000 ;
      LAYER met4 ;
        RECT 15.920000 90.495000 16.240000 90.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 68.065000 16.305000 68.385000 ;
      LAYER met4 ;
        RECT 15.985000 68.065000 16.305000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 68.475000 16.305000 68.795000 ;
      LAYER met4 ;
        RECT 15.985000 68.475000 16.305000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 68.885000 16.305000 69.205000 ;
      LAYER met4 ;
        RECT 15.985000 68.885000 16.305000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 69.295000 16.305000 69.615000 ;
      LAYER met4 ;
        RECT 15.985000 69.295000 16.305000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 69.705000 16.305000 70.025000 ;
      LAYER met4 ;
        RECT 15.985000 69.705000 16.305000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 70.115000 16.305000 70.435000 ;
      LAYER met4 ;
        RECT 15.985000 70.115000 16.305000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 70.525000 16.305000 70.845000 ;
      LAYER met4 ;
        RECT 15.985000 70.525000 16.305000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 70.935000 16.305000 71.255000 ;
      LAYER met4 ;
        RECT 15.985000 70.935000 16.305000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 71.345000 16.305000 71.665000 ;
      LAYER met4 ;
        RECT 15.985000 71.345000 16.305000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 71.755000 16.305000 72.075000 ;
      LAYER met4 ;
        RECT 15.985000 71.755000 16.305000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 72.165000 16.305000 72.485000 ;
      LAYER met4 ;
        RECT 15.985000 72.165000 16.305000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 72.575000 16.305000 72.895000 ;
      LAYER met4 ;
        RECT 15.985000 72.575000 16.305000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 72.985000 16.305000 73.305000 ;
      LAYER met4 ;
        RECT 15.985000 72.985000 16.305000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 73.390000 16.305000 73.710000 ;
      LAYER met4 ;
        RECT 15.985000 73.390000 16.305000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 73.795000 16.305000 74.115000 ;
      LAYER met4 ;
        RECT 15.985000 73.795000 16.305000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 74.200000 16.305000 74.520000 ;
      LAYER met4 ;
        RECT 15.985000 74.200000 16.305000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 74.605000 16.305000 74.925000 ;
      LAYER met4 ;
        RECT 15.985000 74.605000 16.305000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 75.010000 16.305000 75.330000 ;
      LAYER met4 ;
        RECT 15.985000 75.010000 16.305000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 75.415000 16.305000 75.735000 ;
      LAYER met4 ;
        RECT 15.985000 75.415000 16.305000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 75.820000 16.305000 76.140000 ;
      LAYER met4 ;
        RECT 15.985000 75.820000 16.305000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 76.225000 16.305000 76.545000 ;
      LAYER met4 ;
        RECT 15.985000 76.225000 16.305000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 76.630000 16.305000 76.950000 ;
      LAYER met4 ;
        RECT 15.985000 76.630000 16.305000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 77.035000 16.305000 77.355000 ;
      LAYER met4 ;
        RECT 15.985000 77.035000 16.305000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 77.440000 16.305000 77.760000 ;
      LAYER met4 ;
        RECT 15.985000 77.440000 16.305000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 77.845000 16.305000 78.165000 ;
      LAYER met4 ;
        RECT 15.985000 77.845000 16.305000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 78.250000 16.305000 78.570000 ;
      LAYER met4 ;
        RECT 15.985000 78.250000 16.305000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 78.655000 16.305000 78.975000 ;
      LAYER met4 ;
        RECT 15.985000 78.655000 16.305000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 79.060000 16.305000 79.380000 ;
      LAYER met4 ;
        RECT 15.985000 79.060000 16.305000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 79.465000 16.305000 79.785000 ;
      LAYER met4 ;
        RECT 15.985000 79.465000 16.305000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 79.870000 16.305000 80.190000 ;
      LAYER met4 ;
        RECT 15.985000 79.870000 16.305000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 80.275000 16.305000 80.595000 ;
      LAYER met4 ;
        RECT 15.985000 80.275000 16.305000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 80.680000 16.305000 81.000000 ;
      LAYER met4 ;
        RECT 15.985000 80.680000 16.305000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 81.085000 16.305000 81.405000 ;
      LAYER met4 ;
        RECT 15.985000 81.085000 16.305000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 81.490000 16.305000 81.810000 ;
      LAYER met4 ;
        RECT 15.985000 81.490000 16.305000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 81.895000 16.305000 82.215000 ;
      LAYER met4 ;
        RECT 15.985000 81.895000 16.305000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 82.300000 16.305000 82.620000 ;
      LAYER met4 ;
        RECT 15.985000 82.300000 16.305000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020000 17.800000 16.340000 18.120000 ;
      LAYER met4 ;
        RECT 16.020000 17.800000 16.340000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020000 18.230000 16.340000 18.550000 ;
      LAYER met4 ;
        RECT 16.020000 18.230000 16.340000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020000 18.660000 16.340000 18.980000 ;
      LAYER met4 ;
        RECT 16.020000 18.660000 16.340000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020000 19.090000 16.340000 19.410000 ;
      LAYER met4 ;
        RECT 16.020000 19.090000 16.340000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020000 19.520000 16.340000 19.840000 ;
      LAYER met4 ;
        RECT 16.020000 19.520000 16.340000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020000 19.950000 16.340000 20.270000 ;
      LAYER met4 ;
        RECT 16.020000 19.950000 16.340000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020000 20.380000 16.340000 20.700000 ;
      LAYER met4 ;
        RECT 16.020000 20.380000 16.340000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020000 20.810000 16.340000 21.130000 ;
      LAYER met4 ;
        RECT 16.020000 20.810000 16.340000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020000 21.240000 16.340000 21.560000 ;
      LAYER met4 ;
        RECT 16.020000 21.240000 16.340000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020000 21.670000 16.340000 21.990000 ;
      LAYER met4 ;
        RECT 16.020000 21.670000 16.340000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020000 22.100000 16.340000 22.420000 ;
      LAYER met4 ;
        RECT 16.020000 22.100000 16.340000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045000 82.995000 16.365000 83.315000 ;
      LAYER met4 ;
        RECT 16.045000 82.995000 16.365000 83.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045000 83.395000 16.365000 83.715000 ;
      LAYER met4 ;
        RECT 16.045000 83.395000 16.365000 83.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045000 83.795000 16.365000 84.115000 ;
      LAYER met4 ;
        RECT 16.045000 83.795000 16.365000 84.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045000 84.195000 16.365000 84.515000 ;
      LAYER met4 ;
        RECT 16.045000 84.195000 16.365000 84.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045000 84.595000 16.365000 84.915000 ;
      LAYER met4 ;
        RECT 16.045000 84.595000 16.365000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045000 84.995000 16.365000 85.315000 ;
      LAYER met4 ;
        RECT 16.045000 84.995000 16.365000 85.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045000 85.395000 16.365000 85.715000 ;
      LAYER met4 ;
        RECT 16.045000 85.395000 16.365000 85.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045000 85.795000 16.365000 86.115000 ;
      LAYER met4 ;
        RECT 16.045000 85.795000 16.365000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045000 86.195000 16.365000 86.515000 ;
      LAYER met4 ;
        RECT 16.045000 86.195000 16.365000 86.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045000 86.600000 16.365000 86.920000 ;
      LAYER met4 ;
        RECT 16.045000 86.600000 16.365000 86.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045000 87.005000 16.365000 87.325000 ;
      LAYER met4 ;
        RECT 16.045000 87.005000 16.365000 87.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045000 87.410000 16.365000 87.730000 ;
      LAYER met4 ;
        RECT 16.045000 87.410000 16.365000 87.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045000 87.815000 16.365000 88.135000 ;
      LAYER met4 ;
        RECT 16.045000 87.815000 16.365000 88.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 68.065000 16.705000 68.385000 ;
      LAYER met4 ;
        RECT 16.385000 68.065000 16.705000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 68.475000 16.705000 68.795000 ;
      LAYER met4 ;
        RECT 16.385000 68.475000 16.705000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 68.885000 16.705000 69.205000 ;
      LAYER met4 ;
        RECT 16.385000 68.885000 16.705000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 69.295000 16.705000 69.615000 ;
      LAYER met4 ;
        RECT 16.385000 69.295000 16.705000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 69.705000 16.705000 70.025000 ;
      LAYER met4 ;
        RECT 16.385000 69.705000 16.705000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 70.115000 16.705000 70.435000 ;
      LAYER met4 ;
        RECT 16.385000 70.115000 16.705000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 70.525000 16.705000 70.845000 ;
      LAYER met4 ;
        RECT 16.385000 70.525000 16.705000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 70.935000 16.705000 71.255000 ;
      LAYER met4 ;
        RECT 16.385000 70.935000 16.705000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 71.345000 16.705000 71.665000 ;
      LAYER met4 ;
        RECT 16.385000 71.345000 16.705000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 71.755000 16.705000 72.075000 ;
      LAYER met4 ;
        RECT 16.385000 71.755000 16.705000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 72.165000 16.705000 72.485000 ;
      LAYER met4 ;
        RECT 16.385000 72.165000 16.705000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 72.575000 16.705000 72.895000 ;
      LAYER met4 ;
        RECT 16.385000 72.575000 16.705000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 72.985000 16.705000 73.305000 ;
      LAYER met4 ;
        RECT 16.385000 72.985000 16.705000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 73.390000 16.705000 73.710000 ;
      LAYER met4 ;
        RECT 16.385000 73.390000 16.705000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 73.795000 16.705000 74.115000 ;
      LAYER met4 ;
        RECT 16.385000 73.795000 16.705000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 74.200000 16.705000 74.520000 ;
      LAYER met4 ;
        RECT 16.385000 74.200000 16.705000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 74.605000 16.705000 74.925000 ;
      LAYER met4 ;
        RECT 16.385000 74.605000 16.705000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 75.010000 16.705000 75.330000 ;
      LAYER met4 ;
        RECT 16.385000 75.010000 16.705000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 75.415000 16.705000 75.735000 ;
      LAYER met4 ;
        RECT 16.385000 75.415000 16.705000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 75.820000 16.705000 76.140000 ;
      LAYER met4 ;
        RECT 16.385000 75.820000 16.705000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 76.225000 16.705000 76.545000 ;
      LAYER met4 ;
        RECT 16.385000 76.225000 16.705000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 76.630000 16.705000 76.950000 ;
      LAYER met4 ;
        RECT 16.385000 76.630000 16.705000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 77.035000 16.705000 77.355000 ;
      LAYER met4 ;
        RECT 16.385000 77.035000 16.705000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 77.440000 16.705000 77.760000 ;
      LAYER met4 ;
        RECT 16.385000 77.440000 16.705000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 77.845000 16.705000 78.165000 ;
      LAYER met4 ;
        RECT 16.385000 77.845000 16.705000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 78.250000 16.705000 78.570000 ;
      LAYER met4 ;
        RECT 16.385000 78.250000 16.705000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 78.655000 16.705000 78.975000 ;
      LAYER met4 ;
        RECT 16.385000 78.655000 16.705000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 79.060000 16.705000 79.380000 ;
      LAYER met4 ;
        RECT 16.385000 79.060000 16.705000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 79.465000 16.705000 79.785000 ;
      LAYER met4 ;
        RECT 16.385000 79.465000 16.705000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 79.870000 16.705000 80.190000 ;
      LAYER met4 ;
        RECT 16.385000 79.870000 16.705000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 80.275000 16.705000 80.595000 ;
      LAYER met4 ;
        RECT 16.385000 80.275000 16.705000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 80.680000 16.705000 81.000000 ;
      LAYER met4 ;
        RECT 16.385000 80.680000 16.705000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 81.085000 16.705000 81.405000 ;
      LAYER met4 ;
        RECT 16.385000 81.085000 16.705000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 81.490000 16.705000 81.810000 ;
      LAYER met4 ;
        RECT 16.385000 81.490000 16.705000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 81.895000 16.705000 82.215000 ;
      LAYER met4 ;
        RECT 16.385000 81.895000 16.705000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385000 82.300000 16.705000 82.620000 ;
      LAYER met4 ;
        RECT 16.385000 82.300000 16.705000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.420000 88.370000 16.740000 88.690000 ;
      LAYER met4 ;
        RECT 16.420000 88.370000 16.740000 88.690000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.420000 88.785000 16.740000 89.105000 ;
      LAYER met4 ;
        RECT 16.420000 88.785000 16.740000 89.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.420000 89.205000 16.740000 89.525000 ;
      LAYER met4 ;
        RECT 16.420000 89.205000 16.740000 89.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425000 17.800000 16.745000 18.120000 ;
      LAYER met4 ;
        RECT 16.425000 17.800000 16.745000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425000 18.230000 16.745000 18.550000 ;
      LAYER met4 ;
        RECT 16.425000 18.230000 16.745000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425000 18.660000 16.745000 18.980000 ;
      LAYER met4 ;
        RECT 16.425000 18.660000 16.745000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425000 19.090000 16.745000 19.410000 ;
      LAYER met4 ;
        RECT 16.425000 19.090000 16.745000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425000 19.520000 16.745000 19.840000 ;
      LAYER met4 ;
        RECT 16.425000 19.520000 16.745000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425000 19.950000 16.745000 20.270000 ;
      LAYER met4 ;
        RECT 16.425000 19.950000 16.745000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425000 20.380000 16.745000 20.700000 ;
      LAYER met4 ;
        RECT 16.425000 20.380000 16.745000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425000 20.810000 16.745000 21.130000 ;
      LAYER met4 ;
        RECT 16.425000 20.810000 16.745000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425000 21.240000 16.745000 21.560000 ;
      LAYER met4 ;
        RECT 16.425000 21.240000 16.745000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425000 21.670000 16.745000 21.990000 ;
      LAYER met4 ;
        RECT 16.425000 21.670000 16.745000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425000 22.100000 16.745000 22.420000 ;
      LAYER met4 ;
        RECT 16.425000 22.100000 16.745000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 82.995000 16.775000 83.315000 ;
      LAYER met4 ;
        RECT 16.455000 82.995000 16.775000 83.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 83.395000 16.775000 83.715000 ;
      LAYER met4 ;
        RECT 16.455000 83.395000 16.775000 83.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 83.795000 16.775000 84.115000 ;
      LAYER met4 ;
        RECT 16.455000 83.795000 16.775000 84.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 84.195000 16.775000 84.515000 ;
      LAYER met4 ;
        RECT 16.455000 84.195000 16.775000 84.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 84.595000 16.775000 84.915000 ;
      LAYER met4 ;
        RECT 16.455000 84.595000 16.775000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 84.995000 16.775000 85.315000 ;
      LAYER met4 ;
        RECT 16.455000 84.995000 16.775000 85.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 85.395000 16.775000 85.715000 ;
      LAYER met4 ;
        RECT 16.455000 85.395000 16.775000 85.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 85.795000 16.775000 86.115000 ;
      LAYER met4 ;
        RECT 16.455000 85.795000 16.775000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 86.195000 16.775000 86.515000 ;
      LAYER met4 ;
        RECT 16.455000 86.195000 16.775000 86.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 86.600000 16.775000 86.920000 ;
      LAYER met4 ;
        RECT 16.455000 86.600000 16.775000 86.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 87.005000 16.775000 87.325000 ;
      LAYER met4 ;
        RECT 16.455000 87.005000 16.775000 87.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 87.410000 16.775000 87.730000 ;
      LAYER met4 ;
        RECT 16.455000 87.410000 16.775000 87.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 87.815000 16.775000 88.135000 ;
      LAYER met4 ;
        RECT 16.455000 87.815000 16.775000 88.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 68.065000 17.105000 68.385000 ;
      LAYER met4 ;
        RECT 16.785000 68.065000 17.105000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 68.475000 17.105000 68.795000 ;
      LAYER met4 ;
        RECT 16.785000 68.475000 17.105000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 68.885000 17.105000 69.205000 ;
      LAYER met4 ;
        RECT 16.785000 68.885000 17.105000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 69.295000 17.105000 69.615000 ;
      LAYER met4 ;
        RECT 16.785000 69.295000 17.105000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 69.705000 17.105000 70.025000 ;
      LAYER met4 ;
        RECT 16.785000 69.705000 17.105000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 70.115000 17.105000 70.435000 ;
      LAYER met4 ;
        RECT 16.785000 70.115000 17.105000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 70.525000 17.105000 70.845000 ;
      LAYER met4 ;
        RECT 16.785000 70.525000 17.105000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 70.935000 17.105000 71.255000 ;
      LAYER met4 ;
        RECT 16.785000 70.935000 17.105000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 71.345000 17.105000 71.665000 ;
      LAYER met4 ;
        RECT 16.785000 71.345000 17.105000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 71.755000 17.105000 72.075000 ;
      LAYER met4 ;
        RECT 16.785000 71.755000 17.105000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 72.165000 17.105000 72.485000 ;
      LAYER met4 ;
        RECT 16.785000 72.165000 17.105000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 72.575000 17.105000 72.895000 ;
      LAYER met4 ;
        RECT 16.785000 72.575000 17.105000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 72.985000 17.105000 73.305000 ;
      LAYER met4 ;
        RECT 16.785000 72.985000 17.105000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 73.390000 17.105000 73.710000 ;
      LAYER met4 ;
        RECT 16.785000 73.390000 17.105000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 73.795000 17.105000 74.115000 ;
      LAYER met4 ;
        RECT 16.785000 73.795000 17.105000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 74.200000 17.105000 74.520000 ;
      LAYER met4 ;
        RECT 16.785000 74.200000 17.105000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 74.605000 17.105000 74.925000 ;
      LAYER met4 ;
        RECT 16.785000 74.605000 17.105000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 75.010000 17.105000 75.330000 ;
      LAYER met4 ;
        RECT 16.785000 75.010000 17.105000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 75.415000 17.105000 75.735000 ;
      LAYER met4 ;
        RECT 16.785000 75.415000 17.105000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 75.820000 17.105000 76.140000 ;
      LAYER met4 ;
        RECT 16.785000 75.820000 17.105000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 76.225000 17.105000 76.545000 ;
      LAYER met4 ;
        RECT 16.785000 76.225000 17.105000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 76.630000 17.105000 76.950000 ;
      LAYER met4 ;
        RECT 16.785000 76.630000 17.105000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 77.035000 17.105000 77.355000 ;
      LAYER met4 ;
        RECT 16.785000 77.035000 17.105000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 77.440000 17.105000 77.760000 ;
      LAYER met4 ;
        RECT 16.785000 77.440000 17.105000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 77.845000 17.105000 78.165000 ;
      LAYER met4 ;
        RECT 16.785000 77.845000 17.105000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 78.250000 17.105000 78.570000 ;
      LAYER met4 ;
        RECT 16.785000 78.250000 17.105000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 78.655000 17.105000 78.975000 ;
      LAYER met4 ;
        RECT 16.785000 78.655000 17.105000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 79.060000 17.105000 79.380000 ;
      LAYER met4 ;
        RECT 16.785000 79.060000 17.105000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 79.465000 17.105000 79.785000 ;
      LAYER met4 ;
        RECT 16.785000 79.465000 17.105000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 79.870000 17.105000 80.190000 ;
      LAYER met4 ;
        RECT 16.785000 79.870000 17.105000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 80.275000 17.105000 80.595000 ;
      LAYER met4 ;
        RECT 16.785000 80.275000 17.105000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 80.680000 17.105000 81.000000 ;
      LAYER met4 ;
        RECT 16.785000 80.680000 17.105000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 81.085000 17.105000 81.405000 ;
      LAYER met4 ;
        RECT 16.785000 81.085000 17.105000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 81.490000 17.105000 81.810000 ;
      LAYER met4 ;
        RECT 16.785000 81.490000 17.105000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 81.895000 17.105000 82.215000 ;
      LAYER met4 ;
        RECT 16.785000 81.895000 17.105000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785000 82.300000 17.105000 82.620000 ;
      LAYER met4 ;
        RECT 16.785000 82.300000 17.105000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830000 17.800000 17.150000 18.120000 ;
      LAYER met4 ;
        RECT 16.830000 17.800000 17.150000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830000 18.230000 17.150000 18.550000 ;
      LAYER met4 ;
        RECT 16.830000 18.230000 17.150000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830000 18.660000 17.150000 18.980000 ;
      LAYER met4 ;
        RECT 16.830000 18.660000 17.150000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830000 19.090000 17.150000 19.410000 ;
      LAYER met4 ;
        RECT 16.830000 19.090000 17.150000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830000 19.520000 17.150000 19.840000 ;
      LAYER met4 ;
        RECT 16.830000 19.520000 17.150000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830000 19.950000 17.150000 20.270000 ;
      LAYER met4 ;
        RECT 16.830000 19.950000 17.150000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830000 20.380000 17.150000 20.700000 ;
      LAYER met4 ;
        RECT 16.830000 20.380000 17.150000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830000 20.810000 17.150000 21.130000 ;
      LAYER met4 ;
        RECT 16.830000 20.810000 17.150000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830000 21.240000 17.150000 21.560000 ;
      LAYER met4 ;
        RECT 16.830000 21.240000 17.150000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830000 21.670000 17.150000 21.990000 ;
      LAYER met4 ;
        RECT 16.830000 21.670000 17.150000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830000 22.100000 17.150000 22.420000 ;
      LAYER met4 ;
        RECT 16.830000 22.100000 17.150000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865000 82.995000 17.185000 83.315000 ;
      LAYER met4 ;
        RECT 16.865000 82.995000 17.185000 83.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865000 83.395000 17.185000 83.715000 ;
      LAYER met4 ;
        RECT 16.865000 83.395000 17.185000 83.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865000 83.795000 17.185000 84.115000 ;
      LAYER met4 ;
        RECT 16.865000 83.795000 17.185000 84.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865000 84.195000 17.185000 84.515000 ;
      LAYER met4 ;
        RECT 16.865000 84.195000 17.185000 84.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865000 84.595000 17.185000 84.915000 ;
      LAYER met4 ;
        RECT 16.865000 84.595000 17.185000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865000 84.995000 17.185000 85.315000 ;
      LAYER met4 ;
        RECT 16.865000 84.995000 17.185000 85.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865000 85.395000 17.185000 85.715000 ;
      LAYER met4 ;
        RECT 16.865000 85.395000 17.185000 85.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865000 85.795000 17.185000 86.115000 ;
      LAYER met4 ;
        RECT 16.865000 85.795000 17.185000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865000 86.195000 17.185000 86.515000 ;
      LAYER met4 ;
        RECT 16.865000 86.195000 17.185000 86.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865000 86.600000 17.185000 86.920000 ;
      LAYER met4 ;
        RECT 16.865000 86.600000 17.185000 86.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865000 87.005000 17.185000 87.325000 ;
      LAYER met4 ;
        RECT 16.865000 87.005000 17.185000 87.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865000 87.410000 17.185000 87.730000 ;
      LAYER met4 ;
        RECT 16.865000 87.410000 17.185000 87.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865000 87.815000 17.185000 88.135000 ;
      LAYER met4 ;
        RECT 16.865000 87.815000 17.185000 88.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 68.065000 17.505000 68.385000 ;
      LAYER met4 ;
        RECT 17.185000 68.065000 17.505000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 68.475000 17.505000 68.795000 ;
      LAYER met4 ;
        RECT 17.185000 68.475000 17.505000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 68.885000 17.505000 69.205000 ;
      LAYER met4 ;
        RECT 17.185000 68.885000 17.505000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 69.295000 17.505000 69.615000 ;
      LAYER met4 ;
        RECT 17.185000 69.295000 17.505000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 69.705000 17.505000 70.025000 ;
      LAYER met4 ;
        RECT 17.185000 69.705000 17.505000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 70.115000 17.505000 70.435000 ;
      LAYER met4 ;
        RECT 17.185000 70.115000 17.505000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 70.525000 17.505000 70.845000 ;
      LAYER met4 ;
        RECT 17.185000 70.525000 17.505000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 70.935000 17.505000 71.255000 ;
      LAYER met4 ;
        RECT 17.185000 70.935000 17.505000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 71.345000 17.505000 71.665000 ;
      LAYER met4 ;
        RECT 17.185000 71.345000 17.505000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 71.755000 17.505000 72.075000 ;
      LAYER met4 ;
        RECT 17.185000 71.755000 17.505000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 72.165000 17.505000 72.485000 ;
      LAYER met4 ;
        RECT 17.185000 72.165000 17.505000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 72.575000 17.505000 72.895000 ;
      LAYER met4 ;
        RECT 17.185000 72.575000 17.505000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 72.985000 17.505000 73.305000 ;
      LAYER met4 ;
        RECT 17.185000 72.985000 17.505000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 73.390000 17.505000 73.710000 ;
      LAYER met4 ;
        RECT 17.185000 73.390000 17.505000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 73.795000 17.505000 74.115000 ;
      LAYER met4 ;
        RECT 17.185000 73.795000 17.505000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 74.200000 17.505000 74.520000 ;
      LAYER met4 ;
        RECT 17.185000 74.200000 17.505000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 74.605000 17.505000 74.925000 ;
      LAYER met4 ;
        RECT 17.185000 74.605000 17.505000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 75.010000 17.505000 75.330000 ;
      LAYER met4 ;
        RECT 17.185000 75.010000 17.505000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 75.415000 17.505000 75.735000 ;
      LAYER met4 ;
        RECT 17.185000 75.415000 17.505000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 75.820000 17.505000 76.140000 ;
      LAYER met4 ;
        RECT 17.185000 75.820000 17.505000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 76.225000 17.505000 76.545000 ;
      LAYER met4 ;
        RECT 17.185000 76.225000 17.505000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 76.630000 17.505000 76.950000 ;
      LAYER met4 ;
        RECT 17.185000 76.630000 17.505000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 77.035000 17.505000 77.355000 ;
      LAYER met4 ;
        RECT 17.185000 77.035000 17.505000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 77.440000 17.505000 77.760000 ;
      LAYER met4 ;
        RECT 17.185000 77.440000 17.505000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 77.845000 17.505000 78.165000 ;
      LAYER met4 ;
        RECT 17.185000 77.845000 17.505000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 78.250000 17.505000 78.570000 ;
      LAYER met4 ;
        RECT 17.185000 78.250000 17.505000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 78.655000 17.505000 78.975000 ;
      LAYER met4 ;
        RECT 17.185000 78.655000 17.505000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 79.060000 17.505000 79.380000 ;
      LAYER met4 ;
        RECT 17.185000 79.060000 17.505000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 79.465000 17.505000 79.785000 ;
      LAYER met4 ;
        RECT 17.185000 79.465000 17.505000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 79.870000 17.505000 80.190000 ;
      LAYER met4 ;
        RECT 17.185000 79.870000 17.505000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 80.275000 17.505000 80.595000 ;
      LAYER met4 ;
        RECT 17.185000 80.275000 17.505000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 80.680000 17.505000 81.000000 ;
      LAYER met4 ;
        RECT 17.185000 80.680000 17.505000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 81.085000 17.505000 81.405000 ;
      LAYER met4 ;
        RECT 17.185000 81.085000 17.505000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 81.490000 17.505000 81.810000 ;
      LAYER met4 ;
        RECT 17.185000 81.490000 17.505000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 81.895000 17.505000 82.215000 ;
      LAYER met4 ;
        RECT 17.185000 81.895000 17.505000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185000 82.300000 17.505000 82.620000 ;
      LAYER met4 ;
        RECT 17.185000 82.300000 17.505000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200000 88.370000 17.520000 88.690000 ;
      LAYER met4 ;
        RECT 17.200000 88.370000 17.520000 88.690000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200000 88.785000 17.520000 89.105000 ;
      LAYER met4 ;
        RECT 17.200000 88.785000 17.520000 89.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200000 89.205000 17.520000 89.525000 ;
      LAYER met4 ;
        RECT 17.200000 89.205000 17.520000 89.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235000 17.800000 17.555000 18.120000 ;
      LAYER met4 ;
        RECT 17.235000 17.800000 17.555000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235000 18.230000 17.555000 18.550000 ;
      LAYER met4 ;
        RECT 17.235000 18.230000 17.555000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235000 18.660000 17.555000 18.980000 ;
      LAYER met4 ;
        RECT 17.235000 18.660000 17.555000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235000 19.090000 17.555000 19.410000 ;
      LAYER met4 ;
        RECT 17.235000 19.090000 17.555000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235000 19.520000 17.555000 19.840000 ;
      LAYER met4 ;
        RECT 17.235000 19.520000 17.555000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235000 19.950000 17.555000 20.270000 ;
      LAYER met4 ;
        RECT 17.235000 19.950000 17.555000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235000 20.380000 17.555000 20.700000 ;
      LAYER met4 ;
        RECT 17.235000 20.380000 17.555000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235000 20.810000 17.555000 21.130000 ;
      LAYER met4 ;
        RECT 17.235000 20.810000 17.555000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235000 21.240000 17.555000 21.560000 ;
      LAYER met4 ;
        RECT 17.235000 21.240000 17.555000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235000 21.670000 17.555000 21.990000 ;
      LAYER met4 ;
        RECT 17.235000 21.670000 17.555000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235000 22.100000 17.555000 22.420000 ;
      LAYER met4 ;
        RECT 17.235000 22.100000 17.555000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275000 82.995000 17.595000 83.315000 ;
      LAYER met4 ;
        RECT 17.275000 82.995000 17.595000 83.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275000 83.395000 17.595000 83.715000 ;
      LAYER met4 ;
        RECT 17.275000 83.395000 17.595000 83.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275000 83.795000 17.595000 84.115000 ;
      LAYER met4 ;
        RECT 17.275000 83.795000 17.595000 84.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275000 84.195000 17.595000 84.515000 ;
      LAYER met4 ;
        RECT 17.275000 84.195000 17.595000 84.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275000 84.595000 17.595000 84.915000 ;
      LAYER met4 ;
        RECT 17.275000 84.595000 17.595000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275000 84.995000 17.595000 85.315000 ;
      LAYER met4 ;
        RECT 17.275000 84.995000 17.595000 85.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275000 85.395000 17.595000 85.715000 ;
      LAYER met4 ;
        RECT 17.275000 85.395000 17.595000 85.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275000 85.795000 17.595000 86.115000 ;
      LAYER met4 ;
        RECT 17.275000 85.795000 17.595000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275000 86.195000 17.595000 86.515000 ;
      LAYER met4 ;
        RECT 17.275000 86.195000 17.595000 86.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275000 86.600000 17.595000 86.920000 ;
      LAYER met4 ;
        RECT 17.275000 86.600000 17.595000 86.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275000 87.005000 17.595000 87.325000 ;
      LAYER met4 ;
        RECT 17.275000 87.005000 17.595000 87.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275000 87.410000 17.595000 87.730000 ;
      LAYER met4 ;
        RECT 17.275000 87.410000 17.595000 87.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275000 87.815000 17.595000 88.135000 ;
      LAYER met4 ;
        RECT 17.275000 87.815000 17.595000 88.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 68.065000 17.905000 68.385000 ;
      LAYER met4 ;
        RECT 17.585000 68.065000 17.905000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 68.475000 17.905000 68.795000 ;
      LAYER met4 ;
        RECT 17.585000 68.475000 17.905000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 68.885000 17.905000 69.205000 ;
      LAYER met4 ;
        RECT 17.585000 68.885000 17.905000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 69.295000 17.905000 69.615000 ;
      LAYER met4 ;
        RECT 17.585000 69.295000 17.905000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 69.705000 17.905000 70.025000 ;
      LAYER met4 ;
        RECT 17.585000 69.705000 17.905000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 70.115000 17.905000 70.435000 ;
      LAYER met4 ;
        RECT 17.585000 70.115000 17.905000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 70.525000 17.905000 70.845000 ;
      LAYER met4 ;
        RECT 17.585000 70.525000 17.905000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 70.935000 17.905000 71.255000 ;
      LAYER met4 ;
        RECT 17.585000 70.935000 17.905000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 71.345000 17.905000 71.665000 ;
      LAYER met4 ;
        RECT 17.585000 71.345000 17.905000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 71.755000 17.905000 72.075000 ;
      LAYER met4 ;
        RECT 17.585000 71.755000 17.905000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 72.165000 17.905000 72.485000 ;
      LAYER met4 ;
        RECT 17.585000 72.165000 17.905000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 72.575000 17.905000 72.895000 ;
      LAYER met4 ;
        RECT 17.585000 72.575000 17.905000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 72.985000 17.905000 73.305000 ;
      LAYER met4 ;
        RECT 17.585000 72.985000 17.905000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 73.390000 17.905000 73.710000 ;
      LAYER met4 ;
        RECT 17.585000 73.390000 17.905000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 73.795000 17.905000 74.115000 ;
      LAYER met4 ;
        RECT 17.585000 73.795000 17.905000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 74.200000 17.905000 74.520000 ;
      LAYER met4 ;
        RECT 17.585000 74.200000 17.905000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 74.605000 17.905000 74.925000 ;
      LAYER met4 ;
        RECT 17.585000 74.605000 17.905000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 75.010000 17.905000 75.330000 ;
      LAYER met4 ;
        RECT 17.585000 75.010000 17.905000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 75.415000 17.905000 75.735000 ;
      LAYER met4 ;
        RECT 17.585000 75.415000 17.905000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 75.820000 17.905000 76.140000 ;
      LAYER met4 ;
        RECT 17.585000 75.820000 17.905000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 76.225000 17.905000 76.545000 ;
      LAYER met4 ;
        RECT 17.585000 76.225000 17.905000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 76.630000 17.905000 76.950000 ;
      LAYER met4 ;
        RECT 17.585000 76.630000 17.905000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 77.035000 17.905000 77.355000 ;
      LAYER met4 ;
        RECT 17.585000 77.035000 17.905000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 77.440000 17.905000 77.760000 ;
      LAYER met4 ;
        RECT 17.585000 77.440000 17.905000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 77.845000 17.905000 78.165000 ;
      LAYER met4 ;
        RECT 17.585000 77.845000 17.905000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 78.250000 17.905000 78.570000 ;
      LAYER met4 ;
        RECT 17.585000 78.250000 17.905000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 78.655000 17.905000 78.975000 ;
      LAYER met4 ;
        RECT 17.585000 78.655000 17.905000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 79.060000 17.905000 79.380000 ;
      LAYER met4 ;
        RECT 17.585000 79.060000 17.905000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 79.465000 17.905000 79.785000 ;
      LAYER met4 ;
        RECT 17.585000 79.465000 17.905000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 79.870000 17.905000 80.190000 ;
      LAYER met4 ;
        RECT 17.585000 79.870000 17.905000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 80.275000 17.905000 80.595000 ;
      LAYER met4 ;
        RECT 17.585000 80.275000 17.905000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 80.680000 17.905000 81.000000 ;
      LAYER met4 ;
        RECT 17.585000 80.680000 17.905000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 81.085000 17.905000 81.405000 ;
      LAYER met4 ;
        RECT 17.585000 81.085000 17.905000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 81.490000 17.905000 81.810000 ;
      LAYER met4 ;
        RECT 17.585000 81.490000 17.905000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 81.895000 17.905000 82.215000 ;
      LAYER met4 ;
        RECT 17.585000 81.895000 17.905000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585000 82.300000 17.905000 82.620000 ;
      LAYER met4 ;
        RECT 17.585000 82.300000 17.905000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640000 17.800000 17.960000 18.120000 ;
      LAYER met4 ;
        RECT 17.640000 17.800000 17.960000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640000 18.230000 17.960000 18.550000 ;
      LAYER met4 ;
        RECT 17.640000 18.230000 17.960000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640000 18.660000 17.960000 18.980000 ;
      LAYER met4 ;
        RECT 17.640000 18.660000 17.960000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640000 19.090000 17.960000 19.410000 ;
      LAYER met4 ;
        RECT 17.640000 19.090000 17.960000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640000 19.520000 17.960000 19.840000 ;
      LAYER met4 ;
        RECT 17.640000 19.520000 17.960000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640000 19.950000 17.960000 20.270000 ;
      LAYER met4 ;
        RECT 17.640000 19.950000 17.960000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640000 20.380000 17.960000 20.700000 ;
      LAYER met4 ;
        RECT 17.640000 20.380000 17.960000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640000 20.810000 17.960000 21.130000 ;
      LAYER met4 ;
        RECT 17.640000 20.810000 17.960000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640000 21.240000 17.960000 21.560000 ;
      LAYER met4 ;
        RECT 17.640000 21.240000 17.960000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640000 21.670000 17.960000 21.990000 ;
      LAYER met4 ;
        RECT 17.640000 21.670000 17.960000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640000 22.100000 17.960000 22.420000 ;
      LAYER met4 ;
        RECT 17.640000 22.100000 17.960000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685000 82.995000 18.005000 83.315000 ;
      LAYER met4 ;
        RECT 17.685000 82.995000 18.005000 83.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685000 83.395000 18.005000 83.715000 ;
      LAYER met4 ;
        RECT 17.685000 83.395000 18.005000 83.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685000 83.795000 18.005000 84.115000 ;
      LAYER met4 ;
        RECT 17.685000 83.795000 18.005000 84.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685000 84.195000 18.005000 84.515000 ;
      LAYER met4 ;
        RECT 17.685000 84.195000 18.005000 84.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685000 84.595000 18.005000 84.915000 ;
      LAYER met4 ;
        RECT 17.685000 84.595000 18.005000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685000 84.995000 18.005000 85.315000 ;
      LAYER met4 ;
        RECT 17.685000 84.995000 18.005000 85.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685000 85.395000 18.005000 85.715000 ;
      LAYER met4 ;
        RECT 17.685000 85.395000 18.005000 85.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685000 85.795000 18.005000 86.115000 ;
      LAYER met4 ;
        RECT 17.685000 85.795000 18.005000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685000 86.195000 18.005000 86.515000 ;
      LAYER met4 ;
        RECT 17.685000 86.195000 18.005000 86.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685000 86.600000 18.005000 86.920000 ;
      LAYER met4 ;
        RECT 17.685000 86.600000 18.005000 86.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685000 87.005000 18.005000 87.325000 ;
      LAYER met4 ;
        RECT 17.685000 87.005000 18.005000 87.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685000 87.410000 18.005000 87.730000 ;
      LAYER met4 ;
        RECT 17.685000 87.410000 18.005000 87.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685000 87.815000 18.005000 88.135000 ;
      LAYER met4 ;
        RECT 17.685000 87.815000 18.005000 88.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 68.065000 18.305000 68.385000 ;
      LAYER met4 ;
        RECT 17.985000 68.065000 18.305000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 68.475000 18.305000 68.795000 ;
      LAYER met4 ;
        RECT 17.985000 68.475000 18.305000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 68.885000 18.305000 69.205000 ;
      LAYER met4 ;
        RECT 17.985000 68.885000 18.305000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 69.295000 18.305000 69.615000 ;
      LAYER met4 ;
        RECT 17.985000 69.295000 18.305000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 69.705000 18.305000 70.025000 ;
      LAYER met4 ;
        RECT 17.985000 69.705000 18.305000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 70.115000 18.305000 70.435000 ;
      LAYER met4 ;
        RECT 17.985000 70.115000 18.305000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 70.525000 18.305000 70.845000 ;
      LAYER met4 ;
        RECT 17.985000 70.525000 18.305000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 70.935000 18.305000 71.255000 ;
      LAYER met4 ;
        RECT 17.985000 70.935000 18.305000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 71.345000 18.305000 71.665000 ;
      LAYER met4 ;
        RECT 17.985000 71.345000 18.305000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 71.755000 18.305000 72.075000 ;
      LAYER met4 ;
        RECT 17.985000 71.755000 18.305000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 72.165000 18.305000 72.485000 ;
      LAYER met4 ;
        RECT 17.985000 72.165000 18.305000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 72.575000 18.305000 72.895000 ;
      LAYER met4 ;
        RECT 17.985000 72.575000 18.305000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 72.985000 18.305000 73.305000 ;
      LAYER met4 ;
        RECT 17.985000 72.985000 18.305000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 73.390000 18.305000 73.710000 ;
      LAYER met4 ;
        RECT 17.985000 73.390000 18.305000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 73.795000 18.305000 74.115000 ;
      LAYER met4 ;
        RECT 17.985000 73.795000 18.305000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 74.200000 18.305000 74.520000 ;
      LAYER met4 ;
        RECT 17.985000 74.200000 18.305000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 74.605000 18.305000 74.925000 ;
      LAYER met4 ;
        RECT 17.985000 74.605000 18.305000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 75.010000 18.305000 75.330000 ;
      LAYER met4 ;
        RECT 17.985000 75.010000 18.305000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 75.415000 18.305000 75.735000 ;
      LAYER met4 ;
        RECT 17.985000 75.415000 18.305000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 75.820000 18.305000 76.140000 ;
      LAYER met4 ;
        RECT 17.985000 75.820000 18.305000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 76.225000 18.305000 76.545000 ;
      LAYER met4 ;
        RECT 17.985000 76.225000 18.305000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 76.630000 18.305000 76.950000 ;
      LAYER met4 ;
        RECT 17.985000 76.630000 18.305000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 77.035000 18.305000 77.355000 ;
      LAYER met4 ;
        RECT 17.985000 77.035000 18.305000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 77.440000 18.305000 77.760000 ;
      LAYER met4 ;
        RECT 17.985000 77.440000 18.305000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 77.845000 18.305000 78.165000 ;
      LAYER met4 ;
        RECT 17.985000 77.845000 18.305000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 78.250000 18.305000 78.570000 ;
      LAYER met4 ;
        RECT 17.985000 78.250000 18.305000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 78.655000 18.305000 78.975000 ;
      LAYER met4 ;
        RECT 17.985000 78.655000 18.305000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 79.060000 18.305000 79.380000 ;
      LAYER met4 ;
        RECT 17.985000 79.060000 18.305000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 79.465000 18.305000 79.785000 ;
      LAYER met4 ;
        RECT 17.985000 79.465000 18.305000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 79.870000 18.305000 80.190000 ;
      LAYER met4 ;
        RECT 17.985000 79.870000 18.305000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 80.275000 18.305000 80.595000 ;
      LAYER met4 ;
        RECT 17.985000 80.275000 18.305000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 80.680000 18.305000 81.000000 ;
      LAYER met4 ;
        RECT 17.985000 80.680000 18.305000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 81.085000 18.305000 81.405000 ;
      LAYER met4 ;
        RECT 17.985000 81.085000 18.305000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 81.490000 18.305000 81.810000 ;
      LAYER met4 ;
        RECT 17.985000 81.490000 18.305000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 81.895000 18.305000 82.215000 ;
      LAYER met4 ;
        RECT 17.985000 81.895000 18.305000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985000 82.300000 18.305000 82.620000 ;
      LAYER met4 ;
        RECT 17.985000 82.300000 18.305000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 17.800000 18.365000 18.120000 ;
      LAYER met4 ;
        RECT 18.045000 17.800000 18.365000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 18.230000 18.365000 18.550000 ;
      LAYER met4 ;
        RECT 18.045000 18.230000 18.365000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 18.660000 18.365000 18.980000 ;
      LAYER met4 ;
        RECT 18.045000 18.660000 18.365000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 19.090000 18.365000 19.410000 ;
      LAYER met4 ;
        RECT 18.045000 19.090000 18.365000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 19.520000 18.365000 19.840000 ;
      LAYER met4 ;
        RECT 18.045000 19.520000 18.365000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 19.950000 18.365000 20.270000 ;
      LAYER met4 ;
        RECT 18.045000 19.950000 18.365000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 20.380000 18.365000 20.700000 ;
      LAYER met4 ;
        RECT 18.045000 20.380000 18.365000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 20.810000 18.365000 21.130000 ;
      LAYER met4 ;
        RECT 18.045000 20.810000 18.365000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 21.240000 18.365000 21.560000 ;
      LAYER met4 ;
        RECT 18.045000 21.240000 18.365000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 21.670000 18.365000 21.990000 ;
      LAYER met4 ;
        RECT 18.045000 21.670000 18.365000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 22.100000 18.365000 22.420000 ;
      LAYER met4 ;
        RECT 18.045000 22.100000 18.365000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095000 82.995000 18.415000 83.315000 ;
      LAYER met4 ;
        RECT 18.095000 82.995000 18.415000 83.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095000 83.395000 18.415000 83.715000 ;
      LAYER met4 ;
        RECT 18.095000 83.395000 18.415000 83.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095000 83.795000 18.415000 84.115000 ;
      LAYER met4 ;
        RECT 18.095000 83.795000 18.415000 84.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095000 84.195000 18.415000 84.515000 ;
      LAYER met4 ;
        RECT 18.095000 84.195000 18.415000 84.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095000 84.595000 18.415000 84.915000 ;
      LAYER met4 ;
        RECT 18.095000 84.595000 18.415000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095000 84.995000 18.415000 85.315000 ;
      LAYER met4 ;
        RECT 18.095000 84.995000 18.415000 85.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095000 85.395000 18.415000 85.715000 ;
      LAYER met4 ;
        RECT 18.095000 85.395000 18.415000 85.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095000 85.795000 18.415000 86.115000 ;
      LAYER met4 ;
        RECT 18.095000 85.795000 18.415000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095000 86.195000 18.415000 86.515000 ;
      LAYER met4 ;
        RECT 18.095000 86.195000 18.415000 86.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095000 86.600000 18.415000 86.920000 ;
      LAYER met4 ;
        RECT 18.095000 86.600000 18.415000 86.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095000 87.005000 18.415000 87.325000 ;
      LAYER met4 ;
        RECT 18.095000 87.005000 18.415000 87.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095000 87.410000 18.415000 87.730000 ;
      LAYER met4 ;
        RECT 18.095000 87.410000 18.415000 87.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095000 87.815000 18.415000 88.135000 ;
      LAYER met4 ;
        RECT 18.095000 87.815000 18.415000 88.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 68.065000 18.705000 68.385000 ;
      LAYER met4 ;
        RECT 18.385000 68.065000 18.705000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 68.475000 18.705000 68.795000 ;
      LAYER met4 ;
        RECT 18.385000 68.475000 18.705000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 68.885000 18.705000 69.205000 ;
      LAYER met4 ;
        RECT 18.385000 68.885000 18.705000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 69.295000 18.705000 69.615000 ;
      LAYER met4 ;
        RECT 18.385000 69.295000 18.705000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 69.705000 18.705000 70.025000 ;
      LAYER met4 ;
        RECT 18.385000 69.705000 18.705000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 70.115000 18.705000 70.435000 ;
      LAYER met4 ;
        RECT 18.385000 70.115000 18.705000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 70.525000 18.705000 70.845000 ;
      LAYER met4 ;
        RECT 18.385000 70.525000 18.705000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 70.935000 18.705000 71.255000 ;
      LAYER met4 ;
        RECT 18.385000 70.935000 18.705000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 71.345000 18.705000 71.665000 ;
      LAYER met4 ;
        RECT 18.385000 71.345000 18.705000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 71.755000 18.705000 72.075000 ;
      LAYER met4 ;
        RECT 18.385000 71.755000 18.705000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 72.165000 18.705000 72.485000 ;
      LAYER met4 ;
        RECT 18.385000 72.165000 18.705000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 72.575000 18.705000 72.895000 ;
      LAYER met4 ;
        RECT 18.385000 72.575000 18.705000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 72.985000 18.705000 73.305000 ;
      LAYER met4 ;
        RECT 18.385000 72.985000 18.705000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 73.390000 18.705000 73.710000 ;
      LAYER met4 ;
        RECT 18.385000 73.390000 18.705000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 73.795000 18.705000 74.115000 ;
      LAYER met4 ;
        RECT 18.385000 73.795000 18.705000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 74.200000 18.705000 74.520000 ;
      LAYER met4 ;
        RECT 18.385000 74.200000 18.705000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 74.605000 18.705000 74.925000 ;
      LAYER met4 ;
        RECT 18.385000 74.605000 18.705000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 75.010000 18.705000 75.330000 ;
      LAYER met4 ;
        RECT 18.385000 75.010000 18.705000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 75.415000 18.705000 75.735000 ;
      LAYER met4 ;
        RECT 18.385000 75.415000 18.705000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 75.820000 18.705000 76.140000 ;
      LAYER met4 ;
        RECT 18.385000 75.820000 18.705000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 76.225000 18.705000 76.545000 ;
      LAYER met4 ;
        RECT 18.385000 76.225000 18.705000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 76.630000 18.705000 76.950000 ;
      LAYER met4 ;
        RECT 18.385000 76.630000 18.705000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 77.035000 18.705000 77.355000 ;
      LAYER met4 ;
        RECT 18.385000 77.035000 18.705000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 77.440000 18.705000 77.760000 ;
      LAYER met4 ;
        RECT 18.385000 77.440000 18.705000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 77.845000 18.705000 78.165000 ;
      LAYER met4 ;
        RECT 18.385000 77.845000 18.705000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 78.250000 18.705000 78.570000 ;
      LAYER met4 ;
        RECT 18.385000 78.250000 18.705000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 78.655000 18.705000 78.975000 ;
      LAYER met4 ;
        RECT 18.385000 78.655000 18.705000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 79.060000 18.705000 79.380000 ;
      LAYER met4 ;
        RECT 18.385000 79.060000 18.705000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 79.465000 18.705000 79.785000 ;
      LAYER met4 ;
        RECT 18.385000 79.465000 18.705000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 79.870000 18.705000 80.190000 ;
      LAYER met4 ;
        RECT 18.385000 79.870000 18.705000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 80.275000 18.705000 80.595000 ;
      LAYER met4 ;
        RECT 18.385000 80.275000 18.705000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 80.680000 18.705000 81.000000 ;
      LAYER met4 ;
        RECT 18.385000 80.680000 18.705000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 81.085000 18.705000 81.405000 ;
      LAYER met4 ;
        RECT 18.385000 81.085000 18.705000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 81.490000 18.705000 81.810000 ;
      LAYER met4 ;
        RECT 18.385000 81.490000 18.705000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 81.895000 18.705000 82.215000 ;
      LAYER met4 ;
        RECT 18.385000 81.895000 18.705000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385000 82.300000 18.705000 82.620000 ;
      LAYER met4 ;
        RECT 18.385000 82.300000 18.705000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450000 17.800000 18.770000 18.120000 ;
      LAYER met4 ;
        RECT 18.450000 17.800000 18.770000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450000 18.230000 18.770000 18.550000 ;
      LAYER met4 ;
        RECT 18.450000 18.230000 18.770000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450000 18.660000 18.770000 18.980000 ;
      LAYER met4 ;
        RECT 18.450000 18.660000 18.770000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450000 19.090000 18.770000 19.410000 ;
      LAYER met4 ;
        RECT 18.450000 19.090000 18.770000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450000 19.520000 18.770000 19.840000 ;
      LAYER met4 ;
        RECT 18.450000 19.520000 18.770000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450000 19.950000 18.770000 20.270000 ;
      LAYER met4 ;
        RECT 18.450000 19.950000 18.770000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450000 20.380000 18.770000 20.700000 ;
      LAYER met4 ;
        RECT 18.450000 20.380000 18.770000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450000 20.810000 18.770000 21.130000 ;
      LAYER met4 ;
        RECT 18.450000 20.810000 18.770000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450000 21.240000 18.770000 21.560000 ;
      LAYER met4 ;
        RECT 18.450000 21.240000 18.770000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450000 21.670000 18.770000 21.990000 ;
      LAYER met4 ;
        RECT 18.450000 21.670000 18.770000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450000 22.100000 18.770000 22.420000 ;
      LAYER met4 ;
        RECT 18.450000 22.100000 18.770000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505000 82.995000 18.825000 83.315000 ;
      LAYER met4 ;
        RECT 18.505000 82.995000 18.825000 83.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505000 83.395000 18.825000 83.715000 ;
      LAYER met4 ;
        RECT 18.505000 83.395000 18.825000 83.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505000 83.795000 18.825000 84.115000 ;
      LAYER met4 ;
        RECT 18.505000 83.795000 18.825000 84.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505000 84.195000 18.825000 84.515000 ;
      LAYER met4 ;
        RECT 18.505000 84.195000 18.825000 84.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505000 84.595000 18.825000 84.915000 ;
      LAYER met4 ;
        RECT 18.505000 84.595000 18.825000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505000 84.995000 18.825000 85.315000 ;
      LAYER met4 ;
        RECT 18.505000 84.995000 18.825000 85.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505000 85.395000 18.825000 85.715000 ;
      LAYER met4 ;
        RECT 18.505000 85.395000 18.825000 85.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505000 85.795000 18.825000 86.115000 ;
      LAYER met4 ;
        RECT 18.505000 85.795000 18.825000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505000 86.195000 18.825000 86.515000 ;
      LAYER met4 ;
        RECT 18.505000 86.195000 18.825000 86.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505000 86.600000 18.825000 86.920000 ;
      LAYER met4 ;
        RECT 18.505000 86.600000 18.825000 86.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505000 87.005000 18.825000 87.325000 ;
      LAYER met4 ;
        RECT 18.505000 87.005000 18.825000 87.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505000 87.410000 18.825000 87.730000 ;
      LAYER met4 ;
        RECT 18.505000 87.410000 18.825000 87.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505000 87.815000 18.825000 88.135000 ;
      LAYER met4 ;
        RECT 18.505000 87.815000 18.825000 88.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 68.065000 19.105000 68.385000 ;
      LAYER met4 ;
        RECT 18.785000 68.065000 19.105000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 68.475000 19.105000 68.795000 ;
      LAYER met4 ;
        RECT 18.785000 68.475000 19.105000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 68.885000 19.105000 69.205000 ;
      LAYER met4 ;
        RECT 18.785000 68.885000 19.105000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 69.295000 19.105000 69.615000 ;
      LAYER met4 ;
        RECT 18.785000 69.295000 19.105000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 69.705000 19.105000 70.025000 ;
      LAYER met4 ;
        RECT 18.785000 69.705000 19.105000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 70.115000 19.105000 70.435000 ;
      LAYER met4 ;
        RECT 18.785000 70.115000 19.105000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 70.525000 19.105000 70.845000 ;
      LAYER met4 ;
        RECT 18.785000 70.525000 19.105000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 70.935000 19.105000 71.255000 ;
      LAYER met4 ;
        RECT 18.785000 70.935000 19.105000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 71.345000 19.105000 71.665000 ;
      LAYER met4 ;
        RECT 18.785000 71.345000 19.105000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 71.755000 19.105000 72.075000 ;
      LAYER met4 ;
        RECT 18.785000 71.755000 19.105000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 72.165000 19.105000 72.485000 ;
      LAYER met4 ;
        RECT 18.785000 72.165000 19.105000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 72.575000 19.105000 72.895000 ;
      LAYER met4 ;
        RECT 18.785000 72.575000 19.105000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 72.985000 19.105000 73.305000 ;
      LAYER met4 ;
        RECT 18.785000 72.985000 19.105000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 73.390000 19.105000 73.710000 ;
      LAYER met4 ;
        RECT 18.785000 73.390000 19.105000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 73.795000 19.105000 74.115000 ;
      LAYER met4 ;
        RECT 18.785000 73.795000 19.105000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 74.200000 19.105000 74.520000 ;
      LAYER met4 ;
        RECT 18.785000 74.200000 19.105000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 74.605000 19.105000 74.925000 ;
      LAYER met4 ;
        RECT 18.785000 74.605000 19.105000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 75.010000 19.105000 75.330000 ;
      LAYER met4 ;
        RECT 18.785000 75.010000 19.105000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 75.415000 19.105000 75.735000 ;
      LAYER met4 ;
        RECT 18.785000 75.415000 19.105000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 75.820000 19.105000 76.140000 ;
      LAYER met4 ;
        RECT 18.785000 75.820000 19.105000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 76.225000 19.105000 76.545000 ;
      LAYER met4 ;
        RECT 18.785000 76.225000 19.105000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 76.630000 19.105000 76.950000 ;
      LAYER met4 ;
        RECT 18.785000 76.630000 19.105000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 77.035000 19.105000 77.355000 ;
      LAYER met4 ;
        RECT 18.785000 77.035000 19.105000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 77.440000 19.105000 77.760000 ;
      LAYER met4 ;
        RECT 18.785000 77.440000 19.105000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 77.845000 19.105000 78.165000 ;
      LAYER met4 ;
        RECT 18.785000 77.845000 19.105000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 78.250000 19.105000 78.570000 ;
      LAYER met4 ;
        RECT 18.785000 78.250000 19.105000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 78.655000 19.105000 78.975000 ;
      LAYER met4 ;
        RECT 18.785000 78.655000 19.105000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 79.060000 19.105000 79.380000 ;
      LAYER met4 ;
        RECT 18.785000 79.060000 19.105000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 79.465000 19.105000 79.785000 ;
      LAYER met4 ;
        RECT 18.785000 79.465000 19.105000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 79.870000 19.105000 80.190000 ;
      LAYER met4 ;
        RECT 18.785000 79.870000 19.105000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 80.275000 19.105000 80.595000 ;
      LAYER met4 ;
        RECT 18.785000 80.275000 19.105000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 80.680000 19.105000 81.000000 ;
      LAYER met4 ;
        RECT 18.785000 80.680000 19.105000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 81.085000 19.105000 81.405000 ;
      LAYER met4 ;
        RECT 18.785000 81.085000 19.105000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 81.490000 19.105000 81.810000 ;
      LAYER met4 ;
        RECT 18.785000 81.490000 19.105000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 81.895000 19.105000 82.215000 ;
      LAYER met4 ;
        RECT 18.785000 81.895000 19.105000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 82.300000 19.105000 82.620000 ;
      LAYER met4 ;
        RECT 18.785000 82.300000 19.105000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855000 17.800000 19.175000 18.120000 ;
      LAYER met4 ;
        RECT 18.855000 17.800000 19.175000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855000 18.230000 19.175000 18.550000 ;
      LAYER met4 ;
        RECT 18.855000 18.230000 19.175000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855000 18.660000 19.175000 18.980000 ;
      LAYER met4 ;
        RECT 18.855000 18.660000 19.175000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855000 19.090000 19.175000 19.410000 ;
      LAYER met4 ;
        RECT 18.855000 19.090000 19.175000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855000 19.520000 19.175000 19.840000 ;
      LAYER met4 ;
        RECT 18.855000 19.520000 19.175000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855000 19.950000 19.175000 20.270000 ;
      LAYER met4 ;
        RECT 18.855000 19.950000 19.175000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855000 20.380000 19.175000 20.700000 ;
      LAYER met4 ;
        RECT 18.855000 20.380000 19.175000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855000 20.810000 19.175000 21.130000 ;
      LAYER met4 ;
        RECT 18.855000 20.810000 19.175000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855000 21.240000 19.175000 21.560000 ;
      LAYER met4 ;
        RECT 18.855000 21.240000 19.175000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855000 21.670000 19.175000 21.990000 ;
      LAYER met4 ;
        RECT 18.855000 21.670000 19.175000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855000 22.100000 19.175000 22.420000 ;
      LAYER met4 ;
        RECT 18.855000 22.100000 19.175000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.000000 85.815000 19.320000 86.135000 ;
      LAYER met4 ;
        RECT 19.000000 85.815000 19.320000 86.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.000000 86.250000 19.320000 86.570000 ;
      LAYER met4 ;
        RECT 19.000000 86.250000 19.320000 86.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.000000 86.690000 19.320000 87.010000 ;
      LAYER met4 ;
        RECT 19.000000 86.690000 19.320000 87.010000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 68.065000 19.505000 68.385000 ;
      LAYER met4 ;
        RECT 19.185000 68.065000 19.505000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 68.475000 19.505000 68.795000 ;
      LAYER met4 ;
        RECT 19.185000 68.475000 19.505000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 68.885000 19.505000 69.205000 ;
      LAYER met4 ;
        RECT 19.185000 68.885000 19.505000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 69.295000 19.505000 69.615000 ;
      LAYER met4 ;
        RECT 19.185000 69.295000 19.505000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 69.705000 19.505000 70.025000 ;
      LAYER met4 ;
        RECT 19.185000 69.705000 19.505000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 70.115000 19.505000 70.435000 ;
      LAYER met4 ;
        RECT 19.185000 70.115000 19.505000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 70.525000 19.505000 70.845000 ;
      LAYER met4 ;
        RECT 19.185000 70.525000 19.505000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 70.935000 19.505000 71.255000 ;
      LAYER met4 ;
        RECT 19.185000 70.935000 19.505000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 71.345000 19.505000 71.665000 ;
      LAYER met4 ;
        RECT 19.185000 71.345000 19.505000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 71.755000 19.505000 72.075000 ;
      LAYER met4 ;
        RECT 19.185000 71.755000 19.505000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 72.165000 19.505000 72.485000 ;
      LAYER met4 ;
        RECT 19.185000 72.165000 19.505000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 72.575000 19.505000 72.895000 ;
      LAYER met4 ;
        RECT 19.185000 72.575000 19.505000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 72.985000 19.505000 73.305000 ;
      LAYER met4 ;
        RECT 19.185000 72.985000 19.505000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 73.390000 19.505000 73.710000 ;
      LAYER met4 ;
        RECT 19.185000 73.390000 19.505000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 73.795000 19.505000 74.115000 ;
      LAYER met4 ;
        RECT 19.185000 73.795000 19.505000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 74.200000 19.505000 74.520000 ;
      LAYER met4 ;
        RECT 19.185000 74.200000 19.505000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 74.605000 19.505000 74.925000 ;
      LAYER met4 ;
        RECT 19.185000 74.605000 19.505000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 75.010000 19.505000 75.330000 ;
      LAYER met4 ;
        RECT 19.185000 75.010000 19.505000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 75.415000 19.505000 75.735000 ;
      LAYER met4 ;
        RECT 19.185000 75.415000 19.505000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 75.820000 19.505000 76.140000 ;
      LAYER met4 ;
        RECT 19.185000 75.820000 19.505000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 76.225000 19.505000 76.545000 ;
      LAYER met4 ;
        RECT 19.185000 76.225000 19.505000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 76.630000 19.505000 76.950000 ;
      LAYER met4 ;
        RECT 19.185000 76.630000 19.505000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 77.035000 19.505000 77.355000 ;
      LAYER met4 ;
        RECT 19.185000 77.035000 19.505000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 77.440000 19.505000 77.760000 ;
      LAYER met4 ;
        RECT 19.185000 77.440000 19.505000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 77.845000 19.505000 78.165000 ;
      LAYER met4 ;
        RECT 19.185000 77.845000 19.505000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 78.250000 19.505000 78.570000 ;
      LAYER met4 ;
        RECT 19.185000 78.250000 19.505000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 78.655000 19.505000 78.975000 ;
      LAYER met4 ;
        RECT 19.185000 78.655000 19.505000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 79.060000 19.505000 79.380000 ;
      LAYER met4 ;
        RECT 19.185000 79.060000 19.505000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 79.465000 19.505000 79.785000 ;
      LAYER met4 ;
        RECT 19.185000 79.465000 19.505000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 79.870000 19.505000 80.190000 ;
      LAYER met4 ;
        RECT 19.185000 79.870000 19.505000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 80.275000 19.505000 80.595000 ;
      LAYER met4 ;
        RECT 19.185000 80.275000 19.505000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 80.680000 19.505000 81.000000 ;
      LAYER met4 ;
        RECT 19.185000 80.680000 19.505000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 81.085000 19.505000 81.405000 ;
      LAYER met4 ;
        RECT 19.185000 81.085000 19.505000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 81.490000 19.505000 81.810000 ;
      LAYER met4 ;
        RECT 19.185000 81.490000 19.505000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 81.895000 19.505000 82.215000 ;
      LAYER met4 ;
        RECT 19.185000 81.895000 19.505000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 82.300000 19.505000 82.620000 ;
      LAYER met4 ;
        RECT 19.185000 82.300000 19.505000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 82.950000 19.510000 83.270000 ;
      LAYER met4 ;
        RECT 19.190000 82.950000 19.510000 83.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 83.410000 19.510000 83.730000 ;
      LAYER met4 ;
        RECT 19.190000 83.410000 19.510000 83.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 83.870000 19.510000 84.190000 ;
      LAYER met4 ;
        RECT 19.190000 83.870000 19.510000 84.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 84.335000 19.510000 84.655000 ;
      LAYER met4 ;
        RECT 19.190000 84.335000 19.510000 84.655000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 84.800000 19.510000 85.120000 ;
      LAYER met4 ;
        RECT 19.190000 84.800000 19.510000 85.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 85.265000 19.510000 85.585000 ;
      LAYER met4 ;
        RECT 19.190000 85.265000 19.510000 85.585000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260000 17.800000 19.580000 18.120000 ;
      LAYER met4 ;
        RECT 19.260000 17.800000 19.580000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260000 18.230000 19.580000 18.550000 ;
      LAYER met4 ;
        RECT 19.260000 18.230000 19.580000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260000 18.660000 19.580000 18.980000 ;
      LAYER met4 ;
        RECT 19.260000 18.660000 19.580000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260000 19.090000 19.580000 19.410000 ;
      LAYER met4 ;
        RECT 19.260000 19.090000 19.580000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260000 19.520000 19.580000 19.840000 ;
      LAYER met4 ;
        RECT 19.260000 19.520000 19.580000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260000 19.950000 19.580000 20.270000 ;
      LAYER met4 ;
        RECT 19.260000 19.950000 19.580000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260000 20.380000 19.580000 20.700000 ;
      LAYER met4 ;
        RECT 19.260000 20.380000 19.580000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260000 20.810000 19.580000 21.130000 ;
      LAYER met4 ;
        RECT 19.260000 20.810000 19.580000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260000 21.240000 19.580000 21.560000 ;
      LAYER met4 ;
        RECT 19.260000 21.240000 19.580000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260000 21.670000 19.580000 21.990000 ;
      LAYER met4 ;
        RECT 19.260000 21.670000 19.580000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260000 22.100000 19.580000 22.420000 ;
      LAYER met4 ;
        RECT 19.260000 22.100000 19.580000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 68.065000 19.905000 68.385000 ;
      LAYER met4 ;
        RECT 19.585000 68.065000 19.905000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 68.475000 19.905000 68.795000 ;
      LAYER met4 ;
        RECT 19.585000 68.475000 19.905000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 68.885000 19.905000 69.205000 ;
      LAYER met4 ;
        RECT 19.585000 68.885000 19.905000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 69.295000 19.905000 69.615000 ;
      LAYER met4 ;
        RECT 19.585000 69.295000 19.905000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 69.705000 19.905000 70.025000 ;
      LAYER met4 ;
        RECT 19.585000 69.705000 19.905000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 70.115000 19.905000 70.435000 ;
      LAYER met4 ;
        RECT 19.585000 70.115000 19.905000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 70.525000 19.905000 70.845000 ;
      LAYER met4 ;
        RECT 19.585000 70.525000 19.905000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 70.935000 19.905000 71.255000 ;
      LAYER met4 ;
        RECT 19.585000 70.935000 19.905000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 71.345000 19.905000 71.665000 ;
      LAYER met4 ;
        RECT 19.585000 71.345000 19.905000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 71.755000 19.905000 72.075000 ;
      LAYER met4 ;
        RECT 19.585000 71.755000 19.905000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 72.165000 19.905000 72.485000 ;
      LAYER met4 ;
        RECT 19.585000 72.165000 19.905000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 72.575000 19.905000 72.895000 ;
      LAYER met4 ;
        RECT 19.585000 72.575000 19.905000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 72.985000 19.905000 73.305000 ;
      LAYER met4 ;
        RECT 19.585000 72.985000 19.905000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 73.390000 19.905000 73.710000 ;
      LAYER met4 ;
        RECT 19.585000 73.390000 19.905000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 73.795000 19.905000 74.115000 ;
      LAYER met4 ;
        RECT 19.585000 73.795000 19.905000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 74.200000 19.905000 74.520000 ;
      LAYER met4 ;
        RECT 19.585000 74.200000 19.905000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 74.605000 19.905000 74.925000 ;
      LAYER met4 ;
        RECT 19.585000 74.605000 19.905000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 75.010000 19.905000 75.330000 ;
      LAYER met4 ;
        RECT 19.585000 75.010000 19.905000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 75.415000 19.905000 75.735000 ;
      LAYER met4 ;
        RECT 19.585000 75.415000 19.905000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 75.820000 19.905000 76.140000 ;
      LAYER met4 ;
        RECT 19.585000 75.820000 19.905000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 76.225000 19.905000 76.545000 ;
      LAYER met4 ;
        RECT 19.585000 76.225000 19.905000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 76.630000 19.905000 76.950000 ;
      LAYER met4 ;
        RECT 19.585000 76.630000 19.905000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 77.035000 19.905000 77.355000 ;
      LAYER met4 ;
        RECT 19.585000 77.035000 19.905000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 77.440000 19.905000 77.760000 ;
      LAYER met4 ;
        RECT 19.585000 77.440000 19.905000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 77.845000 19.905000 78.165000 ;
      LAYER met4 ;
        RECT 19.585000 77.845000 19.905000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 78.250000 19.905000 78.570000 ;
      LAYER met4 ;
        RECT 19.585000 78.250000 19.905000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 78.655000 19.905000 78.975000 ;
      LAYER met4 ;
        RECT 19.585000 78.655000 19.905000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 79.060000 19.905000 79.380000 ;
      LAYER met4 ;
        RECT 19.585000 79.060000 19.905000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 79.465000 19.905000 79.785000 ;
      LAYER met4 ;
        RECT 19.585000 79.465000 19.905000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 79.870000 19.905000 80.190000 ;
      LAYER met4 ;
        RECT 19.585000 79.870000 19.905000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 80.275000 19.905000 80.595000 ;
      LAYER met4 ;
        RECT 19.585000 80.275000 19.905000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 80.680000 19.905000 81.000000 ;
      LAYER met4 ;
        RECT 19.585000 80.680000 19.905000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 81.085000 19.905000 81.405000 ;
      LAYER met4 ;
        RECT 19.585000 81.085000 19.905000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 81.490000 19.905000 81.810000 ;
      LAYER met4 ;
        RECT 19.585000 81.490000 19.905000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 81.895000 19.905000 82.215000 ;
      LAYER met4 ;
        RECT 19.585000 81.895000 19.905000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585000 82.300000 19.905000 82.620000 ;
      LAYER met4 ;
        RECT 19.585000 82.300000 19.905000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665000 17.800000 19.985000 18.120000 ;
      LAYER met4 ;
        RECT 19.665000 17.800000 19.985000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665000 18.230000 19.985000 18.550000 ;
      LAYER met4 ;
        RECT 19.665000 18.230000 19.985000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665000 18.660000 19.985000 18.980000 ;
      LAYER met4 ;
        RECT 19.665000 18.660000 19.985000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665000 19.090000 19.985000 19.410000 ;
      LAYER met4 ;
        RECT 19.665000 19.090000 19.985000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665000 19.520000 19.985000 19.840000 ;
      LAYER met4 ;
        RECT 19.665000 19.520000 19.985000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665000 19.950000 19.985000 20.270000 ;
      LAYER met4 ;
        RECT 19.665000 19.950000 19.985000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665000 20.380000 19.985000 20.700000 ;
      LAYER met4 ;
        RECT 19.665000 20.380000 19.985000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665000 20.810000 19.985000 21.130000 ;
      LAYER met4 ;
        RECT 19.665000 20.810000 19.985000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665000 21.240000 19.985000 21.560000 ;
      LAYER met4 ;
        RECT 19.665000 21.240000 19.985000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665000 21.670000 19.985000 21.990000 ;
      LAYER met4 ;
        RECT 19.665000 21.670000 19.985000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665000 22.100000 19.985000 22.420000 ;
      LAYER met4 ;
        RECT 19.665000 22.100000 19.985000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.670000 82.950000 19.990000 83.270000 ;
      LAYER met4 ;
        RECT 19.670000 82.950000 19.990000 83.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.670000 83.410000 19.990000 83.730000 ;
      LAYER met4 ;
        RECT 19.670000 83.410000 19.990000 83.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.670000 83.870000 19.990000 84.190000 ;
      LAYER met4 ;
        RECT 19.670000 83.870000 19.990000 84.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.670000 84.335000 19.990000 84.655000 ;
      LAYER met4 ;
        RECT 19.670000 84.335000 19.990000 84.655000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.670000 84.800000 19.990000 85.120000 ;
      LAYER met4 ;
        RECT 19.670000 84.800000 19.990000 85.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.670000 85.265000 19.990000 85.585000 ;
      LAYER met4 ;
        RECT 19.670000 85.265000 19.990000 85.585000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.740000 85.815000 20.060000 86.135000 ;
      LAYER met4 ;
        RECT 19.740000 85.815000 20.060000 86.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.740000 86.250000 20.060000 86.570000 ;
      LAYER met4 ;
        RECT 19.740000 86.250000 20.060000 86.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.740000 86.690000 20.060000 87.010000 ;
      LAYER met4 ;
        RECT 19.740000 86.690000 20.060000 87.010000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 68.065000 20.305000 68.385000 ;
      LAYER met4 ;
        RECT 19.985000 68.065000 20.305000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 68.475000 20.305000 68.795000 ;
      LAYER met4 ;
        RECT 19.985000 68.475000 20.305000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 68.885000 20.305000 69.205000 ;
      LAYER met4 ;
        RECT 19.985000 68.885000 20.305000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 69.295000 20.305000 69.615000 ;
      LAYER met4 ;
        RECT 19.985000 69.295000 20.305000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 69.705000 20.305000 70.025000 ;
      LAYER met4 ;
        RECT 19.985000 69.705000 20.305000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 70.115000 20.305000 70.435000 ;
      LAYER met4 ;
        RECT 19.985000 70.115000 20.305000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 70.525000 20.305000 70.845000 ;
      LAYER met4 ;
        RECT 19.985000 70.525000 20.305000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 70.935000 20.305000 71.255000 ;
      LAYER met4 ;
        RECT 19.985000 70.935000 20.305000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 71.345000 20.305000 71.665000 ;
      LAYER met4 ;
        RECT 19.985000 71.345000 20.305000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 71.755000 20.305000 72.075000 ;
      LAYER met4 ;
        RECT 19.985000 71.755000 20.305000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 72.165000 20.305000 72.485000 ;
      LAYER met4 ;
        RECT 19.985000 72.165000 20.305000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 72.575000 20.305000 72.895000 ;
      LAYER met4 ;
        RECT 19.985000 72.575000 20.305000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 72.985000 20.305000 73.305000 ;
      LAYER met4 ;
        RECT 19.985000 72.985000 20.305000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 73.390000 20.305000 73.710000 ;
      LAYER met4 ;
        RECT 19.985000 73.390000 20.305000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 73.795000 20.305000 74.115000 ;
      LAYER met4 ;
        RECT 19.985000 73.795000 20.305000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 74.200000 20.305000 74.520000 ;
      LAYER met4 ;
        RECT 19.985000 74.200000 20.305000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 74.605000 20.305000 74.925000 ;
      LAYER met4 ;
        RECT 19.985000 74.605000 20.305000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 75.010000 20.305000 75.330000 ;
      LAYER met4 ;
        RECT 19.985000 75.010000 20.305000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 75.415000 20.305000 75.735000 ;
      LAYER met4 ;
        RECT 19.985000 75.415000 20.305000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 75.820000 20.305000 76.140000 ;
      LAYER met4 ;
        RECT 19.985000 75.820000 20.305000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 76.225000 20.305000 76.545000 ;
      LAYER met4 ;
        RECT 19.985000 76.225000 20.305000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 76.630000 20.305000 76.950000 ;
      LAYER met4 ;
        RECT 19.985000 76.630000 20.305000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 77.035000 20.305000 77.355000 ;
      LAYER met4 ;
        RECT 19.985000 77.035000 20.305000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 77.440000 20.305000 77.760000 ;
      LAYER met4 ;
        RECT 19.985000 77.440000 20.305000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 77.845000 20.305000 78.165000 ;
      LAYER met4 ;
        RECT 19.985000 77.845000 20.305000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 78.250000 20.305000 78.570000 ;
      LAYER met4 ;
        RECT 19.985000 78.250000 20.305000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 78.655000 20.305000 78.975000 ;
      LAYER met4 ;
        RECT 19.985000 78.655000 20.305000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 79.060000 20.305000 79.380000 ;
      LAYER met4 ;
        RECT 19.985000 79.060000 20.305000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 79.465000 20.305000 79.785000 ;
      LAYER met4 ;
        RECT 19.985000 79.465000 20.305000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 79.870000 20.305000 80.190000 ;
      LAYER met4 ;
        RECT 19.985000 79.870000 20.305000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 80.275000 20.305000 80.595000 ;
      LAYER met4 ;
        RECT 19.985000 80.275000 20.305000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 80.680000 20.305000 81.000000 ;
      LAYER met4 ;
        RECT 19.985000 80.680000 20.305000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 81.085000 20.305000 81.405000 ;
      LAYER met4 ;
        RECT 19.985000 81.085000 20.305000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 81.490000 20.305000 81.810000 ;
      LAYER met4 ;
        RECT 19.985000 81.490000 20.305000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 81.895000 20.305000 82.215000 ;
      LAYER met4 ;
        RECT 19.985000 81.895000 20.305000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985000 82.300000 20.305000 82.620000 ;
      LAYER met4 ;
        RECT 19.985000 82.300000 20.305000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250000 17.800000 2.570000 18.120000 ;
      LAYER met4 ;
        RECT 2.250000 17.800000 2.570000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250000 18.230000 2.570000 18.550000 ;
      LAYER met4 ;
        RECT 2.250000 18.230000 2.570000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250000 18.660000 2.570000 18.980000 ;
      LAYER met4 ;
        RECT 2.250000 18.660000 2.570000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250000 19.090000 2.570000 19.410000 ;
      LAYER met4 ;
        RECT 2.250000 19.090000 2.570000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250000 19.520000 2.570000 19.840000 ;
      LAYER met4 ;
        RECT 2.250000 19.520000 2.570000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250000 19.950000 2.570000 20.270000 ;
      LAYER met4 ;
        RECT 2.250000 19.950000 2.570000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250000 20.380000 2.570000 20.700000 ;
      LAYER met4 ;
        RECT 2.250000 20.380000 2.570000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250000 20.810000 2.570000 21.130000 ;
      LAYER met4 ;
        RECT 2.250000 20.810000 2.570000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250000 21.240000 2.570000 21.560000 ;
      LAYER met4 ;
        RECT 2.250000 21.240000 2.570000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250000 21.670000 2.570000 21.990000 ;
      LAYER met4 ;
        RECT 2.250000 21.670000 2.570000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250000 22.100000 2.570000 22.420000 ;
      LAYER met4 ;
        RECT 2.250000 22.100000 2.570000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 82.795000 2.635000 83.115000 ;
      LAYER met4 ;
        RECT 2.315000 82.795000 2.635000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 83.205000 2.635000 83.525000 ;
      LAYER met4 ;
        RECT 2.315000 83.205000 2.635000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 83.615000 2.635000 83.935000 ;
      LAYER met4 ;
        RECT 2.315000 83.615000 2.635000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 84.025000 2.635000 84.345000 ;
      LAYER met4 ;
        RECT 2.315000 84.025000 2.635000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 84.435000 2.635000 84.755000 ;
      LAYER met4 ;
        RECT 2.315000 84.435000 2.635000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 84.845000 2.635000 85.165000 ;
      LAYER met4 ;
        RECT 2.315000 84.845000 2.635000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 85.255000 2.635000 85.575000 ;
      LAYER met4 ;
        RECT 2.315000 85.255000 2.635000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 85.665000 2.635000 85.985000 ;
      LAYER met4 ;
        RECT 2.315000 85.665000 2.635000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 86.075000 2.635000 86.395000 ;
      LAYER met4 ;
        RECT 2.315000 86.075000 2.635000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 86.485000 2.635000 86.805000 ;
      LAYER met4 ;
        RECT 2.315000 86.485000 2.635000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 86.895000 2.635000 87.215000 ;
      LAYER met4 ;
        RECT 2.315000 86.895000 2.635000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 87.305000 2.635000 87.625000 ;
      LAYER met4 ;
        RECT 2.315000 87.305000 2.635000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 87.715000 2.635000 88.035000 ;
      LAYER met4 ;
        RECT 2.315000 87.715000 2.635000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 88.125000 2.635000 88.445000 ;
      LAYER met4 ;
        RECT 2.315000 88.125000 2.635000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 88.535000 2.635000 88.855000 ;
      LAYER met4 ;
        RECT 2.315000 88.535000 2.635000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 88.945000 2.635000 89.265000 ;
      LAYER met4 ;
        RECT 2.315000 88.945000 2.635000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 89.355000 2.635000 89.675000 ;
      LAYER met4 ;
        RECT 2.315000 89.355000 2.635000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 89.765000 2.635000 90.085000 ;
      LAYER met4 ;
        RECT 2.315000 89.765000 2.635000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 90.175000 2.635000 90.495000 ;
      LAYER met4 ;
        RECT 2.315000 90.175000 2.635000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 90.585000 2.635000 90.905000 ;
      LAYER met4 ;
        RECT 2.315000 90.585000 2.635000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 90.995000 2.635000 91.315000 ;
      LAYER met4 ;
        RECT 2.315000 90.995000 2.635000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 91.405000 2.635000 91.725000 ;
      LAYER met4 ;
        RECT 2.315000 91.405000 2.635000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 91.815000 2.635000 92.135000 ;
      LAYER met4 ;
        RECT 2.315000 91.815000 2.635000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 92.225000 2.635000 92.545000 ;
      LAYER met4 ;
        RECT 2.315000 92.225000 2.635000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315000 92.635000 2.635000 92.955000 ;
      LAYER met4 ;
        RECT 2.315000 92.635000 2.635000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 68.065000 2.705000 68.385000 ;
      LAYER met4 ;
        RECT 2.385000 68.065000 2.705000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 68.475000 2.705000 68.795000 ;
      LAYER met4 ;
        RECT 2.385000 68.475000 2.705000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 68.885000 2.705000 69.205000 ;
      LAYER met4 ;
        RECT 2.385000 68.885000 2.705000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 69.295000 2.705000 69.615000 ;
      LAYER met4 ;
        RECT 2.385000 69.295000 2.705000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 69.705000 2.705000 70.025000 ;
      LAYER met4 ;
        RECT 2.385000 69.705000 2.705000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 70.115000 2.705000 70.435000 ;
      LAYER met4 ;
        RECT 2.385000 70.115000 2.705000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 70.525000 2.705000 70.845000 ;
      LAYER met4 ;
        RECT 2.385000 70.525000 2.705000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 70.935000 2.705000 71.255000 ;
      LAYER met4 ;
        RECT 2.385000 70.935000 2.705000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 71.345000 2.705000 71.665000 ;
      LAYER met4 ;
        RECT 2.385000 71.345000 2.705000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 71.755000 2.705000 72.075000 ;
      LAYER met4 ;
        RECT 2.385000 71.755000 2.705000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 72.165000 2.705000 72.485000 ;
      LAYER met4 ;
        RECT 2.385000 72.165000 2.705000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 72.575000 2.705000 72.895000 ;
      LAYER met4 ;
        RECT 2.385000 72.575000 2.705000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 72.985000 2.705000 73.305000 ;
      LAYER met4 ;
        RECT 2.385000 72.985000 2.705000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 73.390000 2.705000 73.710000 ;
      LAYER met4 ;
        RECT 2.385000 73.390000 2.705000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 73.795000 2.705000 74.115000 ;
      LAYER met4 ;
        RECT 2.385000 73.795000 2.705000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 74.200000 2.705000 74.520000 ;
      LAYER met4 ;
        RECT 2.385000 74.200000 2.705000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 74.605000 2.705000 74.925000 ;
      LAYER met4 ;
        RECT 2.385000 74.605000 2.705000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 75.010000 2.705000 75.330000 ;
      LAYER met4 ;
        RECT 2.385000 75.010000 2.705000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 75.415000 2.705000 75.735000 ;
      LAYER met4 ;
        RECT 2.385000 75.415000 2.705000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 75.820000 2.705000 76.140000 ;
      LAYER met4 ;
        RECT 2.385000 75.820000 2.705000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 76.225000 2.705000 76.545000 ;
      LAYER met4 ;
        RECT 2.385000 76.225000 2.705000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 76.630000 2.705000 76.950000 ;
      LAYER met4 ;
        RECT 2.385000 76.630000 2.705000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 77.035000 2.705000 77.355000 ;
      LAYER met4 ;
        RECT 2.385000 77.035000 2.705000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 77.440000 2.705000 77.760000 ;
      LAYER met4 ;
        RECT 2.385000 77.440000 2.705000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 77.845000 2.705000 78.165000 ;
      LAYER met4 ;
        RECT 2.385000 77.845000 2.705000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 78.250000 2.705000 78.570000 ;
      LAYER met4 ;
        RECT 2.385000 78.250000 2.705000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 78.655000 2.705000 78.975000 ;
      LAYER met4 ;
        RECT 2.385000 78.655000 2.705000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 79.060000 2.705000 79.380000 ;
      LAYER met4 ;
        RECT 2.385000 79.060000 2.705000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 79.465000 2.705000 79.785000 ;
      LAYER met4 ;
        RECT 2.385000 79.465000 2.705000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 79.870000 2.705000 80.190000 ;
      LAYER met4 ;
        RECT 2.385000 79.870000 2.705000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 80.275000 2.705000 80.595000 ;
      LAYER met4 ;
        RECT 2.385000 80.275000 2.705000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 80.680000 2.705000 81.000000 ;
      LAYER met4 ;
        RECT 2.385000 80.680000 2.705000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 81.085000 2.705000 81.405000 ;
      LAYER met4 ;
        RECT 2.385000 81.085000 2.705000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 81.490000 2.705000 81.810000 ;
      LAYER met4 ;
        RECT 2.385000 81.490000 2.705000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 81.895000 2.705000 82.215000 ;
      LAYER met4 ;
        RECT 2.385000 81.895000 2.705000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385000 82.300000 2.705000 82.620000 ;
      LAYER met4 ;
        RECT 2.385000 82.300000 2.705000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655000 17.800000 2.975000 18.120000 ;
      LAYER met4 ;
        RECT 2.655000 17.800000 2.975000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655000 18.230000 2.975000 18.550000 ;
      LAYER met4 ;
        RECT 2.655000 18.230000 2.975000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655000 18.660000 2.975000 18.980000 ;
      LAYER met4 ;
        RECT 2.655000 18.660000 2.975000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655000 19.090000 2.975000 19.410000 ;
      LAYER met4 ;
        RECT 2.655000 19.090000 2.975000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655000 19.520000 2.975000 19.840000 ;
      LAYER met4 ;
        RECT 2.655000 19.520000 2.975000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655000 19.950000 2.975000 20.270000 ;
      LAYER met4 ;
        RECT 2.655000 19.950000 2.975000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655000 20.380000 2.975000 20.700000 ;
      LAYER met4 ;
        RECT 2.655000 20.380000 2.975000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655000 20.810000 2.975000 21.130000 ;
      LAYER met4 ;
        RECT 2.655000 20.810000 2.975000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655000 21.240000 2.975000 21.560000 ;
      LAYER met4 ;
        RECT 2.655000 21.240000 2.975000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655000 21.670000 2.975000 21.990000 ;
      LAYER met4 ;
        RECT 2.655000 21.670000 2.975000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655000 22.100000 2.975000 22.420000 ;
      LAYER met4 ;
        RECT 2.655000 22.100000 2.975000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 82.795000 3.045000 83.115000 ;
      LAYER met4 ;
        RECT 2.725000 82.795000 3.045000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 83.205000 3.045000 83.525000 ;
      LAYER met4 ;
        RECT 2.725000 83.205000 3.045000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 83.615000 3.045000 83.935000 ;
      LAYER met4 ;
        RECT 2.725000 83.615000 3.045000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 84.025000 3.045000 84.345000 ;
      LAYER met4 ;
        RECT 2.725000 84.025000 3.045000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 84.435000 3.045000 84.755000 ;
      LAYER met4 ;
        RECT 2.725000 84.435000 3.045000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 84.845000 3.045000 85.165000 ;
      LAYER met4 ;
        RECT 2.725000 84.845000 3.045000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 85.255000 3.045000 85.575000 ;
      LAYER met4 ;
        RECT 2.725000 85.255000 3.045000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 85.665000 3.045000 85.985000 ;
      LAYER met4 ;
        RECT 2.725000 85.665000 3.045000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 86.075000 3.045000 86.395000 ;
      LAYER met4 ;
        RECT 2.725000 86.075000 3.045000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 86.485000 3.045000 86.805000 ;
      LAYER met4 ;
        RECT 2.725000 86.485000 3.045000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 86.895000 3.045000 87.215000 ;
      LAYER met4 ;
        RECT 2.725000 86.895000 3.045000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 87.305000 3.045000 87.625000 ;
      LAYER met4 ;
        RECT 2.725000 87.305000 3.045000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 87.715000 3.045000 88.035000 ;
      LAYER met4 ;
        RECT 2.725000 87.715000 3.045000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 88.125000 3.045000 88.445000 ;
      LAYER met4 ;
        RECT 2.725000 88.125000 3.045000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 88.535000 3.045000 88.855000 ;
      LAYER met4 ;
        RECT 2.725000 88.535000 3.045000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 88.945000 3.045000 89.265000 ;
      LAYER met4 ;
        RECT 2.725000 88.945000 3.045000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 89.355000 3.045000 89.675000 ;
      LAYER met4 ;
        RECT 2.725000 89.355000 3.045000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 89.765000 3.045000 90.085000 ;
      LAYER met4 ;
        RECT 2.725000 89.765000 3.045000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 90.175000 3.045000 90.495000 ;
      LAYER met4 ;
        RECT 2.725000 90.175000 3.045000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 90.585000 3.045000 90.905000 ;
      LAYER met4 ;
        RECT 2.725000 90.585000 3.045000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 90.995000 3.045000 91.315000 ;
      LAYER met4 ;
        RECT 2.725000 90.995000 3.045000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 91.405000 3.045000 91.725000 ;
      LAYER met4 ;
        RECT 2.725000 91.405000 3.045000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 91.815000 3.045000 92.135000 ;
      LAYER met4 ;
        RECT 2.725000 91.815000 3.045000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 92.225000 3.045000 92.545000 ;
      LAYER met4 ;
        RECT 2.725000 92.225000 3.045000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725000 92.635000 3.045000 92.955000 ;
      LAYER met4 ;
        RECT 2.725000 92.635000 3.045000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 68.065000 3.105000 68.385000 ;
      LAYER met4 ;
        RECT 2.785000 68.065000 3.105000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 68.475000 3.105000 68.795000 ;
      LAYER met4 ;
        RECT 2.785000 68.475000 3.105000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 68.885000 3.105000 69.205000 ;
      LAYER met4 ;
        RECT 2.785000 68.885000 3.105000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 69.295000 3.105000 69.615000 ;
      LAYER met4 ;
        RECT 2.785000 69.295000 3.105000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 69.705000 3.105000 70.025000 ;
      LAYER met4 ;
        RECT 2.785000 69.705000 3.105000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 70.115000 3.105000 70.435000 ;
      LAYER met4 ;
        RECT 2.785000 70.115000 3.105000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 70.525000 3.105000 70.845000 ;
      LAYER met4 ;
        RECT 2.785000 70.525000 3.105000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 70.935000 3.105000 71.255000 ;
      LAYER met4 ;
        RECT 2.785000 70.935000 3.105000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 71.345000 3.105000 71.665000 ;
      LAYER met4 ;
        RECT 2.785000 71.345000 3.105000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 71.755000 3.105000 72.075000 ;
      LAYER met4 ;
        RECT 2.785000 71.755000 3.105000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 72.165000 3.105000 72.485000 ;
      LAYER met4 ;
        RECT 2.785000 72.165000 3.105000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 72.575000 3.105000 72.895000 ;
      LAYER met4 ;
        RECT 2.785000 72.575000 3.105000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 72.985000 3.105000 73.305000 ;
      LAYER met4 ;
        RECT 2.785000 72.985000 3.105000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 73.390000 3.105000 73.710000 ;
      LAYER met4 ;
        RECT 2.785000 73.390000 3.105000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 73.795000 3.105000 74.115000 ;
      LAYER met4 ;
        RECT 2.785000 73.795000 3.105000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 74.200000 3.105000 74.520000 ;
      LAYER met4 ;
        RECT 2.785000 74.200000 3.105000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 74.605000 3.105000 74.925000 ;
      LAYER met4 ;
        RECT 2.785000 74.605000 3.105000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 75.010000 3.105000 75.330000 ;
      LAYER met4 ;
        RECT 2.785000 75.010000 3.105000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 75.415000 3.105000 75.735000 ;
      LAYER met4 ;
        RECT 2.785000 75.415000 3.105000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 75.820000 3.105000 76.140000 ;
      LAYER met4 ;
        RECT 2.785000 75.820000 3.105000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 76.225000 3.105000 76.545000 ;
      LAYER met4 ;
        RECT 2.785000 76.225000 3.105000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 76.630000 3.105000 76.950000 ;
      LAYER met4 ;
        RECT 2.785000 76.630000 3.105000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 77.035000 3.105000 77.355000 ;
      LAYER met4 ;
        RECT 2.785000 77.035000 3.105000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 77.440000 3.105000 77.760000 ;
      LAYER met4 ;
        RECT 2.785000 77.440000 3.105000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 77.845000 3.105000 78.165000 ;
      LAYER met4 ;
        RECT 2.785000 77.845000 3.105000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 78.250000 3.105000 78.570000 ;
      LAYER met4 ;
        RECT 2.785000 78.250000 3.105000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 78.655000 3.105000 78.975000 ;
      LAYER met4 ;
        RECT 2.785000 78.655000 3.105000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 79.060000 3.105000 79.380000 ;
      LAYER met4 ;
        RECT 2.785000 79.060000 3.105000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 79.465000 3.105000 79.785000 ;
      LAYER met4 ;
        RECT 2.785000 79.465000 3.105000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 79.870000 3.105000 80.190000 ;
      LAYER met4 ;
        RECT 2.785000 79.870000 3.105000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 80.275000 3.105000 80.595000 ;
      LAYER met4 ;
        RECT 2.785000 80.275000 3.105000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 80.680000 3.105000 81.000000 ;
      LAYER met4 ;
        RECT 2.785000 80.680000 3.105000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 81.085000 3.105000 81.405000 ;
      LAYER met4 ;
        RECT 2.785000 81.085000 3.105000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 81.490000 3.105000 81.810000 ;
      LAYER met4 ;
        RECT 2.785000 81.490000 3.105000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 81.895000 3.105000 82.215000 ;
      LAYER met4 ;
        RECT 2.785000 81.895000 3.105000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785000 82.300000 3.105000 82.620000 ;
      LAYER met4 ;
        RECT 2.785000 82.300000 3.105000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070000 17.800000 20.390000 18.120000 ;
      LAYER met4 ;
        RECT 20.070000 17.800000 20.390000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070000 18.230000 20.390000 18.550000 ;
      LAYER met4 ;
        RECT 20.070000 18.230000 20.390000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070000 18.660000 20.390000 18.980000 ;
      LAYER met4 ;
        RECT 20.070000 18.660000 20.390000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070000 19.090000 20.390000 19.410000 ;
      LAYER met4 ;
        RECT 20.070000 19.090000 20.390000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070000 19.520000 20.390000 19.840000 ;
      LAYER met4 ;
        RECT 20.070000 19.520000 20.390000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070000 19.950000 20.390000 20.270000 ;
      LAYER met4 ;
        RECT 20.070000 19.950000 20.390000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070000 20.380000 20.390000 20.700000 ;
      LAYER met4 ;
        RECT 20.070000 20.380000 20.390000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070000 20.810000 20.390000 21.130000 ;
      LAYER met4 ;
        RECT 20.070000 20.810000 20.390000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070000 21.240000 20.390000 21.560000 ;
      LAYER met4 ;
        RECT 20.070000 21.240000 20.390000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070000 21.670000 20.390000 21.990000 ;
      LAYER met4 ;
        RECT 20.070000 21.670000 20.390000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070000 22.100000 20.390000 22.420000 ;
      LAYER met4 ;
        RECT 20.070000 22.100000 20.390000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150000 82.950000 20.470000 83.270000 ;
      LAYER met4 ;
        RECT 20.150000 82.950000 20.470000 83.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150000 83.410000 20.470000 83.730000 ;
      LAYER met4 ;
        RECT 20.150000 83.410000 20.470000 83.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150000 83.870000 20.470000 84.190000 ;
      LAYER met4 ;
        RECT 20.150000 83.870000 20.470000 84.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150000 84.335000 20.470000 84.655000 ;
      LAYER met4 ;
        RECT 20.150000 84.335000 20.470000 84.655000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150000 84.800000 20.470000 85.120000 ;
      LAYER met4 ;
        RECT 20.150000 84.800000 20.470000 85.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150000 85.265000 20.470000 85.585000 ;
      LAYER met4 ;
        RECT 20.150000 85.265000 20.470000 85.585000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 68.065000 20.705000 68.385000 ;
      LAYER met4 ;
        RECT 20.385000 68.065000 20.705000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 68.475000 20.705000 68.795000 ;
      LAYER met4 ;
        RECT 20.385000 68.475000 20.705000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 68.885000 20.705000 69.205000 ;
      LAYER met4 ;
        RECT 20.385000 68.885000 20.705000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 69.295000 20.705000 69.615000 ;
      LAYER met4 ;
        RECT 20.385000 69.295000 20.705000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 69.705000 20.705000 70.025000 ;
      LAYER met4 ;
        RECT 20.385000 69.705000 20.705000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 70.115000 20.705000 70.435000 ;
      LAYER met4 ;
        RECT 20.385000 70.115000 20.705000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 70.525000 20.705000 70.845000 ;
      LAYER met4 ;
        RECT 20.385000 70.525000 20.705000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 70.935000 20.705000 71.255000 ;
      LAYER met4 ;
        RECT 20.385000 70.935000 20.705000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 71.345000 20.705000 71.665000 ;
      LAYER met4 ;
        RECT 20.385000 71.345000 20.705000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 71.755000 20.705000 72.075000 ;
      LAYER met4 ;
        RECT 20.385000 71.755000 20.705000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 72.165000 20.705000 72.485000 ;
      LAYER met4 ;
        RECT 20.385000 72.165000 20.705000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 72.575000 20.705000 72.895000 ;
      LAYER met4 ;
        RECT 20.385000 72.575000 20.705000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 72.985000 20.705000 73.305000 ;
      LAYER met4 ;
        RECT 20.385000 72.985000 20.705000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 73.390000 20.705000 73.710000 ;
      LAYER met4 ;
        RECT 20.385000 73.390000 20.705000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 73.795000 20.705000 74.115000 ;
      LAYER met4 ;
        RECT 20.385000 73.795000 20.705000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 74.200000 20.705000 74.520000 ;
      LAYER met4 ;
        RECT 20.385000 74.200000 20.705000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 74.605000 20.705000 74.925000 ;
      LAYER met4 ;
        RECT 20.385000 74.605000 20.705000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 75.010000 20.705000 75.330000 ;
      LAYER met4 ;
        RECT 20.385000 75.010000 20.705000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 75.415000 20.705000 75.735000 ;
      LAYER met4 ;
        RECT 20.385000 75.415000 20.705000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 75.820000 20.705000 76.140000 ;
      LAYER met4 ;
        RECT 20.385000 75.820000 20.705000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 76.225000 20.705000 76.545000 ;
      LAYER met4 ;
        RECT 20.385000 76.225000 20.705000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 76.630000 20.705000 76.950000 ;
      LAYER met4 ;
        RECT 20.385000 76.630000 20.705000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 77.035000 20.705000 77.355000 ;
      LAYER met4 ;
        RECT 20.385000 77.035000 20.705000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 77.440000 20.705000 77.760000 ;
      LAYER met4 ;
        RECT 20.385000 77.440000 20.705000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 77.845000 20.705000 78.165000 ;
      LAYER met4 ;
        RECT 20.385000 77.845000 20.705000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 78.250000 20.705000 78.570000 ;
      LAYER met4 ;
        RECT 20.385000 78.250000 20.705000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 78.655000 20.705000 78.975000 ;
      LAYER met4 ;
        RECT 20.385000 78.655000 20.705000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 79.060000 20.705000 79.380000 ;
      LAYER met4 ;
        RECT 20.385000 79.060000 20.705000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 79.465000 20.705000 79.785000 ;
      LAYER met4 ;
        RECT 20.385000 79.465000 20.705000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 79.870000 20.705000 80.190000 ;
      LAYER met4 ;
        RECT 20.385000 79.870000 20.705000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 80.275000 20.705000 80.595000 ;
      LAYER met4 ;
        RECT 20.385000 80.275000 20.705000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 80.680000 20.705000 81.000000 ;
      LAYER met4 ;
        RECT 20.385000 80.680000 20.705000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 81.085000 20.705000 81.405000 ;
      LAYER met4 ;
        RECT 20.385000 81.085000 20.705000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 81.490000 20.705000 81.810000 ;
      LAYER met4 ;
        RECT 20.385000 81.490000 20.705000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 81.895000 20.705000 82.215000 ;
      LAYER met4 ;
        RECT 20.385000 81.895000 20.705000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385000 82.300000 20.705000 82.620000 ;
      LAYER met4 ;
        RECT 20.385000 82.300000 20.705000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475000 17.800000 20.795000 18.120000 ;
      LAYER met4 ;
        RECT 20.475000 17.800000 20.795000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475000 18.230000 20.795000 18.550000 ;
      LAYER met4 ;
        RECT 20.475000 18.230000 20.795000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475000 18.660000 20.795000 18.980000 ;
      LAYER met4 ;
        RECT 20.475000 18.660000 20.795000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475000 19.090000 20.795000 19.410000 ;
      LAYER met4 ;
        RECT 20.475000 19.090000 20.795000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475000 19.520000 20.795000 19.840000 ;
      LAYER met4 ;
        RECT 20.475000 19.520000 20.795000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475000 19.950000 20.795000 20.270000 ;
      LAYER met4 ;
        RECT 20.475000 19.950000 20.795000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475000 20.380000 20.795000 20.700000 ;
      LAYER met4 ;
        RECT 20.475000 20.380000 20.795000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475000 20.810000 20.795000 21.130000 ;
      LAYER met4 ;
        RECT 20.475000 20.810000 20.795000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475000 21.240000 20.795000 21.560000 ;
      LAYER met4 ;
        RECT 20.475000 21.240000 20.795000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475000 21.670000 20.795000 21.990000 ;
      LAYER met4 ;
        RECT 20.475000 21.670000 20.795000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475000 22.100000 20.795000 22.420000 ;
      LAYER met4 ;
        RECT 20.475000 22.100000 20.795000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.630000 82.950000 20.950000 83.270000 ;
      LAYER met4 ;
        RECT 20.630000 82.950000 20.950000 83.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.630000 83.410000 20.950000 83.730000 ;
      LAYER met4 ;
        RECT 20.630000 83.410000 20.950000 83.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.630000 83.870000 20.950000 84.190000 ;
      LAYER met4 ;
        RECT 20.630000 83.870000 20.950000 84.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.630000 84.335000 20.950000 84.655000 ;
      LAYER met4 ;
        RECT 20.630000 84.335000 20.950000 84.655000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.630000 84.800000 20.950000 85.120000 ;
      LAYER met4 ;
        RECT 20.630000 84.800000 20.950000 85.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.630000 85.265000 20.950000 85.585000 ;
      LAYER met4 ;
        RECT 20.630000 85.265000 20.950000 85.585000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 68.065000 21.105000 68.385000 ;
      LAYER met4 ;
        RECT 20.785000 68.065000 21.105000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 68.475000 21.105000 68.795000 ;
      LAYER met4 ;
        RECT 20.785000 68.475000 21.105000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 68.885000 21.105000 69.205000 ;
      LAYER met4 ;
        RECT 20.785000 68.885000 21.105000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 69.295000 21.105000 69.615000 ;
      LAYER met4 ;
        RECT 20.785000 69.295000 21.105000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 69.705000 21.105000 70.025000 ;
      LAYER met4 ;
        RECT 20.785000 69.705000 21.105000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 70.115000 21.105000 70.435000 ;
      LAYER met4 ;
        RECT 20.785000 70.115000 21.105000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 70.525000 21.105000 70.845000 ;
      LAYER met4 ;
        RECT 20.785000 70.525000 21.105000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 70.935000 21.105000 71.255000 ;
      LAYER met4 ;
        RECT 20.785000 70.935000 21.105000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 71.345000 21.105000 71.665000 ;
      LAYER met4 ;
        RECT 20.785000 71.345000 21.105000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 71.755000 21.105000 72.075000 ;
      LAYER met4 ;
        RECT 20.785000 71.755000 21.105000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 72.165000 21.105000 72.485000 ;
      LAYER met4 ;
        RECT 20.785000 72.165000 21.105000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 72.575000 21.105000 72.895000 ;
      LAYER met4 ;
        RECT 20.785000 72.575000 21.105000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 72.985000 21.105000 73.305000 ;
      LAYER met4 ;
        RECT 20.785000 72.985000 21.105000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 73.390000 21.105000 73.710000 ;
      LAYER met4 ;
        RECT 20.785000 73.390000 21.105000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 73.795000 21.105000 74.115000 ;
      LAYER met4 ;
        RECT 20.785000 73.795000 21.105000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 74.200000 21.105000 74.520000 ;
      LAYER met4 ;
        RECT 20.785000 74.200000 21.105000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 74.605000 21.105000 74.925000 ;
      LAYER met4 ;
        RECT 20.785000 74.605000 21.105000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 75.010000 21.105000 75.330000 ;
      LAYER met4 ;
        RECT 20.785000 75.010000 21.105000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 75.415000 21.105000 75.735000 ;
      LAYER met4 ;
        RECT 20.785000 75.415000 21.105000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 75.820000 21.105000 76.140000 ;
      LAYER met4 ;
        RECT 20.785000 75.820000 21.105000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 76.225000 21.105000 76.545000 ;
      LAYER met4 ;
        RECT 20.785000 76.225000 21.105000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 76.630000 21.105000 76.950000 ;
      LAYER met4 ;
        RECT 20.785000 76.630000 21.105000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 77.035000 21.105000 77.355000 ;
      LAYER met4 ;
        RECT 20.785000 77.035000 21.105000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 77.440000 21.105000 77.760000 ;
      LAYER met4 ;
        RECT 20.785000 77.440000 21.105000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 77.845000 21.105000 78.165000 ;
      LAYER met4 ;
        RECT 20.785000 77.845000 21.105000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 78.250000 21.105000 78.570000 ;
      LAYER met4 ;
        RECT 20.785000 78.250000 21.105000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 78.655000 21.105000 78.975000 ;
      LAYER met4 ;
        RECT 20.785000 78.655000 21.105000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 79.060000 21.105000 79.380000 ;
      LAYER met4 ;
        RECT 20.785000 79.060000 21.105000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 79.465000 21.105000 79.785000 ;
      LAYER met4 ;
        RECT 20.785000 79.465000 21.105000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 79.870000 21.105000 80.190000 ;
      LAYER met4 ;
        RECT 20.785000 79.870000 21.105000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 80.275000 21.105000 80.595000 ;
      LAYER met4 ;
        RECT 20.785000 80.275000 21.105000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 80.680000 21.105000 81.000000 ;
      LAYER met4 ;
        RECT 20.785000 80.680000 21.105000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 81.085000 21.105000 81.405000 ;
      LAYER met4 ;
        RECT 20.785000 81.085000 21.105000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 81.490000 21.105000 81.810000 ;
      LAYER met4 ;
        RECT 20.785000 81.490000 21.105000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 81.895000 21.105000 82.215000 ;
      LAYER met4 ;
        RECT 20.785000 81.895000 21.105000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785000 82.300000 21.105000 82.620000 ;
      LAYER met4 ;
        RECT 20.785000 82.300000 21.105000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880000 17.800000 21.200000 18.120000 ;
      LAYER met4 ;
        RECT 20.880000 17.800000 21.200000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880000 18.230000 21.200000 18.550000 ;
      LAYER met4 ;
        RECT 20.880000 18.230000 21.200000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880000 18.660000 21.200000 18.980000 ;
      LAYER met4 ;
        RECT 20.880000 18.660000 21.200000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880000 19.090000 21.200000 19.410000 ;
      LAYER met4 ;
        RECT 20.880000 19.090000 21.200000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880000 19.520000 21.200000 19.840000 ;
      LAYER met4 ;
        RECT 20.880000 19.520000 21.200000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880000 19.950000 21.200000 20.270000 ;
      LAYER met4 ;
        RECT 20.880000 19.950000 21.200000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880000 20.380000 21.200000 20.700000 ;
      LAYER met4 ;
        RECT 20.880000 20.380000 21.200000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880000 20.810000 21.200000 21.130000 ;
      LAYER met4 ;
        RECT 20.880000 20.810000 21.200000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880000 21.240000 21.200000 21.560000 ;
      LAYER met4 ;
        RECT 20.880000 21.240000 21.200000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880000 21.670000 21.200000 21.990000 ;
      LAYER met4 ;
        RECT 20.880000 21.670000 21.200000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880000 22.100000 21.200000 22.420000 ;
      LAYER met4 ;
        RECT 20.880000 22.100000 21.200000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.110000 82.950000 21.430000 83.270000 ;
      LAYER met4 ;
        RECT 21.110000 82.950000 21.430000 83.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.110000 83.410000 21.430000 83.730000 ;
      LAYER met4 ;
        RECT 21.110000 83.410000 21.430000 83.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.110000 83.870000 21.430000 84.190000 ;
      LAYER met4 ;
        RECT 21.110000 83.870000 21.430000 84.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.110000 84.335000 21.430000 84.655000 ;
      LAYER met4 ;
        RECT 21.110000 84.335000 21.430000 84.655000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.110000 84.800000 21.430000 85.120000 ;
      LAYER met4 ;
        RECT 21.110000 84.800000 21.430000 85.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.110000 85.265000 21.430000 85.585000 ;
      LAYER met4 ;
        RECT 21.110000 85.265000 21.430000 85.585000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 68.065000 21.505000 68.385000 ;
      LAYER met4 ;
        RECT 21.185000 68.065000 21.505000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 68.475000 21.505000 68.795000 ;
      LAYER met4 ;
        RECT 21.185000 68.475000 21.505000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 68.885000 21.505000 69.205000 ;
      LAYER met4 ;
        RECT 21.185000 68.885000 21.505000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 69.295000 21.505000 69.615000 ;
      LAYER met4 ;
        RECT 21.185000 69.295000 21.505000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 69.705000 21.505000 70.025000 ;
      LAYER met4 ;
        RECT 21.185000 69.705000 21.505000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 70.115000 21.505000 70.435000 ;
      LAYER met4 ;
        RECT 21.185000 70.115000 21.505000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 70.525000 21.505000 70.845000 ;
      LAYER met4 ;
        RECT 21.185000 70.525000 21.505000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 70.935000 21.505000 71.255000 ;
      LAYER met4 ;
        RECT 21.185000 70.935000 21.505000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 71.345000 21.505000 71.665000 ;
      LAYER met4 ;
        RECT 21.185000 71.345000 21.505000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 71.755000 21.505000 72.075000 ;
      LAYER met4 ;
        RECT 21.185000 71.755000 21.505000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 72.165000 21.505000 72.485000 ;
      LAYER met4 ;
        RECT 21.185000 72.165000 21.505000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 72.575000 21.505000 72.895000 ;
      LAYER met4 ;
        RECT 21.185000 72.575000 21.505000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 72.985000 21.505000 73.305000 ;
      LAYER met4 ;
        RECT 21.185000 72.985000 21.505000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 73.390000 21.505000 73.710000 ;
      LAYER met4 ;
        RECT 21.185000 73.390000 21.505000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 73.795000 21.505000 74.115000 ;
      LAYER met4 ;
        RECT 21.185000 73.795000 21.505000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 74.200000 21.505000 74.520000 ;
      LAYER met4 ;
        RECT 21.185000 74.200000 21.505000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 74.605000 21.505000 74.925000 ;
      LAYER met4 ;
        RECT 21.185000 74.605000 21.505000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 75.010000 21.505000 75.330000 ;
      LAYER met4 ;
        RECT 21.185000 75.010000 21.505000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 75.415000 21.505000 75.735000 ;
      LAYER met4 ;
        RECT 21.185000 75.415000 21.505000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 75.820000 21.505000 76.140000 ;
      LAYER met4 ;
        RECT 21.185000 75.820000 21.505000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 76.225000 21.505000 76.545000 ;
      LAYER met4 ;
        RECT 21.185000 76.225000 21.505000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 76.630000 21.505000 76.950000 ;
      LAYER met4 ;
        RECT 21.185000 76.630000 21.505000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 77.035000 21.505000 77.355000 ;
      LAYER met4 ;
        RECT 21.185000 77.035000 21.505000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 77.440000 21.505000 77.760000 ;
      LAYER met4 ;
        RECT 21.185000 77.440000 21.505000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 77.845000 21.505000 78.165000 ;
      LAYER met4 ;
        RECT 21.185000 77.845000 21.505000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 78.250000 21.505000 78.570000 ;
      LAYER met4 ;
        RECT 21.185000 78.250000 21.505000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 78.655000 21.505000 78.975000 ;
      LAYER met4 ;
        RECT 21.185000 78.655000 21.505000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 79.060000 21.505000 79.380000 ;
      LAYER met4 ;
        RECT 21.185000 79.060000 21.505000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 79.465000 21.505000 79.785000 ;
      LAYER met4 ;
        RECT 21.185000 79.465000 21.505000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 79.870000 21.505000 80.190000 ;
      LAYER met4 ;
        RECT 21.185000 79.870000 21.505000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 80.275000 21.505000 80.595000 ;
      LAYER met4 ;
        RECT 21.185000 80.275000 21.505000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 80.680000 21.505000 81.000000 ;
      LAYER met4 ;
        RECT 21.185000 80.680000 21.505000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 81.085000 21.505000 81.405000 ;
      LAYER met4 ;
        RECT 21.185000 81.085000 21.505000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 81.490000 21.505000 81.810000 ;
      LAYER met4 ;
        RECT 21.185000 81.490000 21.505000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 81.895000 21.505000 82.215000 ;
      LAYER met4 ;
        RECT 21.185000 81.895000 21.505000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185000 82.300000 21.505000 82.620000 ;
      LAYER met4 ;
        RECT 21.185000 82.300000 21.505000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285000 17.800000 21.605000 18.120000 ;
      LAYER met4 ;
        RECT 21.285000 17.800000 21.605000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285000 18.230000 21.605000 18.550000 ;
      LAYER met4 ;
        RECT 21.285000 18.230000 21.605000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285000 18.660000 21.605000 18.980000 ;
      LAYER met4 ;
        RECT 21.285000 18.660000 21.605000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285000 19.090000 21.605000 19.410000 ;
      LAYER met4 ;
        RECT 21.285000 19.090000 21.605000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285000 19.520000 21.605000 19.840000 ;
      LAYER met4 ;
        RECT 21.285000 19.520000 21.605000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285000 19.950000 21.605000 20.270000 ;
      LAYER met4 ;
        RECT 21.285000 19.950000 21.605000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285000 20.380000 21.605000 20.700000 ;
      LAYER met4 ;
        RECT 21.285000 20.380000 21.605000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285000 20.810000 21.605000 21.130000 ;
      LAYER met4 ;
        RECT 21.285000 20.810000 21.605000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285000 21.240000 21.605000 21.560000 ;
      LAYER met4 ;
        RECT 21.285000 21.240000 21.605000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285000 21.670000 21.605000 21.990000 ;
      LAYER met4 ;
        RECT 21.285000 21.670000 21.605000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285000 22.100000 21.605000 22.420000 ;
      LAYER met4 ;
        RECT 21.285000 22.100000 21.605000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 68.065000 21.905000 68.385000 ;
      LAYER met4 ;
        RECT 21.585000 68.065000 21.905000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 68.475000 21.905000 68.795000 ;
      LAYER met4 ;
        RECT 21.585000 68.475000 21.905000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 68.885000 21.905000 69.205000 ;
      LAYER met4 ;
        RECT 21.585000 68.885000 21.905000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 69.295000 21.905000 69.615000 ;
      LAYER met4 ;
        RECT 21.585000 69.295000 21.905000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 69.705000 21.905000 70.025000 ;
      LAYER met4 ;
        RECT 21.585000 69.705000 21.905000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 70.115000 21.905000 70.435000 ;
      LAYER met4 ;
        RECT 21.585000 70.115000 21.905000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 70.525000 21.905000 70.845000 ;
      LAYER met4 ;
        RECT 21.585000 70.525000 21.905000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 70.935000 21.905000 71.255000 ;
      LAYER met4 ;
        RECT 21.585000 70.935000 21.905000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 71.345000 21.905000 71.665000 ;
      LAYER met4 ;
        RECT 21.585000 71.345000 21.905000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 71.755000 21.905000 72.075000 ;
      LAYER met4 ;
        RECT 21.585000 71.755000 21.905000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 72.165000 21.905000 72.485000 ;
      LAYER met4 ;
        RECT 21.585000 72.165000 21.905000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 72.575000 21.905000 72.895000 ;
      LAYER met4 ;
        RECT 21.585000 72.575000 21.905000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 72.985000 21.905000 73.305000 ;
      LAYER met4 ;
        RECT 21.585000 72.985000 21.905000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 73.390000 21.905000 73.710000 ;
      LAYER met4 ;
        RECT 21.585000 73.390000 21.905000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 73.795000 21.905000 74.115000 ;
      LAYER met4 ;
        RECT 21.585000 73.795000 21.905000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 74.200000 21.905000 74.520000 ;
      LAYER met4 ;
        RECT 21.585000 74.200000 21.905000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 74.605000 21.905000 74.925000 ;
      LAYER met4 ;
        RECT 21.585000 74.605000 21.905000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 75.010000 21.905000 75.330000 ;
      LAYER met4 ;
        RECT 21.585000 75.010000 21.905000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 75.415000 21.905000 75.735000 ;
      LAYER met4 ;
        RECT 21.585000 75.415000 21.905000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 75.820000 21.905000 76.140000 ;
      LAYER met4 ;
        RECT 21.585000 75.820000 21.905000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 76.225000 21.905000 76.545000 ;
      LAYER met4 ;
        RECT 21.585000 76.225000 21.905000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 76.630000 21.905000 76.950000 ;
      LAYER met4 ;
        RECT 21.585000 76.630000 21.905000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 77.035000 21.905000 77.355000 ;
      LAYER met4 ;
        RECT 21.585000 77.035000 21.905000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 77.440000 21.905000 77.760000 ;
      LAYER met4 ;
        RECT 21.585000 77.440000 21.905000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 77.845000 21.905000 78.165000 ;
      LAYER met4 ;
        RECT 21.585000 77.845000 21.905000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 78.250000 21.905000 78.570000 ;
      LAYER met4 ;
        RECT 21.585000 78.250000 21.905000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 78.655000 21.905000 78.975000 ;
      LAYER met4 ;
        RECT 21.585000 78.655000 21.905000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 79.060000 21.905000 79.380000 ;
      LAYER met4 ;
        RECT 21.585000 79.060000 21.905000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 79.465000 21.905000 79.785000 ;
      LAYER met4 ;
        RECT 21.585000 79.465000 21.905000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 79.870000 21.905000 80.190000 ;
      LAYER met4 ;
        RECT 21.585000 79.870000 21.905000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 80.275000 21.905000 80.595000 ;
      LAYER met4 ;
        RECT 21.585000 80.275000 21.905000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 80.680000 21.905000 81.000000 ;
      LAYER met4 ;
        RECT 21.585000 80.680000 21.905000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 81.085000 21.905000 81.405000 ;
      LAYER met4 ;
        RECT 21.585000 81.085000 21.905000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 81.490000 21.905000 81.810000 ;
      LAYER met4 ;
        RECT 21.585000 81.490000 21.905000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 81.895000 21.905000 82.215000 ;
      LAYER met4 ;
        RECT 21.585000 81.895000 21.905000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585000 82.300000 21.905000 82.620000 ;
      LAYER met4 ;
        RECT 21.585000 82.300000 21.905000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.655000 82.860000 21.975000 83.180000 ;
      LAYER met4 ;
        RECT 21.655000 82.860000 21.975000 83.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.655000 83.410000 21.975000 83.730000 ;
      LAYER met4 ;
        RECT 21.655000 83.410000 21.975000 83.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.655000 83.960000 21.975000 84.280000 ;
      LAYER met4 ;
        RECT 21.655000 83.960000 21.975000 84.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690000 17.800000 22.010000 18.120000 ;
      LAYER met4 ;
        RECT 21.690000 17.800000 22.010000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690000 18.230000 22.010000 18.550000 ;
      LAYER met4 ;
        RECT 21.690000 18.230000 22.010000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690000 18.660000 22.010000 18.980000 ;
      LAYER met4 ;
        RECT 21.690000 18.660000 22.010000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690000 19.090000 22.010000 19.410000 ;
      LAYER met4 ;
        RECT 21.690000 19.090000 22.010000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690000 19.520000 22.010000 19.840000 ;
      LAYER met4 ;
        RECT 21.690000 19.520000 22.010000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690000 19.950000 22.010000 20.270000 ;
      LAYER met4 ;
        RECT 21.690000 19.950000 22.010000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690000 20.380000 22.010000 20.700000 ;
      LAYER met4 ;
        RECT 21.690000 20.380000 22.010000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690000 20.810000 22.010000 21.130000 ;
      LAYER met4 ;
        RECT 21.690000 20.810000 22.010000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690000 21.240000 22.010000 21.560000 ;
      LAYER met4 ;
        RECT 21.690000 21.240000 22.010000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690000 21.670000 22.010000 21.990000 ;
      LAYER met4 ;
        RECT 21.690000 21.670000 22.010000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690000 22.100000 22.010000 22.420000 ;
      LAYER met4 ;
        RECT 21.690000 22.100000 22.010000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 68.065000 22.305000 68.385000 ;
      LAYER met4 ;
        RECT 21.985000 68.065000 22.305000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 68.475000 22.305000 68.795000 ;
      LAYER met4 ;
        RECT 21.985000 68.475000 22.305000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 68.885000 22.305000 69.205000 ;
      LAYER met4 ;
        RECT 21.985000 68.885000 22.305000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 69.295000 22.305000 69.615000 ;
      LAYER met4 ;
        RECT 21.985000 69.295000 22.305000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 69.705000 22.305000 70.025000 ;
      LAYER met4 ;
        RECT 21.985000 69.705000 22.305000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 70.115000 22.305000 70.435000 ;
      LAYER met4 ;
        RECT 21.985000 70.115000 22.305000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 70.525000 22.305000 70.845000 ;
      LAYER met4 ;
        RECT 21.985000 70.525000 22.305000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 70.935000 22.305000 71.255000 ;
      LAYER met4 ;
        RECT 21.985000 70.935000 22.305000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 71.345000 22.305000 71.665000 ;
      LAYER met4 ;
        RECT 21.985000 71.345000 22.305000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 71.755000 22.305000 72.075000 ;
      LAYER met4 ;
        RECT 21.985000 71.755000 22.305000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 72.165000 22.305000 72.485000 ;
      LAYER met4 ;
        RECT 21.985000 72.165000 22.305000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 72.575000 22.305000 72.895000 ;
      LAYER met4 ;
        RECT 21.985000 72.575000 22.305000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 72.985000 22.305000 73.305000 ;
      LAYER met4 ;
        RECT 21.985000 72.985000 22.305000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 73.390000 22.305000 73.710000 ;
      LAYER met4 ;
        RECT 21.985000 73.390000 22.305000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 73.795000 22.305000 74.115000 ;
      LAYER met4 ;
        RECT 21.985000 73.795000 22.305000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 74.200000 22.305000 74.520000 ;
      LAYER met4 ;
        RECT 21.985000 74.200000 22.305000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 74.605000 22.305000 74.925000 ;
      LAYER met4 ;
        RECT 21.985000 74.605000 22.305000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 75.010000 22.305000 75.330000 ;
      LAYER met4 ;
        RECT 21.985000 75.010000 22.305000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 75.415000 22.305000 75.735000 ;
      LAYER met4 ;
        RECT 21.985000 75.415000 22.305000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 75.820000 22.305000 76.140000 ;
      LAYER met4 ;
        RECT 21.985000 75.820000 22.305000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 76.225000 22.305000 76.545000 ;
      LAYER met4 ;
        RECT 21.985000 76.225000 22.305000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 76.630000 22.305000 76.950000 ;
      LAYER met4 ;
        RECT 21.985000 76.630000 22.305000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 77.035000 22.305000 77.355000 ;
      LAYER met4 ;
        RECT 21.985000 77.035000 22.305000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 77.440000 22.305000 77.760000 ;
      LAYER met4 ;
        RECT 21.985000 77.440000 22.305000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 77.845000 22.305000 78.165000 ;
      LAYER met4 ;
        RECT 21.985000 77.845000 22.305000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 78.250000 22.305000 78.570000 ;
      LAYER met4 ;
        RECT 21.985000 78.250000 22.305000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 78.655000 22.305000 78.975000 ;
      LAYER met4 ;
        RECT 21.985000 78.655000 22.305000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 79.060000 22.305000 79.380000 ;
      LAYER met4 ;
        RECT 21.985000 79.060000 22.305000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 79.465000 22.305000 79.785000 ;
      LAYER met4 ;
        RECT 21.985000 79.465000 22.305000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 79.870000 22.305000 80.190000 ;
      LAYER met4 ;
        RECT 21.985000 79.870000 22.305000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 80.275000 22.305000 80.595000 ;
      LAYER met4 ;
        RECT 21.985000 80.275000 22.305000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 80.680000 22.305000 81.000000 ;
      LAYER met4 ;
        RECT 21.985000 80.680000 22.305000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 81.085000 22.305000 81.405000 ;
      LAYER met4 ;
        RECT 21.985000 81.085000 22.305000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 81.490000 22.305000 81.810000 ;
      LAYER met4 ;
        RECT 21.985000 81.490000 22.305000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 81.895000 22.305000 82.215000 ;
      LAYER met4 ;
        RECT 21.985000 81.895000 22.305000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985000 82.300000 22.305000 82.620000 ;
      LAYER met4 ;
        RECT 21.985000 82.300000 22.305000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100000 17.800000 22.420000 18.120000 ;
      LAYER met4 ;
        RECT 22.100000 17.800000 22.420000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100000 18.230000 22.420000 18.550000 ;
      LAYER met4 ;
        RECT 22.100000 18.230000 22.420000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100000 18.660000 22.420000 18.980000 ;
      LAYER met4 ;
        RECT 22.100000 18.660000 22.420000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100000 19.090000 22.420000 19.410000 ;
      LAYER met4 ;
        RECT 22.100000 19.090000 22.420000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100000 19.520000 22.420000 19.840000 ;
      LAYER met4 ;
        RECT 22.100000 19.520000 22.420000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100000 19.950000 22.420000 20.270000 ;
      LAYER met4 ;
        RECT 22.100000 19.950000 22.420000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100000 20.380000 22.420000 20.700000 ;
      LAYER met4 ;
        RECT 22.100000 20.380000 22.420000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100000 20.810000 22.420000 21.130000 ;
      LAYER met4 ;
        RECT 22.100000 20.810000 22.420000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100000 21.240000 22.420000 21.560000 ;
      LAYER met4 ;
        RECT 22.100000 21.240000 22.420000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100000 21.670000 22.420000 21.990000 ;
      LAYER met4 ;
        RECT 22.100000 21.670000 22.420000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100000 22.100000 22.420000 22.420000 ;
      LAYER met4 ;
        RECT 22.100000 22.100000 22.420000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 68.065000 22.705000 68.385000 ;
      LAYER met4 ;
        RECT 22.385000 68.065000 22.705000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 68.475000 22.705000 68.795000 ;
      LAYER met4 ;
        RECT 22.385000 68.475000 22.705000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 68.885000 22.705000 69.205000 ;
      LAYER met4 ;
        RECT 22.385000 68.885000 22.705000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 69.295000 22.705000 69.615000 ;
      LAYER met4 ;
        RECT 22.385000 69.295000 22.705000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 69.705000 22.705000 70.025000 ;
      LAYER met4 ;
        RECT 22.385000 69.705000 22.705000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 70.115000 22.705000 70.435000 ;
      LAYER met4 ;
        RECT 22.385000 70.115000 22.705000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 70.525000 22.705000 70.845000 ;
      LAYER met4 ;
        RECT 22.385000 70.525000 22.705000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 70.935000 22.705000 71.255000 ;
      LAYER met4 ;
        RECT 22.385000 70.935000 22.705000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 71.345000 22.705000 71.665000 ;
      LAYER met4 ;
        RECT 22.385000 71.345000 22.705000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 71.755000 22.705000 72.075000 ;
      LAYER met4 ;
        RECT 22.385000 71.755000 22.705000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 72.165000 22.705000 72.485000 ;
      LAYER met4 ;
        RECT 22.385000 72.165000 22.705000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 72.575000 22.705000 72.895000 ;
      LAYER met4 ;
        RECT 22.385000 72.575000 22.705000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 72.985000 22.705000 73.305000 ;
      LAYER met4 ;
        RECT 22.385000 72.985000 22.705000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 73.390000 22.705000 73.710000 ;
      LAYER met4 ;
        RECT 22.385000 73.390000 22.705000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 73.795000 22.705000 74.115000 ;
      LAYER met4 ;
        RECT 22.385000 73.795000 22.705000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 74.200000 22.705000 74.520000 ;
      LAYER met4 ;
        RECT 22.385000 74.200000 22.705000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 74.605000 22.705000 74.925000 ;
      LAYER met4 ;
        RECT 22.385000 74.605000 22.705000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 75.010000 22.705000 75.330000 ;
      LAYER met4 ;
        RECT 22.385000 75.010000 22.705000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 75.415000 22.705000 75.735000 ;
      LAYER met4 ;
        RECT 22.385000 75.415000 22.705000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 75.820000 22.705000 76.140000 ;
      LAYER met4 ;
        RECT 22.385000 75.820000 22.705000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 76.225000 22.705000 76.545000 ;
      LAYER met4 ;
        RECT 22.385000 76.225000 22.705000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 76.630000 22.705000 76.950000 ;
      LAYER met4 ;
        RECT 22.385000 76.630000 22.705000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 77.035000 22.705000 77.355000 ;
      LAYER met4 ;
        RECT 22.385000 77.035000 22.705000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 77.440000 22.705000 77.760000 ;
      LAYER met4 ;
        RECT 22.385000 77.440000 22.705000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 77.845000 22.705000 78.165000 ;
      LAYER met4 ;
        RECT 22.385000 77.845000 22.705000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 78.250000 22.705000 78.570000 ;
      LAYER met4 ;
        RECT 22.385000 78.250000 22.705000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 78.655000 22.705000 78.975000 ;
      LAYER met4 ;
        RECT 22.385000 78.655000 22.705000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 79.060000 22.705000 79.380000 ;
      LAYER met4 ;
        RECT 22.385000 79.060000 22.705000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 79.465000 22.705000 79.785000 ;
      LAYER met4 ;
        RECT 22.385000 79.465000 22.705000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 79.870000 22.705000 80.190000 ;
      LAYER met4 ;
        RECT 22.385000 79.870000 22.705000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 80.275000 22.705000 80.595000 ;
      LAYER met4 ;
        RECT 22.385000 80.275000 22.705000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 80.680000 22.705000 81.000000 ;
      LAYER met4 ;
        RECT 22.385000 80.680000 22.705000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 81.085000 22.705000 81.405000 ;
      LAYER met4 ;
        RECT 22.385000 81.085000 22.705000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 81.490000 22.705000 81.810000 ;
      LAYER met4 ;
        RECT 22.385000 81.490000 22.705000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 81.895000 22.705000 82.215000 ;
      LAYER met4 ;
        RECT 22.385000 81.895000 22.705000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385000 82.300000 22.705000 82.620000 ;
      LAYER met4 ;
        RECT 22.385000 82.300000 22.705000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445000 82.860000 22.765000 83.180000 ;
      LAYER met4 ;
        RECT 22.445000 82.860000 22.765000 83.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445000 83.410000 22.765000 83.730000 ;
      LAYER met4 ;
        RECT 22.445000 83.410000 22.765000 83.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445000 83.960000 22.765000 84.280000 ;
      LAYER met4 ;
        RECT 22.445000 83.960000 22.765000 84.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510000 17.800000 22.830000 18.120000 ;
      LAYER met4 ;
        RECT 22.510000 17.800000 22.830000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510000 18.230000 22.830000 18.550000 ;
      LAYER met4 ;
        RECT 22.510000 18.230000 22.830000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510000 18.660000 22.830000 18.980000 ;
      LAYER met4 ;
        RECT 22.510000 18.660000 22.830000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510000 19.090000 22.830000 19.410000 ;
      LAYER met4 ;
        RECT 22.510000 19.090000 22.830000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510000 19.520000 22.830000 19.840000 ;
      LAYER met4 ;
        RECT 22.510000 19.520000 22.830000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510000 19.950000 22.830000 20.270000 ;
      LAYER met4 ;
        RECT 22.510000 19.950000 22.830000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510000 20.380000 22.830000 20.700000 ;
      LAYER met4 ;
        RECT 22.510000 20.380000 22.830000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510000 20.810000 22.830000 21.130000 ;
      LAYER met4 ;
        RECT 22.510000 20.810000 22.830000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510000 21.240000 22.830000 21.560000 ;
      LAYER met4 ;
        RECT 22.510000 21.240000 22.830000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510000 21.670000 22.830000 21.990000 ;
      LAYER met4 ;
        RECT 22.510000 21.670000 22.830000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510000 22.100000 22.830000 22.420000 ;
      LAYER met4 ;
        RECT 22.510000 22.100000 22.830000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 68.065000 23.105000 68.385000 ;
      LAYER met4 ;
        RECT 22.785000 68.065000 23.105000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 68.475000 23.105000 68.795000 ;
      LAYER met4 ;
        RECT 22.785000 68.475000 23.105000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 68.885000 23.105000 69.205000 ;
      LAYER met4 ;
        RECT 22.785000 68.885000 23.105000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 69.295000 23.105000 69.615000 ;
      LAYER met4 ;
        RECT 22.785000 69.295000 23.105000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 69.705000 23.105000 70.025000 ;
      LAYER met4 ;
        RECT 22.785000 69.705000 23.105000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 70.115000 23.105000 70.435000 ;
      LAYER met4 ;
        RECT 22.785000 70.115000 23.105000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 70.525000 23.105000 70.845000 ;
      LAYER met4 ;
        RECT 22.785000 70.525000 23.105000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 70.935000 23.105000 71.255000 ;
      LAYER met4 ;
        RECT 22.785000 70.935000 23.105000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 71.345000 23.105000 71.665000 ;
      LAYER met4 ;
        RECT 22.785000 71.345000 23.105000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 71.755000 23.105000 72.075000 ;
      LAYER met4 ;
        RECT 22.785000 71.755000 23.105000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 72.165000 23.105000 72.485000 ;
      LAYER met4 ;
        RECT 22.785000 72.165000 23.105000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 72.575000 23.105000 72.895000 ;
      LAYER met4 ;
        RECT 22.785000 72.575000 23.105000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 72.985000 23.105000 73.305000 ;
      LAYER met4 ;
        RECT 22.785000 72.985000 23.105000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 73.390000 23.105000 73.710000 ;
      LAYER met4 ;
        RECT 22.785000 73.390000 23.105000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 73.795000 23.105000 74.115000 ;
      LAYER met4 ;
        RECT 22.785000 73.795000 23.105000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 74.200000 23.105000 74.520000 ;
      LAYER met4 ;
        RECT 22.785000 74.200000 23.105000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 74.605000 23.105000 74.925000 ;
      LAYER met4 ;
        RECT 22.785000 74.605000 23.105000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 75.010000 23.105000 75.330000 ;
      LAYER met4 ;
        RECT 22.785000 75.010000 23.105000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 75.415000 23.105000 75.735000 ;
      LAYER met4 ;
        RECT 22.785000 75.415000 23.105000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 75.820000 23.105000 76.140000 ;
      LAYER met4 ;
        RECT 22.785000 75.820000 23.105000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 76.225000 23.105000 76.545000 ;
      LAYER met4 ;
        RECT 22.785000 76.225000 23.105000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 76.630000 23.105000 76.950000 ;
      LAYER met4 ;
        RECT 22.785000 76.630000 23.105000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 77.035000 23.105000 77.355000 ;
      LAYER met4 ;
        RECT 22.785000 77.035000 23.105000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 77.440000 23.105000 77.760000 ;
      LAYER met4 ;
        RECT 22.785000 77.440000 23.105000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 77.845000 23.105000 78.165000 ;
      LAYER met4 ;
        RECT 22.785000 77.845000 23.105000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 78.250000 23.105000 78.570000 ;
      LAYER met4 ;
        RECT 22.785000 78.250000 23.105000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 78.655000 23.105000 78.975000 ;
      LAYER met4 ;
        RECT 22.785000 78.655000 23.105000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 79.060000 23.105000 79.380000 ;
      LAYER met4 ;
        RECT 22.785000 79.060000 23.105000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 79.465000 23.105000 79.785000 ;
      LAYER met4 ;
        RECT 22.785000 79.465000 23.105000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 79.870000 23.105000 80.190000 ;
      LAYER met4 ;
        RECT 22.785000 79.870000 23.105000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 80.275000 23.105000 80.595000 ;
      LAYER met4 ;
        RECT 22.785000 80.275000 23.105000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 80.680000 23.105000 81.000000 ;
      LAYER met4 ;
        RECT 22.785000 80.680000 23.105000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 81.085000 23.105000 81.405000 ;
      LAYER met4 ;
        RECT 22.785000 81.085000 23.105000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 81.490000 23.105000 81.810000 ;
      LAYER met4 ;
        RECT 22.785000 81.490000 23.105000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 81.895000 23.105000 82.215000 ;
      LAYER met4 ;
        RECT 22.785000 81.895000 23.105000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785000 82.300000 23.105000 82.620000 ;
      LAYER met4 ;
        RECT 22.785000 82.300000 23.105000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920000 17.800000 23.240000 18.120000 ;
      LAYER met4 ;
        RECT 22.920000 17.800000 23.240000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920000 18.230000 23.240000 18.550000 ;
      LAYER met4 ;
        RECT 22.920000 18.230000 23.240000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920000 18.660000 23.240000 18.980000 ;
      LAYER met4 ;
        RECT 22.920000 18.660000 23.240000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920000 19.090000 23.240000 19.410000 ;
      LAYER met4 ;
        RECT 22.920000 19.090000 23.240000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920000 19.520000 23.240000 19.840000 ;
      LAYER met4 ;
        RECT 22.920000 19.520000 23.240000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920000 19.950000 23.240000 20.270000 ;
      LAYER met4 ;
        RECT 22.920000 19.950000 23.240000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920000 20.380000 23.240000 20.700000 ;
      LAYER met4 ;
        RECT 22.920000 20.380000 23.240000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920000 20.810000 23.240000 21.130000 ;
      LAYER met4 ;
        RECT 22.920000 20.810000 23.240000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920000 21.240000 23.240000 21.560000 ;
      LAYER met4 ;
        RECT 22.920000 21.240000 23.240000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920000 21.670000 23.240000 21.990000 ;
      LAYER met4 ;
        RECT 22.920000 21.670000 23.240000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920000 22.100000 23.240000 22.420000 ;
      LAYER met4 ;
        RECT 22.920000 22.100000 23.240000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 68.065000 23.505000 68.385000 ;
      LAYER met4 ;
        RECT 23.185000 68.065000 23.505000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 68.475000 23.505000 68.795000 ;
      LAYER met4 ;
        RECT 23.185000 68.475000 23.505000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 68.885000 23.505000 69.205000 ;
      LAYER met4 ;
        RECT 23.185000 68.885000 23.505000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 69.295000 23.505000 69.615000 ;
      LAYER met4 ;
        RECT 23.185000 69.295000 23.505000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 69.705000 23.505000 70.025000 ;
      LAYER met4 ;
        RECT 23.185000 69.705000 23.505000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 70.115000 23.505000 70.435000 ;
      LAYER met4 ;
        RECT 23.185000 70.115000 23.505000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 70.525000 23.505000 70.845000 ;
      LAYER met4 ;
        RECT 23.185000 70.525000 23.505000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 70.935000 23.505000 71.255000 ;
      LAYER met4 ;
        RECT 23.185000 70.935000 23.505000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 71.345000 23.505000 71.665000 ;
      LAYER met4 ;
        RECT 23.185000 71.345000 23.505000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 71.755000 23.505000 72.075000 ;
      LAYER met4 ;
        RECT 23.185000 71.755000 23.505000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 72.165000 23.505000 72.485000 ;
      LAYER met4 ;
        RECT 23.185000 72.165000 23.505000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 72.575000 23.505000 72.895000 ;
      LAYER met4 ;
        RECT 23.185000 72.575000 23.505000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 72.985000 23.505000 73.305000 ;
      LAYER met4 ;
        RECT 23.185000 72.985000 23.505000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 73.390000 23.505000 73.710000 ;
      LAYER met4 ;
        RECT 23.185000 73.390000 23.505000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 73.795000 23.505000 74.115000 ;
      LAYER met4 ;
        RECT 23.185000 73.795000 23.505000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 74.200000 23.505000 74.520000 ;
      LAYER met4 ;
        RECT 23.185000 74.200000 23.505000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 74.605000 23.505000 74.925000 ;
      LAYER met4 ;
        RECT 23.185000 74.605000 23.505000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 75.010000 23.505000 75.330000 ;
      LAYER met4 ;
        RECT 23.185000 75.010000 23.505000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 75.415000 23.505000 75.735000 ;
      LAYER met4 ;
        RECT 23.185000 75.415000 23.505000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 75.820000 23.505000 76.140000 ;
      LAYER met4 ;
        RECT 23.185000 75.820000 23.505000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 76.225000 23.505000 76.545000 ;
      LAYER met4 ;
        RECT 23.185000 76.225000 23.505000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 76.630000 23.505000 76.950000 ;
      LAYER met4 ;
        RECT 23.185000 76.630000 23.505000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 77.035000 23.505000 77.355000 ;
      LAYER met4 ;
        RECT 23.185000 77.035000 23.505000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 77.440000 23.505000 77.760000 ;
      LAYER met4 ;
        RECT 23.185000 77.440000 23.505000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 77.845000 23.505000 78.165000 ;
      LAYER met4 ;
        RECT 23.185000 77.845000 23.505000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 78.250000 23.505000 78.570000 ;
      LAYER met4 ;
        RECT 23.185000 78.250000 23.505000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 78.655000 23.505000 78.975000 ;
      LAYER met4 ;
        RECT 23.185000 78.655000 23.505000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 79.060000 23.505000 79.380000 ;
      LAYER met4 ;
        RECT 23.185000 79.060000 23.505000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 79.465000 23.505000 79.785000 ;
      LAYER met4 ;
        RECT 23.185000 79.465000 23.505000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 79.870000 23.505000 80.190000 ;
      LAYER met4 ;
        RECT 23.185000 79.870000 23.505000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 80.275000 23.505000 80.595000 ;
      LAYER met4 ;
        RECT 23.185000 80.275000 23.505000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 80.680000 23.505000 81.000000 ;
      LAYER met4 ;
        RECT 23.185000 80.680000 23.505000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 81.085000 23.505000 81.405000 ;
      LAYER met4 ;
        RECT 23.185000 81.085000 23.505000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 81.490000 23.505000 81.810000 ;
      LAYER met4 ;
        RECT 23.185000 81.490000 23.505000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 81.895000 23.505000 82.215000 ;
      LAYER met4 ;
        RECT 23.185000 81.895000 23.505000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185000 82.300000 23.505000 82.620000 ;
      LAYER met4 ;
        RECT 23.185000 82.300000 23.505000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330000 17.800000 23.650000 18.120000 ;
      LAYER met4 ;
        RECT 23.330000 17.800000 23.650000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330000 18.230000 23.650000 18.550000 ;
      LAYER met4 ;
        RECT 23.330000 18.230000 23.650000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330000 18.660000 23.650000 18.980000 ;
      LAYER met4 ;
        RECT 23.330000 18.660000 23.650000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330000 19.090000 23.650000 19.410000 ;
      LAYER met4 ;
        RECT 23.330000 19.090000 23.650000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330000 19.520000 23.650000 19.840000 ;
      LAYER met4 ;
        RECT 23.330000 19.520000 23.650000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330000 19.950000 23.650000 20.270000 ;
      LAYER met4 ;
        RECT 23.330000 19.950000 23.650000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330000 20.380000 23.650000 20.700000 ;
      LAYER met4 ;
        RECT 23.330000 20.380000 23.650000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330000 20.810000 23.650000 21.130000 ;
      LAYER met4 ;
        RECT 23.330000 20.810000 23.650000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330000 21.240000 23.650000 21.560000 ;
      LAYER met4 ;
        RECT 23.330000 21.240000 23.650000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330000 21.670000 23.650000 21.990000 ;
      LAYER met4 ;
        RECT 23.330000 21.670000 23.650000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330000 22.100000 23.650000 22.420000 ;
      LAYER met4 ;
        RECT 23.330000 22.100000 23.650000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 68.065000 23.905000 68.385000 ;
      LAYER met4 ;
        RECT 23.585000 68.065000 23.905000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 68.475000 23.905000 68.795000 ;
      LAYER met4 ;
        RECT 23.585000 68.475000 23.905000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 68.885000 23.905000 69.205000 ;
      LAYER met4 ;
        RECT 23.585000 68.885000 23.905000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 69.295000 23.905000 69.615000 ;
      LAYER met4 ;
        RECT 23.585000 69.295000 23.905000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 69.705000 23.905000 70.025000 ;
      LAYER met4 ;
        RECT 23.585000 69.705000 23.905000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 70.115000 23.905000 70.435000 ;
      LAYER met4 ;
        RECT 23.585000 70.115000 23.905000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 70.525000 23.905000 70.845000 ;
      LAYER met4 ;
        RECT 23.585000 70.525000 23.905000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 70.935000 23.905000 71.255000 ;
      LAYER met4 ;
        RECT 23.585000 70.935000 23.905000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 71.345000 23.905000 71.665000 ;
      LAYER met4 ;
        RECT 23.585000 71.345000 23.905000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 71.755000 23.905000 72.075000 ;
      LAYER met4 ;
        RECT 23.585000 71.755000 23.905000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 72.165000 23.905000 72.485000 ;
      LAYER met4 ;
        RECT 23.585000 72.165000 23.905000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 72.575000 23.905000 72.895000 ;
      LAYER met4 ;
        RECT 23.585000 72.575000 23.905000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 72.985000 23.905000 73.305000 ;
      LAYER met4 ;
        RECT 23.585000 72.985000 23.905000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 73.390000 23.905000 73.710000 ;
      LAYER met4 ;
        RECT 23.585000 73.390000 23.905000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 73.795000 23.905000 74.115000 ;
      LAYER met4 ;
        RECT 23.585000 73.795000 23.905000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 74.200000 23.905000 74.520000 ;
      LAYER met4 ;
        RECT 23.585000 74.200000 23.905000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 74.605000 23.905000 74.925000 ;
      LAYER met4 ;
        RECT 23.585000 74.605000 23.905000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 75.010000 23.905000 75.330000 ;
      LAYER met4 ;
        RECT 23.585000 75.010000 23.905000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 75.415000 23.905000 75.735000 ;
      LAYER met4 ;
        RECT 23.585000 75.415000 23.905000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 75.820000 23.905000 76.140000 ;
      LAYER met4 ;
        RECT 23.585000 75.820000 23.905000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 76.225000 23.905000 76.545000 ;
      LAYER met4 ;
        RECT 23.585000 76.225000 23.905000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 76.630000 23.905000 76.950000 ;
      LAYER met4 ;
        RECT 23.585000 76.630000 23.905000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 77.035000 23.905000 77.355000 ;
      LAYER met4 ;
        RECT 23.585000 77.035000 23.905000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 77.440000 23.905000 77.760000 ;
      LAYER met4 ;
        RECT 23.585000 77.440000 23.905000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 77.845000 23.905000 78.165000 ;
      LAYER met4 ;
        RECT 23.585000 77.845000 23.905000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 78.250000 23.905000 78.570000 ;
      LAYER met4 ;
        RECT 23.585000 78.250000 23.905000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 78.655000 23.905000 78.975000 ;
      LAYER met4 ;
        RECT 23.585000 78.655000 23.905000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 79.060000 23.905000 79.380000 ;
      LAYER met4 ;
        RECT 23.585000 79.060000 23.905000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 79.465000 23.905000 79.785000 ;
      LAYER met4 ;
        RECT 23.585000 79.465000 23.905000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 79.870000 23.905000 80.190000 ;
      LAYER met4 ;
        RECT 23.585000 79.870000 23.905000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 80.275000 23.905000 80.595000 ;
      LAYER met4 ;
        RECT 23.585000 80.275000 23.905000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 80.680000 23.905000 81.000000 ;
      LAYER met4 ;
        RECT 23.585000 80.680000 23.905000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 81.085000 23.905000 81.405000 ;
      LAYER met4 ;
        RECT 23.585000 81.085000 23.905000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 81.490000 23.905000 81.810000 ;
      LAYER met4 ;
        RECT 23.585000 81.490000 23.905000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 81.895000 23.905000 82.215000 ;
      LAYER met4 ;
        RECT 23.585000 81.895000 23.905000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585000 82.300000 23.905000 82.620000 ;
      LAYER met4 ;
        RECT 23.585000 82.300000 23.905000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740000 17.800000 24.060000 18.120000 ;
      LAYER met4 ;
        RECT 23.740000 17.800000 24.060000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740000 18.230000 24.060000 18.550000 ;
      LAYER met4 ;
        RECT 23.740000 18.230000 24.060000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740000 18.660000 24.060000 18.980000 ;
      LAYER met4 ;
        RECT 23.740000 18.660000 24.060000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740000 19.090000 24.060000 19.410000 ;
      LAYER met4 ;
        RECT 23.740000 19.090000 24.060000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740000 19.520000 24.060000 19.840000 ;
      LAYER met4 ;
        RECT 23.740000 19.520000 24.060000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740000 19.950000 24.060000 20.270000 ;
      LAYER met4 ;
        RECT 23.740000 19.950000 24.060000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740000 20.380000 24.060000 20.700000 ;
      LAYER met4 ;
        RECT 23.740000 20.380000 24.060000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740000 20.810000 24.060000 21.130000 ;
      LAYER met4 ;
        RECT 23.740000 20.810000 24.060000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740000 21.240000 24.060000 21.560000 ;
      LAYER met4 ;
        RECT 23.740000 21.240000 24.060000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740000 21.670000 24.060000 21.990000 ;
      LAYER met4 ;
        RECT 23.740000 21.670000 24.060000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740000 22.100000 24.060000 22.420000 ;
      LAYER met4 ;
        RECT 23.740000 22.100000 24.060000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 68.065000 24.305000 68.385000 ;
      LAYER met4 ;
        RECT 23.985000 68.065000 24.305000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 68.475000 24.305000 68.795000 ;
      LAYER met4 ;
        RECT 23.985000 68.475000 24.305000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 68.885000 24.305000 69.205000 ;
      LAYER met4 ;
        RECT 23.985000 68.885000 24.305000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 69.295000 24.305000 69.615000 ;
      LAYER met4 ;
        RECT 23.985000 69.295000 24.305000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 69.705000 24.305000 70.025000 ;
      LAYER met4 ;
        RECT 23.985000 69.705000 24.305000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 70.115000 24.305000 70.435000 ;
      LAYER met4 ;
        RECT 23.985000 70.115000 24.305000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 70.525000 24.305000 70.845000 ;
      LAYER met4 ;
        RECT 23.985000 70.525000 24.305000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 70.935000 24.305000 71.255000 ;
      LAYER met4 ;
        RECT 23.985000 70.935000 24.305000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 71.345000 24.305000 71.665000 ;
      LAYER met4 ;
        RECT 23.985000 71.345000 24.305000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 71.755000 24.305000 72.075000 ;
      LAYER met4 ;
        RECT 23.985000 71.755000 24.305000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 72.165000 24.305000 72.485000 ;
      LAYER met4 ;
        RECT 23.985000 72.165000 24.305000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 72.575000 24.305000 72.895000 ;
      LAYER met4 ;
        RECT 23.985000 72.575000 24.305000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 72.985000 24.305000 73.305000 ;
      LAYER met4 ;
        RECT 23.985000 72.985000 24.305000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 73.390000 24.305000 73.710000 ;
      LAYER met4 ;
        RECT 23.985000 73.390000 24.305000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 73.795000 24.305000 74.115000 ;
      LAYER met4 ;
        RECT 23.985000 73.795000 24.305000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 74.200000 24.305000 74.520000 ;
      LAYER met4 ;
        RECT 23.985000 74.200000 24.305000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 74.605000 24.305000 74.925000 ;
      LAYER met4 ;
        RECT 23.985000 74.605000 24.305000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 75.010000 24.305000 75.330000 ;
      LAYER met4 ;
        RECT 23.985000 75.010000 24.305000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 75.415000 24.305000 75.735000 ;
      LAYER met4 ;
        RECT 23.985000 75.415000 24.305000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 75.820000 24.305000 76.140000 ;
      LAYER met4 ;
        RECT 23.985000 75.820000 24.305000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 76.225000 24.305000 76.545000 ;
      LAYER met4 ;
        RECT 23.985000 76.225000 24.305000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 76.630000 24.305000 76.950000 ;
      LAYER met4 ;
        RECT 23.985000 76.630000 24.305000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 77.035000 24.305000 77.355000 ;
      LAYER met4 ;
        RECT 23.985000 77.035000 24.305000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 77.440000 24.305000 77.760000 ;
      LAYER met4 ;
        RECT 23.985000 77.440000 24.305000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 77.845000 24.305000 78.165000 ;
      LAYER met4 ;
        RECT 23.985000 77.845000 24.305000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 78.250000 24.305000 78.570000 ;
      LAYER met4 ;
        RECT 23.985000 78.250000 24.305000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 78.655000 24.305000 78.975000 ;
      LAYER met4 ;
        RECT 23.985000 78.655000 24.305000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 79.060000 24.305000 79.380000 ;
      LAYER met4 ;
        RECT 23.985000 79.060000 24.305000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 79.465000 24.305000 79.785000 ;
      LAYER met4 ;
        RECT 23.985000 79.465000 24.305000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 79.870000 24.305000 80.190000 ;
      LAYER met4 ;
        RECT 23.985000 79.870000 24.305000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 80.275000 24.305000 80.595000 ;
      LAYER met4 ;
        RECT 23.985000 80.275000 24.305000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 80.680000 24.305000 81.000000 ;
      LAYER met4 ;
        RECT 23.985000 80.680000 24.305000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 81.085000 24.305000 81.405000 ;
      LAYER met4 ;
        RECT 23.985000 81.085000 24.305000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 81.490000 24.305000 81.810000 ;
      LAYER met4 ;
        RECT 23.985000 81.490000 24.305000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 81.895000 24.305000 82.215000 ;
      LAYER met4 ;
        RECT 23.985000 81.895000 24.305000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985000 82.300000 24.305000 82.620000 ;
      LAYER met4 ;
        RECT 23.985000 82.300000 24.305000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 17.800000 24.470000 18.120000 ;
      LAYER met4 ;
        RECT 24.150000 17.800000 24.470000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 18.230000 24.470000 18.550000 ;
      LAYER met4 ;
        RECT 24.150000 18.230000 24.470000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 18.660000 24.470000 18.980000 ;
      LAYER met4 ;
        RECT 24.150000 18.660000 24.470000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 19.090000 24.470000 19.410000 ;
      LAYER met4 ;
        RECT 24.150000 19.090000 24.470000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 19.520000 24.470000 19.840000 ;
      LAYER met4 ;
        RECT 24.150000 19.520000 24.470000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 19.950000 24.470000 20.270000 ;
      LAYER met4 ;
        RECT 24.150000 19.950000 24.470000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 20.380000 24.470000 20.700000 ;
      LAYER met4 ;
        RECT 24.150000 20.380000 24.470000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 20.810000 24.470000 21.130000 ;
      LAYER met4 ;
        RECT 24.150000 20.810000 24.470000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 21.240000 24.470000 21.560000 ;
      LAYER met4 ;
        RECT 24.150000 21.240000 24.470000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 21.670000 24.470000 21.990000 ;
      LAYER met4 ;
        RECT 24.150000 21.670000 24.470000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 22.100000 24.470000 22.420000 ;
      LAYER met4 ;
        RECT 24.150000 22.100000 24.470000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060000 17.800000 3.380000 18.120000 ;
      LAYER met4 ;
        RECT 3.060000 17.800000 3.380000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060000 18.230000 3.380000 18.550000 ;
      LAYER met4 ;
        RECT 3.060000 18.230000 3.380000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060000 18.660000 3.380000 18.980000 ;
      LAYER met4 ;
        RECT 3.060000 18.660000 3.380000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060000 19.090000 3.380000 19.410000 ;
      LAYER met4 ;
        RECT 3.060000 19.090000 3.380000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060000 19.520000 3.380000 19.840000 ;
      LAYER met4 ;
        RECT 3.060000 19.520000 3.380000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060000 19.950000 3.380000 20.270000 ;
      LAYER met4 ;
        RECT 3.060000 19.950000 3.380000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060000 20.380000 3.380000 20.700000 ;
      LAYER met4 ;
        RECT 3.060000 20.380000 3.380000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060000 20.810000 3.380000 21.130000 ;
      LAYER met4 ;
        RECT 3.060000 20.810000 3.380000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060000 21.240000 3.380000 21.560000 ;
      LAYER met4 ;
        RECT 3.060000 21.240000 3.380000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060000 21.670000 3.380000 21.990000 ;
      LAYER met4 ;
        RECT 3.060000 21.670000 3.380000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060000 22.100000 3.380000 22.420000 ;
      LAYER met4 ;
        RECT 3.060000 22.100000 3.380000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 82.795000 3.455000 83.115000 ;
      LAYER met4 ;
        RECT 3.135000 82.795000 3.455000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 83.205000 3.455000 83.525000 ;
      LAYER met4 ;
        RECT 3.135000 83.205000 3.455000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 83.615000 3.455000 83.935000 ;
      LAYER met4 ;
        RECT 3.135000 83.615000 3.455000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 84.025000 3.455000 84.345000 ;
      LAYER met4 ;
        RECT 3.135000 84.025000 3.455000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 84.435000 3.455000 84.755000 ;
      LAYER met4 ;
        RECT 3.135000 84.435000 3.455000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 84.845000 3.455000 85.165000 ;
      LAYER met4 ;
        RECT 3.135000 84.845000 3.455000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 85.255000 3.455000 85.575000 ;
      LAYER met4 ;
        RECT 3.135000 85.255000 3.455000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 85.665000 3.455000 85.985000 ;
      LAYER met4 ;
        RECT 3.135000 85.665000 3.455000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 86.075000 3.455000 86.395000 ;
      LAYER met4 ;
        RECT 3.135000 86.075000 3.455000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 86.485000 3.455000 86.805000 ;
      LAYER met4 ;
        RECT 3.135000 86.485000 3.455000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 86.895000 3.455000 87.215000 ;
      LAYER met4 ;
        RECT 3.135000 86.895000 3.455000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 87.305000 3.455000 87.625000 ;
      LAYER met4 ;
        RECT 3.135000 87.305000 3.455000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 87.715000 3.455000 88.035000 ;
      LAYER met4 ;
        RECT 3.135000 87.715000 3.455000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 88.125000 3.455000 88.445000 ;
      LAYER met4 ;
        RECT 3.135000 88.125000 3.455000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 88.535000 3.455000 88.855000 ;
      LAYER met4 ;
        RECT 3.135000 88.535000 3.455000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 88.945000 3.455000 89.265000 ;
      LAYER met4 ;
        RECT 3.135000 88.945000 3.455000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 89.355000 3.455000 89.675000 ;
      LAYER met4 ;
        RECT 3.135000 89.355000 3.455000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 89.765000 3.455000 90.085000 ;
      LAYER met4 ;
        RECT 3.135000 89.765000 3.455000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 90.175000 3.455000 90.495000 ;
      LAYER met4 ;
        RECT 3.135000 90.175000 3.455000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 90.585000 3.455000 90.905000 ;
      LAYER met4 ;
        RECT 3.135000 90.585000 3.455000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 90.995000 3.455000 91.315000 ;
      LAYER met4 ;
        RECT 3.135000 90.995000 3.455000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 91.405000 3.455000 91.725000 ;
      LAYER met4 ;
        RECT 3.135000 91.405000 3.455000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 91.815000 3.455000 92.135000 ;
      LAYER met4 ;
        RECT 3.135000 91.815000 3.455000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 92.225000 3.455000 92.545000 ;
      LAYER met4 ;
        RECT 3.135000 92.225000 3.455000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135000 92.635000 3.455000 92.955000 ;
      LAYER met4 ;
        RECT 3.135000 92.635000 3.455000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 68.065000 3.505000 68.385000 ;
      LAYER met4 ;
        RECT 3.185000 68.065000 3.505000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 68.475000 3.505000 68.795000 ;
      LAYER met4 ;
        RECT 3.185000 68.475000 3.505000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 68.885000 3.505000 69.205000 ;
      LAYER met4 ;
        RECT 3.185000 68.885000 3.505000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 69.295000 3.505000 69.615000 ;
      LAYER met4 ;
        RECT 3.185000 69.295000 3.505000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 69.705000 3.505000 70.025000 ;
      LAYER met4 ;
        RECT 3.185000 69.705000 3.505000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 70.115000 3.505000 70.435000 ;
      LAYER met4 ;
        RECT 3.185000 70.115000 3.505000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 70.525000 3.505000 70.845000 ;
      LAYER met4 ;
        RECT 3.185000 70.525000 3.505000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 70.935000 3.505000 71.255000 ;
      LAYER met4 ;
        RECT 3.185000 70.935000 3.505000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 71.345000 3.505000 71.665000 ;
      LAYER met4 ;
        RECT 3.185000 71.345000 3.505000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 71.755000 3.505000 72.075000 ;
      LAYER met4 ;
        RECT 3.185000 71.755000 3.505000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 72.165000 3.505000 72.485000 ;
      LAYER met4 ;
        RECT 3.185000 72.165000 3.505000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 72.575000 3.505000 72.895000 ;
      LAYER met4 ;
        RECT 3.185000 72.575000 3.505000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 72.985000 3.505000 73.305000 ;
      LAYER met4 ;
        RECT 3.185000 72.985000 3.505000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 73.390000 3.505000 73.710000 ;
      LAYER met4 ;
        RECT 3.185000 73.390000 3.505000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 73.795000 3.505000 74.115000 ;
      LAYER met4 ;
        RECT 3.185000 73.795000 3.505000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 74.200000 3.505000 74.520000 ;
      LAYER met4 ;
        RECT 3.185000 74.200000 3.505000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 74.605000 3.505000 74.925000 ;
      LAYER met4 ;
        RECT 3.185000 74.605000 3.505000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 75.010000 3.505000 75.330000 ;
      LAYER met4 ;
        RECT 3.185000 75.010000 3.505000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 75.415000 3.505000 75.735000 ;
      LAYER met4 ;
        RECT 3.185000 75.415000 3.505000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 75.820000 3.505000 76.140000 ;
      LAYER met4 ;
        RECT 3.185000 75.820000 3.505000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 76.225000 3.505000 76.545000 ;
      LAYER met4 ;
        RECT 3.185000 76.225000 3.505000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 76.630000 3.505000 76.950000 ;
      LAYER met4 ;
        RECT 3.185000 76.630000 3.505000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 77.035000 3.505000 77.355000 ;
      LAYER met4 ;
        RECT 3.185000 77.035000 3.505000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 77.440000 3.505000 77.760000 ;
      LAYER met4 ;
        RECT 3.185000 77.440000 3.505000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 77.845000 3.505000 78.165000 ;
      LAYER met4 ;
        RECT 3.185000 77.845000 3.505000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 78.250000 3.505000 78.570000 ;
      LAYER met4 ;
        RECT 3.185000 78.250000 3.505000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 78.655000 3.505000 78.975000 ;
      LAYER met4 ;
        RECT 3.185000 78.655000 3.505000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 79.060000 3.505000 79.380000 ;
      LAYER met4 ;
        RECT 3.185000 79.060000 3.505000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 79.465000 3.505000 79.785000 ;
      LAYER met4 ;
        RECT 3.185000 79.465000 3.505000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 79.870000 3.505000 80.190000 ;
      LAYER met4 ;
        RECT 3.185000 79.870000 3.505000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 80.275000 3.505000 80.595000 ;
      LAYER met4 ;
        RECT 3.185000 80.275000 3.505000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 80.680000 3.505000 81.000000 ;
      LAYER met4 ;
        RECT 3.185000 80.680000 3.505000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 81.085000 3.505000 81.405000 ;
      LAYER met4 ;
        RECT 3.185000 81.085000 3.505000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 81.490000 3.505000 81.810000 ;
      LAYER met4 ;
        RECT 3.185000 81.490000 3.505000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 81.895000 3.505000 82.215000 ;
      LAYER met4 ;
        RECT 3.185000 81.895000 3.505000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185000 82.300000 3.505000 82.620000 ;
      LAYER met4 ;
        RECT 3.185000 82.300000 3.505000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465000 17.800000 3.785000 18.120000 ;
      LAYER met4 ;
        RECT 3.465000 17.800000 3.785000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465000 18.230000 3.785000 18.550000 ;
      LAYER met4 ;
        RECT 3.465000 18.230000 3.785000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465000 18.660000 3.785000 18.980000 ;
      LAYER met4 ;
        RECT 3.465000 18.660000 3.785000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465000 19.090000 3.785000 19.410000 ;
      LAYER met4 ;
        RECT 3.465000 19.090000 3.785000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465000 19.520000 3.785000 19.840000 ;
      LAYER met4 ;
        RECT 3.465000 19.520000 3.785000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465000 19.950000 3.785000 20.270000 ;
      LAYER met4 ;
        RECT 3.465000 19.950000 3.785000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465000 20.380000 3.785000 20.700000 ;
      LAYER met4 ;
        RECT 3.465000 20.380000 3.785000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465000 20.810000 3.785000 21.130000 ;
      LAYER met4 ;
        RECT 3.465000 20.810000 3.785000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465000 21.240000 3.785000 21.560000 ;
      LAYER met4 ;
        RECT 3.465000 21.240000 3.785000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465000 21.670000 3.785000 21.990000 ;
      LAYER met4 ;
        RECT 3.465000 21.670000 3.785000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465000 22.100000 3.785000 22.420000 ;
      LAYER met4 ;
        RECT 3.465000 22.100000 3.785000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 82.795000 3.865000 83.115000 ;
      LAYER met4 ;
        RECT 3.545000 82.795000 3.865000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 83.205000 3.865000 83.525000 ;
      LAYER met4 ;
        RECT 3.545000 83.205000 3.865000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 83.615000 3.865000 83.935000 ;
      LAYER met4 ;
        RECT 3.545000 83.615000 3.865000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 84.025000 3.865000 84.345000 ;
      LAYER met4 ;
        RECT 3.545000 84.025000 3.865000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 84.435000 3.865000 84.755000 ;
      LAYER met4 ;
        RECT 3.545000 84.435000 3.865000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 84.845000 3.865000 85.165000 ;
      LAYER met4 ;
        RECT 3.545000 84.845000 3.865000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 85.255000 3.865000 85.575000 ;
      LAYER met4 ;
        RECT 3.545000 85.255000 3.865000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 85.665000 3.865000 85.985000 ;
      LAYER met4 ;
        RECT 3.545000 85.665000 3.865000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 86.075000 3.865000 86.395000 ;
      LAYER met4 ;
        RECT 3.545000 86.075000 3.865000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 86.485000 3.865000 86.805000 ;
      LAYER met4 ;
        RECT 3.545000 86.485000 3.865000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 86.895000 3.865000 87.215000 ;
      LAYER met4 ;
        RECT 3.545000 86.895000 3.865000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 87.305000 3.865000 87.625000 ;
      LAYER met4 ;
        RECT 3.545000 87.305000 3.865000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 87.715000 3.865000 88.035000 ;
      LAYER met4 ;
        RECT 3.545000 87.715000 3.865000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 88.125000 3.865000 88.445000 ;
      LAYER met4 ;
        RECT 3.545000 88.125000 3.865000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 88.535000 3.865000 88.855000 ;
      LAYER met4 ;
        RECT 3.545000 88.535000 3.865000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 88.945000 3.865000 89.265000 ;
      LAYER met4 ;
        RECT 3.545000 88.945000 3.865000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 89.355000 3.865000 89.675000 ;
      LAYER met4 ;
        RECT 3.545000 89.355000 3.865000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 89.765000 3.865000 90.085000 ;
      LAYER met4 ;
        RECT 3.545000 89.765000 3.865000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 90.175000 3.865000 90.495000 ;
      LAYER met4 ;
        RECT 3.545000 90.175000 3.865000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 90.585000 3.865000 90.905000 ;
      LAYER met4 ;
        RECT 3.545000 90.585000 3.865000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 90.995000 3.865000 91.315000 ;
      LAYER met4 ;
        RECT 3.545000 90.995000 3.865000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 91.405000 3.865000 91.725000 ;
      LAYER met4 ;
        RECT 3.545000 91.405000 3.865000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 91.815000 3.865000 92.135000 ;
      LAYER met4 ;
        RECT 3.545000 91.815000 3.865000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 92.225000 3.865000 92.545000 ;
      LAYER met4 ;
        RECT 3.545000 92.225000 3.865000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545000 92.635000 3.865000 92.955000 ;
      LAYER met4 ;
        RECT 3.545000 92.635000 3.865000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 68.065000 3.905000 68.385000 ;
      LAYER met4 ;
        RECT 3.585000 68.065000 3.905000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 68.475000 3.905000 68.795000 ;
      LAYER met4 ;
        RECT 3.585000 68.475000 3.905000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 68.885000 3.905000 69.205000 ;
      LAYER met4 ;
        RECT 3.585000 68.885000 3.905000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 69.295000 3.905000 69.615000 ;
      LAYER met4 ;
        RECT 3.585000 69.295000 3.905000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 69.705000 3.905000 70.025000 ;
      LAYER met4 ;
        RECT 3.585000 69.705000 3.905000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 70.115000 3.905000 70.435000 ;
      LAYER met4 ;
        RECT 3.585000 70.115000 3.905000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 70.525000 3.905000 70.845000 ;
      LAYER met4 ;
        RECT 3.585000 70.525000 3.905000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 70.935000 3.905000 71.255000 ;
      LAYER met4 ;
        RECT 3.585000 70.935000 3.905000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 71.345000 3.905000 71.665000 ;
      LAYER met4 ;
        RECT 3.585000 71.345000 3.905000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 71.755000 3.905000 72.075000 ;
      LAYER met4 ;
        RECT 3.585000 71.755000 3.905000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 72.165000 3.905000 72.485000 ;
      LAYER met4 ;
        RECT 3.585000 72.165000 3.905000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 72.575000 3.905000 72.895000 ;
      LAYER met4 ;
        RECT 3.585000 72.575000 3.905000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 72.985000 3.905000 73.305000 ;
      LAYER met4 ;
        RECT 3.585000 72.985000 3.905000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 73.390000 3.905000 73.710000 ;
      LAYER met4 ;
        RECT 3.585000 73.390000 3.905000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 73.795000 3.905000 74.115000 ;
      LAYER met4 ;
        RECT 3.585000 73.795000 3.905000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 74.200000 3.905000 74.520000 ;
      LAYER met4 ;
        RECT 3.585000 74.200000 3.905000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 74.605000 3.905000 74.925000 ;
      LAYER met4 ;
        RECT 3.585000 74.605000 3.905000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 75.010000 3.905000 75.330000 ;
      LAYER met4 ;
        RECT 3.585000 75.010000 3.905000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 75.415000 3.905000 75.735000 ;
      LAYER met4 ;
        RECT 3.585000 75.415000 3.905000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 75.820000 3.905000 76.140000 ;
      LAYER met4 ;
        RECT 3.585000 75.820000 3.905000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 76.225000 3.905000 76.545000 ;
      LAYER met4 ;
        RECT 3.585000 76.225000 3.905000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 76.630000 3.905000 76.950000 ;
      LAYER met4 ;
        RECT 3.585000 76.630000 3.905000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 77.035000 3.905000 77.355000 ;
      LAYER met4 ;
        RECT 3.585000 77.035000 3.905000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 77.440000 3.905000 77.760000 ;
      LAYER met4 ;
        RECT 3.585000 77.440000 3.905000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 77.845000 3.905000 78.165000 ;
      LAYER met4 ;
        RECT 3.585000 77.845000 3.905000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 78.250000 3.905000 78.570000 ;
      LAYER met4 ;
        RECT 3.585000 78.250000 3.905000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 78.655000 3.905000 78.975000 ;
      LAYER met4 ;
        RECT 3.585000 78.655000 3.905000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 79.060000 3.905000 79.380000 ;
      LAYER met4 ;
        RECT 3.585000 79.060000 3.905000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 79.465000 3.905000 79.785000 ;
      LAYER met4 ;
        RECT 3.585000 79.465000 3.905000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 79.870000 3.905000 80.190000 ;
      LAYER met4 ;
        RECT 3.585000 79.870000 3.905000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 80.275000 3.905000 80.595000 ;
      LAYER met4 ;
        RECT 3.585000 80.275000 3.905000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 80.680000 3.905000 81.000000 ;
      LAYER met4 ;
        RECT 3.585000 80.680000 3.905000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 81.085000 3.905000 81.405000 ;
      LAYER met4 ;
        RECT 3.585000 81.085000 3.905000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 81.490000 3.905000 81.810000 ;
      LAYER met4 ;
        RECT 3.585000 81.490000 3.905000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 81.895000 3.905000 82.215000 ;
      LAYER met4 ;
        RECT 3.585000 81.895000 3.905000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585000 82.300000 3.905000 82.620000 ;
      LAYER met4 ;
        RECT 3.585000 82.300000 3.905000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870000 17.800000 4.190000 18.120000 ;
      LAYER met4 ;
        RECT 3.870000 17.800000 4.190000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870000 18.230000 4.190000 18.550000 ;
      LAYER met4 ;
        RECT 3.870000 18.230000 4.190000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870000 18.660000 4.190000 18.980000 ;
      LAYER met4 ;
        RECT 3.870000 18.660000 4.190000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870000 19.090000 4.190000 19.410000 ;
      LAYER met4 ;
        RECT 3.870000 19.090000 4.190000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870000 19.520000 4.190000 19.840000 ;
      LAYER met4 ;
        RECT 3.870000 19.520000 4.190000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870000 19.950000 4.190000 20.270000 ;
      LAYER met4 ;
        RECT 3.870000 19.950000 4.190000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870000 20.380000 4.190000 20.700000 ;
      LAYER met4 ;
        RECT 3.870000 20.380000 4.190000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870000 20.810000 4.190000 21.130000 ;
      LAYER met4 ;
        RECT 3.870000 20.810000 4.190000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870000 21.240000 4.190000 21.560000 ;
      LAYER met4 ;
        RECT 3.870000 21.240000 4.190000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870000 21.670000 4.190000 21.990000 ;
      LAYER met4 ;
        RECT 3.870000 21.670000 4.190000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870000 22.100000 4.190000 22.420000 ;
      LAYER met4 ;
        RECT 3.870000 22.100000 4.190000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 82.795000 4.275000 83.115000 ;
      LAYER met4 ;
        RECT 3.955000 82.795000 4.275000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 83.205000 4.275000 83.525000 ;
      LAYER met4 ;
        RECT 3.955000 83.205000 4.275000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 83.615000 4.275000 83.935000 ;
      LAYER met4 ;
        RECT 3.955000 83.615000 4.275000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 84.025000 4.275000 84.345000 ;
      LAYER met4 ;
        RECT 3.955000 84.025000 4.275000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 84.435000 4.275000 84.755000 ;
      LAYER met4 ;
        RECT 3.955000 84.435000 4.275000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 84.845000 4.275000 85.165000 ;
      LAYER met4 ;
        RECT 3.955000 84.845000 4.275000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 85.255000 4.275000 85.575000 ;
      LAYER met4 ;
        RECT 3.955000 85.255000 4.275000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 85.665000 4.275000 85.985000 ;
      LAYER met4 ;
        RECT 3.955000 85.665000 4.275000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 86.075000 4.275000 86.395000 ;
      LAYER met4 ;
        RECT 3.955000 86.075000 4.275000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 86.485000 4.275000 86.805000 ;
      LAYER met4 ;
        RECT 3.955000 86.485000 4.275000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 86.895000 4.275000 87.215000 ;
      LAYER met4 ;
        RECT 3.955000 86.895000 4.275000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 87.305000 4.275000 87.625000 ;
      LAYER met4 ;
        RECT 3.955000 87.305000 4.275000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 87.715000 4.275000 88.035000 ;
      LAYER met4 ;
        RECT 3.955000 87.715000 4.275000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 88.125000 4.275000 88.445000 ;
      LAYER met4 ;
        RECT 3.955000 88.125000 4.275000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 88.535000 4.275000 88.855000 ;
      LAYER met4 ;
        RECT 3.955000 88.535000 4.275000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 88.945000 4.275000 89.265000 ;
      LAYER met4 ;
        RECT 3.955000 88.945000 4.275000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 89.355000 4.275000 89.675000 ;
      LAYER met4 ;
        RECT 3.955000 89.355000 4.275000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 89.765000 4.275000 90.085000 ;
      LAYER met4 ;
        RECT 3.955000 89.765000 4.275000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 90.175000 4.275000 90.495000 ;
      LAYER met4 ;
        RECT 3.955000 90.175000 4.275000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 90.585000 4.275000 90.905000 ;
      LAYER met4 ;
        RECT 3.955000 90.585000 4.275000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 90.995000 4.275000 91.315000 ;
      LAYER met4 ;
        RECT 3.955000 90.995000 4.275000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 91.405000 4.275000 91.725000 ;
      LAYER met4 ;
        RECT 3.955000 91.405000 4.275000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 91.815000 4.275000 92.135000 ;
      LAYER met4 ;
        RECT 3.955000 91.815000 4.275000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 92.225000 4.275000 92.545000 ;
      LAYER met4 ;
        RECT 3.955000 92.225000 4.275000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955000 92.635000 4.275000 92.955000 ;
      LAYER met4 ;
        RECT 3.955000 92.635000 4.275000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 68.065000 4.305000 68.385000 ;
      LAYER met4 ;
        RECT 3.985000 68.065000 4.305000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 68.475000 4.305000 68.795000 ;
      LAYER met4 ;
        RECT 3.985000 68.475000 4.305000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 68.885000 4.305000 69.205000 ;
      LAYER met4 ;
        RECT 3.985000 68.885000 4.305000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 69.295000 4.305000 69.615000 ;
      LAYER met4 ;
        RECT 3.985000 69.295000 4.305000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 69.705000 4.305000 70.025000 ;
      LAYER met4 ;
        RECT 3.985000 69.705000 4.305000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 70.115000 4.305000 70.435000 ;
      LAYER met4 ;
        RECT 3.985000 70.115000 4.305000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 70.525000 4.305000 70.845000 ;
      LAYER met4 ;
        RECT 3.985000 70.525000 4.305000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 70.935000 4.305000 71.255000 ;
      LAYER met4 ;
        RECT 3.985000 70.935000 4.305000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 71.345000 4.305000 71.665000 ;
      LAYER met4 ;
        RECT 3.985000 71.345000 4.305000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 71.755000 4.305000 72.075000 ;
      LAYER met4 ;
        RECT 3.985000 71.755000 4.305000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 72.165000 4.305000 72.485000 ;
      LAYER met4 ;
        RECT 3.985000 72.165000 4.305000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 72.575000 4.305000 72.895000 ;
      LAYER met4 ;
        RECT 3.985000 72.575000 4.305000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 72.985000 4.305000 73.305000 ;
      LAYER met4 ;
        RECT 3.985000 72.985000 4.305000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 73.390000 4.305000 73.710000 ;
      LAYER met4 ;
        RECT 3.985000 73.390000 4.305000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 73.795000 4.305000 74.115000 ;
      LAYER met4 ;
        RECT 3.985000 73.795000 4.305000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 74.200000 4.305000 74.520000 ;
      LAYER met4 ;
        RECT 3.985000 74.200000 4.305000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 74.605000 4.305000 74.925000 ;
      LAYER met4 ;
        RECT 3.985000 74.605000 4.305000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 75.010000 4.305000 75.330000 ;
      LAYER met4 ;
        RECT 3.985000 75.010000 4.305000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 75.415000 4.305000 75.735000 ;
      LAYER met4 ;
        RECT 3.985000 75.415000 4.305000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 75.820000 4.305000 76.140000 ;
      LAYER met4 ;
        RECT 3.985000 75.820000 4.305000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 76.225000 4.305000 76.545000 ;
      LAYER met4 ;
        RECT 3.985000 76.225000 4.305000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 76.630000 4.305000 76.950000 ;
      LAYER met4 ;
        RECT 3.985000 76.630000 4.305000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 77.035000 4.305000 77.355000 ;
      LAYER met4 ;
        RECT 3.985000 77.035000 4.305000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 77.440000 4.305000 77.760000 ;
      LAYER met4 ;
        RECT 3.985000 77.440000 4.305000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 77.845000 4.305000 78.165000 ;
      LAYER met4 ;
        RECT 3.985000 77.845000 4.305000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 78.250000 4.305000 78.570000 ;
      LAYER met4 ;
        RECT 3.985000 78.250000 4.305000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 78.655000 4.305000 78.975000 ;
      LAYER met4 ;
        RECT 3.985000 78.655000 4.305000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 79.060000 4.305000 79.380000 ;
      LAYER met4 ;
        RECT 3.985000 79.060000 4.305000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 79.465000 4.305000 79.785000 ;
      LAYER met4 ;
        RECT 3.985000 79.465000 4.305000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 79.870000 4.305000 80.190000 ;
      LAYER met4 ;
        RECT 3.985000 79.870000 4.305000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 80.275000 4.305000 80.595000 ;
      LAYER met4 ;
        RECT 3.985000 80.275000 4.305000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 80.680000 4.305000 81.000000 ;
      LAYER met4 ;
        RECT 3.985000 80.680000 4.305000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 81.085000 4.305000 81.405000 ;
      LAYER met4 ;
        RECT 3.985000 81.085000 4.305000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 81.490000 4.305000 81.810000 ;
      LAYER met4 ;
        RECT 3.985000 81.490000 4.305000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 81.895000 4.305000 82.215000 ;
      LAYER met4 ;
        RECT 3.985000 81.895000 4.305000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985000 82.300000 4.305000 82.620000 ;
      LAYER met4 ;
        RECT 3.985000 82.300000 4.305000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275000 17.800000 4.595000 18.120000 ;
      LAYER met4 ;
        RECT 4.275000 17.800000 4.595000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275000 18.230000 4.595000 18.550000 ;
      LAYER met4 ;
        RECT 4.275000 18.230000 4.595000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275000 18.660000 4.595000 18.980000 ;
      LAYER met4 ;
        RECT 4.275000 18.660000 4.595000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275000 19.090000 4.595000 19.410000 ;
      LAYER met4 ;
        RECT 4.275000 19.090000 4.595000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275000 19.520000 4.595000 19.840000 ;
      LAYER met4 ;
        RECT 4.275000 19.520000 4.595000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275000 19.950000 4.595000 20.270000 ;
      LAYER met4 ;
        RECT 4.275000 19.950000 4.595000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275000 20.380000 4.595000 20.700000 ;
      LAYER met4 ;
        RECT 4.275000 20.380000 4.595000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275000 20.810000 4.595000 21.130000 ;
      LAYER met4 ;
        RECT 4.275000 20.810000 4.595000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275000 21.240000 4.595000 21.560000 ;
      LAYER met4 ;
        RECT 4.275000 21.240000 4.595000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275000 21.670000 4.595000 21.990000 ;
      LAYER met4 ;
        RECT 4.275000 21.670000 4.595000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275000 22.100000 4.595000 22.420000 ;
      LAYER met4 ;
        RECT 4.275000 22.100000 4.595000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 82.795000 4.685000 83.115000 ;
      LAYER met4 ;
        RECT 4.365000 82.795000 4.685000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 83.205000 4.685000 83.525000 ;
      LAYER met4 ;
        RECT 4.365000 83.205000 4.685000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 83.615000 4.685000 83.935000 ;
      LAYER met4 ;
        RECT 4.365000 83.615000 4.685000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 84.025000 4.685000 84.345000 ;
      LAYER met4 ;
        RECT 4.365000 84.025000 4.685000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 84.435000 4.685000 84.755000 ;
      LAYER met4 ;
        RECT 4.365000 84.435000 4.685000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 84.845000 4.685000 85.165000 ;
      LAYER met4 ;
        RECT 4.365000 84.845000 4.685000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 85.255000 4.685000 85.575000 ;
      LAYER met4 ;
        RECT 4.365000 85.255000 4.685000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 85.665000 4.685000 85.985000 ;
      LAYER met4 ;
        RECT 4.365000 85.665000 4.685000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 86.075000 4.685000 86.395000 ;
      LAYER met4 ;
        RECT 4.365000 86.075000 4.685000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 86.485000 4.685000 86.805000 ;
      LAYER met4 ;
        RECT 4.365000 86.485000 4.685000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 86.895000 4.685000 87.215000 ;
      LAYER met4 ;
        RECT 4.365000 86.895000 4.685000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 87.305000 4.685000 87.625000 ;
      LAYER met4 ;
        RECT 4.365000 87.305000 4.685000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 87.715000 4.685000 88.035000 ;
      LAYER met4 ;
        RECT 4.365000 87.715000 4.685000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 88.125000 4.685000 88.445000 ;
      LAYER met4 ;
        RECT 4.365000 88.125000 4.685000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 88.535000 4.685000 88.855000 ;
      LAYER met4 ;
        RECT 4.365000 88.535000 4.685000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 88.945000 4.685000 89.265000 ;
      LAYER met4 ;
        RECT 4.365000 88.945000 4.685000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 89.355000 4.685000 89.675000 ;
      LAYER met4 ;
        RECT 4.365000 89.355000 4.685000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 89.765000 4.685000 90.085000 ;
      LAYER met4 ;
        RECT 4.365000 89.765000 4.685000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 90.175000 4.685000 90.495000 ;
      LAYER met4 ;
        RECT 4.365000 90.175000 4.685000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 90.585000 4.685000 90.905000 ;
      LAYER met4 ;
        RECT 4.365000 90.585000 4.685000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 90.995000 4.685000 91.315000 ;
      LAYER met4 ;
        RECT 4.365000 90.995000 4.685000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 91.405000 4.685000 91.725000 ;
      LAYER met4 ;
        RECT 4.365000 91.405000 4.685000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 91.815000 4.685000 92.135000 ;
      LAYER met4 ;
        RECT 4.365000 91.815000 4.685000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 92.225000 4.685000 92.545000 ;
      LAYER met4 ;
        RECT 4.365000 92.225000 4.685000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365000 92.635000 4.685000 92.955000 ;
      LAYER met4 ;
        RECT 4.365000 92.635000 4.685000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 68.065000 4.705000 68.385000 ;
      LAYER met4 ;
        RECT 4.385000 68.065000 4.705000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 68.475000 4.705000 68.795000 ;
      LAYER met4 ;
        RECT 4.385000 68.475000 4.705000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 68.885000 4.705000 69.205000 ;
      LAYER met4 ;
        RECT 4.385000 68.885000 4.705000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 69.295000 4.705000 69.615000 ;
      LAYER met4 ;
        RECT 4.385000 69.295000 4.705000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 69.705000 4.705000 70.025000 ;
      LAYER met4 ;
        RECT 4.385000 69.705000 4.705000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 70.115000 4.705000 70.435000 ;
      LAYER met4 ;
        RECT 4.385000 70.115000 4.705000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 70.525000 4.705000 70.845000 ;
      LAYER met4 ;
        RECT 4.385000 70.525000 4.705000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 70.935000 4.705000 71.255000 ;
      LAYER met4 ;
        RECT 4.385000 70.935000 4.705000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 71.345000 4.705000 71.665000 ;
      LAYER met4 ;
        RECT 4.385000 71.345000 4.705000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 71.755000 4.705000 72.075000 ;
      LAYER met4 ;
        RECT 4.385000 71.755000 4.705000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 72.165000 4.705000 72.485000 ;
      LAYER met4 ;
        RECT 4.385000 72.165000 4.705000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 72.575000 4.705000 72.895000 ;
      LAYER met4 ;
        RECT 4.385000 72.575000 4.705000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 72.985000 4.705000 73.305000 ;
      LAYER met4 ;
        RECT 4.385000 72.985000 4.705000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 73.390000 4.705000 73.710000 ;
      LAYER met4 ;
        RECT 4.385000 73.390000 4.705000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 73.795000 4.705000 74.115000 ;
      LAYER met4 ;
        RECT 4.385000 73.795000 4.705000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 74.200000 4.705000 74.520000 ;
      LAYER met4 ;
        RECT 4.385000 74.200000 4.705000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 74.605000 4.705000 74.925000 ;
      LAYER met4 ;
        RECT 4.385000 74.605000 4.705000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 75.010000 4.705000 75.330000 ;
      LAYER met4 ;
        RECT 4.385000 75.010000 4.705000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 75.415000 4.705000 75.735000 ;
      LAYER met4 ;
        RECT 4.385000 75.415000 4.705000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 75.820000 4.705000 76.140000 ;
      LAYER met4 ;
        RECT 4.385000 75.820000 4.705000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 76.225000 4.705000 76.545000 ;
      LAYER met4 ;
        RECT 4.385000 76.225000 4.705000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 76.630000 4.705000 76.950000 ;
      LAYER met4 ;
        RECT 4.385000 76.630000 4.705000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 77.035000 4.705000 77.355000 ;
      LAYER met4 ;
        RECT 4.385000 77.035000 4.705000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 77.440000 4.705000 77.760000 ;
      LAYER met4 ;
        RECT 4.385000 77.440000 4.705000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 77.845000 4.705000 78.165000 ;
      LAYER met4 ;
        RECT 4.385000 77.845000 4.705000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 78.250000 4.705000 78.570000 ;
      LAYER met4 ;
        RECT 4.385000 78.250000 4.705000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 78.655000 4.705000 78.975000 ;
      LAYER met4 ;
        RECT 4.385000 78.655000 4.705000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 79.060000 4.705000 79.380000 ;
      LAYER met4 ;
        RECT 4.385000 79.060000 4.705000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 79.465000 4.705000 79.785000 ;
      LAYER met4 ;
        RECT 4.385000 79.465000 4.705000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 79.870000 4.705000 80.190000 ;
      LAYER met4 ;
        RECT 4.385000 79.870000 4.705000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 80.275000 4.705000 80.595000 ;
      LAYER met4 ;
        RECT 4.385000 80.275000 4.705000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 80.680000 4.705000 81.000000 ;
      LAYER met4 ;
        RECT 4.385000 80.680000 4.705000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 81.085000 4.705000 81.405000 ;
      LAYER met4 ;
        RECT 4.385000 81.085000 4.705000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 81.490000 4.705000 81.810000 ;
      LAYER met4 ;
        RECT 4.385000 81.490000 4.705000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 81.895000 4.705000 82.215000 ;
      LAYER met4 ;
        RECT 4.385000 81.895000 4.705000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385000 82.300000 4.705000 82.620000 ;
      LAYER met4 ;
        RECT 4.385000 82.300000 4.705000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680000 17.800000 5.000000 18.120000 ;
      LAYER met4 ;
        RECT 4.680000 17.800000 5.000000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680000 18.230000 5.000000 18.550000 ;
      LAYER met4 ;
        RECT 4.680000 18.230000 5.000000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680000 18.660000 5.000000 18.980000 ;
      LAYER met4 ;
        RECT 4.680000 18.660000 5.000000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680000 19.090000 5.000000 19.410000 ;
      LAYER met4 ;
        RECT 4.680000 19.090000 5.000000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680000 19.520000 5.000000 19.840000 ;
      LAYER met4 ;
        RECT 4.680000 19.520000 5.000000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680000 19.950000 5.000000 20.270000 ;
      LAYER met4 ;
        RECT 4.680000 19.950000 5.000000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680000 20.380000 5.000000 20.700000 ;
      LAYER met4 ;
        RECT 4.680000 20.380000 5.000000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680000 20.810000 5.000000 21.130000 ;
      LAYER met4 ;
        RECT 4.680000 20.810000 5.000000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680000 21.240000 5.000000 21.560000 ;
      LAYER met4 ;
        RECT 4.680000 21.240000 5.000000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680000 21.670000 5.000000 21.990000 ;
      LAYER met4 ;
        RECT 4.680000 21.670000 5.000000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680000 22.100000 5.000000 22.420000 ;
      LAYER met4 ;
        RECT 4.680000 22.100000 5.000000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 82.795000 5.095000 83.115000 ;
      LAYER met4 ;
        RECT 4.775000 82.795000 5.095000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 83.205000 5.095000 83.525000 ;
      LAYER met4 ;
        RECT 4.775000 83.205000 5.095000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 83.615000 5.095000 83.935000 ;
      LAYER met4 ;
        RECT 4.775000 83.615000 5.095000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 84.025000 5.095000 84.345000 ;
      LAYER met4 ;
        RECT 4.775000 84.025000 5.095000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 84.435000 5.095000 84.755000 ;
      LAYER met4 ;
        RECT 4.775000 84.435000 5.095000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 84.845000 5.095000 85.165000 ;
      LAYER met4 ;
        RECT 4.775000 84.845000 5.095000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 85.255000 5.095000 85.575000 ;
      LAYER met4 ;
        RECT 4.775000 85.255000 5.095000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 85.665000 5.095000 85.985000 ;
      LAYER met4 ;
        RECT 4.775000 85.665000 5.095000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 86.075000 5.095000 86.395000 ;
      LAYER met4 ;
        RECT 4.775000 86.075000 5.095000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 86.485000 5.095000 86.805000 ;
      LAYER met4 ;
        RECT 4.775000 86.485000 5.095000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 86.895000 5.095000 87.215000 ;
      LAYER met4 ;
        RECT 4.775000 86.895000 5.095000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 87.305000 5.095000 87.625000 ;
      LAYER met4 ;
        RECT 4.775000 87.305000 5.095000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 87.715000 5.095000 88.035000 ;
      LAYER met4 ;
        RECT 4.775000 87.715000 5.095000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 88.125000 5.095000 88.445000 ;
      LAYER met4 ;
        RECT 4.775000 88.125000 5.095000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 88.535000 5.095000 88.855000 ;
      LAYER met4 ;
        RECT 4.775000 88.535000 5.095000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 88.945000 5.095000 89.265000 ;
      LAYER met4 ;
        RECT 4.775000 88.945000 5.095000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 89.355000 5.095000 89.675000 ;
      LAYER met4 ;
        RECT 4.775000 89.355000 5.095000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 89.765000 5.095000 90.085000 ;
      LAYER met4 ;
        RECT 4.775000 89.765000 5.095000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 90.175000 5.095000 90.495000 ;
      LAYER met4 ;
        RECT 4.775000 90.175000 5.095000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 90.585000 5.095000 90.905000 ;
      LAYER met4 ;
        RECT 4.775000 90.585000 5.095000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 90.995000 5.095000 91.315000 ;
      LAYER met4 ;
        RECT 4.775000 90.995000 5.095000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 91.405000 5.095000 91.725000 ;
      LAYER met4 ;
        RECT 4.775000 91.405000 5.095000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 91.815000 5.095000 92.135000 ;
      LAYER met4 ;
        RECT 4.775000 91.815000 5.095000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 92.225000 5.095000 92.545000 ;
      LAYER met4 ;
        RECT 4.775000 92.225000 5.095000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775000 92.635000 5.095000 92.955000 ;
      LAYER met4 ;
        RECT 4.775000 92.635000 5.095000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 68.065000 5.105000 68.385000 ;
      LAYER met4 ;
        RECT 4.785000 68.065000 5.105000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 68.475000 5.105000 68.795000 ;
      LAYER met4 ;
        RECT 4.785000 68.475000 5.105000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 68.885000 5.105000 69.205000 ;
      LAYER met4 ;
        RECT 4.785000 68.885000 5.105000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 69.295000 5.105000 69.615000 ;
      LAYER met4 ;
        RECT 4.785000 69.295000 5.105000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 69.705000 5.105000 70.025000 ;
      LAYER met4 ;
        RECT 4.785000 69.705000 5.105000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 70.115000 5.105000 70.435000 ;
      LAYER met4 ;
        RECT 4.785000 70.115000 5.105000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 70.525000 5.105000 70.845000 ;
      LAYER met4 ;
        RECT 4.785000 70.525000 5.105000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 70.935000 5.105000 71.255000 ;
      LAYER met4 ;
        RECT 4.785000 70.935000 5.105000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 71.345000 5.105000 71.665000 ;
      LAYER met4 ;
        RECT 4.785000 71.345000 5.105000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 71.755000 5.105000 72.075000 ;
      LAYER met4 ;
        RECT 4.785000 71.755000 5.105000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 72.165000 5.105000 72.485000 ;
      LAYER met4 ;
        RECT 4.785000 72.165000 5.105000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 72.575000 5.105000 72.895000 ;
      LAYER met4 ;
        RECT 4.785000 72.575000 5.105000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 72.985000 5.105000 73.305000 ;
      LAYER met4 ;
        RECT 4.785000 72.985000 5.105000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 73.390000 5.105000 73.710000 ;
      LAYER met4 ;
        RECT 4.785000 73.390000 5.105000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 73.795000 5.105000 74.115000 ;
      LAYER met4 ;
        RECT 4.785000 73.795000 5.105000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 74.200000 5.105000 74.520000 ;
      LAYER met4 ;
        RECT 4.785000 74.200000 5.105000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 74.605000 5.105000 74.925000 ;
      LAYER met4 ;
        RECT 4.785000 74.605000 5.105000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 75.010000 5.105000 75.330000 ;
      LAYER met4 ;
        RECT 4.785000 75.010000 5.105000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 75.415000 5.105000 75.735000 ;
      LAYER met4 ;
        RECT 4.785000 75.415000 5.105000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 75.820000 5.105000 76.140000 ;
      LAYER met4 ;
        RECT 4.785000 75.820000 5.105000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 76.225000 5.105000 76.545000 ;
      LAYER met4 ;
        RECT 4.785000 76.225000 5.105000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 76.630000 5.105000 76.950000 ;
      LAYER met4 ;
        RECT 4.785000 76.630000 5.105000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 77.035000 5.105000 77.355000 ;
      LAYER met4 ;
        RECT 4.785000 77.035000 5.105000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 77.440000 5.105000 77.760000 ;
      LAYER met4 ;
        RECT 4.785000 77.440000 5.105000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 77.845000 5.105000 78.165000 ;
      LAYER met4 ;
        RECT 4.785000 77.845000 5.105000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 78.250000 5.105000 78.570000 ;
      LAYER met4 ;
        RECT 4.785000 78.250000 5.105000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 78.655000 5.105000 78.975000 ;
      LAYER met4 ;
        RECT 4.785000 78.655000 5.105000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 79.060000 5.105000 79.380000 ;
      LAYER met4 ;
        RECT 4.785000 79.060000 5.105000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 79.465000 5.105000 79.785000 ;
      LAYER met4 ;
        RECT 4.785000 79.465000 5.105000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 79.870000 5.105000 80.190000 ;
      LAYER met4 ;
        RECT 4.785000 79.870000 5.105000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 80.275000 5.105000 80.595000 ;
      LAYER met4 ;
        RECT 4.785000 80.275000 5.105000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 80.680000 5.105000 81.000000 ;
      LAYER met4 ;
        RECT 4.785000 80.680000 5.105000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 81.085000 5.105000 81.405000 ;
      LAYER met4 ;
        RECT 4.785000 81.085000 5.105000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 81.490000 5.105000 81.810000 ;
      LAYER met4 ;
        RECT 4.785000 81.490000 5.105000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 81.895000 5.105000 82.215000 ;
      LAYER met4 ;
        RECT 4.785000 81.895000 5.105000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785000 82.300000 5.105000 82.620000 ;
      LAYER met4 ;
        RECT 4.785000 82.300000 5.105000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 17.800000 5.405000 18.120000 ;
      LAYER met4 ;
        RECT 5.085000 17.800000 5.405000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 18.230000 5.405000 18.550000 ;
      LAYER met4 ;
        RECT 5.085000 18.230000 5.405000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 18.660000 5.405000 18.980000 ;
      LAYER met4 ;
        RECT 5.085000 18.660000 5.405000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 19.090000 5.405000 19.410000 ;
      LAYER met4 ;
        RECT 5.085000 19.090000 5.405000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 19.520000 5.405000 19.840000 ;
      LAYER met4 ;
        RECT 5.085000 19.520000 5.405000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 19.950000 5.405000 20.270000 ;
      LAYER met4 ;
        RECT 5.085000 19.950000 5.405000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 20.380000 5.405000 20.700000 ;
      LAYER met4 ;
        RECT 5.085000 20.380000 5.405000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 20.810000 5.405000 21.130000 ;
      LAYER met4 ;
        RECT 5.085000 20.810000 5.405000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 21.240000 5.405000 21.560000 ;
      LAYER met4 ;
        RECT 5.085000 21.240000 5.405000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 21.670000 5.405000 21.990000 ;
      LAYER met4 ;
        RECT 5.085000 21.670000 5.405000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 22.100000 5.405000 22.420000 ;
      LAYER met4 ;
        RECT 5.085000 22.100000 5.405000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 68.065000 5.505000 68.385000 ;
      LAYER met4 ;
        RECT 5.185000 68.065000 5.505000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 68.475000 5.505000 68.795000 ;
      LAYER met4 ;
        RECT 5.185000 68.475000 5.505000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 68.885000 5.505000 69.205000 ;
      LAYER met4 ;
        RECT 5.185000 68.885000 5.505000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 69.295000 5.505000 69.615000 ;
      LAYER met4 ;
        RECT 5.185000 69.295000 5.505000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 69.705000 5.505000 70.025000 ;
      LAYER met4 ;
        RECT 5.185000 69.705000 5.505000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 70.115000 5.505000 70.435000 ;
      LAYER met4 ;
        RECT 5.185000 70.115000 5.505000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 70.525000 5.505000 70.845000 ;
      LAYER met4 ;
        RECT 5.185000 70.525000 5.505000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 70.935000 5.505000 71.255000 ;
      LAYER met4 ;
        RECT 5.185000 70.935000 5.505000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 71.345000 5.505000 71.665000 ;
      LAYER met4 ;
        RECT 5.185000 71.345000 5.505000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 71.755000 5.505000 72.075000 ;
      LAYER met4 ;
        RECT 5.185000 71.755000 5.505000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 72.165000 5.505000 72.485000 ;
      LAYER met4 ;
        RECT 5.185000 72.165000 5.505000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 72.575000 5.505000 72.895000 ;
      LAYER met4 ;
        RECT 5.185000 72.575000 5.505000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 72.985000 5.505000 73.305000 ;
      LAYER met4 ;
        RECT 5.185000 72.985000 5.505000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 73.390000 5.505000 73.710000 ;
      LAYER met4 ;
        RECT 5.185000 73.390000 5.505000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 73.795000 5.505000 74.115000 ;
      LAYER met4 ;
        RECT 5.185000 73.795000 5.505000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 74.200000 5.505000 74.520000 ;
      LAYER met4 ;
        RECT 5.185000 74.200000 5.505000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 74.605000 5.505000 74.925000 ;
      LAYER met4 ;
        RECT 5.185000 74.605000 5.505000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 75.010000 5.505000 75.330000 ;
      LAYER met4 ;
        RECT 5.185000 75.010000 5.505000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 75.415000 5.505000 75.735000 ;
      LAYER met4 ;
        RECT 5.185000 75.415000 5.505000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 75.820000 5.505000 76.140000 ;
      LAYER met4 ;
        RECT 5.185000 75.820000 5.505000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 76.225000 5.505000 76.545000 ;
      LAYER met4 ;
        RECT 5.185000 76.225000 5.505000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 76.630000 5.505000 76.950000 ;
      LAYER met4 ;
        RECT 5.185000 76.630000 5.505000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 77.035000 5.505000 77.355000 ;
      LAYER met4 ;
        RECT 5.185000 77.035000 5.505000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 77.440000 5.505000 77.760000 ;
      LAYER met4 ;
        RECT 5.185000 77.440000 5.505000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 77.845000 5.505000 78.165000 ;
      LAYER met4 ;
        RECT 5.185000 77.845000 5.505000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 78.250000 5.505000 78.570000 ;
      LAYER met4 ;
        RECT 5.185000 78.250000 5.505000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 78.655000 5.505000 78.975000 ;
      LAYER met4 ;
        RECT 5.185000 78.655000 5.505000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 79.060000 5.505000 79.380000 ;
      LAYER met4 ;
        RECT 5.185000 79.060000 5.505000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 79.465000 5.505000 79.785000 ;
      LAYER met4 ;
        RECT 5.185000 79.465000 5.505000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 79.870000 5.505000 80.190000 ;
      LAYER met4 ;
        RECT 5.185000 79.870000 5.505000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 80.275000 5.505000 80.595000 ;
      LAYER met4 ;
        RECT 5.185000 80.275000 5.505000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 80.680000 5.505000 81.000000 ;
      LAYER met4 ;
        RECT 5.185000 80.680000 5.505000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 81.085000 5.505000 81.405000 ;
      LAYER met4 ;
        RECT 5.185000 81.085000 5.505000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 81.490000 5.505000 81.810000 ;
      LAYER met4 ;
        RECT 5.185000 81.490000 5.505000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 81.895000 5.505000 82.215000 ;
      LAYER met4 ;
        RECT 5.185000 81.895000 5.505000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 82.300000 5.505000 82.620000 ;
      LAYER met4 ;
        RECT 5.185000 82.300000 5.505000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 82.795000 5.505000 83.115000 ;
      LAYER met4 ;
        RECT 5.185000 82.795000 5.505000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 83.205000 5.505000 83.525000 ;
      LAYER met4 ;
        RECT 5.185000 83.205000 5.505000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 83.615000 5.505000 83.935000 ;
      LAYER met4 ;
        RECT 5.185000 83.615000 5.505000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 84.025000 5.505000 84.345000 ;
      LAYER met4 ;
        RECT 5.185000 84.025000 5.505000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 84.435000 5.505000 84.755000 ;
      LAYER met4 ;
        RECT 5.185000 84.435000 5.505000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 84.845000 5.505000 85.165000 ;
      LAYER met4 ;
        RECT 5.185000 84.845000 5.505000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 85.255000 5.505000 85.575000 ;
      LAYER met4 ;
        RECT 5.185000 85.255000 5.505000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 85.665000 5.505000 85.985000 ;
      LAYER met4 ;
        RECT 5.185000 85.665000 5.505000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 86.075000 5.505000 86.395000 ;
      LAYER met4 ;
        RECT 5.185000 86.075000 5.505000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 86.485000 5.505000 86.805000 ;
      LAYER met4 ;
        RECT 5.185000 86.485000 5.505000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 86.895000 5.505000 87.215000 ;
      LAYER met4 ;
        RECT 5.185000 86.895000 5.505000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 87.305000 5.505000 87.625000 ;
      LAYER met4 ;
        RECT 5.185000 87.305000 5.505000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 87.715000 5.505000 88.035000 ;
      LAYER met4 ;
        RECT 5.185000 87.715000 5.505000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 88.125000 5.505000 88.445000 ;
      LAYER met4 ;
        RECT 5.185000 88.125000 5.505000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 88.535000 5.505000 88.855000 ;
      LAYER met4 ;
        RECT 5.185000 88.535000 5.505000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 88.945000 5.505000 89.265000 ;
      LAYER met4 ;
        RECT 5.185000 88.945000 5.505000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 89.355000 5.505000 89.675000 ;
      LAYER met4 ;
        RECT 5.185000 89.355000 5.505000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 89.765000 5.505000 90.085000 ;
      LAYER met4 ;
        RECT 5.185000 89.765000 5.505000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 90.175000 5.505000 90.495000 ;
      LAYER met4 ;
        RECT 5.185000 90.175000 5.505000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 90.585000 5.505000 90.905000 ;
      LAYER met4 ;
        RECT 5.185000 90.585000 5.505000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 90.995000 5.505000 91.315000 ;
      LAYER met4 ;
        RECT 5.185000 90.995000 5.505000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 91.405000 5.505000 91.725000 ;
      LAYER met4 ;
        RECT 5.185000 91.405000 5.505000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 91.815000 5.505000 92.135000 ;
      LAYER met4 ;
        RECT 5.185000 91.815000 5.505000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 92.225000 5.505000 92.545000 ;
      LAYER met4 ;
        RECT 5.185000 92.225000 5.505000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185000 92.635000 5.505000 92.955000 ;
      LAYER met4 ;
        RECT 5.185000 92.635000 5.505000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490000 17.800000 5.810000 18.120000 ;
      LAYER met4 ;
        RECT 5.490000 17.800000 5.810000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490000 18.230000 5.810000 18.550000 ;
      LAYER met4 ;
        RECT 5.490000 18.230000 5.810000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490000 18.660000 5.810000 18.980000 ;
      LAYER met4 ;
        RECT 5.490000 18.660000 5.810000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490000 19.090000 5.810000 19.410000 ;
      LAYER met4 ;
        RECT 5.490000 19.090000 5.810000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490000 19.520000 5.810000 19.840000 ;
      LAYER met4 ;
        RECT 5.490000 19.520000 5.810000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490000 19.950000 5.810000 20.270000 ;
      LAYER met4 ;
        RECT 5.490000 19.950000 5.810000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490000 20.380000 5.810000 20.700000 ;
      LAYER met4 ;
        RECT 5.490000 20.380000 5.810000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490000 20.810000 5.810000 21.130000 ;
      LAYER met4 ;
        RECT 5.490000 20.810000 5.810000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490000 21.240000 5.810000 21.560000 ;
      LAYER met4 ;
        RECT 5.490000 21.240000 5.810000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490000 21.670000 5.810000 21.990000 ;
      LAYER met4 ;
        RECT 5.490000 21.670000 5.810000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490000 22.100000 5.810000 22.420000 ;
      LAYER met4 ;
        RECT 5.490000 22.100000 5.810000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 68.065000 5.905000 68.385000 ;
      LAYER met4 ;
        RECT 5.585000 68.065000 5.905000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 68.475000 5.905000 68.795000 ;
      LAYER met4 ;
        RECT 5.585000 68.475000 5.905000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 68.885000 5.905000 69.205000 ;
      LAYER met4 ;
        RECT 5.585000 68.885000 5.905000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 69.295000 5.905000 69.615000 ;
      LAYER met4 ;
        RECT 5.585000 69.295000 5.905000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 69.705000 5.905000 70.025000 ;
      LAYER met4 ;
        RECT 5.585000 69.705000 5.905000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 70.115000 5.905000 70.435000 ;
      LAYER met4 ;
        RECT 5.585000 70.115000 5.905000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 70.525000 5.905000 70.845000 ;
      LAYER met4 ;
        RECT 5.585000 70.525000 5.905000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 70.935000 5.905000 71.255000 ;
      LAYER met4 ;
        RECT 5.585000 70.935000 5.905000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 71.345000 5.905000 71.665000 ;
      LAYER met4 ;
        RECT 5.585000 71.345000 5.905000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 71.755000 5.905000 72.075000 ;
      LAYER met4 ;
        RECT 5.585000 71.755000 5.905000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 72.165000 5.905000 72.485000 ;
      LAYER met4 ;
        RECT 5.585000 72.165000 5.905000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 72.575000 5.905000 72.895000 ;
      LAYER met4 ;
        RECT 5.585000 72.575000 5.905000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 72.985000 5.905000 73.305000 ;
      LAYER met4 ;
        RECT 5.585000 72.985000 5.905000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 73.390000 5.905000 73.710000 ;
      LAYER met4 ;
        RECT 5.585000 73.390000 5.905000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 73.795000 5.905000 74.115000 ;
      LAYER met4 ;
        RECT 5.585000 73.795000 5.905000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 74.200000 5.905000 74.520000 ;
      LAYER met4 ;
        RECT 5.585000 74.200000 5.905000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 74.605000 5.905000 74.925000 ;
      LAYER met4 ;
        RECT 5.585000 74.605000 5.905000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 75.010000 5.905000 75.330000 ;
      LAYER met4 ;
        RECT 5.585000 75.010000 5.905000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 75.415000 5.905000 75.735000 ;
      LAYER met4 ;
        RECT 5.585000 75.415000 5.905000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 75.820000 5.905000 76.140000 ;
      LAYER met4 ;
        RECT 5.585000 75.820000 5.905000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 76.225000 5.905000 76.545000 ;
      LAYER met4 ;
        RECT 5.585000 76.225000 5.905000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 76.630000 5.905000 76.950000 ;
      LAYER met4 ;
        RECT 5.585000 76.630000 5.905000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 77.035000 5.905000 77.355000 ;
      LAYER met4 ;
        RECT 5.585000 77.035000 5.905000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 77.440000 5.905000 77.760000 ;
      LAYER met4 ;
        RECT 5.585000 77.440000 5.905000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 77.845000 5.905000 78.165000 ;
      LAYER met4 ;
        RECT 5.585000 77.845000 5.905000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 78.250000 5.905000 78.570000 ;
      LAYER met4 ;
        RECT 5.585000 78.250000 5.905000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 78.655000 5.905000 78.975000 ;
      LAYER met4 ;
        RECT 5.585000 78.655000 5.905000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 79.060000 5.905000 79.380000 ;
      LAYER met4 ;
        RECT 5.585000 79.060000 5.905000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 79.465000 5.905000 79.785000 ;
      LAYER met4 ;
        RECT 5.585000 79.465000 5.905000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 79.870000 5.905000 80.190000 ;
      LAYER met4 ;
        RECT 5.585000 79.870000 5.905000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 80.275000 5.905000 80.595000 ;
      LAYER met4 ;
        RECT 5.585000 80.275000 5.905000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 80.680000 5.905000 81.000000 ;
      LAYER met4 ;
        RECT 5.585000 80.680000 5.905000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 81.085000 5.905000 81.405000 ;
      LAYER met4 ;
        RECT 5.585000 81.085000 5.905000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 81.490000 5.905000 81.810000 ;
      LAYER met4 ;
        RECT 5.585000 81.490000 5.905000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 81.895000 5.905000 82.215000 ;
      LAYER met4 ;
        RECT 5.585000 81.895000 5.905000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585000 82.300000 5.905000 82.620000 ;
      LAYER met4 ;
        RECT 5.585000 82.300000 5.905000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 82.795000 5.915000 83.115000 ;
      LAYER met4 ;
        RECT 5.595000 82.795000 5.915000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 83.205000 5.915000 83.525000 ;
      LAYER met4 ;
        RECT 5.595000 83.205000 5.915000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 83.615000 5.915000 83.935000 ;
      LAYER met4 ;
        RECT 5.595000 83.615000 5.915000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 84.025000 5.915000 84.345000 ;
      LAYER met4 ;
        RECT 5.595000 84.025000 5.915000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 84.435000 5.915000 84.755000 ;
      LAYER met4 ;
        RECT 5.595000 84.435000 5.915000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 84.845000 5.915000 85.165000 ;
      LAYER met4 ;
        RECT 5.595000 84.845000 5.915000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 85.255000 5.915000 85.575000 ;
      LAYER met4 ;
        RECT 5.595000 85.255000 5.915000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 85.665000 5.915000 85.985000 ;
      LAYER met4 ;
        RECT 5.595000 85.665000 5.915000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 86.075000 5.915000 86.395000 ;
      LAYER met4 ;
        RECT 5.595000 86.075000 5.915000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 86.485000 5.915000 86.805000 ;
      LAYER met4 ;
        RECT 5.595000 86.485000 5.915000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 86.895000 5.915000 87.215000 ;
      LAYER met4 ;
        RECT 5.595000 86.895000 5.915000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 87.305000 5.915000 87.625000 ;
      LAYER met4 ;
        RECT 5.595000 87.305000 5.915000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 87.715000 5.915000 88.035000 ;
      LAYER met4 ;
        RECT 5.595000 87.715000 5.915000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 88.125000 5.915000 88.445000 ;
      LAYER met4 ;
        RECT 5.595000 88.125000 5.915000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 88.535000 5.915000 88.855000 ;
      LAYER met4 ;
        RECT 5.595000 88.535000 5.915000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 88.945000 5.915000 89.265000 ;
      LAYER met4 ;
        RECT 5.595000 88.945000 5.915000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 89.355000 5.915000 89.675000 ;
      LAYER met4 ;
        RECT 5.595000 89.355000 5.915000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 89.765000 5.915000 90.085000 ;
      LAYER met4 ;
        RECT 5.595000 89.765000 5.915000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 90.175000 5.915000 90.495000 ;
      LAYER met4 ;
        RECT 5.595000 90.175000 5.915000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 90.585000 5.915000 90.905000 ;
      LAYER met4 ;
        RECT 5.595000 90.585000 5.915000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 90.995000 5.915000 91.315000 ;
      LAYER met4 ;
        RECT 5.595000 90.995000 5.915000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 91.405000 5.915000 91.725000 ;
      LAYER met4 ;
        RECT 5.595000 91.405000 5.915000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 91.815000 5.915000 92.135000 ;
      LAYER met4 ;
        RECT 5.595000 91.815000 5.915000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 92.225000 5.915000 92.545000 ;
      LAYER met4 ;
        RECT 5.595000 92.225000 5.915000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595000 92.635000 5.915000 92.955000 ;
      LAYER met4 ;
        RECT 5.595000 92.635000 5.915000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895000 17.800000 6.215000 18.120000 ;
      LAYER met4 ;
        RECT 5.895000 17.800000 6.215000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895000 18.230000 6.215000 18.550000 ;
      LAYER met4 ;
        RECT 5.895000 18.230000 6.215000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895000 18.660000 6.215000 18.980000 ;
      LAYER met4 ;
        RECT 5.895000 18.660000 6.215000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895000 19.090000 6.215000 19.410000 ;
      LAYER met4 ;
        RECT 5.895000 19.090000 6.215000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895000 19.520000 6.215000 19.840000 ;
      LAYER met4 ;
        RECT 5.895000 19.520000 6.215000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895000 19.950000 6.215000 20.270000 ;
      LAYER met4 ;
        RECT 5.895000 19.950000 6.215000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895000 20.380000 6.215000 20.700000 ;
      LAYER met4 ;
        RECT 5.895000 20.380000 6.215000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895000 20.810000 6.215000 21.130000 ;
      LAYER met4 ;
        RECT 5.895000 20.810000 6.215000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895000 21.240000 6.215000 21.560000 ;
      LAYER met4 ;
        RECT 5.895000 21.240000 6.215000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895000 21.670000 6.215000 21.990000 ;
      LAYER met4 ;
        RECT 5.895000 21.670000 6.215000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895000 22.100000 6.215000 22.420000 ;
      LAYER met4 ;
        RECT 5.895000 22.100000 6.215000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 68.065000 6.305000 68.385000 ;
      LAYER met4 ;
        RECT 5.985000 68.065000 6.305000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 68.475000 6.305000 68.795000 ;
      LAYER met4 ;
        RECT 5.985000 68.475000 6.305000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 68.885000 6.305000 69.205000 ;
      LAYER met4 ;
        RECT 5.985000 68.885000 6.305000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 69.295000 6.305000 69.615000 ;
      LAYER met4 ;
        RECT 5.985000 69.295000 6.305000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 69.705000 6.305000 70.025000 ;
      LAYER met4 ;
        RECT 5.985000 69.705000 6.305000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 70.115000 6.305000 70.435000 ;
      LAYER met4 ;
        RECT 5.985000 70.115000 6.305000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 70.525000 6.305000 70.845000 ;
      LAYER met4 ;
        RECT 5.985000 70.525000 6.305000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 70.935000 6.305000 71.255000 ;
      LAYER met4 ;
        RECT 5.985000 70.935000 6.305000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 71.345000 6.305000 71.665000 ;
      LAYER met4 ;
        RECT 5.985000 71.345000 6.305000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 71.755000 6.305000 72.075000 ;
      LAYER met4 ;
        RECT 5.985000 71.755000 6.305000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 72.165000 6.305000 72.485000 ;
      LAYER met4 ;
        RECT 5.985000 72.165000 6.305000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 72.575000 6.305000 72.895000 ;
      LAYER met4 ;
        RECT 5.985000 72.575000 6.305000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 72.985000 6.305000 73.305000 ;
      LAYER met4 ;
        RECT 5.985000 72.985000 6.305000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 73.390000 6.305000 73.710000 ;
      LAYER met4 ;
        RECT 5.985000 73.390000 6.305000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 73.795000 6.305000 74.115000 ;
      LAYER met4 ;
        RECT 5.985000 73.795000 6.305000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 74.200000 6.305000 74.520000 ;
      LAYER met4 ;
        RECT 5.985000 74.200000 6.305000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 74.605000 6.305000 74.925000 ;
      LAYER met4 ;
        RECT 5.985000 74.605000 6.305000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 75.010000 6.305000 75.330000 ;
      LAYER met4 ;
        RECT 5.985000 75.010000 6.305000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 75.415000 6.305000 75.735000 ;
      LAYER met4 ;
        RECT 5.985000 75.415000 6.305000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 75.820000 6.305000 76.140000 ;
      LAYER met4 ;
        RECT 5.985000 75.820000 6.305000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 76.225000 6.305000 76.545000 ;
      LAYER met4 ;
        RECT 5.985000 76.225000 6.305000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 76.630000 6.305000 76.950000 ;
      LAYER met4 ;
        RECT 5.985000 76.630000 6.305000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 77.035000 6.305000 77.355000 ;
      LAYER met4 ;
        RECT 5.985000 77.035000 6.305000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 77.440000 6.305000 77.760000 ;
      LAYER met4 ;
        RECT 5.985000 77.440000 6.305000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 77.845000 6.305000 78.165000 ;
      LAYER met4 ;
        RECT 5.985000 77.845000 6.305000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 78.250000 6.305000 78.570000 ;
      LAYER met4 ;
        RECT 5.985000 78.250000 6.305000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 78.655000 6.305000 78.975000 ;
      LAYER met4 ;
        RECT 5.985000 78.655000 6.305000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 79.060000 6.305000 79.380000 ;
      LAYER met4 ;
        RECT 5.985000 79.060000 6.305000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 79.465000 6.305000 79.785000 ;
      LAYER met4 ;
        RECT 5.985000 79.465000 6.305000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 79.870000 6.305000 80.190000 ;
      LAYER met4 ;
        RECT 5.985000 79.870000 6.305000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 80.275000 6.305000 80.595000 ;
      LAYER met4 ;
        RECT 5.985000 80.275000 6.305000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 80.680000 6.305000 81.000000 ;
      LAYER met4 ;
        RECT 5.985000 80.680000 6.305000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 81.085000 6.305000 81.405000 ;
      LAYER met4 ;
        RECT 5.985000 81.085000 6.305000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 81.490000 6.305000 81.810000 ;
      LAYER met4 ;
        RECT 5.985000 81.490000 6.305000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 81.895000 6.305000 82.215000 ;
      LAYER met4 ;
        RECT 5.985000 81.895000 6.305000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985000 82.300000 6.305000 82.620000 ;
      LAYER met4 ;
        RECT 5.985000 82.300000 6.305000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 17.800000 51.105000 18.120000 ;
      LAYER met4 ;
        RECT 50.785000 17.800000 51.105000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 18.230000 51.105000 18.550000 ;
      LAYER met4 ;
        RECT 50.785000 18.230000 51.105000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 18.660000 51.105000 18.980000 ;
      LAYER met4 ;
        RECT 50.785000 18.660000 51.105000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 19.090000 51.105000 19.410000 ;
      LAYER met4 ;
        RECT 50.785000 19.090000 51.105000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 19.520000 51.105000 19.840000 ;
      LAYER met4 ;
        RECT 50.785000 19.520000 51.105000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 19.950000 51.105000 20.270000 ;
      LAYER met4 ;
        RECT 50.785000 19.950000 51.105000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 20.380000 51.105000 20.700000 ;
      LAYER met4 ;
        RECT 50.785000 20.380000 51.105000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 20.810000 51.105000 21.130000 ;
      LAYER met4 ;
        RECT 50.785000 20.810000 51.105000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 21.240000 51.105000 21.560000 ;
      LAYER met4 ;
        RECT 50.785000 21.240000 51.105000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 21.670000 51.105000 21.990000 ;
      LAYER met4 ;
        RECT 50.785000 21.670000 51.105000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 22.100000 51.105000 22.420000 ;
      LAYER met4 ;
        RECT 50.785000 22.100000 51.105000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 68.065000 51.270000 68.385000 ;
      LAYER met4 ;
        RECT 50.950000 68.065000 51.270000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 68.475000 51.270000 68.795000 ;
      LAYER met4 ;
        RECT 50.950000 68.475000 51.270000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 68.885000 51.270000 69.205000 ;
      LAYER met4 ;
        RECT 50.950000 68.885000 51.270000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 69.295000 51.270000 69.615000 ;
      LAYER met4 ;
        RECT 50.950000 69.295000 51.270000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 69.705000 51.270000 70.025000 ;
      LAYER met4 ;
        RECT 50.950000 69.705000 51.270000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 70.115000 51.270000 70.435000 ;
      LAYER met4 ;
        RECT 50.950000 70.115000 51.270000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 70.525000 51.270000 70.845000 ;
      LAYER met4 ;
        RECT 50.950000 70.525000 51.270000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 70.935000 51.270000 71.255000 ;
      LAYER met4 ;
        RECT 50.950000 70.935000 51.270000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 71.345000 51.270000 71.665000 ;
      LAYER met4 ;
        RECT 50.950000 71.345000 51.270000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 71.755000 51.270000 72.075000 ;
      LAYER met4 ;
        RECT 50.950000 71.755000 51.270000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 72.165000 51.270000 72.485000 ;
      LAYER met4 ;
        RECT 50.950000 72.165000 51.270000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 72.575000 51.270000 72.895000 ;
      LAYER met4 ;
        RECT 50.950000 72.575000 51.270000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 72.985000 51.270000 73.305000 ;
      LAYER met4 ;
        RECT 50.950000 72.985000 51.270000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 73.390000 51.270000 73.710000 ;
      LAYER met4 ;
        RECT 50.950000 73.390000 51.270000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 73.795000 51.270000 74.115000 ;
      LAYER met4 ;
        RECT 50.950000 73.795000 51.270000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 74.200000 51.270000 74.520000 ;
      LAYER met4 ;
        RECT 50.950000 74.200000 51.270000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 74.605000 51.270000 74.925000 ;
      LAYER met4 ;
        RECT 50.950000 74.605000 51.270000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 75.010000 51.270000 75.330000 ;
      LAYER met4 ;
        RECT 50.950000 75.010000 51.270000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 75.415000 51.270000 75.735000 ;
      LAYER met4 ;
        RECT 50.950000 75.415000 51.270000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 75.820000 51.270000 76.140000 ;
      LAYER met4 ;
        RECT 50.950000 75.820000 51.270000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 76.225000 51.270000 76.545000 ;
      LAYER met4 ;
        RECT 50.950000 76.225000 51.270000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 76.630000 51.270000 76.950000 ;
      LAYER met4 ;
        RECT 50.950000 76.630000 51.270000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 77.035000 51.270000 77.355000 ;
      LAYER met4 ;
        RECT 50.950000 77.035000 51.270000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 77.440000 51.270000 77.760000 ;
      LAYER met4 ;
        RECT 50.950000 77.440000 51.270000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 77.845000 51.270000 78.165000 ;
      LAYER met4 ;
        RECT 50.950000 77.845000 51.270000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 78.250000 51.270000 78.570000 ;
      LAYER met4 ;
        RECT 50.950000 78.250000 51.270000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 78.655000 51.270000 78.975000 ;
      LAYER met4 ;
        RECT 50.950000 78.655000 51.270000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 79.060000 51.270000 79.380000 ;
      LAYER met4 ;
        RECT 50.950000 79.060000 51.270000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 79.465000 51.270000 79.785000 ;
      LAYER met4 ;
        RECT 50.950000 79.465000 51.270000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 79.870000 51.270000 80.190000 ;
      LAYER met4 ;
        RECT 50.950000 79.870000 51.270000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 80.275000 51.270000 80.595000 ;
      LAYER met4 ;
        RECT 50.950000 80.275000 51.270000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 80.680000 51.270000 81.000000 ;
      LAYER met4 ;
        RECT 50.950000 80.680000 51.270000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 81.085000 51.270000 81.405000 ;
      LAYER met4 ;
        RECT 50.950000 81.085000 51.270000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 81.490000 51.270000 81.810000 ;
      LAYER met4 ;
        RECT 50.950000 81.490000 51.270000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 81.895000 51.270000 82.215000 ;
      LAYER met4 ;
        RECT 50.950000 81.895000 51.270000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.950000 82.300000 51.270000 82.620000 ;
      LAYER met4 ;
        RECT 50.950000 82.300000 51.270000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.190000 17.800000 51.510000 18.120000 ;
      LAYER met4 ;
        RECT 51.190000 17.800000 51.510000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.190000 18.230000 51.510000 18.550000 ;
      LAYER met4 ;
        RECT 51.190000 18.230000 51.510000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.190000 18.660000 51.510000 18.980000 ;
      LAYER met4 ;
        RECT 51.190000 18.660000 51.510000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.190000 19.090000 51.510000 19.410000 ;
      LAYER met4 ;
        RECT 51.190000 19.090000 51.510000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.190000 19.520000 51.510000 19.840000 ;
      LAYER met4 ;
        RECT 51.190000 19.520000 51.510000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.190000 19.950000 51.510000 20.270000 ;
      LAYER met4 ;
        RECT 51.190000 19.950000 51.510000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.190000 20.380000 51.510000 20.700000 ;
      LAYER met4 ;
        RECT 51.190000 20.380000 51.510000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.190000 20.810000 51.510000 21.130000 ;
      LAYER met4 ;
        RECT 51.190000 20.810000 51.510000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.190000 21.240000 51.510000 21.560000 ;
      LAYER met4 ;
        RECT 51.190000 21.240000 51.510000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.190000 21.670000 51.510000 21.990000 ;
      LAYER met4 ;
        RECT 51.190000 21.670000 51.510000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.190000 22.100000 51.510000 22.420000 ;
      LAYER met4 ;
        RECT 51.190000 22.100000 51.510000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 68.065000 51.670000 68.385000 ;
      LAYER met4 ;
        RECT 51.350000 68.065000 51.670000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 68.475000 51.670000 68.795000 ;
      LAYER met4 ;
        RECT 51.350000 68.475000 51.670000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 68.885000 51.670000 69.205000 ;
      LAYER met4 ;
        RECT 51.350000 68.885000 51.670000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 69.295000 51.670000 69.615000 ;
      LAYER met4 ;
        RECT 51.350000 69.295000 51.670000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 69.705000 51.670000 70.025000 ;
      LAYER met4 ;
        RECT 51.350000 69.705000 51.670000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 70.115000 51.670000 70.435000 ;
      LAYER met4 ;
        RECT 51.350000 70.115000 51.670000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 70.525000 51.670000 70.845000 ;
      LAYER met4 ;
        RECT 51.350000 70.525000 51.670000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 70.935000 51.670000 71.255000 ;
      LAYER met4 ;
        RECT 51.350000 70.935000 51.670000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 71.345000 51.670000 71.665000 ;
      LAYER met4 ;
        RECT 51.350000 71.345000 51.670000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 71.755000 51.670000 72.075000 ;
      LAYER met4 ;
        RECT 51.350000 71.755000 51.670000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 72.165000 51.670000 72.485000 ;
      LAYER met4 ;
        RECT 51.350000 72.165000 51.670000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 72.575000 51.670000 72.895000 ;
      LAYER met4 ;
        RECT 51.350000 72.575000 51.670000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 72.985000 51.670000 73.305000 ;
      LAYER met4 ;
        RECT 51.350000 72.985000 51.670000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 73.390000 51.670000 73.710000 ;
      LAYER met4 ;
        RECT 51.350000 73.390000 51.670000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 73.795000 51.670000 74.115000 ;
      LAYER met4 ;
        RECT 51.350000 73.795000 51.670000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 74.200000 51.670000 74.520000 ;
      LAYER met4 ;
        RECT 51.350000 74.200000 51.670000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 74.605000 51.670000 74.925000 ;
      LAYER met4 ;
        RECT 51.350000 74.605000 51.670000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 75.010000 51.670000 75.330000 ;
      LAYER met4 ;
        RECT 51.350000 75.010000 51.670000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 75.415000 51.670000 75.735000 ;
      LAYER met4 ;
        RECT 51.350000 75.415000 51.670000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 75.820000 51.670000 76.140000 ;
      LAYER met4 ;
        RECT 51.350000 75.820000 51.670000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 76.225000 51.670000 76.545000 ;
      LAYER met4 ;
        RECT 51.350000 76.225000 51.670000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 76.630000 51.670000 76.950000 ;
      LAYER met4 ;
        RECT 51.350000 76.630000 51.670000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 77.035000 51.670000 77.355000 ;
      LAYER met4 ;
        RECT 51.350000 77.035000 51.670000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 77.440000 51.670000 77.760000 ;
      LAYER met4 ;
        RECT 51.350000 77.440000 51.670000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 77.845000 51.670000 78.165000 ;
      LAYER met4 ;
        RECT 51.350000 77.845000 51.670000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 78.250000 51.670000 78.570000 ;
      LAYER met4 ;
        RECT 51.350000 78.250000 51.670000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 78.655000 51.670000 78.975000 ;
      LAYER met4 ;
        RECT 51.350000 78.655000 51.670000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 79.060000 51.670000 79.380000 ;
      LAYER met4 ;
        RECT 51.350000 79.060000 51.670000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 79.465000 51.670000 79.785000 ;
      LAYER met4 ;
        RECT 51.350000 79.465000 51.670000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 79.870000 51.670000 80.190000 ;
      LAYER met4 ;
        RECT 51.350000 79.870000 51.670000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 80.275000 51.670000 80.595000 ;
      LAYER met4 ;
        RECT 51.350000 80.275000 51.670000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 80.680000 51.670000 81.000000 ;
      LAYER met4 ;
        RECT 51.350000 80.680000 51.670000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 81.085000 51.670000 81.405000 ;
      LAYER met4 ;
        RECT 51.350000 81.085000 51.670000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 81.490000 51.670000 81.810000 ;
      LAYER met4 ;
        RECT 51.350000 81.490000 51.670000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 81.895000 51.670000 82.215000 ;
      LAYER met4 ;
        RECT 51.350000 81.895000 51.670000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.350000 82.300000 51.670000 82.620000 ;
      LAYER met4 ;
        RECT 51.350000 82.300000 51.670000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.595000 17.800000 51.915000 18.120000 ;
      LAYER met4 ;
        RECT 51.595000 17.800000 51.915000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.595000 18.230000 51.915000 18.550000 ;
      LAYER met4 ;
        RECT 51.595000 18.230000 51.915000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.595000 18.660000 51.915000 18.980000 ;
      LAYER met4 ;
        RECT 51.595000 18.660000 51.915000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.595000 19.090000 51.915000 19.410000 ;
      LAYER met4 ;
        RECT 51.595000 19.090000 51.915000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.595000 19.520000 51.915000 19.840000 ;
      LAYER met4 ;
        RECT 51.595000 19.520000 51.915000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.595000 19.950000 51.915000 20.270000 ;
      LAYER met4 ;
        RECT 51.595000 19.950000 51.915000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.595000 20.380000 51.915000 20.700000 ;
      LAYER met4 ;
        RECT 51.595000 20.380000 51.915000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.595000 20.810000 51.915000 21.130000 ;
      LAYER met4 ;
        RECT 51.595000 20.810000 51.915000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.595000 21.240000 51.915000 21.560000 ;
      LAYER met4 ;
        RECT 51.595000 21.240000 51.915000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.595000 21.670000 51.915000 21.990000 ;
      LAYER met4 ;
        RECT 51.595000 21.670000 51.915000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.595000 22.100000 51.915000 22.420000 ;
      LAYER met4 ;
        RECT 51.595000 22.100000 51.915000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 68.065000 52.070000 68.385000 ;
      LAYER met4 ;
        RECT 51.750000 68.065000 52.070000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 68.475000 52.070000 68.795000 ;
      LAYER met4 ;
        RECT 51.750000 68.475000 52.070000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 68.885000 52.070000 69.205000 ;
      LAYER met4 ;
        RECT 51.750000 68.885000 52.070000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 69.295000 52.070000 69.615000 ;
      LAYER met4 ;
        RECT 51.750000 69.295000 52.070000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 69.705000 52.070000 70.025000 ;
      LAYER met4 ;
        RECT 51.750000 69.705000 52.070000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 70.115000 52.070000 70.435000 ;
      LAYER met4 ;
        RECT 51.750000 70.115000 52.070000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 70.525000 52.070000 70.845000 ;
      LAYER met4 ;
        RECT 51.750000 70.525000 52.070000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 70.935000 52.070000 71.255000 ;
      LAYER met4 ;
        RECT 51.750000 70.935000 52.070000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 71.345000 52.070000 71.665000 ;
      LAYER met4 ;
        RECT 51.750000 71.345000 52.070000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 71.755000 52.070000 72.075000 ;
      LAYER met4 ;
        RECT 51.750000 71.755000 52.070000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 72.165000 52.070000 72.485000 ;
      LAYER met4 ;
        RECT 51.750000 72.165000 52.070000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 72.575000 52.070000 72.895000 ;
      LAYER met4 ;
        RECT 51.750000 72.575000 52.070000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 72.985000 52.070000 73.305000 ;
      LAYER met4 ;
        RECT 51.750000 72.985000 52.070000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 73.390000 52.070000 73.710000 ;
      LAYER met4 ;
        RECT 51.750000 73.390000 52.070000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 73.795000 52.070000 74.115000 ;
      LAYER met4 ;
        RECT 51.750000 73.795000 52.070000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 74.200000 52.070000 74.520000 ;
      LAYER met4 ;
        RECT 51.750000 74.200000 52.070000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 74.605000 52.070000 74.925000 ;
      LAYER met4 ;
        RECT 51.750000 74.605000 52.070000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 75.010000 52.070000 75.330000 ;
      LAYER met4 ;
        RECT 51.750000 75.010000 52.070000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 75.415000 52.070000 75.735000 ;
      LAYER met4 ;
        RECT 51.750000 75.415000 52.070000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 75.820000 52.070000 76.140000 ;
      LAYER met4 ;
        RECT 51.750000 75.820000 52.070000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 76.225000 52.070000 76.545000 ;
      LAYER met4 ;
        RECT 51.750000 76.225000 52.070000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 76.630000 52.070000 76.950000 ;
      LAYER met4 ;
        RECT 51.750000 76.630000 52.070000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 77.035000 52.070000 77.355000 ;
      LAYER met4 ;
        RECT 51.750000 77.035000 52.070000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 77.440000 52.070000 77.760000 ;
      LAYER met4 ;
        RECT 51.750000 77.440000 52.070000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 77.845000 52.070000 78.165000 ;
      LAYER met4 ;
        RECT 51.750000 77.845000 52.070000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 78.250000 52.070000 78.570000 ;
      LAYER met4 ;
        RECT 51.750000 78.250000 52.070000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 78.655000 52.070000 78.975000 ;
      LAYER met4 ;
        RECT 51.750000 78.655000 52.070000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 79.060000 52.070000 79.380000 ;
      LAYER met4 ;
        RECT 51.750000 79.060000 52.070000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 79.465000 52.070000 79.785000 ;
      LAYER met4 ;
        RECT 51.750000 79.465000 52.070000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 79.870000 52.070000 80.190000 ;
      LAYER met4 ;
        RECT 51.750000 79.870000 52.070000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 80.275000 52.070000 80.595000 ;
      LAYER met4 ;
        RECT 51.750000 80.275000 52.070000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 80.680000 52.070000 81.000000 ;
      LAYER met4 ;
        RECT 51.750000 80.680000 52.070000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 81.085000 52.070000 81.405000 ;
      LAYER met4 ;
        RECT 51.750000 81.085000 52.070000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 81.490000 52.070000 81.810000 ;
      LAYER met4 ;
        RECT 51.750000 81.490000 52.070000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 81.895000 52.070000 82.215000 ;
      LAYER met4 ;
        RECT 51.750000 81.895000 52.070000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.750000 82.300000 52.070000 82.620000 ;
      LAYER met4 ;
        RECT 51.750000 82.300000 52.070000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.000000 17.800000 52.320000 18.120000 ;
      LAYER met4 ;
        RECT 52.000000 17.800000 52.320000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.000000 18.230000 52.320000 18.550000 ;
      LAYER met4 ;
        RECT 52.000000 18.230000 52.320000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.000000 18.660000 52.320000 18.980000 ;
      LAYER met4 ;
        RECT 52.000000 18.660000 52.320000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.000000 19.090000 52.320000 19.410000 ;
      LAYER met4 ;
        RECT 52.000000 19.090000 52.320000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.000000 19.520000 52.320000 19.840000 ;
      LAYER met4 ;
        RECT 52.000000 19.520000 52.320000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.000000 19.950000 52.320000 20.270000 ;
      LAYER met4 ;
        RECT 52.000000 19.950000 52.320000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.000000 20.380000 52.320000 20.700000 ;
      LAYER met4 ;
        RECT 52.000000 20.380000 52.320000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.000000 20.810000 52.320000 21.130000 ;
      LAYER met4 ;
        RECT 52.000000 20.810000 52.320000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.000000 21.240000 52.320000 21.560000 ;
      LAYER met4 ;
        RECT 52.000000 21.240000 52.320000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.000000 21.670000 52.320000 21.990000 ;
      LAYER met4 ;
        RECT 52.000000 21.670000 52.320000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.000000 22.100000 52.320000 22.420000 ;
      LAYER met4 ;
        RECT 52.000000 22.100000 52.320000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 68.065000 52.470000 68.385000 ;
      LAYER met4 ;
        RECT 52.150000 68.065000 52.470000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 68.475000 52.470000 68.795000 ;
      LAYER met4 ;
        RECT 52.150000 68.475000 52.470000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 68.885000 52.470000 69.205000 ;
      LAYER met4 ;
        RECT 52.150000 68.885000 52.470000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 69.295000 52.470000 69.615000 ;
      LAYER met4 ;
        RECT 52.150000 69.295000 52.470000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 69.705000 52.470000 70.025000 ;
      LAYER met4 ;
        RECT 52.150000 69.705000 52.470000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 70.115000 52.470000 70.435000 ;
      LAYER met4 ;
        RECT 52.150000 70.115000 52.470000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 70.525000 52.470000 70.845000 ;
      LAYER met4 ;
        RECT 52.150000 70.525000 52.470000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 70.935000 52.470000 71.255000 ;
      LAYER met4 ;
        RECT 52.150000 70.935000 52.470000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 71.345000 52.470000 71.665000 ;
      LAYER met4 ;
        RECT 52.150000 71.345000 52.470000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 71.755000 52.470000 72.075000 ;
      LAYER met4 ;
        RECT 52.150000 71.755000 52.470000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 72.165000 52.470000 72.485000 ;
      LAYER met4 ;
        RECT 52.150000 72.165000 52.470000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 72.575000 52.470000 72.895000 ;
      LAYER met4 ;
        RECT 52.150000 72.575000 52.470000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 72.985000 52.470000 73.305000 ;
      LAYER met4 ;
        RECT 52.150000 72.985000 52.470000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 73.390000 52.470000 73.710000 ;
      LAYER met4 ;
        RECT 52.150000 73.390000 52.470000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 73.795000 52.470000 74.115000 ;
      LAYER met4 ;
        RECT 52.150000 73.795000 52.470000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 74.200000 52.470000 74.520000 ;
      LAYER met4 ;
        RECT 52.150000 74.200000 52.470000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 74.605000 52.470000 74.925000 ;
      LAYER met4 ;
        RECT 52.150000 74.605000 52.470000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 75.010000 52.470000 75.330000 ;
      LAYER met4 ;
        RECT 52.150000 75.010000 52.470000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 75.415000 52.470000 75.735000 ;
      LAYER met4 ;
        RECT 52.150000 75.415000 52.470000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 75.820000 52.470000 76.140000 ;
      LAYER met4 ;
        RECT 52.150000 75.820000 52.470000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 76.225000 52.470000 76.545000 ;
      LAYER met4 ;
        RECT 52.150000 76.225000 52.470000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 76.630000 52.470000 76.950000 ;
      LAYER met4 ;
        RECT 52.150000 76.630000 52.470000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 77.035000 52.470000 77.355000 ;
      LAYER met4 ;
        RECT 52.150000 77.035000 52.470000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 77.440000 52.470000 77.760000 ;
      LAYER met4 ;
        RECT 52.150000 77.440000 52.470000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 77.845000 52.470000 78.165000 ;
      LAYER met4 ;
        RECT 52.150000 77.845000 52.470000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 78.250000 52.470000 78.570000 ;
      LAYER met4 ;
        RECT 52.150000 78.250000 52.470000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 78.655000 52.470000 78.975000 ;
      LAYER met4 ;
        RECT 52.150000 78.655000 52.470000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 79.060000 52.470000 79.380000 ;
      LAYER met4 ;
        RECT 52.150000 79.060000 52.470000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 79.465000 52.470000 79.785000 ;
      LAYER met4 ;
        RECT 52.150000 79.465000 52.470000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 79.870000 52.470000 80.190000 ;
      LAYER met4 ;
        RECT 52.150000 79.870000 52.470000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 80.275000 52.470000 80.595000 ;
      LAYER met4 ;
        RECT 52.150000 80.275000 52.470000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 80.680000 52.470000 81.000000 ;
      LAYER met4 ;
        RECT 52.150000 80.680000 52.470000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 81.085000 52.470000 81.405000 ;
      LAYER met4 ;
        RECT 52.150000 81.085000 52.470000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 81.490000 52.470000 81.810000 ;
      LAYER met4 ;
        RECT 52.150000 81.490000 52.470000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 81.895000 52.470000 82.215000 ;
      LAYER met4 ;
        RECT 52.150000 81.895000 52.470000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.150000 82.300000 52.470000 82.620000 ;
      LAYER met4 ;
        RECT 52.150000 82.300000 52.470000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 17.800000 52.725000 18.120000 ;
      LAYER met4 ;
        RECT 52.405000 17.800000 52.725000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 18.230000 52.725000 18.550000 ;
      LAYER met4 ;
        RECT 52.405000 18.230000 52.725000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 18.660000 52.725000 18.980000 ;
      LAYER met4 ;
        RECT 52.405000 18.660000 52.725000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 19.090000 52.725000 19.410000 ;
      LAYER met4 ;
        RECT 52.405000 19.090000 52.725000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 19.520000 52.725000 19.840000 ;
      LAYER met4 ;
        RECT 52.405000 19.520000 52.725000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 19.950000 52.725000 20.270000 ;
      LAYER met4 ;
        RECT 52.405000 19.950000 52.725000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 20.380000 52.725000 20.700000 ;
      LAYER met4 ;
        RECT 52.405000 20.380000 52.725000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 20.810000 52.725000 21.130000 ;
      LAYER met4 ;
        RECT 52.405000 20.810000 52.725000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 21.240000 52.725000 21.560000 ;
      LAYER met4 ;
        RECT 52.405000 21.240000 52.725000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 21.670000 52.725000 21.990000 ;
      LAYER met4 ;
        RECT 52.405000 21.670000 52.725000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 22.100000 52.725000 22.420000 ;
      LAYER met4 ;
        RECT 52.405000 22.100000 52.725000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.490000 82.860000 52.810000 83.180000 ;
      LAYER met4 ;
        RECT 52.490000 82.860000 52.810000 83.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.490000 83.410000 52.810000 83.730000 ;
      LAYER met4 ;
        RECT 52.490000 83.410000 52.810000 83.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.490000 83.960000 52.810000 84.280000 ;
      LAYER met4 ;
        RECT 52.490000 83.960000 52.810000 84.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 68.065000 52.870000 68.385000 ;
      LAYER met4 ;
        RECT 52.550000 68.065000 52.870000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 68.475000 52.870000 68.795000 ;
      LAYER met4 ;
        RECT 52.550000 68.475000 52.870000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 68.885000 52.870000 69.205000 ;
      LAYER met4 ;
        RECT 52.550000 68.885000 52.870000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 69.295000 52.870000 69.615000 ;
      LAYER met4 ;
        RECT 52.550000 69.295000 52.870000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 69.705000 52.870000 70.025000 ;
      LAYER met4 ;
        RECT 52.550000 69.705000 52.870000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 70.115000 52.870000 70.435000 ;
      LAYER met4 ;
        RECT 52.550000 70.115000 52.870000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 70.525000 52.870000 70.845000 ;
      LAYER met4 ;
        RECT 52.550000 70.525000 52.870000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 70.935000 52.870000 71.255000 ;
      LAYER met4 ;
        RECT 52.550000 70.935000 52.870000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 71.345000 52.870000 71.665000 ;
      LAYER met4 ;
        RECT 52.550000 71.345000 52.870000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 71.755000 52.870000 72.075000 ;
      LAYER met4 ;
        RECT 52.550000 71.755000 52.870000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 72.165000 52.870000 72.485000 ;
      LAYER met4 ;
        RECT 52.550000 72.165000 52.870000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 72.575000 52.870000 72.895000 ;
      LAYER met4 ;
        RECT 52.550000 72.575000 52.870000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 72.985000 52.870000 73.305000 ;
      LAYER met4 ;
        RECT 52.550000 72.985000 52.870000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 73.390000 52.870000 73.710000 ;
      LAYER met4 ;
        RECT 52.550000 73.390000 52.870000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 73.795000 52.870000 74.115000 ;
      LAYER met4 ;
        RECT 52.550000 73.795000 52.870000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 74.200000 52.870000 74.520000 ;
      LAYER met4 ;
        RECT 52.550000 74.200000 52.870000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 74.605000 52.870000 74.925000 ;
      LAYER met4 ;
        RECT 52.550000 74.605000 52.870000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 75.010000 52.870000 75.330000 ;
      LAYER met4 ;
        RECT 52.550000 75.010000 52.870000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 75.415000 52.870000 75.735000 ;
      LAYER met4 ;
        RECT 52.550000 75.415000 52.870000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 75.820000 52.870000 76.140000 ;
      LAYER met4 ;
        RECT 52.550000 75.820000 52.870000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 76.225000 52.870000 76.545000 ;
      LAYER met4 ;
        RECT 52.550000 76.225000 52.870000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 76.630000 52.870000 76.950000 ;
      LAYER met4 ;
        RECT 52.550000 76.630000 52.870000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 77.035000 52.870000 77.355000 ;
      LAYER met4 ;
        RECT 52.550000 77.035000 52.870000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 77.440000 52.870000 77.760000 ;
      LAYER met4 ;
        RECT 52.550000 77.440000 52.870000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 77.845000 52.870000 78.165000 ;
      LAYER met4 ;
        RECT 52.550000 77.845000 52.870000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 78.250000 52.870000 78.570000 ;
      LAYER met4 ;
        RECT 52.550000 78.250000 52.870000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 78.655000 52.870000 78.975000 ;
      LAYER met4 ;
        RECT 52.550000 78.655000 52.870000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 79.060000 52.870000 79.380000 ;
      LAYER met4 ;
        RECT 52.550000 79.060000 52.870000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 79.465000 52.870000 79.785000 ;
      LAYER met4 ;
        RECT 52.550000 79.465000 52.870000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 79.870000 52.870000 80.190000 ;
      LAYER met4 ;
        RECT 52.550000 79.870000 52.870000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 80.275000 52.870000 80.595000 ;
      LAYER met4 ;
        RECT 52.550000 80.275000 52.870000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 80.680000 52.870000 81.000000 ;
      LAYER met4 ;
        RECT 52.550000 80.680000 52.870000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 81.085000 52.870000 81.405000 ;
      LAYER met4 ;
        RECT 52.550000 81.085000 52.870000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 81.490000 52.870000 81.810000 ;
      LAYER met4 ;
        RECT 52.550000 81.490000 52.870000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 81.895000 52.870000 82.215000 ;
      LAYER met4 ;
        RECT 52.550000 81.895000 52.870000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.550000 82.300000 52.870000 82.620000 ;
      LAYER met4 ;
        RECT 52.550000 82.300000 52.870000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.810000 17.800000 53.130000 18.120000 ;
      LAYER met4 ;
        RECT 52.810000 17.800000 53.130000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.810000 18.230000 53.130000 18.550000 ;
      LAYER met4 ;
        RECT 52.810000 18.230000 53.130000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.810000 18.660000 53.130000 18.980000 ;
      LAYER met4 ;
        RECT 52.810000 18.660000 53.130000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.810000 19.090000 53.130000 19.410000 ;
      LAYER met4 ;
        RECT 52.810000 19.090000 53.130000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.810000 19.520000 53.130000 19.840000 ;
      LAYER met4 ;
        RECT 52.810000 19.520000 53.130000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.810000 19.950000 53.130000 20.270000 ;
      LAYER met4 ;
        RECT 52.810000 19.950000 53.130000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.810000 20.380000 53.130000 20.700000 ;
      LAYER met4 ;
        RECT 52.810000 20.380000 53.130000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.810000 20.810000 53.130000 21.130000 ;
      LAYER met4 ;
        RECT 52.810000 20.810000 53.130000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.810000 21.240000 53.130000 21.560000 ;
      LAYER met4 ;
        RECT 52.810000 21.240000 53.130000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.810000 21.670000 53.130000 21.990000 ;
      LAYER met4 ;
        RECT 52.810000 21.670000 53.130000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.810000 22.100000 53.130000 22.420000 ;
      LAYER met4 ;
        RECT 52.810000 22.100000 53.130000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 68.065000 53.270000 68.385000 ;
      LAYER met4 ;
        RECT 52.950000 68.065000 53.270000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 68.475000 53.270000 68.795000 ;
      LAYER met4 ;
        RECT 52.950000 68.475000 53.270000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 68.885000 53.270000 69.205000 ;
      LAYER met4 ;
        RECT 52.950000 68.885000 53.270000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 69.295000 53.270000 69.615000 ;
      LAYER met4 ;
        RECT 52.950000 69.295000 53.270000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 69.705000 53.270000 70.025000 ;
      LAYER met4 ;
        RECT 52.950000 69.705000 53.270000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 70.115000 53.270000 70.435000 ;
      LAYER met4 ;
        RECT 52.950000 70.115000 53.270000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 70.525000 53.270000 70.845000 ;
      LAYER met4 ;
        RECT 52.950000 70.525000 53.270000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 70.935000 53.270000 71.255000 ;
      LAYER met4 ;
        RECT 52.950000 70.935000 53.270000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 71.345000 53.270000 71.665000 ;
      LAYER met4 ;
        RECT 52.950000 71.345000 53.270000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 71.755000 53.270000 72.075000 ;
      LAYER met4 ;
        RECT 52.950000 71.755000 53.270000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 72.165000 53.270000 72.485000 ;
      LAYER met4 ;
        RECT 52.950000 72.165000 53.270000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 72.575000 53.270000 72.895000 ;
      LAYER met4 ;
        RECT 52.950000 72.575000 53.270000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 72.985000 53.270000 73.305000 ;
      LAYER met4 ;
        RECT 52.950000 72.985000 53.270000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 73.390000 53.270000 73.710000 ;
      LAYER met4 ;
        RECT 52.950000 73.390000 53.270000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 73.795000 53.270000 74.115000 ;
      LAYER met4 ;
        RECT 52.950000 73.795000 53.270000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 74.200000 53.270000 74.520000 ;
      LAYER met4 ;
        RECT 52.950000 74.200000 53.270000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 74.605000 53.270000 74.925000 ;
      LAYER met4 ;
        RECT 52.950000 74.605000 53.270000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 75.010000 53.270000 75.330000 ;
      LAYER met4 ;
        RECT 52.950000 75.010000 53.270000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 75.415000 53.270000 75.735000 ;
      LAYER met4 ;
        RECT 52.950000 75.415000 53.270000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 75.820000 53.270000 76.140000 ;
      LAYER met4 ;
        RECT 52.950000 75.820000 53.270000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 76.225000 53.270000 76.545000 ;
      LAYER met4 ;
        RECT 52.950000 76.225000 53.270000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 76.630000 53.270000 76.950000 ;
      LAYER met4 ;
        RECT 52.950000 76.630000 53.270000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 77.035000 53.270000 77.355000 ;
      LAYER met4 ;
        RECT 52.950000 77.035000 53.270000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 77.440000 53.270000 77.760000 ;
      LAYER met4 ;
        RECT 52.950000 77.440000 53.270000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 77.845000 53.270000 78.165000 ;
      LAYER met4 ;
        RECT 52.950000 77.845000 53.270000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 78.250000 53.270000 78.570000 ;
      LAYER met4 ;
        RECT 52.950000 78.250000 53.270000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 78.655000 53.270000 78.975000 ;
      LAYER met4 ;
        RECT 52.950000 78.655000 53.270000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 79.060000 53.270000 79.380000 ;
      LAYER met4 ;
        RECT 52.950000 79.060000 53.270000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 79.465000 53.270000 79.785000 ;
      LAYER met4 ;
        RECT 52.950000 79.465000 53.270000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 79.870000 53.270000 80.190000 ;
      LAYER met4 ;
        RECT 52.950000 79.870000 53.270000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 80.275000 53.270000 80.595000 ;
      LAYER met4 ;
        RECT 52.950000 80.275000 53.270000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 80.680000 53.270000 81.000000 ;
      LAYER met4 ;
        RECT 52.950000 80.680000 53.270000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 81.085000 53.270000 81.405000 ;
      LAYER met4 ;
        RECT 52.950000 81.085000 53.270000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 81.490000 53.270000 81.810000 ;
      LAYER met4 ;
        RECT 52.950000 81.490000 53.270000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 81.895000 53.270000 82.215000 ;
      LAYER met4 ;
        RECT 52.950000 81.895000 53.270000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.950000 82.300000 53.270000 82.620000 ;
      LAYER met4 ;
        RECT 52.950000 82.300000 53.270000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.215000 17.800000 53.535000 18.120000 ;
      LAYER met4 ;
        RECT 53.215000 17.800000 53.535000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.215000 18.230000 53.535000 18.550000 ;
      LAYER met4 ;
        RECT 53.215000 18.230000 53.535000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.215000 18.660000 53.535000 18.980000 ;
      LAYER met4 ;
        RECT 53.215000 18.660000 53.535000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.215000 19.090000 53.535000 19.410000 ;
      LAYER met4 ;
        RECT 53.215000 19.090000 53.535000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.215000 19.520000 53.535000 19.840000 ;
      LAYER met4 ;
        RECT 53.215000 19.520000 53.535000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.215000 19.950000 53.535000 20.270000 ;
      LAYER met4 ;
        RECT 53.215000 19.950000 53.535000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.215000 20.380000 53.535000 20.700000 ;
      LAYER met4 ;
        RECT 53.215000 20.380000 53.535000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.215000 20.810000 53.535000 21.130000 ;
      LAYER met4 ;
        RECT 53.215000 20.810000 53.535000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.215000 21.240000 53.535000 21.560000 ;
      LAYER met4 ;
        RECT 53.215000 21.240000 53.535000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.215000 21.670000 53.535000 21.990000 ;
      LAYER met4 ;
        RECT 53.215000 21.670000 53.535000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.215000 22.100000 53.535000 22.420000 ;
      LAYER met4 ;
        RECT 53.215000 22.100000 53.535000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.280000 82.860000 53.600000 83.180000 ;
      LAYER met4 ;
        RECT 53.280000 82.860000 53.600000 83.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.280000 83.410000 53.600000 83.730000 ;
      LAYER met4 ;
        RECT 53.280000 83.410000 53.600000 83.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.280000 83.960000 53.600000 84.280000 ;
      LAYER met4 ;
        RECT 53.280000 83.960000 53.600000 84.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 68.065000 53.670000 68.385000 ;
      LAYER met4 ;
        RECT 53.350000 68.065000 53.670000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 68.475000 53.670000 68.795000 ;
      LAYER met4 ;
        RECT 53.350000 68.475000 53.670000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 68.885000 53.670000 69.205000 ;
      LAYER met4 ;
        RECT 53.350000 68.885000 53.670000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 69.295000 53.670000 69.615000 ;
      LAYER met4 ;
        RECT 53.350000 69.295000 53.670000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 69.705000 53.670000 70.025000 ;
      LAYER met4 ;
        RECT 53.350000 69.705000 53.670000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 70.115000 53.670000 70.435000 ;
      LAYER met4 ;
        RECT 53.350000 70.115000 53.670000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 70.525000 53.670000 70.845000 ;
      LAYER met4 ;
        RECT 53.350000 70.525000 53.670000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 70.935000 53.670000 71.255000 ;
      LAYER met4 ;
        RECT 53.350000 70.935000 53.670000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 71.345000 53.670000 71.665000 ;
      LAYER met4 ;
        RECT 53.350000 71.345000 53.670000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 71.755000 53.670000 72.075000 ;
      LAYER met4 ;
        RECT 53.350000 71.755000 53.670000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 72.165000 53.670000 72.485000 ;
      LAYER met4 ;
        RECT 53.350000 72.165000 53.670000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 72.575000 53.670000 72.895000 ;
      LAYER met4 ;
        RECT 53.350000 72.575000 53.670000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 72.985000 53.670000 73.305000 ;
      LAYER met4 ;
        RECT 53.350000 72.985000 53.670000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 73.390000 53.670000 73.710000 ;
      LAYER met4 ;
        RECT 53.350000 73.390000 53.670000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 73.795000 53.670000 74.115000 ;
      LAYER met4 ;
        RECT 53.350000 73.795000 53.670000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 74.200000 53.670000 74.520000 ;
      LAYER met4 ;
        RECT 53.350000 74.200000 53.670000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 74.605000 53.670000 74.925000 ;
      LAYER met4 ;
        RECT 53.350000 74.605000 53.670000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 75.010000 53.670000 75.330000 ;
      LAYER met4 ;
        RECT 53.350000 75.010000 53.670000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 75.415000 53.670000 75.735000 ;
      LAYER met4 ;
        RECT 53.350000 75.415000 53.670000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 75.820000 53.670000 76.140000 ;
      LAYER met4 ;
        RECT 53.350000 75.820000 53.670000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 76.225000 53.670000 76.545000 ;
      LAYER met4 ;
        RECT 53.350000 76.225000 53.670000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 76.630000 53.670000 76.950000 ;
      LAYER met4 ;
        RECT 53.350000 76.630000 53.670000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 77.035000 53.670000 77.355000 ;
      LAYER met4 ;
        RECT 53.350000 77.035000 53.670000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 77.440000 53.670000 77.760000 ;
      LAYER met4 ;
        RECT 53.350000 77.440000 53.670000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 77.845000 53.670000 78.165000 ;
      LAYER met4 ;
        RECT 53.350000 77.845000 53.670000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 78.250000 53.670000 78.570000 ;
      LAYER met4 ;
        RECT 53.350000 78.250000 53.670000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 78.655000 53.670000 78.975000 ;
      LAYER met4 ;
        RECT 53.350000 78.655000 53.670000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 79.060000 53.670000 79.380000 ;
      LAYER met4 ;
        RECT 53.350000 79.060000 53.670000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 79.465000 53.670000 79.785000 ;
      LAYER met4 ;
        RECT 53.350000 79.465000 53.670000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 79.870000 53.670000 80.190000 ;
      LAYER met4 ;
        RECT 53.350000 79.870000 53.670000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 80.275000 53.670000 80.595000 ;
      LAYER met4 ;
        RECT 53.350000 80.275000 53.670000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 80.680000 53.670000 81.000000 ;
      LAYER met4 ;
        RECT 53.350000 80.680000 53.670000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 81.085000 53.670000 81.405000 ;
      LAYER met4 ;
        RECT 53.350000 81.085000 53.670000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 81.490000 53.670000 81.810000 ;
      LAYER met4 ;
        RECT 53.350000 81.490000 53.670000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 81.895000 53.670000 82.215000 ;
      LAYER met4 ;
        RECT 53.350000 81.895000 53.670000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.350000 82.300000 53.670000 82.620000 ;
      LAYER met4 ;
        RECT 53.350000 82.300000 53.670000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.620000 17.800000 53.940000 18.120000 ;
      LAYER met4 ;
        RECT 53.620000 17.800000 53.940000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.620000 18.230000 53.940000 18.550000 ;
      LAYER met4 ;
        RECT 53.620000 18.230000 53.940000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.620000 18.660000 53.940000 18.980000 ;
      LAYER met4 ;
        RECT 53.620000 18.660000 53.940000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.620000 19.090000 53.940000 19.410000 ;
      LAYER met4 ;
        RECT 53.620000 19.090000 53.940000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.620000 19.520000 53.940000 19.840000 ;
      LAYER met4 ;
        RECT 53.620000 19.520000 53.940000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.620000 19.950000 53.940000 20.270000 ;
      LAYER met4 ;
        RECT 53.620000 19.950000 53.940000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.620000 20.380000 53.940000 20.700000 ;
      LAYER met4 ;
        RECT 53.620000 20.380000 53.940000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.620000 20.810000 53.940000 21.130000 ;
      LAYER met4 ;
        RECT 53.620000 20.810000 53.940000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.620000 21.240000 53.940000 21.560000 ;
      LAYER met4 ;
        RECT 53.620000 21.240000 53.940000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.620000 21.670000 53.940000 21.990000 ;
      LAYER met4 ;
        RECT 53.620000 21.670000 53.940000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.620000 22.100000 53.940000 22.420000 ;
      LAYER met4 ;
        RECT 53.620000 22.100000 53.940000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 68.065000 54.070000 68.385000 ;
      LAYER met4 ;
        RECT 53.750000 68.065000 54.070000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 68.475000 54.070000 68.795000 ;
      LAYER met4 ;
        RECT 53.750000 68.475000 54.070000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 68.885000 54.070000 69.205000 ;
      LAYER met4 ;
        RECT 53.750000 68.885000 54.070000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 69.295000 54.070000 69.615000 ;
      LAYER met4 ;
        RECT 53.750000 69.295000 54.070000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 69.705000 54.070000 70.025000 ;
      LAYER met4 ;
        RECT 53.750000 69.705000 54.070000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 70.115000 54.070000 70.435000 ;
      LAYER met4 ;
        RECT 53.750000 70.115000 54.070000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 70.525000 54.070000 70.845000 ;
      LAYER met4 ;
        RECT 53.750000 70.525000 54.070000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 70.935000 54.070000 71.255000 ;
      LAYER met4 ;
        RECT 53.750000 70.935000 54.070000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 71.345000 54.070000 71.665000 ;
      LAYER met4 ;
        RECT 53.750000 71.345000 54.070000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 71.755000 54.070000 72.075000 ;
      LAYER met4 ;
        RECT 53.750000 71.755000 54.070000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 72.165000 54.070000 72.485000 ;
      LAYER met4 ;
        RECT 53.750000 72.165000 54.070000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 72.575000 54.070000 72.895000 ;
      LAYER met4 ;
        RECT 53.750000 72.575000 54.070000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 72.985000 54.070000 73.305000 ;
      LAYER met4 ;
        RECT 53.750000 72.985000 54.070000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 73.390000 54.070000 73.710000 ;
      LAYER met4 ;
        RECT 53.750000 73.390000 54.070000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 73.795000 54.070000 74.115000 ;
      LAYER met4 ;
        RECT 53.750000 73.795000 54.070000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 74.200000 54.070000 74.520000 ;
      LAYER met4 ;
        RECT 53.750000 74.200000 54.070000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 74.605000 54.070000 74.925000 ;
      LAYER met4 ;
        RECT 53.750000 74.605000 54.070000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 75.010000 54.070000 75.330000 ;
      LAYER met4 ;
        RECT 53.750000 75.010000 54.070000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 75.415000 54.070000 75.735000 ;
      LAYER met4 ;
        RECT 53.750000 75.415000 54.070000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 75.820000 54.070000 76.140000 ;
      LAYER met4 ;
        RECT 53.750000 75.820000 54.070000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 76.225000 54.070000 76.545000 ;
      LAYER met4 ;
        RECT 53.750000 76.225000 54.070000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 76.630000 54.070000 76.950000 ;
      LAYER met4 ;
        RECT 53.750000 76.630000 54.070000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 77.035000 54.070000 77.355000 ;
      LAYER met4 ;
        RECT 53.750000 77.035000 54.070000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 77.440000 54.070000 77.760000 ;
      LAYER met4 ;
        RECT 53.750000 77.440000 54.070000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 77.845000 54.070000 78.165000 ;
      LAYER met4 ;
        RECT 53.750000 77.845000 54.070000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 78.250000 54.070000 78.570000 ;
      LAYER met4 ;
        RECT 53.750000 78.250000 54.070000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 78.655000 54.070000 78.975000 ;
      LAYER met4 ;
        RECT 53.750000 78.655000 54.070000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 79.060000 54.070000 79.380000 ;
      LAYER met4 ;
        RECT 53.750000 79.060000 54.070000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 79.465000 54.070000 79.785000 ;
      LAYER met4 ;
        RECT 53.750000 79.465000 54.070000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 79.870000 54.070000 80.190000 ;
      LAYER met4 ;
        RECT 53.750000 79.870000 54.070000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 80.275000 54.070000 80.595000 ;
      LAYER met4 ;
        RECT 53.750000 80.275000 54.070000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 80.680000 54.070000 81.000000 ;
      LAYER met4 ;
        RECT 53.750000 80.680000 54.070000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 81.085000 54.070000 81.405000 ;
      LAYER met4 ;
        RECT 53.750000 81.085000 54.070000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 81.490000 54.070000 81.810000 ;
      LAYER met4 ;
        RECT 53.750000 81.490000 54.070000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 81.895000 54.070000 82.215000 ;
      LAYER met4 ;
        RECT 53.750000 81.895000 54.070000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750000 82.300000 54.070000 82.620000 ;
      LAYER met4 ;
        RECT 53.750000 82.300000 54.070000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.825000 82.950000 54.145000 83.270000 ;
      LAYER met4 ;
        RECT 53.825000 82.950000 54.145000 83.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.825000 83.410000 54.145000 83.730000 ;
      LAYER met4 ;
        RECT 53.825000 83.410000 54.145000 83.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.825000 83.870000 54.145000 84.190000 ;
      LAYER met4 ;
        RECT 53.825000 83.870000 54.145000 84.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.825000 84.335000 54.145000 84.655000 ;
      LAYER met4 ;
        RECT 53.825000 84.335000 54.145000 84.655000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.825000 84.800000 54.145000 85.120000 ;
      LAYER met4 ;
        RECT 53.825000 84.800000 54.145000 85.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.825000 85.265000 54.145000 85.585000 ;
      LAYER met4 ;
        RECT 53.825000 85.265000 54.145000 85.585000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.025000 17.800000 54.345000 18.120000 ;
      LAYER met4 ;
        RECT 54.025000 17.800000 54.345000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.025000 18.230000 54.345000 18.550000 ;
      LAYER met4 ;
        RECT 54.025000 18.230000 54.345000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.025000 18.660000 54.345000 18.980000 ;
      LAYER met4 ;
        RECT 54.025000 18.660000 54.345000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.025000 19.090000 54.345000 19.410000 ;
      LAYER met4 ;
        RECT 54.025000 19.090000 54.345000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.025000 19.520000 54.345000 19.840000 ;
      LAYER met4 ;
        RECT 54.025000 19.520000 54.345000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.025000 19.950000 54.345000 20.270000 ;
      LAYER met4 ;
        RECT 54.025000 19.950000 54.345000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.025000 20.380000 54.345000 20.700000 ;
      LAYER met4 ;
        RECT 54.025000 20.380000 54.345000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.025000 20.810000 54.345000 21.130000 ;
      LAYER met4 ;
        RECT 54.025000 20.810000 54.345000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.025000 21.240000 54.345000 21.560000 ;
      LAYER met4 ;
        RECT 54.025000 21.240000 54.345000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.025000 21.670000 54.345000 21.990000 ;
      LAYER met4 ;
        RECT 54.025000 21.670000 54.345000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.025000 22.100000 54.345000 22.420000 ;
      LAYER met4 ;
        RECT 54.025000 22.100000 54.345000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 68.065000 54.470000 68.385000 ;
      LAYER met4 ;
        RECT 54.150000 68.065000 54.470000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 68.475000 54.470000 68.795000 ;
      LAYER met4 ;
        RECT 54.150000 68.475000 54.470000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 68.885000 54.470000 69.205000 ;
      LAYER met4 ;
        RECT 54.150000 68.885000 54.470000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 69.295000 54.470000 69.615000 ;
      LAYER met4 ;
        RECT 54.150000 69.295000 54.470000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 69.705000 54.470000 70.025000 ;
      LAYER met4 ;
        RECT 54.150000 69.705000 54.470000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 70.115000 54.470000 70.435000 ;
      LAYER met4 ;
        RECT 54.150000 70.115000 54.470000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 70.525000 54.470000 70.845000 ;
      LAYER met4 ;
        RECT 54.150000 70.525000 54.470000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 70.935000 54.470000 71.255000 ;
      LAYER met4 ;
        RECT 54.150000 70.935000 54.470000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 71.345000 54.470000 71.665000 ;
      LAYER met4 ;
        RECT 54.150000 71.345000 54.470000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 71.755000 54.470000 72.075000 ;
      LAYER met4 ;
        RECT 54.150000 71.755000 54.470000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 72.165000 54.470000 72.485000 ;
      LAYER met4 ;
        RECT 54.150000 72.165000 54.470000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 72.575000 54.470000 72.895000 ;
      LAYER met4 ;
        RECT 54.150000 72.575000 54.470000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 72.985000 54.470000 73.305000 ;
      LAYER met4 ;
        RECT 54.150000 72.985000 54.470000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 73.390000 54.470000 73.710000 ;
      LAYER met4 ;
        RECT 54.150000 73.390000 54.470000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 73.795000 54.470000 74.115000 ;
      LAYER met4 ;
        RECT 54.150000 73.795000 54.470000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 74.200000 54.470000 74.520000 ;
      LAYER met4 ;
        RECT 54.150000 74.200000 54.470000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 74.605000 54.470000 74.925000 ;
      LAYER met4 ;
        RECT 54.150000 74.605000 54.470000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 75.010000 54.470000 75.330000 ;
      LAYER met4 ;
        RECT 54.150000 75.010000 54.470000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 75.415000 54.470000 75.735000 ;
      LAYER met4 ;
        RECT 54.150000 75.415000 54.470000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 75.820000 54.470000 76.140000 ;
      LAYER met4 ;
        RECT 54.150000 75.820000 54.470000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 76.225000 54.470000 76.545000 ;
      LAYER met4 ;
        RECT 54.150000 76.225000 54.470000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 76.630000 54.470000 76.950000 ;
      LAYER met4 ;
        RECT 54.150000 76.630000 54.470000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 77.035000 54.470000 77.355000 ;
      LAYER met4 ;
        RECT 54.150000 77.035000 54.470000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 77.440000 54.470000 77.760000 ;
      LAYER met4 ;
        RECT 54.150000 77.440000 54.470000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 77.845000 54.470000 78.165000 ;
      LAYER met4 ;
        RECT 54.150000 77.845000 54.470000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 78.250000 54.470000 78.570000 ;
      LAYER met4 ;
        RECT 54.150000 78.250000 54.470000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 78.655000 54.470000 78.975000 ;
      LAYER met4 ;
        RECT 54.150000 78.655000 54.470000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 79.060000 54.470000 79.380000 ;
      LAYER met4 ;
        RECT 54.150000 79.060000 54.470000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 79.465000 54.470000 79.785000 ;
      LAYER met4 ;
        RECT 54.150000 79.465000 54.470000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 79.870000 54.470000 80.190000 ;
      LAYER met4 ;
        RECT 54.150000 79.870000 54.470000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 80.275000 54.470000 80.595000 ;
      LAYER met4 ;
        RECT 54.150000 80.275000 54.470000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 80.680000 54.470000 81.000000 ;
      LAYER met4 ;
        RECT 54.150000 80.680000 54.470000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 81.085000 54.470000 81.405000 ;
      LAYER met4 ;
        RECT 54.150000 81.085000 54.470000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 81.490000 54.470000 81.810000 ;
      LAYER met4 ;
        RECT 54.150000 81.490000 54.470000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 81.895000 54.470000 82.215000 ;
      LAYER met4 ;
        RECT 54.150000 81.895000 54.470000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.150000 82.300000 54.470000 82.620000 ;
      LAYER met4 ;
        RECT 54.150000 82.300000 54.470000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.305000 82.950000 54.625000 83.270000 ;
      LAYER met4 ;
        RECT 54.305000 82.950000 54.625000 83.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.305000 83.410000 54.625000 83.730000 ;
      LAYER met4 ;
        RECT 54.305000 83.410000 54.625000 83.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.305000 83.870000 54.625000 84.190000 ;
      LAYER met4 ;
        RECT 54.305000 83.870000 54.625000 84.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.305000 84.335000 54.625000 84.655000 ;
      LAYER met4 ;
        RECT 54.305000 84.335000 54.625000 84.655000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.305000 84.800000 54.625000 85.120000 ;
      LAYER met4 ;
        RECT 54.305000 84.800000 54.625000 85.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.305000 85.265000 54.625000 85.585000 ;
      LAYER met4 ;
        RECT 54.305000 85.265000 54.625000 85.585000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.430000 17.800000 54.750000 18.120000 ;
      LAYER met4 ;
        RECT 54.430000 17.800000 54.750000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.430000 18.230000 54.750000 18.550000 ;
      LAYER met4 ;
        RECT 54.430000 18.230000 54.750000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.430000 18.660000 54.750000 18.980000 ;
      LAYER met4 ;
        RECT 54.430000 18.660000 54.750000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.430000 19.090000 54.750000 19.410000 ;
      LAYER met4 ;
        RECT 54.430000 19.090000 54.750000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.430000 19.520000 54.750000 19.840000 ;
      LAYER met4 ;
        RECT 54.430000 19.520000 54.750000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.430000 19.950000 54.750000 20.270000 ;
      LAYER met4 ;
        RECT 54.430000 19.950000 54.750000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.430000 20.380000 54.750000 20.700000 ;
      LAYER met4 ;
        RECT 54.430000 20.380000 54.750000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.430000 20.810000 54.750000 21.130000 ;
      LAYER met4 ;
        RECT 54.430000 20.810000 54.750000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.430000 21.240000 54.750000 21.560000 ;
      LAYER met4 ;
        RECT 54.430000 21.240000 54.750000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.430000 21.670000 54.750000 21.990000 ;
      LAYER met4 ;
        RECT 54.430000 21.670000 54.750000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.430000 22.100000 54.750000 22.420000 ;
      LAYER met4 ;
        RECT 54.430000 22.100000 54.750000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 68.065000 54.870000 68.385000 ;
      LAYER met4 ;
        RECT 54.550000 68.065000 54.870000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 68.475000 54.870000 68.795000 ;
      LAYER met4 ;
        RECT 54.550000 68.475000 54.870000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 68.885000 54.870000 69.205000 ;
      LAYER met4 ;
        RECT 54.550000 68.885000 54.870000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 69.295000 54.870000 69.615000 ;
      LAYER met4 ;
        RECT 54.550000 69.295000 54.870000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 69.705000 54.870000 70.025000 ;
      LAYER met4 ;
        RECT 54.550000 69.705000 54.870000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 70.115000 54.870000 70.435000 ;
      LAYER met4 ;
        RECT 54.550000 70.115000 54.870000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 70.525000 54.870000 70.845000 ;
      LAYER met4 ;
        RECT 54.550000 70.525000 54.870000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 70.935000 54.870000 71.255000 ;
      LAYER met4 ;
        RECT 54.550000 70.935000 54.870000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 71.345000 54.870000 71.665000 ;
      LAYER met4 ;
        RECT 54.550000 71.345000 54.870000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 71.755000 54.870000 72.075000 ;
      LAYER met4 ;
        RECT 54.550000 71.755000 54.870000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 72.165000 54.870000 72.485000 ;
      LAYER met4 ;
        RECT 54.550000 72.165000 54.870000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 72.575000 54.870000 72.895000 ;
      LAYER met4 ;
        RECT 54.550000 72.575000 54.870000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 72.985000 54.870000 73.305000 ;
      LAYER met4 ;
        RECT 54.550000 72.985000 54.870000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 73.390000 54.870000 73.710000 ;
      LAYER met4 ;
        RECT 54.550000 73.390000 54.870000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 73.795000 54.870000 74.115000 ;
      LAYER met4 ;
        RECT 54.550000 73.795000 54.870000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 74.200000 54.870000 74.520000 ;
      LAYER met4 ;
        RECT 54.550000 74.200000 54.870000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 74.605000 54.870000 74.925000 ;
      LAYER met4 ;
        RECT 54.550000 74.605000 54.870000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 75.010000 54.870000 75.330000 ;
      LAYER met4 ;
        RECT 54.550000 75.010000 54.870000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 75.415000 54.870000 75.735000 ;
      LAYER met4 ;
        RECT 54.550000 75.415000 54.870000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 75.820000 54.870000 76.140000 ;
      LAYER met4 ;
        RECT 54.550000 75.820000 54.870000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 76.225000 54.870000 76.545000 ;
      LAYER met4 ;
        RECT 54.550000 76.225000 54.870000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 76.630000 54.870000 76.950000 ;
      LAYER met4 ;
        RECT 54.550000 76.630000 54.870000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 77.035000 54.870000 77.355000 ;
      LAYER met4 ;
        RECT 54.550000 77.035000 54.870000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 77.440000 54.870000 77.760000 ;
      LAYER met4 ;
        RECT 54.550000 77.440000 54.870000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 77.845000 54.870000 78.165000 ;
      LAYER met4 ;
        RECT 54.550000 77.845000 54.870000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 78.250000 54.870000 78.570000 ;
      LAYER met4 ;
        RECT 54.550000 78.250000 54.870000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 78.655000 54.870000 78.975000 ;
      LAYER met4 ;
        RECT 54.550000 78.655000 54.870000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 79.060000 54.870000 79.380000 ;
      LAYER met4 ;
        RECT 54.550000 79.060000 54.870000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 79.465000 54.870000 79.785000 ;
      LAYER met4 ;
        RECT 54.550000 79.465000 54.870000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 79.870000 54.870000 80.190000 ;
      LAYER met4 ;
        RECT 54.550000 79.870000 54.870000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 80.275000 54.870000 80.595000 ;
      LAYER met4 ;
        RECT 54.550000 80.275000 54.870000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 80.680000 54.870000 81.000000 ;
      LAYER met4 ;
        RECT 54.550000 80.680000 54.870000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 81.085000 54.870000 81.405000 ;
      LAYER met4 ;
        RECT 54.550000 81.085000 54.870000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 81.490000 54.870000 81.810000 ;
      LAYER met4 ;
        RECT 54.550000 81.490000 54.870000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 81.895000 54.870000 82.215000 ;
      LAYER met4 ;
        RECT 54.550000 81.895000 54.870000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.550000 82.300000 54.870000 82.620000 ;
      LAYER met4 ;
        RECT 54.550000 82.300000 54.870000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.785000 82.950000 55.105000 83.270000 ;
      LAYER met4 ;
        RECT 54.785000 82.950000 55.105000 83.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.785000 83.410000 55.105000 83.730000 ;
      LAYER met4 ;
        RECT 54.785000 83.410000 55.105000 83.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.785000 83.870000 55.105000 84.190000 ;
      LAYER met4 ;
        RECT 54.785000 83.870000 55.105000 84.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.785000 84.335000 55.105000 84.655000 ;
      LAYER met4 ;
        RECT 54.785000 84.335000 55.105000 84.655000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.785000 84.800000 55.105000 85.120000 ;
      LAYER met4 ;
        RECT 54.785000 84.800000 55.105000 85.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.785000 85.265000 55.105000 85.585000 ;
      LAYER met4 ;
        RECT 54.785000 85.265000 55.105000 85.585000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.835000 17.800000 55.155000 18.120000 ;
      LAYER met4 ;
        RECT 54.835000 17.800000 55.155000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.835000 18.230000 55.155000 18.550000 ;
      LAYER met4 ;
        RECT 54.835000 18.230000 55.155000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.835000 18.660000 55.155000 18.980000 ;
      LAYER met4 ;
        RECT 54.835000 18.660000 55.155000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.835000 19.090000 55.155000 19.410000 ;
      LAYER met4 ;
        RECT 54.835000 19.090000 55.155000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.835000 19.520000 55.155000 19.840000 ;
      LAYER met4 ;
        RECT 54.835000 19.520000 55.155000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.835000 19.950000 55.155000 20.270000 ;
      LAYER met4 ;
        RECT 54.835000 19.950000 55.155000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.835000 20.380000 55.155000 20.700000 ;
      LAYER met4 ;
        RECT 54.835000 20.380000 55.155000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.835000 20.810000 55.155000 21.130000 ;
      LAYER met4 ;
        RECT 54.835000 20.810000 55.155000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.835000 21.240000 55.155000 21.560000 ;
      LAYER met4 ;
        RECT 54.835000 21.240000 55.155000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.835000 21.670000 55.155000 21.990000 ;
      LAYER met4 ;
        RECT 54.835000 21.670000 55.155000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.835000 22.100000 55.155000 22.420000 ;
      LAYER met4 ;
        RECT 54.835000 22.100000 55.155000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 68.065000 55.270000 68.385000 ;
      LAYER met4 ;
        RECT 54.950000 68.065000 55.270000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 68.475000 55.270000 68.795000 ;
      LAYER met4 ;
        RECT 54.950000 68.475000 55.270000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 68.885000 55.270000 69.205000 ;
      LAYER met4 ;
        RECT 54.950000 68.885000 55.270000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 69.295000 55.270000 69.615000 ;
      LAYER met4 ;
        RECT 54.950000 69.295000 55.270000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 69.705000 55.270000 70.025000 ;
      LAYER met4 ;
        RECT 54.950000 69.705000 55.270000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 70.115000 55.270000 70.435000 ;
      LAYER met4 ;
        RECT 54.950000 70.115000 55.270000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 70.525000 55.270000 70.845000 ;
      LAYER met4 ;
        RECT 54.950000 70.525000 55.270000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 70.935000 55.270000 71.255000 ;
      LAYER met4 ;
        RECT 54.950000 70.935000 55.270000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 71.345000 55.270000 71.665000 ;
      LAYER met4 ;
        RECT 54.950000 71.345000 55.270000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 71.755000 55.270000 72.075000 ;
      LAYER met4 ;
        RECT 54.950000 71.755000 55.270000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 72.165000 55.270000 72.485000 ;
      LAYER met4 ;
        RECT 54.950000 72.165000 55.270000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 72.575000 55.270000 72.895000 ;
      LAYER met4 ;
        RECT 54.950000 72.575000 55.270000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 72.985000 55.270000 73.305000 ;
      LAYER met4 ;
        RECT 54.950000 72.985000 55.270000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 73.390000 55.270000 73.710000 ;
      LAYER met4 ;
        RECT 54.950000 73.390000 55.270000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 73.795000 55.270000 74.115000 ;
      LAYER met4 ;
        RECT 54.950000 73.795000 55.270000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 74.200000 55.270000 74.520000 ;
      LAYER met4 ;
        RECT 54.950000 74.200000 55.270000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 74.605000 55.270000 74.925000 ;
      LAYER met4 ;
        RECT 54.950000 74.605000 55.270000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 75.010000 55.270000 75.330000 ;
      LAYER met4 ;
        RECT 54.950000 75.010000 55.270000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 75.415000 55.270000 75.735000 ;
      LAYER met4 ;
        RECT 54.950000 75.415000 55.270000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 75.820000 55.270000 76.140000 ;
      LAYER met4 ;
        RECT 54.950000 75.820000 55.270000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 76.225000 55.270000 76.545000 ;
      LAYER met4 ;
        RECT 54.950000 76.225000 55.270000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 76.630000 55.270000 76.950000 ;
      LAYER met4 ;
        RECT 54.950000 76.630000 55.270000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 77.035000 55.270000 77.355000 ;
      LAYER met4 ;
        RECT 54.950000 77.035000 55.270000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 77.440000 55.270000 77.760000 ;
      LAYER met4 ;
        RECT 54.950000 77.440000 55.270000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 77.845000 55.270000 78.165000 ;
      LAYER met4 ;
        RECT 54.950000 77.845000 55.270000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 78.250000 55.270000 78.570000 ;
      LAYER met4 ;
        RECT 54.950000 78.250000 55.270000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 78.655000 55.270000 78.975000 ;
      LAYER met4 ;
        RECT 54.950000 78.655000 55.270000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 79.060000 55.270000 79.380000 ;
      LAYER met4 ;
        RECT 54.950000 79.060000 55.270000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 79.465000 55.270000 79.785000 ;
      LAYER met4 ;
        RECT 54.950000 79.465000 55.270000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 79.870000 55.270000 80.190000 ;
      LAYER met4 ;
        RECT 54.950000 79.870000 55.270000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 80.275000 55.270000 80.595000 ;
      LAYER met4 ;
        RECT 54.950000 80.275000 55.270000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 80.680000 55.270000 81.000000 ;
      LAYER met4 ;
        RECT 54.950000 80.680000 55.270000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 81.085000 55.270000 81.405000 ;
      LAYER met4 ;
        RECT 54.950000 81.085000 55.270000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 81.490000 55.270000 81.810000 ;
      LAYER met4 ;
        RECT 54.950000 81.490000 55.270000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 81.895000 55.270000 82.215000 ;
      LAYER met4 ;
        RECT 54.950000 81.895000 55.270000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.950000 82.300000 55.270000 82.620000 ;
      LAYER met4 ;
        RECT 54.950000 82.300000 55.270000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.195000 85.815000 55.515000 86.135000 ;
      LAYER met4 ;
        RECT 55.195000 85.815000 55.515000 86.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.195000 86.250000 55.515000 86.570000 ;
      LAYER met4 ;
        RECT 55.195000 86.250000 55.515000 86.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.195000 86.690000 55.515000 87.010000 ;
      LAYER met4 ;
        RECT 55.195000 86.690000 55.515000 87.010000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.240000 17.800000 55.560000 18.120000 ;
      LAYER met4 ;
        RECT 55.240000 17.800000 55.560000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.240000 18.230000 55.560000 18.550000 ;
      LAYER met4 ;
        RECT 55.240000 18.230000 55.560000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.240000 18.660000 55.560000 18.980000 ;
      LAYER met4 ;
        RECT 55.240000 18.660000 55.560000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.240000 19.090000 55.560000 19.410000 ;
      LAYER met4 ;
        RECT 55.240000 19.090000 55.560000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.240000 19.520000 55.560000 19.840000 ;
      LAYER met4 ;
        RECT 55.240000 19.520000 55.560000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.240000 19.950000 55.560000 20.270000 ;
      LAYER met4 ;
        RECT 55.240000 19.950000 55.560000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.240000 20.380000 55.560000 20.700000 ;
      LAYER met4 ;
        RECT 55.240000 20.380000 55.560000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.240000 20.810000 55.560000 21.130000 ;
      LAYER met4 ;
        RECT 55.240000 20.810000 55.560000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.240000 21.240000 55.560000 21.560000 ;
      LAYER met4 ;
        RECT 55.240000 21.240000 55.560000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.240000 21.670000 55.560000 21.990000 ;
      LAYER met4 ;
        RECT 55.240000 21.670000 55.560000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.240000 22.100000 55.560000 22.420000 ;
      LAYER met4 ;
        RECT 55.240000 22.100000 55.560000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.265000 82.950000 55.585000 83.270000 ;
      LAYER met4 ;
        RECT 55.265000 82.950000 55.585000 83.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.265000 83.410000 55.585000 83.730000 ;
      LAYER met4 ;
        RECT 55.265000 83.410000 55.585000 83.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.265000 83.870000 55.585000 84.190000 ;
      LAYER met4 ;
        RECT 55.265000 83.870000 55.585000 84.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.265000 84.335000 55.585000 84.655000 ;
      LAYER met4 ;
        RECT 55.265000 84.335000 55.585000 84.655000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.265000 84.800000 55.585000 85.120000 ;
      LAYER met4 ;
        RECT 55.265000 84.800000 55.585000 85.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.265000 85.265000 55.585000 85.585000 ;
      LAYER met4 ;
        RECT 55.265000 85.265000 55.585000 85.585000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 68.065000 55.670000 68.385000 ;
      LAYER met4 ;
        RECT 55.350000 68.065000 55.670000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 68.475000 55.670000 68.795000 ;
      LAYER met4 ;
        RECT 55.350000 68.475000 55.670000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 68.885000 55.670000 69.205000 ;
      LAYER met4 ;
        RECT 55.350000 68.885000 55.670000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 69.295000 55.670000 69.615000 ;
      LAYER met4 ;
        RECT 55.350000 69.295000 55.670000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 69.705000 55.670000 70.025000 ;
      LAYER met4 ;
        RECT 55.350000 69.705000 55.670000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 70.115000 55.670000 70.435000 ;
      LAYER met4 ;
        RECT 55.350000 70.115000 55.670000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 70.525000 55.670000 70.845000 ;
      LAYER met4 ;
        RECT 55.350000 70.525000 55.670000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 70.935000 55.670000 71.255000 ;
      LAYER met4 ;
        RECT 55.350000 70.935000 55.670000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 71.345000 55.670000 71.665000 ;
      LAYER met4 ;
        RECT 55.350000 71.345000 55.670000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 71.755000 55.670000 72.075000 ;
      LAYER met4 ;
        RECT 55.350000 71.755000 55.670000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 72.165000 55.670000 72.485000 ;
      LAYER met4 ;
        RECT 55.350000 72.165000 55.670000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 72.575000 55.670000 72.895000 ;
      LAYER met4 ;
        RECT 55.350000 72.575000 55.670000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 72.985000 55.670000 73.305000 ;
      LAYER met4 ;
        RECT 55.350000 72.985000 55.670000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 73.390000 55.670000 73.710000 ;
      LAYER met4 ;
        RECT 55.350000 73.390000 55.670000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 73.795000 55.670000 74.115000 ;
      LAYER met4 ;
        RECT 55.350000 73.795000 55.670000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 74.200000 55.670000 74.520000 ;
      LAYER met4 ;
        RECT 55.350000 74.200000 55.670000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 74.605000 55.670000 74.925000 ;
      LAYER met4 ;
        RECT 55.350000 74.605000 55.670000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 75.010000 55.670000 75.330000 ;
      LAYER met4 ;
        RECT 55.350000 75.010000 55.670000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 75.415000 55.670000 75.735000 ;
      LAYER met4 ;
        RECT 55.350000 75.415000 55.670000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 75.820000 55.670000 76.140000 ;
      LAYER met4 ;
        RECT 55.350000 75.820000 55.670000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 76.225000 55.670000 76.545000 ;
      LAYER met4 ;
        RECT 55.350000 76.225000 55.670000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 76.630000 55.670000 76.950000 ;
      LAYER met4 ;
        RECT 55.350000 76.630000 55.670000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 77.035000 55.670000 77.355000 ;
      LAYER met4 ;
        RECT 55.350000 77.035000 55.670000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 77.440000 55.670000 77.760000 ;
      LAYER met4 ;
        RECT 55.350000 77.440000 55.670000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 77.845000 55.670000 78.165000 ;
      LAYER met4 ;
        RECT 55.350000 77.845000 55.670000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 78.250000 55.670000 78.570000 ;
      LAYER met4 ;
        RECT 55.350000 78.250000 55.670000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 78.655000 55.670000 78.975000 ;
      LAYER met4 ;
        RECT 55.350000 78.655000 55.670000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 79.060000 55.670000 79.380000 ;
      LAYER met4 ;
        RECT 55.350000 79.060000 55.670000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 79.465000 55.670000 79.785000 ;
      LAYER met4 ;
        RECT 55.350000 79.465000 55.670000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 79.870000 55.670000 80.190000 ;
      LAYER met4 ;
        RECT 55.350000 79.870000 55.670000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 80.275000 55.670000 80.595000 ;
      LAYER met4 ;
        RECT 55.350000 80.275000 55.670000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 80.680000 55.670000 81.000000 ;
      LAYER met4 ;
        RECT 55.350000 80.680000 55.670000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 81.085000 55.670000 81.405000 ;
      LAYER met4 ;
        RECT 55.350000 81.085000 55.670000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 81.490000 55.670000 81.810000 ;
      LAYER met4 ;
        RECT 55.350000 81.490000 55.670000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 81.895000 55.670000 82.215000 ;
      LAYER met4 ;
        RECT 55.350000 81.895000 55.670000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.350000 82.300000 55.670000 82.620000 ;
      LAYER met4 ;
        RECT 55.350000 82.300000 55.670000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.645000 17.800000 55.965000 18.120000 ;
      LAYER met4 ;
        RECT 55.645000 17.800000 55.965000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.645000 18.230000 55.965000 18.550000 ;
      LAYER met4 ;
        RECT 55.645000 18.230000 55.965000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.645000 18.660000 55.965000 18.980000 ;
      LAYER met4 ;
        RECT 55.645000 18.660000 55.965000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.645000 19.090000 55.965000 19.410000 ;
      LAYER met4 ;
        RECT 55.645000 19.090000 55.965000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.645000 19.520000 55.965000 19.840000 ;
      LAYER met4 ;
        RECT 55.645000 19.520000 55.965000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.645000 19.950000 55.965000 20.270000 ;
      LAYER met4 ;
        RECT 55.645000 19.950000 55.965000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.645000 20.380000 55.965000 20.700000 ;
      LAYER met4 ;
        RECT 55.645000 20.380000 55.965000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.645000 20.810000 55.965000 21.130000 ;
      LAYER met4 ;
        RECT 55.645000 20.810000 55.965000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.645000 21.240000 55.965000 21.560000 ;
      LAYER met4 ;
        RECT 55.645000 21.240000 55.965000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.645000 21.670000 55.965000 21.990000 ;
      LAYER met4 ;
        RECT 55.645000 21.670000 55.965000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.645000 22.100000 55.965000 22.420000 ;
      LAYER met4 ;
        RECT 55.645000 22.100000 55.965000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.745000 82.950000 56.065000 83.270000 ;
      LAYER met4 ;
        RECT 55.745000 82.950000 56.065000 83.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.745000 83.410000 56.065000 83.730000 ;
      LAYER met4 ;
        RECT 55.745000 83.410000 56.065000 83.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.745000 83.870000 56.065000 84.190000 ;
      LAYER met4 ;
        RECT 55.745000 83.870000 56.065000 84.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.745000 84.335000 56.065000 84.655000 ;
      LAYER met4 ;
        RECT 55.745000 84.335000 56.065000 84.655000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.745000 84.800000 56.065000 85.120000 ;
      LAYER met4 ;
        RECT 55.745000 84.800000 56.065000 85.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.745000 85.265000 56.065000 85.585000 ;
      LAYER met4 ;
        RECT 55.745000 85.265000 56.065000 85.585000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 68.065000 56.070000 68.385000 ;
      LAYER met4 ;
        RECT 55.750000 68.065000 56.070000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 68.475000 56.070000 68.795000 ;
      LAYER met4 ;
        RECT 55.750000 68.475000 56.070000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 68.885000 56.070000 69.205000 ;
      LAYER met4 ;
        RECT 55.750000 68.885000 56.070000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 69.295000 56.070000 69.615000 ;
      LAYER met4 ;
        RECT 55.750000 69.295000 56.070000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 69.705000 56.070000 70.025000 ;
      LAYER met4 ;
        RECT 55.750000 69.705000 56.070000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 70.115000 56.070000 70.435000 ;
      LAYER met4 ;
        RECT 55.750000 70.115000 56.070000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 70.525000 56.070000 70.845000 ;
      LAYER met4 ;
        RECT 55.750000 70.525000 56.070000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 70.935000 56.070000 71.255000 ;
      LAYER met4 ;
        RECT 55.750000 70.935000 56.070000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 71.345000 56.070000 71.665000 ;
      LAYER met4 ;
        RECT 55.750000 71.345000 56.070000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 71.755000 56.070000 72.075000 ;
      LAYER met4 ;
        RECT 55.750000 71.755000 56.070000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 72.165000 56.070000 72.485000 ;
      LAYER met4 ;
        RECT 55.750000 72.165000 56.070000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 72.575000 56.070000 72.895000 ;
      LAYER met4 ;
        RECT 55.750000 72.575000 56.070000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 72.985000 56.070000 73.305000 ;
      LAYER met4 ;
        RECT 55.750000 72.985000 56.070000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 73.390000 56.070000 73.710000 ;
      LAYER met4 ;
        RECT 55.750000 73.390000 56.070000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 73.795000 56.070000 74.115000 ;
      LAYER met4 ;
        RECT 55.750000 73.795000 56.070000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 74.200000 56.070000 74.520000 ;
      LAYER met4 ;
        RECT 55.750000 74.200000 56.070000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 74.605000 56.070000 74.925000 ;
      LAYER met4 ;
        RECT 55.750000 74.605000 56.070000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 75.010000 56.070000 75.330000 ;
      LAYER met4 ;
        RECT 55.750000 75.010000 56.070000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 75.415000 56.070000 75.735000 ;
      LAYER met4 ;
        RECT 55.750000 75.415000 56.070000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 75.820000 56.070000 76.140000 ;
      LAYER met4 ;
        RECT 55.750000 75.820000 56.070000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 76.225000 56.070000 76.545000 ;
      LAYER met4 ;
        RECT 55.750000 76.225000 56.070000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 76.630000 56.070000 76.950000 ;
      LAYER met4 ;
        RECT 55.750000 76.630000 56.070000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 77.035000 56.070000 77.355000 ;
      LAYER met4 ;
        RECT 55.750000 77.035000 56.070000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 77.440000 56.070000 77.760000 ;
      LAYER met4 ;
        RECT 55.750000 77.440000 56.070000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 77.845000 56.070000 78.165000 ;
      LAYER met4 ;
        RECT 55.750000 77.845000 56.070000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 78.250000 56.070000 78.570000 ;
      LAYER met4 ;
        RECT 55.750000 78.250000 56.070000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 78.655000 56.070000 78.975000 ;
      LAYER met4 ;
        RECT 55.750000 78.655000 56.070000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 79.060000 56.070000 79.380000 ;
      LAYER met4 ;
        RECT 55.750000 79.060000 56.070000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 79.465000 56.070000 79.785000 ;
      LAYER met4 ;
        RECT 55.750000 79.465000 56.070000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 79.870000 56.070000 80.190000 ;
      LAYER met4 ;
        RECT 55.750000 79.870000 56.070000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 80.275000 56.070000 80.595000 ;
      LAYER met4 ;
        RECT 55.750000 80.275000 56.070000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 80.680000 56.070000 81.000000 ;
      LAYER met4 ;
        RECT 55.750000 80.680000 56.070000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 81.085000 56.070000 81.405000 ;
      LAYER met4 ;
        RECT 55.750000 81.085000 56.070000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 81.490000 56.070000 81.810000 ;
      LAYER met4 ;
        RECT 55.750000 81.490000 56.070000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 81.895000 56.070000 82.215000 ;
      LAYER met4 ;
        RECT 55.750000 81.895000 56.070000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.750000 82.300000 56.070000 82.620000 ;
      LAYER met4 ;
        RECT 55.750000 82.300000 56.070000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.935000 85.815000 56.255000 86.135000 ;
      LAYER met4 ;
        RECT 55.935000 85.815000 56.255000 86.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.935000 86.250000 56.255000 86.570000 ;
      LAYER met4 ;
        RECT 55.935000 86.250000 56.255000 86.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.935000 86.690000 56.255000 87.010000 ;
      LAYER met4 ;
        RECT 55.935000 86.690000 56.255000 87.010000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.050000 17.800000 56.370000 18.120000 ;
      LAYER met4 ;
        RECT 56.050000 17.800000 56.370000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.050000 18.230000 56.370000 18.550000 ;
      LAYER met4 ;
        RECT 56.050000 18.230000 56.370000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.050000 18.660000 56.370000 18.980000 ;
      LAYER met4 ;
        RECT 56.050000 18.660000 56.370000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.050000 19.090000 56.370000 19.410000 ;
      LAYER met4 ;
        RECT 56.050000 19.090000 56.370000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.050000 19.520000 56.370000 19.840000 ;
      LAYER met4 ;
        RECT 56.050000 19.520000 56.370000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.050000 19.950000 56.370000 20.270000 ;
      LAYER met4 ;
        RECT 56.050000 19.950000 56.370000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.050000 20.380000 56.370000 20.700000 ;
      LAYER met4 ;
        RECT 56.050000 20.380000 56.370000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.050000 20.810000 56.370000 21.130000 ;
      LAYER met4 ;
        RECT 56.050000 20.810000 56.370000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.050000 21.240000 56.370000 21.560000 ;
      LAYER met4 ;
        RECT 56.050000 21.240000 56.370000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.050000 21.670000 56.370000 21.990000 ;
      LAYER met4 ;
        RECT 56.050000 21.670000 56.370000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.050000 22.100000 56.370000 22.420000 ;
      LAYER met4 ;
        RECT 56.050000 22.100000 56.370000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 68.065000 56.470000 68.385000 ;
      LAYER met4 ;
        RECT 56.150000 68.065000 56.470000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 68.475000 56.470000 68.795000 ;
      LAYER met4 ;
        RECT 56.150000 68.475000 56.470000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 68.885000 56.470000 69.205000 ;
      LAYER met4 ;
        RECT 56.150000 68.885000 56.470000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 69.295000 56.470000 69.615000 ;
      LAYER met4 ;
        RECT 56.150000 69.295000 56.470000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 69.705000 56.470000 70.025000 ;
      LAYER met4 ;
        RECT 56.150000 69.705000 56.470000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 70.115000 56.470000 70.435000 ;
      LAYER met4 ;
        RECT 56.150000 70.115000 56.470000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 70.525000 56.470000 70.845000 ;
      LAYER met4 ;
        RECT 56.150000 70.525000 56.470000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 70.935000 56.470000 71.255000 ;
      LAYER met4 ;
        RECT 56.150000 70.935000 56.470000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 71.345000 56.470000 71.665000 ;
      LAYER met4 ;
        RECT 56.150000 71.345000 56.470000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 71.755000 56.470000 72.075000 ;
      LAYER met4 ;
        RECT 56.150000 71.755000 56.470000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 72.165000 56.470000 72.485000 ;
      LAYER met4 ;
        RECT 56.150000 72.165000 56.470000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 72.575000 56.470000 72.895000 ;
      LAYER met4 ;
        RECT 56.150000 72.575000 56.470000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 72.985000 56.470000 73.305000 ;
      LAYER met4 ;
        RECT 56.150000 72.985000 56.470000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 73.390000 56.470000 73.710000 ;
      LAYER met4 ;
        RECT 56.150000 73.390000 56.470000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 73.795000 56.470000 74.115000 ;
      LAYER met4 ;
        RECT 56.150000 73.795000 56.470000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 74.200000 56.470000 74.520000 ;
      LAYER met4 ;
        RECT 56.150000 74.200000 56.470000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 74.605000 56.470000 74.925000 ;
      LAYER met4 ;
        RECT 56.150000 74.605000 56.470000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 75.010000 56.470000 75.330000 ;
      LAYER met4 ;
        RECT 56.150000 75.010000 56.470000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 75.415000 56.470000 75.735000 ;
      LAYER met4 ;
        RECT 56.150000 75.415000 56.470000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 75.820000 56.470000 76.140000 ;
      LAYER met4 ;
        RECT 56.150000 75.820000 56.470000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 76.225000 56.470000 76.545000 ;
      LAYER met4 ;
        RECT 56.150000 76.225000 56.470000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 76.630000 56.470000 76.950000 ;
      LAYER met4 ;
        RECT 56.150000 76.630000 56.470000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 77.035000 56.470000 77.355000 ;
      LAYER met4 ;
        RECT 56.150000 77.035000 56.470000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 77.440000 56.470000 77.760000 ;
      LAYER met4 ;
        RECT 56.150000 77.440000 56.470000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 77.845000 56.470000 78.165000 ;
      LAYER met4 ;
        RECT 56.150000 77.845000 56.470000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 78.250000 56.470000 78.570000 ;
      LAYER met4 ;
        RECT 56.150000 78.250000 56.470000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 78.655000 56.470000 78.975000 ;
      LAYER met4 ;
        RECT 56.150000 78.655000 56.470000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 79.060000 56.470000 79.380000 ;
      LAYER met4 ;
        RECT 56.150000 79.060000 56.470000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 79.465000 56.470000 79.785000 ;
      LAYER met4 ;
        RECT 56.150000 79.465000 56.470000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 79.870000 56.470000 80.190000 ;
      LAYER met4 ;
        RECT 56.150000 79.870000 56.470000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 80.275000 56.470000 80.595000 ;
      LAYER met4 ;
        RECT 56.150000 80.275000 56.470000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 80.680000 56.470000 81.000000 ;
      LAYER met4 ;
        RECT 56.150000 80.680000 56.470000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 81.085000 56.470000 81.405000 ;
      LAYER met4 ;
        RECT 56.150000 81.085000 56.470000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 81.490000 56.470000 81.810000 ;
      LAYER met4 ;
        RECT 56.150000 81.490000 56.470000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 81.895000 56.470000 82.215000 ;
      LAYER met4 ;
        RECT 56.150000 81.895000 56.470000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150000 82.300000 56.470000 82.620000 ;
      LAYER met4 ;
        RECT 56.150000 82.300000 56.470000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430000 82.995000 56.750000 83.315000 ;
      LAYER met4 ;
        RECT 56.430000 82.995000 56.750000 83.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430000 83.395000 56.750000 83.715000 ;
      LAYER met4 ;
        RECT 56.430000 83.395000 56.750000 83.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430000 83.795000 56.750000 84.115000 ;
      LAYER met4 ;
        RECT 56.430000 83.795000 56.750000 84.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430000 84.195000 56.750000 84.515000 ;
      LAYER met4 ;
        RECT 56.430000 84.195000 56.750000 84.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430000 84.595000 56.750000 84.915000 ;
      LAYER met4 ;
        RECT 56.430000 84.595000 56.750000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430000 84.995000 56.750000 85.315000 ;
      LAYER met4 ;
        RECT 56.430000 84.995000 56.750000 85.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430000 85.395000 56.750000 85.715000 ;
      LAYER met4 ;
        RECT 56.430000 85.395000 56.750000 85.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430000 85.795000 56.750000 86.115000 ;
      LAYER met4 ;
        RECT 56.430000 85.795000 56.750000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430000 86.195000 56.750000 86.515000 ;
      LAYER met4 ;
        RECT 56.430000 86.195000 56.750000 86.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430000 86.600000 56.750000 86.920000 ;
      LAYER met4 ;
        RECT 56.430000 86.600000 56.750000 86.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430000 87.005000 56.750000 87.325000 ;
      LAYER met4 ;
        RECT 56.430000 87.005000 56.750000 87.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430000 87.410000 56.750000 87.730000 ;
      LAYER met4 ;
        RECT 56.430000 87.410000 56.750000 87.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430000 87.815000 56.750000 88.135000 ;
      LAYER met4 ;
        RECT 56.430000 87.815000 56.750000 88.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 17.800000 56.775000 18.120000 ;
      LAYER met4 ;
        RECT 56.455000 17.800000 56.775000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 18.230000 56.775000 18.550000 ;
      LAYER met4 ;
        RECT 56.455000 18.230000 56.775000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 18.660000 56.775000 18.980000 ;
      LAYER met4 ;
        RECT 56.455000 18.660000 56.775000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 19.090000 56.775000 19.410000 ;
      LAYER met4 ;
        RECT 56.455000 19.090000 56.775000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 19.520000 56.775000 19.840000 ;
      LAYER met4 ;
        RECT 56.455000 19.520000 56.775000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 19.950000 56.775000 20.270000 ;
      LAYER met4 ;
        RECT 56.455000 19.950000 56.775000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 20.380000 56.775000 20.700000 ;
      LAYER met4 ;
        RECT 56.455000 20.380000 56.775000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 20.810000 56.775000 21.130000 ;
      LAYER met4 ;
        RECT 56.455000 20.810000 56.775000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 21.240000 56.775000 21.560000 ;
      LAYER met4 ;
        RECT 56.455000 21.240000 56.775000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 21.670000 56.775000 21.990000 ;
      LAYER met4 ;
        RECT 56.455000 21.670000 56.775000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 22.100000 56.775000 22.420000 ;
      LAYER met4 ;
        RECT 56.455000 22.100000 56.775000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 68.065000 56.870000 68.385000 ;
      LAYER met4 ;
        RECT 56.550000 68.065000 56.870000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 68.475000 56.870000 68.795000 ;
      LAYER met4 ;
        RECT 56.550000 68.475000 56.870000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 68.885000 56.870000 69.205000 ;
      LAYER met4 ;
        RECT 56.550000 68.885000 56.870000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 69.295000 56.870000 69.615000 ;
      LAYER met4 ;
        RECT 56.550000 69.295000 56.870000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 69.705000 56.870000 70.025000 ;
      LAYER met4 ;
        RECT 56.550000 69.705000 56.870000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 70.115000 56.870000 70.435000 ;
      LAYER met4 ;
        RECT 56.550000 70.115000 56.870000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 70.525000 56.870000 70.845000 ;
      LAYER met4 ;
        RECT 56.550000 70.525000 56.870000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 70.935000 56.870000 71.255000 ;
      LAYER met4 ;
        RECT 56.550000 70.935000 56.870000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 71.345000 56.870000 71.665000 ;
      LAYER met4 ;
        RECT 56.550000 71.345000 56.870000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 71.755000 56.870000 72.075000 ;
      LAYER met4 ;
        RECT 56.550000 71.755000 56.870000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 72.165000 56.870000 72.485000 ;
      LAYER met4 ;
        RECT 56.550000 72.165000 56.870000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 72.575000 56.870000 72.895000 ;
      LAYER met4 ;
        RECT 56.550000 72.575000 56.870000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 72.985000 56.870000 73.305000 ;
      LAYER met4 ;
        RECT 56.550000 72.985000 56.870000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 73.390000 56.870000 73.710000 ;
      LAYER met4 ;
        RECT 56.550000 73.390000 56.870000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 73.795000 56.870000 74.115000 ;
      LAYER met4 ;
        RECT 56.550000 73.795000 56.870000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 74.200000 56.870000 74.520000 ;
      LAYER met4 ;
        RECT 56.550000 74.200000 56.870000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 74.605000 56.870000 74.925000 ;
      LAYER met4 ;
        RECT 56.550000 74.605000 56.870000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 75.010000 56.870000 75.330000 ;
      LAYER met4 ;
        RECT 56.550000 75.010000 56.870000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 75.415000 56.870000 75.735000 ;
      LAYER met4 ;
        RECT 56.550000 75.415000 56.870000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 75.820000 56.870000 76.140000 ;
      LAYER met4 ;
        RECT 56.550000 75.820000 56.870000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 76.225000 56.870000 76.545000 ;
      LAYER met4 ;
        RECT 56.550000 76.225000 56.870000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 76.630000 56.870000 76.950000 ;
      LAYER met4 ;
        RECT 56.550000 76.630000 56.870000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 77.035000 56.870000 77.355000 ;
      LAYER met4 ;
        RECT 56.550000 77.035000 56.870000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 77.440000 56.870000 77.760000 ;
      LAYER met4 ;
        RECT 56.550000 77.440000 56.870000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 77.845000 56.870000 78.165000 ;
      LAYER met4 ;
        RECT 56.550000 77.845000 56.870000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 78.250000 56.870000 78.570000 ;
      LAYER met4 ;
        RECT 56.550000 78.250000 56.870000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 78.655000 56.870000 78.975000 ;
      LAYER met4 ;
        RECT 56.550000 78.655000 56.870000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 79.060000 56.870000 79.380000 ;
      LAYER met4 ;
        RECT 56.550000 79.060000 56.870000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 79.465000 56.870000 79.785000 ;
      LAYER met4 ;
        RECT 56.550000 79.465000 56.870000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 79.870000 56.870000 80.190000 ;
      LAYER met4 ;
        RECT 56.550000 79.870000 56.870000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 80.275000 56.870000 80.595000 ;
      LAYER met4 ;
        RECT 56.550000 80.275000 56.870000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 80.680000 56.870000 81.000000 ;
      LAYER met4 ;
        RECT 56.550000 80.680000 56.870000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 81.085000 56.870000 81.405000 ;
      LAYER met4 ;
        RECT 56.550000 81.085000 56.870000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 81.490000 56.870000 81.810000 ;
      LAYER met4 ;
        RECT 56.550000 81.490000 56.870000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 81.895000 56.870000 82.215000 ;
      LAYER met4 ;
        RECT 56.550000 81.895000 56.870000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.550000 82.300000 56.870000 82.620000 ;
      LAYER met4 ;
        RECT 56.550000 82.300000 56.870000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840000 82.995000 57.160000 83.315000 ;
      LAYER met4 ;
        RECT 56.840000 82.995000 57.160000 83.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840000 83.395000 57.160000 83.715000 ;
      LAYER met4 ;
        RECT 56.840000 83.395000 57.160000 83.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840000 83.795000 57.160000 84.115000 ;
      LAYER met4 ;
        RECT 56.840000 83.795000 57.160000 84.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840000 84.195000 57.160000 84.515000 ;
      LAYER met4 ;
        RECT 56.840000 84.195000 57.160000 84.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840000 84.595000 57.160000 84.915000 ;
      LAYER met4 ;
        RECT 56.840000 84.595000 57.160000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840000 84.995000 57.160000 85.315000 ;
      LAYER met4 ;
        RECT 56.840000 84.995000 57.160000 85.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840000 85.395000 57.160000 85.715000 ;
      LAYER met4 ;
        RECT 56.840000 85.395000 57.160000 85.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840000 85.795000 57.160000 86.115000 ;
      LAYER met4 ;
        RECT 56.840000 85.795000 57.160000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840000 86.195000 57.160000 86.515000 ;
      LAYER met4 ;
        RECT 56.840000 86.195000 57.160000 86.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840000 86.600000 57.160000 86.920000 ;
      LAYER met4 ;
        RECT 56.840000 86.600000 57.160000 86.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840000 87.005000 57.160000 87.325000 ;
      LAYER met4 ;
        RECT 56.840000 87.005000 57.160000 87.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840000 87.410000 57.160000 87.730000 ;
      LAYER met4 ;
        RECT 56.840000 87.410000 57.160000 87.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840000 87.815000 57.160000 88.135000 ;
      LAYER met4 ;
        RECT 56.840000 87.815000 57.160000 88.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.860000 17.800000 57.180000 18.120000 ;
      LAYER met4 ;
        RECT 56.860000 17.800000 57.180000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.860000 18.230000 57.180000 18.550000 ;
      LAYER met4 ;
        RECT 56.860000 18.230000 57.180000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.860000 18.660000 57.180000 18.980000 ;
      LAYER met4 ;
        RECT 56.860000 18.660000 57.180000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.860000 19.090000 57.180000 19.410000 ;
      LAYER met4 ;
        RECT 56.860000 19.090000 57.180000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.860000 19.520000 57.180000 19.840000 ;
      LAYER met4 ;
        RECT 56.860000 19.520000 57.180000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.860000 19.950000 57.180000 20.270000 ;
      LAYER met4 ;
        RECT 56.860000 19.950000 57.180000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.860000 20.380000 57.180000 20.700000 ;
      LAYER met4 ;
        RECT 56.860000 20.380000 57.180000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.860000 20.810000 57.180000 21.130000 ;
      LAYER met4 ;
        RECT 56.860000 20.810000 57.180000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.860000 21.240000 57.180000 21.560000 ;
      LAYER met4 ;
        RECT 56.860000 21.240000 57.180000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.860000 21.670000 57.180000 21.990000 ;
      LAYER met4 ;
        RECT 56.860000 21.670000 57.180000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.860000 22.100000 57.180000 22.420000 ;
      LAYER met4 ;
        RECT 56.860000 22.100000 57.180000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 68.065000 57.270000 68.385000 ;
      LAYER met4 ;
        RECT 56.950000 68.065000 57.270000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 68.475000 57.270000 68.795000 ;
      LAYER met4 ;
        RECT 56.950000 68.475000 57.270000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 68.885000 57.270000 69.205000 ;
      LAYER met4 ;
        RECT 56.950000 68.885000 57.270000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 69.295000 57.270000 69.615000 ;
      LAYER met4 ;
        RECT 56.950000 69.295000 57.270000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 69.705000 57.270000 70.025000 ;
      LAYER met4 ;
        RECT 56.950000 69.705000 57.270000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 70.115000 57.270000 70.435000 ;
      LAYER met4 ;
        RECT 56.950000 70.115000 57.270000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 70.525000 57.270000 70.845000 ;
      LAYER met4 ;
        RECT 56.950000 70.525000 57.270000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 70.935000 57.270000 71.255000 ;
      LAYER met4 ;
        RECT 56.950000 70.935000 57.270000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 71.345000 57.270000 71.665000 ;
      LAYER met4 ;
        RECT 56.950000 71.345000 57.270000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 71.755000 57.270000 72.075000 ;
      LAYER met4 ;
        RECT 56.950000 71.755000 57.270000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 72.165000 57.270000 72.485000 ;
      LAYER met4 ;
        RECT 56.950000 72.165000 57.270000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 72.575000 57.270000 72.895000 ;
      LAYER met4 ;
        RECT 56.950000 72.575000 57.270000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 72.985000 57.270000 73.305000 ;
      LAYER met4 ;
        RECT 56.950000 72.985000 57.270000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 73.390000 57.270000 73.710000 ;
      LAYER met4 ;
        RECT 56.950000 73.390000 57.270000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 73.795000 57.270000 74.115000 ;
      LAYER met4 ;
        RECT 56.950000 73.795000 57.270000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 74.200000 57.270000 74.520000 ;
      LAYER met4 ;
        RECT 56.950000 74.200000 57.270000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 74.605000 57.270000 74.925000 ;
      LAYER met4 ;
        RECT 56.950000 74.605000 57.270000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 75.010000 57.270000 75.330000 ;
      LAYER met4 ;
        RECT 56.950000 75.010000 57.270000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 75.415000 57.270000 75.735000 ;
      LAYER met4 ;
        RECT 56.950000 75.415000 57.270000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 75.820000 57.270000 76.140000 ;
      LAYER met4 ;
        RECT 56.950000 75.820000 57.270000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 76.225000 57.270000 76.545000 ;
      LAYER met4 ;
        RECT 56.950000 76.225000 57.270000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 76.630000 57.270000 76.950000 ;
      LAYER met4 ;
        RECT 56.950000 76.630000 57.270000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 77.035000 57.270000 77.355000 ;
      LAYER met4 ;
        RECT 56.950000 77.035000 57.270000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 77.440000 57.270000 77.760000 ;
      LAYER met4 ;
        RECT 56.950000 77.440000 57.270000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 77.845000 57.270000 78.165000 ;
      LAYER met4 ;
        RECT 56.950000 77.845000 57.270000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 78.250000 57.270000 78.570000 ;
      LAYER met4 ;
        RECT 56.950000 78.250000 57.270000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 78.655000 57.270000 78.975000 ;
      LAYER met4 ;
        RECT 56.950000 78.655000 57.270000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 79.060000 57.270000 79.380000 ;
      LAYER met4 ;
        RECT 56.950000 79.060000 57.270000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 79.465000 57.270000 79.785000 ;
      LAYER met4 ;
        RECT 56.950000 79.465000 57.270000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 79.870000 57.270000 80.190000 ;
      LAYER met4 ;
        RECT 56.950000 79.870000 57.270000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 80.275000 57.270000 80.595000 ;
      LAYER met4 ;
        RECT 56.950000 80.275000 57.270000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 80.680000 57.270000 81.000000 ;
      LAYER met4 ;
        RECT 56.950000 80.680000 57.270000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 81.085000 57.270000 81.405000 ;
      LAYER met4 ;
        RECT 56.950000 81.085000 57.270000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 81.490000 57.270000 81.810000 ;
      LAYER met4 ;
        RECT 56.950000 81.490000 57.270000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 81.895000 57.270000 82.215000 ;
      LAYER met4 ;
        RECT 56.950000 81.895000 57.270000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950000 82.300000 57.270000 82.620000 ;
      LAYER met4 ;
        RECT 56.950000 82.300000 57.270000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250000 82.995000 57.570000 83.315000 ;
      LAYER met4 ;
        RECT 57.250000 82.995000 57.570000 83.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250000 83.395000 57.570000 83.715000 ;
      LAYER met4 ;
        RECT 57.250000 83.395000 57.570000 83.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250000 83.795000 57.570000 84.115000 ;
      LAYER met4 ;
        RECT 57.250000 83.795000 57.570000 84.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250000 84.195000 57.570000 84.515000 ;
      LAYER met4 ;
        RECT 57.250000 84.195000 57.570000 84.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250000 84.595000 57.570000 84.915000 ;
      LAYER met4 ;
        RECT 57.250000 84.595000 57.570000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250000 84.995000 57.570000 85.315000 ;
      LAYER met4 ;
        RECT 57.250000 84.995000 57.570000 85.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250000 85.395000 57.570000 85.715000 ;
      LAYER met4 ;
        RECT 57.250000 85.395000 57.570000 85.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250000 85.795000 57.570000 86.115000 ;
      LAYER met4 ;
        RECT 57.250000 85.795000 57.570000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250000 86.195000 57.570000 86.515000 ;
      LAYER met4 ;
        RECT 57.250000 86.195000 57.570000 86.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250000 86.600000 57.570000 86.920000 ;
      LAYER met4 ;
        RECT 57.250000 86.600000 57.570000 86.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250000 87.005000 57.570000 87.325000 ;
      LAYER met4 ;
        RECT 57.250000 87.005000 57.570000 87.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250000 87.410000 57.570000 87.730000 ;
      LAYER met4 ;
        RECT 57.250000 87.410000 57.570000 87.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250000 87.815000 57.570000 88.135000 ;
      LAYER met4 ;
        RECT 57.250000 87.815000 57.570000 88.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.265000 17.800000 57.585000 18.120000 ;
      LAYER met4 ;
        RECT 57.265000 17.800000 57.585000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.265000 18.230000 57.585000 18.550000 ;
      LAYER met4 ;
        RECT 57.265000 18.230000 57.585000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.265000 18.660000 57.585000 18.980000 ;
      LAYER met4 ;
        RECT 57.265000 18.660000 57.585000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.265000 19.090000 57.585000 19.410000 ;
      LAYER met4 ;
        RECT 57.265000 19.090000 57.585000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.265000 19.520000 57.585000 19.840000 ;
      LAYER met4 ;
        RECT 57.265000 19.520000 57.585000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.265000 19.950000 57.585000 20.270000 ;
      LAYER met4 ;
        RECT 57.265000 19.950000 57.585000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.265000 20.380000 57.585000 20.700000 ;
      LAYER met4 ;
        RECT 57.265000 20.380000 57.585000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.265000 20.810000 57.585000 21.130000 ;
      LAYER met4 ;
        RECT 57.265000 20.810000 57.585000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.265000 21.240000 57.585000 21.560000 ;
      LAYER met4 ;
        RECT 57.265000 21.240000 57.585000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.265000 21.670000 57.585000 21.990000 ;
      LAYER met4 ;
        RECT 57.265000 21.670000 57.585000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.265000 22.100000 57.585000 22.420000 ;
      LAYER met4 ;
        RECT 57.265000 22.100000 57.585000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 68.065000 57.670000 68.385000 ;
      LAYER met4 ;
        RECT 57.350000 68.065000 57.670000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 68.475000 57.670000 68.795000 ;
      LAYER met4 ;
        RECT 57.350000 68.475000 57.670000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 68.885000 57.670000 69.205000 ;
      LAYER met4 ;
        RECT 57.350000 68.885000 57.670000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 69.295000 57.670000 69.615000 ;
      LAYER met4 ;
        RECT 57.350000 69.295000 57.670000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 69.705000 57.670000 70.025000 ;
      LAYER met4 ;
        RECT 57.350000 69.705000 57.670000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 70.115000 57.670000 70.435000 ;
      LAYER met4 ;
        RECT 57.350000 70.115000 57.670000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 70.525000 57.670000 70.845000 ;
      LAYER met4 ;
        RECT 57.350000 70.525000 57.670000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 70.935000 57.670000 71.255000 ;
      LAYER met4 ;
        RECT 57.350000 70.935000 57.670000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 71.345000 57.670000 71.665000 ;
      LAYER met4 ;
        RECT 57.350000 71.345000 57.670000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 71.755000 57.670000 72.075000 ;
      LAYER met4 ;
        RECT 57.350000 71.755000 57.670000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 72.165000 57.670000 72.485000 ;
      LAYER met4 ;
        RECT 57.350000 72.165000 57.670000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 72.575000 57.670000 72.895000 ;
      LAYER met4 ;
        RECT 57.350000 72.575000 57.670000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 72.985000 57.670000 73.305000 ;
      LAYER met4 ;
        RECT 57.350000 72.985000 57.670000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 73.390000 57.670000 73.710000 ;
      LAYER met4 ;
        RECT 57.350000 73.390000 57.670000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 73.795000 57.670000 74.115000 ;
      LAYER met4 ;
        RECT 57.350000 73.795000 57.670000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 74.200000 57.670000 74.520000 ;
      LAYER met4 ;
        RECT 57.350000 74.200000 57.670000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 74.605000 57.670000 74.925000 ;
      LAYER met4 ;
        RECT 57.350000 74.605000 57.670000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 75.010000 57.670000 75.330000 ;
      LAYER met4 ;
        RECT 57.350000 75.010000 57.670000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 75.415000 57.670000 75.735000 ;
      LAYER met4 ;
        RECT 57.350000 75.415000 57.670000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 75.820000 57.670000 76.140000 ;
      LAYER met4 ;
        RECT 57.350000 75.820000 57.670000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 76.225000 57.670000 76.545000 ;
      LAYER met4 ;
        RECT 57.350000 76.225000 57.670000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 76.630000 57.670000 76.950000 ;
      LAYER met4 ;
        RECT 57.350000 76.630000 57.670000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 77.035000 57.670000 77.355000 ;
      LAYER met4 ;
        RECT 57.350000 77.035000 57.670000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 77.440000 57.670000 77.760000 ;
      LAYER met4 ;
        RECT 57.350000 77.440000 57.670000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 77.845000 57.670000 78.165000 ;
      LAYER met4 ;
        RECT 57.350000 77.845000 57.670000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 78.250000 57.670000 78.570000 ;
      LAYER met4 ;
        RECT 57.350000 78.250000 57.670000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 78.655000 57.670000 78.975000 ;
      LAYER met4 ;
        RECT 57.350000 78.655000 57.670000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 79.060000 57.670000 79.380000 ;
      LAYER met4 ;
        RECT 57.350000 79.060000 57.670000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 79.465000 57.670000 79.785000 ;
      LAYER met4 ;
        RECT 57.350000 79.465000 57.670000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 79.870000 57.670000 80.190000 ;
      LAYER met4 ;
        RECT 57.350000 79.870000 57.670000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 80.275000 57.670000 80.595000 ;
      LAYER met4 ;
        RECT 57.350000 80.275000 57.670000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 80.680000 57.670000 81.000000 ;
      LAYER met4 ;
        RECT 57.350000 80.680000 57.670000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 81.085000 57.670000 81.405000 ;
      LAYER met4 ;
        RECT 57.350000 81.085000 57.670000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 81.490000 57.670000 81.810000 ;
      LAYER met4 ;
        RECT 57.350000 81.490000 57.670000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 81.895000 57.670000 82.215000 ;
      LAYER met4 ;
        RECT 57.350000 81.895000 57.670000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.350000 82.300000 57.670000 82.620000 ;
      LAYER met4 ;
        RECT 57.350000 82.300000 57.670000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660000 82.995000 57.980000 83.315000 ;
      LAYER met4 ;
        RECT 57.660000 82.995000 57.980000 83.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660000 83.395000 57.980000 83.715000 ;
      LAYER met4 ;
        RECT 57.660000 83.395000 57.980000 83.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660000 83.795000 57.980000 84.115000 ;
      LAYER met4 ;
        RECT 57.660000 83.795000 57.980000 84.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660000 84.195000 57.980000 84.515000 ;
      LAYER met4 ;
        RECT 57.660000 84.195000 57.980000 84.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660000 84.595000 57.980000 84.915000 ;
      LAYER met4 ;
        RECT 57.660000 84.595000 57.980000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660000 84.995000 57.980000 85.315000 ;
      LAYER met4 ;
        RECT 57.660000 84.995000 57.980000 85.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660000 85.395000 57.980000 85.715000 ;
      LAYER met4 ;
        RECT 57.660000 85.395000 57.980000 85.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660000 85.795000 57.980000 86.115000 ;
      LAYER met4 ;
        RECT 57.660000 85.795000 57.980000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660000 86.195000 57.980000 86.515000 ;
      LAYER met4 ;
        RECT 57.660000 86.195000 57.980000 86.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660000 86.600000 57.980000 86.920000 ;
      LAYER met4 ;
        RECT 57.660000 86.600000 57.980000 86.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660000 87.005000 57.980000 87.325000 ;
      LAYER met4 ;
        RECT 57.660000 87.005000 57.980000 87.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660000 87.410000 57.980000 87.730000 ;
      LAYER met4 ;
        RECT 57.660000 87.410000 57.980000 87.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660000 87.815000 57.980000 88.135000 ;
      LAYER met4 ;
        RECT 57.660000 87.815000 57.980000 88.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.670000 17.800000 57.990000 18.120000 ;
      LAYER met4 ;
        RECT 57.670000 17.800000 57.990000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.670000 18.230000 57.990000 18.550000 ;
      LAYER met4 ;
        RECT 57.670000 18.230000 57.990000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.670000 18.660000 57.990000 18.980000 ;
      LAYER met4 ;
        RECT 57.670000 18.660000 57.990000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.670000 19.090000 57.990000 19.410000 ;
      LAYER met4 ;
        RECT 57.670000 19.090000 57.990000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.670000 19.520000 57.990000 19.840000 ;
      LAYER met4 ;
        RECT 57.670000 19.520000 57.990000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.670000 19.950000 57.990000 20.270000 ;
      LAYER met4 ;
        RECT 57.670000 19.950000 57.990000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.670000 20.380000 57.990000 20.700000 ;
      LAYER met4 ;
        RECT 57.670000 20.380000 57.990000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.670000 20.810000 57.990000 21.130000 ;
      LAYER met4 ;
        RECT 57.670000 20.810000 57.990000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.670000 21.240000 57.990000 21.560000 ;
      LAYER met4 ;
        RECT 57.670000 21.240000 57.990000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.670000 21.670000 57.990000 21.990000 ;
      LAYER met4 ;
        RECT 57.670000 21.670000 57.990000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.670000 22.100000 57.990000 22.420000 ;
      LAYER met4 ;
        RECT 57.670000 22.100000 57.990000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.735000 88.370000 58.055000 88.690000 ;
      LAYER met4 ;
        RECT 57.735000 88.370000 58.055000 88.690000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.735000 88.785000 58.055000 89.105000 ;
      LAYER met4 ;
        RECT 57.735000 88.785000 58.055000 89.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.735000 89.205000 58.055000 89.525000 ;
      LAYER met4 ;
        RECT 57.735000 89.205000 58.055000 89.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 68.065000 58.070000 68.385000 ;
      LAYER met4 ;
        RECT 57.750000 68.065000 58.070000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 68.475000 58.070000 68.795000 ;
      LAYER met4 ;
        RECT 57.750000 68.475000 58.070000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 68.885000 58.070000 69.205000 ;
      LAYER met4 ;
        RECT 57.750000 68.885000 58.070000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 69.295000 58.070000 69.615000 ;
      LAYER met4 ;
        RECT 57.750000 69.295000 58.070000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 69.705000 58.070000 70.025000 ;
      LAYER met4 ;
        RECT 57.750000 69.705000 58.070000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 70.115000 58.070000 70.435000 ;
      LAYER met4 ;
        RECT 57.750000 70.115000 58.070000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 70.525000 58.070000 70.845000 ;
      LAYER met4 ;
        RECT 57.750000 70.525000 58.070000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 70.935000 58.070000 71.255000 ;
      LAYER met4 ;
        RECT 57.750000 70.935000 58.070000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 71.345000 58.070000 71.665000 ;
      LAYER met4 ;
        RECT 57.750000 71.345000 58.070000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 71.755000 58.070000 72.075000 ;
      LAYER met4 ;
        RECT 57.750000 71.755000 58.070000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 72.165000 58.070000 72.485000 ;
      LAYER met4 ;
        RECT 57.750000 72.165000 58.070000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 72.575000 58.070000 72.895000 ;
      LAYER met4 ;
        RECT 57.750000 72.575000 58.070000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 72.985000 58.070000 73.305000 ;
      LAYER met4 ;
        RECT 57.750000 72.985000 58.070000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 73.390000 58.070000 73.710000 ;
      LAYER met4 ;
        RECT 57.750000 73.390000 58.070000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 73.795000 58.070000 74.115000 ;
      LAYER met4 ;
        RECT 57.750000 73.795000 58.070000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 74.200000 58.070000 74.520000 ;
      LAYER met4 ;
        RECT 57.750000 74.200000 58.070000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 74.605000 58.070000 74.925000 ;
      LAYER met4 ;
        RECT 57.750000 74.605000 58.070000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 75.010000 58.070000 75.330000 ;
      LAYER met4 ;
        RECT 57.750000 75.010000 58.070000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 75.415000 58.070000 75.735000 ;
      LAYER met4 ;
        RECT 57.750000 75.415000 58.070000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 75.820000 58.070000 76.140000 ;
      LAYER met4 ;
        RECT 57.750000 75.820000 58.070000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 76.225000 58.070000 76.545000 ;
      LAYER met4 ;
        RECT 57.750000 76.225000 58.070000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 76.630000 58.070000 76.950000 ;
      LAYER met4 ;
        RECT 57.750000 76.630000 58.070000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 77.035000 58.070000 77.355000 ;
      LAYER met4 ;
        RECT 57.750000 77.035000 58.070000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 77.440000 58.070000 77.760000 ;
      LAYER met4 ;
        RECT 57.750000 77.440000 58.070000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 77.845000 58.070000 78.165000 ;
      LAYER met4 ;
        RECT 57.750000 77.845000 58.070000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 78.250000 58.070000 78.570000 ;
      LAYER met4 ;
        RECT 57.750000 78.250000 58.070000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 78.655000 58.070000 78.975000 ;
      LAYER met4 ;
        RECT 57.750000 78.655000 58.070000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 79.060000 58.070000 79.380000 ;
      LAYER met4 ;
        RECT 57.750000 79.060000 58.070000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 79.465000 58.070000 79.785000 ;
      LAYER met4 ;
        RECT 57.750000 79.465000 58.070000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 79.870000 58.070000 80.190000 ;
      LAYER met4 ;
        RECT 57.750000 79.870000 58.070000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 80.275000 58.070000 80.595000 ;
      LAYER met4 ;
        RECT 57.750000 80.275000 58.070000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 80.680000 58.070000 81.000000 ;
      LAYER met4 ;
        RECT 57.750000 80.680000 58.070000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 81.085000 58.070000 81.405000 ;
      LAYER met4 ;
        RECT 57.750000 81.085000 58.070000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 81.490000 58.070000 81.810000 ;
      LAYER met4 ;
        RECT 57.750000 81.490000 58.070000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 81.895000 58.070000 82.215000 ;
      LAYER met4 ;
        RECT 57.750000 81.895000 58.070000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.750000 82.300000 58.070000 82.620000 ;
      LAYER met4 ;
        RECT 57.750000 82.300000 58.070000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070000 82.995000 58.390000 83.315000 ;
      LAYER met4 ;
        RECT 58.070000 82.995000 58.390000 83.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070000 83.395000 58.390000 83.715000 ;
      LAYER met4 ;
        RECT 58.070000 83.395000 58.390000 83.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070000 83.795000 58.390000 84.115000 ;
      LAYER met4 ;
        RECT 58.070000 83.795000 58.390000 84.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070000 84.195000 58.390000 84.515000 ;
      LAYER met4 ;
        RECT 58.070000 84.195000 58.390000 84.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070000 84.595000 58.390000 84.915000 ;
      LAYER met4 ;
        RECT 58.070000 84.595000 58.390000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070000 84.995000 58.390000 85.315000 ;
      LAYER met4 ;
        RECT 58.070000 84.995000 58.390000 85.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070000 85.395000 58.390000 85.715000 ;
      LAYER met4 ;
        RECT 58.070000 85.395000 58.390000 85.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070000 85.795000 58.390000 86.115000 ;
      LAYER met4 ;
        RECT 58.070000 85.795000 58.390000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070000 86.195000 58.390000 86.515000 ;
      LAYER met4 ;
        RECT 58.070000 86.195000 58.390000 86.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070000 86.600000 58.390000 86.920000 ;
      LAYER met4 ;
        RECT 58.070000 86.600000 58.390000 86.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070000 87.005000 58.390000 87.325000 ;
      LAYER met4 ;
        RECT 58.070000 87.005000 58.390000 87.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070000 87.410000 58.390000 87.730000 ;
      LAYER met4 ;
        RECT 58.070000 87.410000 58.390000 87.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070000 87.815000 58.390000 88.135000 ;
      LAYER met4 ;
        RECT 58.070000 87.815000 58.390000 88.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.075000 17.800000 58.395000 18.120000 ;
      LAYER met4 ;
        RECT 58.075000 17.800000 58.395000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.075000 18.230000 58.395000 18.550000 ;
      LAYER met4 ;
        RECT 58.075000 18.230000 58.395000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.075000 18.660000 58.395000 18.980000 ;
      LAYER met4 ;
        RECT 58.075000 18.660000 58.395000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.075000 19.090000 58.395000 19.410000 ;
      LAYER met4 ;
        RECT 58.075000 19.090000 58.395000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.075000 19.520000 58.395000 19.840000 ;
      LAYER met4 ;
        RECT 58.075000 19.520000 58.395000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.075000 19.950000 58.395000 20.270000 ;
      LAYER met4 ;
        RECT 58.075000 19.950000 58.395000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.075000 20.380000 58.395000 20.700000 ;
      LAYER met4 ;
        RECT 58.075000 20.380000 58.395000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.075000 20.810000 58.395000 21.130000 ;
      LAYER met4 ;
        RECT 58.075000 20.810000 58.395000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.075000 21.240000 58.395000 21.560000 ;
      LAYER met4 ;
        RECT 58.075000 21.240000 58.395000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.075000 21.670000 58.395000 21.990000 ;
      LAYER met4 ;
        RECT 58.075000 21.670000 58.395000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.075000 22.100000 58.395000 22.420000 ;
      LAYER met4 ;
        RECT 58.075000 22.100000 58.395000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 68.065000 58.470000 68.385000 ;
      LAYER met4 ;
        RECT 58.150000 68.065000 58.470000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 68.475000 58.470000 68.795000 ;
      LAYER met4 ;
        RECT 58.150000 68.475000 58.470000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 68.885000 58.470000 69.205000 ;
      LAYER met4 ;
        RECT 58.150000 68.885000 58.470000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 69.295000 58.470000 69.615000 ;
      LAYER met4 ;
        RECT 58.150000 69.295000 58.470000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 69.705000 58.470000 70.025000 ;
      LAYER met4 ;
        RECT 58.150000 69.705000 58.470000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 70.115000 58.470000 70.435000 ;
      LAYER met4 ;
        RECT 58.150000 70.115000 58.470000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 70.525000 58.470000 70.845000 ;
      LAYER met4 ;
        RECT 58.150000 70.525000 58.470000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 70.935000 58.470000 71.255000 ;
      LAYER met4 ;
        RECT 58.150000 70.935000 58.470000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 71.345000 58.470000 71.665000 ;
      LAYER met4 ;
        RECT 58.150000 71.345000 58.470000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 71.755000 58.470000 72.075000 ;
      LAYER met4 ;
        RECT 58.150000 71.755000 58.470000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 72.165000 58.470000 72.485000 ;
      LAYER met4 ;
        RECT 58.150000 72.165000 58.470000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 72.575000 58.470000 72.895000 ;
      LAYER met4 ;
        RECT 58.150000 72.575000 58.470000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 72.985000 58.470000 73.305000 ;
      LAYER met4 ;
        RECT 58.150000 72.985000 58.470000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 73.390000 58.470000 73.710000 ;
      LAYER met4 ;
        RECT 58.150000 73.390000 58.470000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 73.795000 58.470000 74.115000 ;
      LAYER met4 ;
        RECT 58.150000 73.795000 58.470000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 74.200000 58.470000 74.520000 ;
      LAYER met4 ;
        RECT 58.150000 74.200000 58.470000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 74.605000 58.470000 74.925000 ;
      LAYER met4 ;
        RECT 58.150000 74.605000 58.470000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 75.010000 58.470000 75.330000 ;
      LAYER met4 ;
        RECT 58.150000 75.010000 58.470000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 75.415000 58.470000 75.735000 ;
      LAYER met4 ;
        RECT 58.150000 75.415000 58.470000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 75.820000 58.470000 76.140000 ;
      LAYER met4 ;
        RECT 58.150000 75.820000 58.470000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 76.225000 58.470000 76.545000 ;
      LAYER met4 ;
        RECT 58.150000 76.225000 58.470000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 76.630000 58.470000 76.950000 ;
      LAYER met4 ;
        RECT 58.150000 76.630000 58.470000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 77.035000 58.470000 77.355000 ;
      LAYER met4 ;
        RECT 58.150000 77.035000 58.470000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 77.440000 58.470000 77.760000 ;
      LAYER met4 ;
        RECT 58.150000 77.440000 58.470000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 77.845000 58.470000 78.165000 ;
      LAYER met4 ;
        RECT 58.150000 77.845000 58.470000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 78.250000 58.470000 78.570000 ;
      LAYER met4 ;
        RECT 58.150000 78.250000 58.470000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 78.655000 58.470000 78.975000 ;
      LAYER met4 ;
        RECT 58.150000 78.655000 58.470000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 79.060000 58.470000 79.380000 ;
      LAYER met4 ;
        RECT 58.150000 79.060000 58.470000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 79.465000 58.470000 79.785000 ;
      LAYER met4 ;
        RECT 58.150000 79.465000 58.470000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 79.870000 58.470000 80.190000 ;
      LAYER met4 ;
        RECT 58.150000 79.870000 58.470000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 80.275000 58.470000 80.595000 ;
      LAYER met4 ;
        RECT 58.150000 80.275000 58.470000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 80.680000 58.470000 81.000000 ;
      LAYER met4 ;
        RECT 58.150000 80.680000 58.470000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 81.085000 58.470000 81.405000 ;
      LAYER met4 ;
        RECT 58.150000 81.085000 58.470000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 81.490000 58.470000 81.810000 ;
      LAYER met4 ;
        RECT 58.150000 81.490000 58.470000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 81.895000 58.470000 82.215000 ;
      LAYER met4 ;
        RECT 58.150000 81.895000 58.470000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.150000 82.300000 58.470000 82.620000 ;
      LAYER met4 ;
        RECT 58.150000 82.300000 58.470000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 17.800000 58.800000 18.120000 ;
      LAYER met4 ;
        RECT 58.480000 17.800000 58.800000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 18.230000 58.800000 18.550000 ;
      LAYER met4 ;
        RECT 58.480000 18.230000 58.800000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 18.660000 58.800000 18.980000 ;
      LAYER met4 ;
        RECT 58.480000 18.660000 58.800000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 19.090000 58.800000 19.410000 ;
      LAYER met4 ;
        RECT 58.480000 19.090000 58.800000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 19.520000 58.800000 19.840000 ;
      LAYER met4 ;
        RECT 58.480000 19.520000 58.800000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 19.950000 58.800000 20.270000 ;
      LAYER met4 ;
        RECT 58.480000 19.950000 58.800000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 20.380000 58.800000 20.700000 ;
      LAYER met4 ;
        RECT 58.480000 20.380000 58.800000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 20.810000 58.800000 21.130000 ;
      LAYER met4 ;
        RECT 58.480000 20.810000 58.800000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 21.240000 58.800000 21.560000 ;
      LAYER met4 ;
        RECT 58.480000 21.240000 58.800000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 21.670000 58.800000 21.990000 ;
      LAYER met4 ;
        RECT 58.480000 21.670000 58.800000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 22.100000 58.800000 22.420000 ;
      LAYER met4 ;
        RECT 58.480000 22.100000 58.800000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 82.995000 58.800000 83.315000 ;
      LAYER met4 ;
        RECT 58.480000 82.995000 58.800000 83.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 83.395000 58.800000 83.715000 ;
      LAYER met4 ;
        RECT 58.480000 83.395000 58.800000 83.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 83.795000 58.800000 84.115000 ;
      LAYER met4 ;
        RECT 58.480000 83.795000 58.800000 84.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 84.195000 58.800000 84.515000 ;
      LAYER met4 ;
        RECT 58.480000 84.195000 58.800000 84.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 84.595000 58.800000 84.915000 ;
      LAYER met4 ;
        RECT 58.480000 84.595000 58.800000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 84.995000 58.800000 85.315000 ;
      LAYER met4 ;
        RECT 58.480000 84.995000 58.800000 85.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 85.395000 58.800000 85.715000 ;
      LAYER met4 ;
        RECT 58.480000 85.395000 58.800000 85.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 85.795000 58.800000 86.115000 ;
      LAYER met4 ;
        RECT 58.480000 85.795000 58.800000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 86.195000 58.800000 86.515000 ;
      LAYER met4 ;
        RECT 58.480000 86.195000 58.800000 86.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 86.600000 58.800000 86.920000 ;
      LAYER met4 ;
        RECT 58.480000 86.600000 58.800000 86.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 87.005000 58.800000 87.325000 ;
      LAYER met4 ;
        RECT 58.480000 87.005000 58.800000 87.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 87.410000 58.800000 87.730000 ;
      LAYER met4 ;
        RECT 58.480000 87.410000 58.800000 87.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 87.815000 58.800000 88.135000 ;
      LAYER met4 ;
        RECT 58.480000 87.815000 58.800000 88.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.515000 88.370000 58.835000 88.690000 ;
      LAYER met4 ;
        RECT 58.515000 88.370000 58.835000 88.690000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.515000 88.785000 58.835000 89.105000 ;
      LAYER met4 ;
        RECT 58.515000 88.785000 58.835000 89.105000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.515000 89.205000 58.835000 89.525000 ;
      LAYER met4 ;
        RECT 58.515000 89.205000 58.835000 89.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 68.065000 58.870000 68.385000 ;
      LAYER met4 ;
        RECT 58.550000 68.065000 58.870000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 68.475000 58.870000 68.795000 ;
      LAYER met4 ;
        RECT 58.550000 68.475000 58.870000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 68.885000 58.870000 69.205000 ;
      LAYER met4 ;
        RECT 58.550000 68.885000 58.870000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 69.295000 58.870000 69.615000 ;
      LAYER met4 ;
        RECT 58.550000 69.295000 58.870000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 69.705000 58.870000 70.025000 ;
      LAYER met4 ;
        RECT 58.550000 69.705000 58.870000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 70.115000 58.870000 70.435000 ;
      LAYER met4 ;
        RECT 58.550000 70.115000 58.870000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 70.525000 58.870000 70.845000 ;
      LAYER met4 ;
        RECT 58.550000 70.525000 58.870000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 70.935000 58.870000 71.255000 ;
      LAYER met4 ;
        RECT 58.550000 70.935000 58.870000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 71.345000 58.870000 71.665000 ;
      LAYER met4 ;
        RECT 58.550000 71.345000 58.870000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 71.755000 58.870000 72.075000 ;
      LAYER met4 ;
        RECT 58.550000 71.755000 58.870000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 72.165000 58.870000 72.485000 ;
      LAYER met4 ;
        RECT 58.550000 72.165000 58.870000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 72.575000 58.870000 72.895000 ;
      LAYER met4 ;
        RECT 58.550000 72.575000 58.870000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 72.985000 58.870000 73.305000 ;
      LAYER met4 ;
        RECT 58.550000 72.985000 58.870000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 73.390000 58.870000 73.710000 ;
      LAYER met4 ;
        RECT 58.550000 73.390000 58.870000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 73.795000 58.870000 74.115000 ;
      LAYER met4 ;
        RECT 58.550000 73.795000 58.870000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 74.200000 58.870000 74.520000 ;
      LAYER met4 ;
        RECT 58.550000 74.200000 58.870000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 74.605000 58.870000 74.925000 ;
      LAYER met4 ;
        RECT 58.550000 74.605000 58.870000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 75.010000 58.870000 75.330000 ;
      LAYER met4 ;
        RECT 58.550000 75.010000 58.870000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 75.415000 58.870000 75.735000 ;
      LAYER met4 ;
        RECT 58.550000 75.415000 58.870000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 75.820000 58.870000 76.140000 ;
      LAYER met4 ;
        RECT 58.550000 75.820000 58.870000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 76.225000 58.870000 76.545000 ;
      LAYER met4 ;
        RECT 58.550000 76.225000 58.870000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 76.630000 58.870000 76.950000 ;
      LAYER met4 ;
        RECT 58.550000 76.630000 58.870000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 77.035000 58.870000 77.355000 ;
      LAYER met4 ;
        RECT 58.550000 77.035000 58.870000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 77.440000 58.870000 77.760000 ;
      LAYER met4 ;
        RECT 58.550000 77.440000 58.870000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 77.845000 58.870000 78.165000 ;
      LAYER met4 ;
        RECT 58.550000 77.845000 58.870000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 78.250000 58.870000 78.570000 ;
      LAYER met4 ;
        RECT 58.550000 78.250000 58.870000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 78.655000 58.870000 78.975000 ;
      LAYER met4 ;
        RECT 58.550000 78.655000 58.870000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 79.060000 58.870000 79.380000 ;
      LAYER met4 ;
        RECT 58.550000 79.060000 58.870000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 79.465000 58.870000 79.785000 ;
      LAYER met4 ;
        RECT 58.550000 79.465000 58.870000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 79.870000 58.870000 80.190000 ;
      LAYER met4 ;
        RECT 58.550000 79.870000 58.870000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 80.275000 58.870000 80.595000 ;
      LAYER met4 ;
        RECT 58.550000 80.275000 58.870000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 80.680000 58.870000 81.000000 ;
      LAYER met4 ;
        RECT 58.550000 80.680000 58.870000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 81.085000 58.870000 81.405000 ;
      LAYER met4 ;
        RECT 58.550000 81.085000 58.870000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 81.490000 58.870000 81.810000 ;
      LAYER met4 ;
        RECT 58.550000 81.490000 58.870000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 81.895000 58.870000 82.215000 ;
      LAYER met4 ;
        RECT 58.550000 81.895000 58.870000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 82.300000 58.870000 82.620000 ;
      LAYER met4 ;
        RECT 58.550000 82.300000 58.870000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.885000 17.800000 59.205000 18.120000 ;
      LAYER met4 ;
        RECT 58.885000 17.800000 59.205000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.885000 18.230000 59.205000 18.550000 ;
      LAYER met4 ;
        RECT 58.885000 18.230000 59.205000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.885000 18.660000 59.205000 18.980000 ;
      LAYER met4 ;
        RECT 58.885000 18.660000 59.205000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.885000 19.090000 59.205000 19.410000 ;
      LAYER met4 ;
        RECT 58.885000 19.090000 59.205000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.885000 19.520000 59.205000 19.840000 ;
      LAYER met4 ;
        RECT 58.885000 19.520000 59.205000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.885000 19.950000 59.205000 20.270000 ;
      LAYER met4 ;
        RECT 58.885000 19.950000 59.205000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.885000 20.380000 59.205000 20.700000 ;
      LAYER met4 ;
        RECT 58.885000 20.380000 59.205000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.885000 20.810000 59.205000 21.130000 ;
      LAYER met4 ;
        RECT 58.885000 20.810000 59.205000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.885000 21.240000 59.205000 21.560000 ;
      LAYER met4 ;
        RECT 58.885000 21.240000 59.205000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.885000 21.670000 59.205000 21.990000 ;
      LAYER met4 ;
        RECT 58.885000 21.670000 59.205000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.885000 22.100000 59.205000 22.420000 ;
      LAYER met4 ;
        RECT 58.885000 22.100000 59.205000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890000 82.995000 59.210000 83.315000 ;
      LAYER met4 ;
        RECT 58.890000 82.995000 59.210000 83.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890000 83.395000 59.210000 83.715000 ;
      LAYER met4 ;
        RECT 58.890000 83.395000 59.210000 83.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890000 83.795000 59.210000 84.115000 ;
      LAYER met4 ;
        RECT 58.890000 83.795000 59.210000 84.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890000 84.195000 59.210000 84.515000 ;
      LAYER met4 ;
        RECT 58.890000 84.195000 59.210000 84.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890000 84.595000 59.210000 84.915000 ;
      LAYER met4 ;
        RECT 58.890000 84.595000 59.210000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890000 84.995000 59.210000 85.315000 ;
      LAYER met4 ;
        RECT 58.890000 84.995000 59.210000 85.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890000 85.395000 59.210000 85.715000 ;
      LAYER met4 ;
        RECT 58.890000 85.395000 59.210000 85.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890000 85.795000 59.210000 86.115000 ;
      LAYER met4 ;
        RECT 58.890000 85.795000 59.210000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890000 86.195000 59.210000 86.515000 ;
      LAYER met4 ;
        RECT 58.890000 86.195000 59.210000 86.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890000 86.600000 59.210000 86.920000 ;
      LAYER met4 ;
        RECT 58.890000 86.600000 59.210000 86.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890000 87.005000 59.210000 87.325000 ;
      LAYER met4 ;
        RECT 58.890000 87.005000 59.210000 87.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890000 87.410000 59.210000 87.730000 ;
      LAYER met4 ;
        RECT 58.890000 87.410000 59.210000 87.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890000 87.815000 59.210000 88.135000 ;
      LAYER met4 ;
        RECT 58.890000 87.815000 59.210000 88.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 68.065000 59.270000 68.385000 ;
      LAYER met4 ;
        RECT 58.950000 68.065000 59.270000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 68.475000 59.270000 68.795000 ;
      LAYER met4 ;
        RECT 58.950000 68.475000 59.270000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 68.885000 59.270000 69.205000 ;
      LAYER met4 ;
        RECT 58.950000 68.885000 59.270000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 69.295000 59.270000 69.615000 ;
      LAYER met4 ;
        RECT 58.950000 69.295000 59.270000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 69.705000 59.270000 70.025000 ;
      LAYER met4 ;
        RECT 58.950000 69.705000 59.270000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 70.115000 59.270000 70.435000 ;
      LAYER met4 ;
        RECT 58.950000 70.115000 59.270000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 70.525000 59.270000 70.845000 ;
      LAYER met4 ;
        RECT 58.950000 70.525000 59.270000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 70.935000 59.270000 71.255000 ;
      LAYER met4 ;
        RECT 58.950000 70.935000 59.270000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 71.345000 59.270000 71.665000 ;
      LAYER met4 ;
        RECT 58.950000 71.345000 59.270000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 71.755000 59.270000 72.075000 ;
      LAYER met4 ;
        RECT 58.950000 71.755000 59.270000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 72.165000 59.270000 72.485000 ;
      LAYER met4 ;
        RECT 58.950000 72.165000 59.270000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 72.575000 59.270000 72.895000 ;
      LAYER met4 ;
        RECT 58.950000 72.575000 59.270000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 72.985000 59.270000 73.305000 ;
      LAYER met4 ;
        RECT 58.950000 72.985000 59.270000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 73.390000 59.270000 73.710000 ;
      LAYER met4 ;
        RECT 58.950000 73.390000 59.270000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 73.795000 59.270000 74.115000 ;
      LAYER met4 ;
        RECT 58.950000 73.795000 59.270000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 74.200000 59.270000 74.520000 ;
      LAYER met4 ;
        RECT 58.950000 74.200000 59.270000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 74.605000 59.270000 74.925000 ;
      LAYER met4 ;
        RECT 58.950000 74.605000 59.270000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 75.010000 59.270000 75.330000 ;
      LAYER met4 ;
        RECT 58.950000 75.010000 59.270000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 75.415000 59.270000 75.735000 ;
      LAYER met4 ;
        RECT 58.950000 75.415000 59.270000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 75.820000 59.270000 76.140000 ;
      LAYER met4 ;
        RECT 58.950000 75.820000 59.270000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 76.225000 59.270000 76.545000 ;
      LAYER met4 ;
        RECT 58.950000 76.225000 59.270000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 76.630000 59.270000 76.950000 ;
      LAYER met4 ;
        RECT 58.950000 76.630000 59.270000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 77.035000 59.270000 77.355000 ;
      LAYER met4 ;
        RECT 58.950000 77.035000 59.270000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 77.440000 59.270000 77.760000 ;
      LAYER met4 ;
        RECT 58.950000 77.440000 59.270000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 77.845000 59.270000 78.165000 ;
      LAYER met4 ;
        RECT 58.950000 77.845000 59.270000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 78.250000 59.270000 78.570000 ;
      LAYER met4 ;
        RECT 58.950000 78.250000 59.270000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 78.655000 59.270000 78.975000 ;
      LAYER met4 ;
        RECT 58.950000 78.655000 59.270000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 79.060000 59.270000 79.380000 ;
      LAYER met4 ;
        RECT 58.950000 79.060000 59.270000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 79.465000 59.270000 79.785000 ;
      LAYER met4 ;
        RECT 58.950000 79.465000 59.270000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 79.870000 59.270000 80.190000 ;
      LAYER met4 ;
        RECT 58.950000 79.870000 59.270000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 80.275000 59.270000 80.595000 ;
      LAYER met4 ;
        RECT 58.950000 80.275000 59.270000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 80.680000 59.270000 81.000000 ;
      LAYER met4 ;
        RECT 58.950000 80.680000 59.270000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 81.085000 59.270000 81.405000 ;
      LAYER met4 ;
        RECT 58.950000 81.085000 59.270000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 81.490000 59.270000 81.810000 ;
      LAYER met4 ;
        RECT 58.950000 81.490000 59.270000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 81.895000 59.270000 82.215000 ;
      LAYER met4 ;
        RECT 58.950000 81.895000 59.270000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950000 82.300000 59.270000 82.620000 ;
      LAYER met4 ;
        RECT 58.950000 82.300000 59.270000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015000 88.350000 59.335000 88.670000 ;
      LAYER met4 ;
        RECT 59.015000 88.350000 59.335000 88.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015000 88.775000 59.335000 89.095000 ;
      LAYER met4 ;
        RECT 59.015000 88.775000 59.335000 89.095000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015000 89.205000 59.335000 89.525000 ;
      LAYER met4 ;
        RECT 59.015000 89.205000 59.335000 89.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015000 89.635000 59.335000 89.955000 ;
      LAYER met4 ;
        RECT 59.015000 89.635000 59.335000 89.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015000 90.065000 59.335000 90.385000 ;
      LAYER met4 ;
        RECT 59.015000 90.065000 59.335000 90.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015000 90.495000 59.335000 90.815000 ;
      LAYER met4 ;
        RECT 59.015000 90.495000 59.335000 90.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.290000 17.800000 59.610000 18.120000 ;
      LAYER met4 ;
        RECT 59.290000 17.800000 59.610000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.290000 18.230000 59.610000 18.550000 ;
      LAYER met4 ;
        RECT 59.290000 18.230000 59.610000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.290000 18.660000 59.610000 18.980000 ;
      LAYER met4 ;
        RECT 59.290000 18.660000 59.610000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.290000 19.090000 59.610000 19.410000 ;
      LAYER met4 ;
        RECT 59.290000 19.090000 59.610000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.290000 19.520000 59.610000 19.840000 ;
      LAYER met4 ;
        RECT 59.290000 19.520000 59.610000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.290000 19.950000 59.610000 20.270000 ;
      LAYER met4 ;
        RECT 59.290000 19.950000 59.610000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.290000 20.380000 59.610000 20.700000 ;
      LAYER met4 ;
        RECT 59.290000 20.380000 59.610000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.290000 20.810000 59.610000 21.130000 ;
      LAYER met4 ;
        RECT 59.290000 20.810000 59.610000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.290000 21.240000 59.610000 21.560000 ;
      LAYER met4 ;
        RECT 59.290000 21.240000 59.610000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.290000 21.670000 59.610000 21.990000 ;
      LAYER met4 ;
        RECT 59.290000 21.670000 59.610000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.290000 22.100000 59.610000 22.420000 ;
      LAYER met4 ;
        RECT 59.290000 22.100000 59.610000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300000 82.995000 59.620000 83.315000 ;
      LAYER met4 ;
        RECT 59.300000 82.995000 59.620000 83.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300000 83.395000 59.620000 83.715000 ;
      LAYER met4 ;
        RECT 59.300000 83.395000 59.620000 83.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300000 83.795000 59.620000 84.115000 ;
      LAYER met4 ;
        RECT 59.300000 83.795000 59.620000 84.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300000 84.195000 59.620000 84.515000 ;
      LAYER met4 ;
        RECT 59.300000 84.195000 59.620000 84.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300000 84.595000 59.620000 84.915000 ;
      LAYER met4 ;
        RECT 59.300000 84.595000 59.620000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300000 84.995000 59.620000 85.315000 ;
      LAYER met4 ;
        RECT 59.300000 84.995000 59.620000 85.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300000 85.395000 59.620000 85.715000 ;
      LAYER met4 ;
        RECT 59.300000 85.395000 59.620000 85.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300000 85.795000 59.620000 86.115000 ;
      LAYER met4 ;
        RECT 59.300000 85.795000 59.620000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300000 86.195000 59.620000 86.515000 ;
      LAYER met4 ;
        RECT 59.300000 86.195000 59.620000 86.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300000 86.600000 59.620000 86.920000 ;
      LAYER met4 ;
        RECT 59.300000 86.600000 59.620000 86.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300000 87.005000 59.620000 87.325000 ;
      LAYER met4 ;
        RECT 59.300000 87.005000 59.620000 87.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300000 87.410000 59.620000 87.730000 ;
      LAYER met4 ;
        RECT 59.300000 87.410000 59.620000 87.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300000 87.815000 59.620000 88.135000 ;
      LAYER met4 ;
        RECT 59.300000 87.815000 59.620000 88.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 68.065000 59.670000 68.385000 ;
      LAYER met4 ;
        RECT 59.350000 68.065000 59.670000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 68.475000 59.670000 68.795000 ;
      LAYER met4 ;
        RECT 59.350000 68.475000 59.670000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 68.885000 59.670000 69.205000 ;
      LAYER met4 ;
        RECT 59.350000 68.885000 59.670000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 69.295000 59.670000 69.615000 ;
      LAYER met4 ;
        RECT 59.350000 69.295000 59.670000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 69.705000 59.670000 70.025000 ;
      LAYER met4 ;
        RECT 59.350000 69.705000 59.670000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 70.115000 59.670000 70.435000 ;
      LAYER met4 ;
        RECT 59.350000 70.115000 59.670000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 70.525000 59.670000 70.845000 ;
      LAYER met4 ;
        RECT 59.350000 70.525000 59.670000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 70.935000 59.670000 71.255000 ;
      LAYER met4 ;
        RECT 59.350000 70.935000 59.670000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 71.345000 59.670000 71.665000 ;
      LAYER met4 ;
        RECT 59.350000 71.345000 59.670000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 71.755000 59.670000 72.075000 ;
      LAYER met4 ;
        RECT 59.350000 71.755000 59.670000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 72.165000 59.670000 72.485000 ;
      LAYER met4 ;
        RECT 59.350000 72.165000 59.670000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 72.575000 59.670000 72.895000 ;
      LAYER met4 ;
        RECT 59.350000 72.575000 59.670000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 72.985000 59.670000 73.305000 ;
      LAYER met4 ;
        RECT 59.350000 72.985000 59.670000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 73.390000 59.670000 73.710000 ;
      LAYER met4 ;
        RECT 59.350000 73.390000 59.670000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 73.795000 59.670000 74.115000 ;
      LAYER met4 ;
        RECT 59.350000 73.795000 59.670000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 74.200000 59.670000 74.520000 ;
      LAYER met4 ;
        RECT 59.350000 74.200000 59.670000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 74.605000 59.670000 74.925000 ;
      LAYER met4 ;
        RECT 59.350000 74.605000 59.670000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 75.010000 59.670000 75.330000 ;
      LAYER met4 ;
        RECT 59.350000 75.010000 59.670000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 75.415000 59.670000 75.735000 ;
      LAYER met4 ;
        RECT 59.350000 75.415000 59.670000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 75.820000 59.670000 76.140000 ;
      LAYER met4 ;
        RECT 59.350000 75.820000 59.670000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 76.225000 59.670000 76.545000 ;
      LAYER met4 ;
        RECT 59.350000 76.225000 59.670000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 76.630000 59.670000 76.950000 ;
      LAYER met4 ;
        RECT 59.350000 76.630000 59.670000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 77.035000 59.670000 77.355000 ;
      LAYER met4 ;
        RECT 59.350000 77.035000 59.670000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 77.440000 59.670000 77.760000 ;
      LAYER met4 ;
        RECT 59.350000 77.440000 59.670000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 77.845000 59.670000 78.165000 ;
      LAYER met4 ;
        RECT 59.350000 77.845000 59.670000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 78.250000 59.670000 78.570000 ;
      LAYER met4 ;
        RECT 59.350000 78.250000 59.670000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 78.655000 59.670000 78.975000 ;
      LAYER met4 ;
        RECT 59.350000 78.655000 59.670000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 79.060000 59.670000 79.380000 ;
      LAYER met4 ;
        RECT 59.350000 79.060000 59.670000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 79.465000 59.670000 79.785000 ;
      LAYER met4 ;
        RECT 59.350000 79.465000 59.670000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 79.870000 59.670000 80.190000 ;
      LAYER met4 ;
        RECT 59.350000 79.870000 59.670000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 80.275000 59.670000 80.595000 ;
      LAYER met4 ;
        RECT 59.350000 80.275000 59.670000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 80.680000 59.670000 81.000000 ;
      LAYER met4 ;
        RECT 59.350000 80.680000 59.670000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 81.085000 59.670000 81.405000 ;
      LAYER met4 ;
        RECT 59.350000 81.085000 59.670000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 81.490000 59.670000 81.810000 ;
      LAYER met4 ;
        RECT 59.350000 81.490000 59.670000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 81.895000 59.670000 82.215000 ;
      LAYER met4 ;
        RECT 59.350000 81.895000 59.670000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350000 82.300000 59.670000 82.620000 ;
      LAYER met4 ;
        RECT 59.350000 82.300000 59.670000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425000 88.350000 59.745000 88.670000 ;
      LAYER met4 ;
        RECT 59.425000 88.350000 59.745000 88.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425000 88.775000 59.745000 89.095000 ;
      LAYER met4 ;
        RECT 59.425000 88.775000 59.745000 89.095000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425000 89.205000 59.745000 89.525000 ;
      LAYER met4 ;
        RECT 59.425000 89.205000 59.745000 89.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425000 89.635000 59.745000 89.955000 ;
      LAYER met4 ;
        RECT 59.425000 89.635000 59.745000 89.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425000 90.065000 59.745000 90.385000 ;
      LAYER met4 ;
        RECT 59.425000 90.065000 59.745000 90.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425000 90.495000 59.745000 90.815000 ;
      LAYER met4 ;
        RECT 59.425000 90.495000 59.745000 90.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.695000 17.800000 60.015000 18.120000 ;
      LAYER met4 ;
        RECT 59.695000 17.800000 60.015000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.695000 18.230000 60.015000 18.550000 ;
      LAYER met4 ;
        RECT 59.695000 18.230000 60.015000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.695000 18.660000 60.015000 18.980000 ;
      LAYER met4 ;
        RECT 59.695000 18.660000 60.015000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.695000 19.090000 60.015000 19.410000 ;
      LAYER met4 ;
        RECT 59.695000 19.090000 60.015000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.695000 19.520000 60.015000 19.840000 ;
      LAYER met4 ;
        RECT 59.695000 19.520000 60.015000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.695000 19.950000 60.015000 20.270000 ;
      LAYER met4 ;
        RECT 59.695000 19.950000 60.015000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.695000 20.380000 60.015000 20.700000 ;
      LAYER met4 ;
        RECT 59.695000 20.380000 60.015000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.695000 20.810000 60.015000 21.130000 ;
      LAYER met4 ;
        RECT 59.695000 20.810000 60.015000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.695000 21.240000 60.015000 21.560000 ;
      LAYER met4 ;
        RECT 59.695000 21.240000 60.015000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.695000 21.670000 60.015000 21.990000 ;
      LAYER met4 ;
        RECT 59.695000 21.670000 60.015000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.695000 22.100000 60.015000 22.420000 ;
      LAYER met4 ;
        RECT 59.695000 22.100000 60.015000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710000 82.995000 60.030000 83.315000 ;
      LAYER met4 ;
        RECT 59.710000 82.995000 60.030000 83.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710000 83.395000 60.030000 83.715000 ;
      LAYER met4 ;
        RECT 59.710000 83.395000 60.030000 83.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710000 83.795000 60.030000 84.115000 ;
      LAYER met4 ;
        RECT 59.710000 83.795000 60.030000 84.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710000 84.195000 60.030000 84.515000 ;
      LAYER met4 ;
        RECT 59.710000 84.195000 60.030000 84.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710000 84.595000 60.030000 84.915000 ;
      LAYER met4 ;
        RECT 59.710000 84.595000 60.030000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710000 84.995000 60.030000 85.315000 ;
      LAYER met4 ;
        RECT 59.710000 84.995000 60.030000 85.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710000 85.395000 60.030000 85.715000 ;
      LAYER met4 ;
        RECT 59.710000 85.395000 60.030000 85.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710000 85.795000 60.030000 86.115000 ;
      LAYER met4 ;
        RECT 59.710000 85.795000 60.030000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710000 86.195000 60.030000 86.515000 ;
      LAYER met4 ;
        RECT 59.710000 86.195000 60.030000 86.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710000 86.600000 60.030000 86.920000 ;
      LAYER met4 ;
        RECT 59.710000 86.600000 60.030000 86.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710000 87.005000 60.030000 87.325000 ;
      LAYER met4 ;
        RECT 59.710000 87.005000 60.030000 87.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710000 87.410000 60.030000 87.730000 ;
      LAYER met4 ;
        RECT 59.710000 87.410000 60.030000 87.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710000 87.815000 60.030000 88.135000 ;
      LAYER met4 ;
        RECT 59.710000 87.815000 60.030000 88.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 68.065000 60.070000 68.385000 ;
      LAYER met4 ;
        RECT 59.750000 68.065000 60.070000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 68.475000 60.070000 68.795000 ;
      LAYER met4 ;
        RECT 59.750000 68.475000 60.070000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 68.885000 60.070000 69.205000 ;
      LAYER met4 ;
        RECT 59.750000 68.885000 60.070000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 69.295000 60.070000 69.615000 ;
      LAYER met4 ;
        RECT 59.750000 69.295000 60.070000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 69.705000 60.070000 70.025000 ;
      LAYER met4 ;
        RECT 59.750000 69.705000 60.070000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 70.115000 60.070000 70.435000 ;
      LAYER met4 ;
        RECT 59.750000 70.115000 60.070000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 70.525000 60.070000 70.845000 ;
      LAYER met4 ;
        RECT 59.750000 70.525000 60.070000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 70.935000 60.070000 71.255000 ;
      LAYER met4 ;
        RECT 59.750000 70.935000 60.070000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 71.345000 60.070000 71.665000 ;
      LAYER met4 ;
        RECT 59.750000 71.345000 60.070000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 71.755000 60.070000 72.075000 ;
      LAYER met4 ;
        RECT 59.750000 71.755000 60.070000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 72.165000 60.070000 72.485000 ;
      LAYER met4 ;
        RECT 59.750000 72.165000 60.070000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 72.575000 60.070000 72.895000 ;
      LAYER met4 ;
        RECT 59.750000 72.575000 60.070000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 72.985000 60.070000 73.305000 ;
      LAYER met4 ;
        RECT 59.750000 72.985000 60.070000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 73.390000 60.070000 73.710000 ;
      LAYER met4 ;
        RECT 59.750000 73.390000 60.070000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 73.795000 60.070000 74.115000 ;
      LAYER met4 ;
        RECT 59.750000 73.795000 60.070000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 74.200000 60.070000 74.520000 ;
      LAYER met4 ;
        RECT 59.750000 74.200000 60.070000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 74.605000 60.070000 74.925000 ;
      LAYER met4 ;
        RECT 59.750000 74.605000 60.070000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 75.010000 60.070000 75.330000 ;
      LAYER met4 ;
        RECT 59.750000 75.010000 60.070000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 75.415000 60.070000 75.735000 ;
      LAYER met4 ;
        RECT 59.750000 75.415000 60.070000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 75.820000 60.070000 76.140000 ;
      LAYER met4 ;
        RECT 59.750000 75.820000 60.070000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 76.225000 60.070000 76.545000 ;
      LAYER met4 ;
        RECT 59.750000 76.225000 60.070000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 76.630000 60.070000 76.950000 ;
      LAYER met4 ;
        RECT 59.750000 76.630000 60.070000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 77.035000 60.070000 77.355000 ;
      LAYER met4 ;
        RECT 59.750000 77.035000 60.070000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 77.440000 60.070000 77.760000 ;
      LAYER met4 ;
        RECT 59.750000 77.440000 60.070000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 77.845000 60.070000 78.165000 ;
      LAYER met4 ;
        RECT 59.750000 77.845000 60.070000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 78.250000 60.070000 78.570000 ;
      LAYER met4 ;
        RECT 59.750000 78.250000 60.070000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 78.655000 60.070000 78.975000 ;
      LAYER met4 ;
        RECT 59.750000 78.655000 60.070000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 79.060000 60.070000 79.380000 ;
      LAYER met4 ;
        RECT 59.750000 79.060000 60.070000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 79.465000 60.070000 79.785000 ;
      LAYER met4 ;
        RECT 59.750000 79.465000 60.070000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 79.870000 60.070000 80.190000 ;
      LAYER met4 ;
        RECT 59.750000 79.870000 60.070000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 80.275000 60.070000 80.595000 ;
      LAYER met4 ;
        RECT 59.750000 80.275000 60.070000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 80.680000 60.070000 81.000000 ;
      LAYER met4 ;
        RECT 59.750000 80.680000 60.070000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 81.085000 60.070000 81.405000 ;
      LAYER met4 ;
        RECT 59.750000 81.085000 60.070000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 81.490000 60.070000 81.810000 ;
      LAYER met4 ;
        RECT 59.750000 81.490000 60.070000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 81.895000 60.070000 82.215000 ;
      LAYER met4 ;
        RECT 59.750000 81.895000 60.070000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.750000 82.300000 60.070000 82.620000 ;
      LAYER met4 ;
        RECT 59.750000 82.300000 60.070000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.835000 88.350000 60.155000 88.670000 ;
      LAYER met4 ;
        RECT 59.835000 88.350000 60.155000 88.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.835000 88.775000 60.155000 89.095000 ;
      LAYER met4 ;
        RECT 59.835000 88.775000 60.155000 89.095000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.835000 89.205000 60.155000 89.525000 ;
      LAYER met4 ;
        RECT 59.835000 89.205000 60.155000 89.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.835000 89.635000 60.155000 89.955000 ;
      LAYER met4 ;
        RECT 59.835000 89.635000 60.155000 89.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.835000 90.065000 60.155000 90.385000 ;
      LAYER met4 ;
        RECT 59.835000 90.065000 60.155000 90.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.835000 90.495000 60.155000 90.815000 ;
      LAYER met4 ;
        RECT 59.835000 90.495000 60.155000 90.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.895000 90.955000 60.215000 91.275000 ;
      LAYER met4 ;
        RECT 59.895000 90.955000 60.215000 91.275000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.895000 91.385000 60.215000 91.705000 ;
      LAYER met4 ;
        RECT 59.895000 91.385000 60.215000 91.705000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 82.795000 6.325000 83.115000 ;
      LAYER met4 ;
        RECT 6.005000 82.795000 6.325000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 83.205000 6.325000 83.525000 ;
      LAYER met4 ;
        RECT 6.005000 83.205000 6.325000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 83.615000 6.325000 83.935000 ;
      LAYER met4 ;
        RECT 6.005000 83.615000 6.325000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 84.025000 6.325000 84.345000 ;
      LAYER met4 ;
        RECT 6.005000 84.025000 6.325000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 84.435000 6.325000 84.755000 ;
      LAYER met4 ;
        RECT 6.005000 84.435000 6.325000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 84.845000 6.325000 85.165000 ;
      LAYER met4 ;
        RECT 6.005000 84.845000 6.325000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 85.255000 6.325000 85.575000 ;
      LAYER met4 ;
        RECT 6.005000 85.255000 6.325000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 85.665000 6.325000 85.985000 ;
      LAYER met4 ;
        RECT 6.005000 85.665000 6.325000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 86.075000 6.325000 86.395000 ;
      LAYER met4 ;
        RECT 6.005000 86.075000 6.325000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 86.485000 6.325000 86.805000 ;
      LAYER met4 ;
        RECT 6.005000 86.485000 6.325000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 86.895000 6.325000 87.215000 ;
      LAYER met4 ;
        RECT 6.005000 86.895000 6.325000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 87.305000 6.325000 87.625000 ;
      LAYER met4 ;
        RECT 6.005000 87.305000 6.325000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 87.715000 6.325000 88.035000 ;
      LAYER met4 ;
        RECT 6.005000 87.715000 6.325000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 88.125000 6.325000 88.445000 ;
      LAYER met4 ;
        RECT 6.005000 88.125000 6.325000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 88.535000 6.325000 88.855000 ;
      LAYER met4 ;
        RECT 6.005000 88.535000 6.325000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 88.945000 6.325000 89.265000 ;
      LAYER met4 ;
        RECT 6.005000 88.945000 6.325000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 89.355000 6.325000 89.675000 ;
      LAYER met4 ;
        RECT 6.005000 89.355000 6.325000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 89.765000 6.325000 90.085000 ;
      LAYER met4 ;
        RECT 6.005000 89.765000 6.325000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 90.175000 6.325000 90.495000 ;
      LAYER met4 ;
        RECT 6.005000 90.175000 6.325000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 90.585000 6.325000 90.905000 ;
      LAYER met4 ;
        RECT 6.005000 90.585000 6.325000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 90.995000 6.325000 91.315000 ;
      LAYER met4 ;
        RECT 6.005000 90.995000 6.325000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 91.405000 6.325000 91.725000 ;
      LAYER met4 ;
        RECT 6.005000 91.405000 6.325000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 91.815000 6.325000 92.135000 ;
      LAYER met4 ;
        RECT 6.005000 91.815000 6.325000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 92.225000 6.325000 92.545000 ;
      LAYER met4 ;
        RECT 6.005000 92.225000 6.325000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005000 92.635000 6.325000 92.955000 ;
      LAYER met4 ;
        RECT 6.005000 92.635000 6.325000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300000 17.800000 6.620000 18.120000 ;
      LAYER met4 ;
        RECT 6.300000 17.800000 6.620000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300000 18.230000 6.620000 18.550000 ;
      LAYER met4 ;
        RECT 6.300000 18.230000 6.620000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300000 18.660000 6.620000 18.980000 ;
      LAYER met4 ;
        RECT 6.300000 18.660000 6.620000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300000 19.090000 6.620000 19.410000 ;
      LAYER met4 ;
        RECT 6.300000 19.090000 6.620000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300000 19.520000 6.620000 19.840000 ;
      LAYER met4 ;
        RECT 6.300000 19.520000 6.620000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300000 19.950000 6.620000 20.270000 ;
      LAYER met4 ;
        RECT 6.300000 19.950000 6.620000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300000 20.380000 6.620000 20.700000 ;
      LAYER met4 ;
        RECT 6.300000 20.380000 6.620000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300000 20.810000 6.620000 21.130000 ;
      LAYER met4 ;
        RECT 6.300000 20.810000 6.620000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300000 21.240000 6.620000 21.560000 ;
      LAYER met4 ;
        RECT 6.300000 21.240000 6.620000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300000 21.670000 6.620000 21.990000 ;
      LAYER met4 ;
        RECT 6.300000 21.670000 6.620000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300000 22.100000 6.620000 22.420000 ;
      LAYER met4 ;
        RECT 6.300000 22.100000 6.620000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 68.065000 6.705000 68.385000 ;
      LAYER met4 ;
        RECT 6.385000 68.065000 6.705000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 68.475000 6.705000 68.795000 ;
      LAYER met4 ;
        RECT 6.385000 68.475000 6.705000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 68.885000 6.705000 69.205000 ;
      LAYER met4 ;
        RECT 6.385000 68.885000 6.705000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 69.295000 6.705000 69.615000 ;
      LAYER met4 ;
        RECT 6.385000 69.295000 6.705000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 69.705000 6.705000 70.025000 ;
      LAYER met4 ;
        RECT 6.385000 69.705000 6.705000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 70.115000 6.705000 70.435000 ;
      LAYER met4 ;
        RECT 6.385000 70.115000 6.705000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 70.525000 6.705000 70.845000 ;
      LAYER met4 ;
        RECT 6.385000 70.525000 6.705000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 70.935000 6.705000 71.255000 ;
      LAYER met4 ;
        RECT 6.385000 70.935000 6.705000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 71.345000 6.705000 71.665000 ;
      LAYER met4 ;
        RECT 6.385000 71.345000 6.705000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 71.755000 6.705000 72.075000 ;
      LAYER met4 ;
        RECT 6.385000 71.755000 6.705000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 72.165000 6.705000 72.485000 ;
      LAYER met4 ;
        RECT 6.385000 72.165000 6.705000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 72.575000 6.705000 72.895000 ;
      LAYER met4 ;
        RECT 6.385000 72.575000 6.705000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 72.985000 6.705000 73.305000 ;
      LAYER met4 ;
        RECT 6.385000 72.985000 6.705000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 73.390000 6.705000 73.710000 ;
      LAYER met4 ;
        RECT 6.385000 73.390000 6.705000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 73.795000 6.705000 74.115000 ;
      LAYER met4 ;
        RECT 6.385000 73.795000 6.705000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 74.200000 6.705000 74.520000 ;
      LAYER met4 ;
        RECT 6.385000 74.200000 6.705000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 74.605000 6.705000 74.925000 ;
      LAYER met4 ;
        RECT 6.385000 74.605000 6.705000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 75.010000 6.705000 75.330000 ;
      LAYER met4 ;
        RECT 6.385000 75.010000 6.705000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 75.415000 6.705000 75.735000 ;
      LAYER met4 ;
        RECT 6.385000 75.415000 6.705000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 75.820000 6.705000 76.140000 ;
      LAYER met4 ;
        RECT 6.385000 75.820000 6.705000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 76.225000 6.705000 76.545000 ;
      LAYER met4 ;
        RECT 6.385000 76.225000 6.705000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 76.630000 6.705000 76.950000 ;
      LAYER met4 ;
        RECT 6.385000 76.630000 6.705000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 77.035000 6.705000 77.355000 ;
      LAYER met4 ;
        RECT 6.385000 77.035000 6.705000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 77.440000 6.705000 77.760000 ;
      LAYER met4 ;
        RECT 6.385000 77.440000 6.705000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 77.845000 6.705000 78.165000 ;
      LAYER met4 ;
        RECT 6.385000 77.845000 6.705000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 78.250000 6.705000 78.570000 ;
      LAYER met4 ;
        RECT 6.385000 78.250000 6.705000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 78.655000 6.705000 78.975000 ;
      LAYER met4 ;
        RECT 6.385000 78.655000 6.705000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 79.060000 6.705000 79.380000 ;
      LAYER met4 ;
        RECT 6.385000 79.060000 6.705000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 79.465000 6.705000 79.785000 ;
      LAYER met4 ;
        RECT 6.385000 79.465000 6.705000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 79.870000 6.705000 80.190000 ;
      LAYER met4 ;
        RECT 6.385000 79.870000 6.705000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 80.275000 6.705000 80.595000 ;
      LAYER met4 ;
        RECT 6.385000 80.275000 6.705000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 80.680000 6.705000 81.000000 ;
      LAYER met4 ;
        RECT 6.385000 80.680000 6.705000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 81.085000 6.705000 81.405000 ;
      LAYER met4 ;
        RECT 6.385000 81.085000 6.705000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 81.490000 6.705000 81.810000 ;
      LAYER met4 ;
        RECT 6.385000 81.490000 6.705000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 81.895000 6.705000 82.215000 ;
      LAYER met4 ;
        RECT 6.385000 81.895000 6.705000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385000 82.300000 6.705000 82.620000 ;
      LAYER met4 ;
        RECT 6.385000 82.300000 6.705000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 82.795000 6.735000 83.115000 ;
      LAYER met4 ;
        RECT 6.415000 82.795000 6.735000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 83.205000 6.735000 83.525000 ;
      LAYER met4 ;
        RECT 6.415000 83.205000 6.735000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 83.615000 6.735000 83.935000 ;
      LAYER met4 ;
        RECT 6.415000 83.615000 6.735000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 84.025000 6.735000 84.345000 ;
      LAYER met4 ;
        RECT 6.415000 84.025000 6.735000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 84.435000 6.735000 84.755000 ;
      LAYER met4 ;
        RECT 6.415000 84.435000 6.735000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 84.845000 6.735000 85.165000 ;
      LAYER met4 ;
        RECT 6.415000 84.845000 6.735000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 85.255000 6.735000 85.575000 ;
      LAYER met4 ;
        RECT 6.415000 85.255000 6.735000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 85.665000 6.735000 85.985000 ;
      LAYER met4 ;
        RECT 6.415000 85.665000 6.735000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 86.075000 6.735000 86.395000 ;
      LAYER met4 ;
        RECT 6.415000 86.075000 6.735000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 86.485000 6.735000 86.805000 ;
      LAYER met4 ;
        RECT 6.415000 86.485000 6.735000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 86.895000 6.735000 87.215000 ;
      LAYER met4 ;
        RECT 6.415000 86.895000 6.735000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 87.305000 6.735000 87.625000 ;
      LAYER met4 ;
        RECT 6.415000 87.305000 6.735000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 87.715000 6.735000 88.035000 ;
      LAYER met4 ;
        RECT 6.415000 87.715000 6.735000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 88.125000 6.735000 88.445000 ;
      LAYER met4 ;
        RECT 6.415000 88.125000 6.735000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 88.535000 6.735000 88.855000 ;
      LAYER met4 ;
        RECT 6.415000 88.535000 6.735000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 88.945000 6.735000 89.265000 ;
      LAYER met4 ;
        RECT 6.415000 88.945000 6.735000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 89.355000 6.735000 89.675000 ;
      LAYER met4 ;
        RECT 6.415000 89.355000 6.735000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 89.765000 6.735000 90.085000 ;
      LAYER met4 ;
        RECT 6.415000 89.765000 6.735000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 90.175000 6.735000 90.495000 ;
      LAYER met4 ;
        RECT 6.415000 90.175000 6.735000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 90.585000 6.735000 90.905000 ;
      LAYER met4 ;
        RECT 6.415000 90.585000 6.735000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 90.995000 6.735000 91.315000 ;
      LAYER met4 ;
        RECT 6.415000 90.995000 6.735000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 91.405000 6.735000 91.725000 ;
      LAYER met4 ;
        RECT 6.415000 91.405000 6.735000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 91.815000 6.735000 92.135000 ;
      LAYER met4 ;
        RECT 6.415000 91.815000 6.735000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 92.225000 6.735000 92.545000 ;
      LAYER met4 ;
        RECT 6.415000 92.225000 6.735000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415000 92.635000 6.735000 92.955000 ;
      LAYER met4 ;
        RECT 6.415000 92.635000 6.735000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705000 17.800000 7.025000 18.120000 ;
      LAYER met4 ;
        RECT 6.705000 17.800000 7.025000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705000 18.230000 7.025000 18.550000 ;
      LAYER met4 ;
        RECT 6.705000 18.230000 7.025000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705000 18.660000 7.025000 18.980000 ;
      LAYER met4 ;
        RECT 6.705000 18.660000 7.025000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705000 19.090000 7.025000 19.410000 ;
      LAYER met4 ;
        RECT 6.705000 19.090000 7.025000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705000 19.520000 7.025000 19.840000 ;
      LAYER met4 ;
        RECT 6.705000 19.520000 7.025000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705000 19.950000 7.025000 20.270000 ;
      LAYER met4 ;
        RECT 6.705000 19.950000 7.025000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705000 20.380000 7.025000 20.700000 ;
      LAYER met4 ;
        RECT 6.705000 20.380000 7.025000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705000 20.810000 7.025000 21.130000 ;
      LAYER met4 ;
        RECT 6.705000 20.810000 7.025000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705000 21.240000 7.025000 21.560000 ;
      LAYER met4 ;
        RECT 6.705000 21.240000 7.025000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705000 21.670000 7.025000 21.990000 ;
      LAYER met4 ;
        RECT 6.705000 21.670000 7.025000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705000 22.100000 7.025000 22.420000 ;
      LAYER met4 ;
        RECT 6.705000 22.100000 7.025000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 68.065000 7.105000 68.385000 ;
      LAYER met4 ;
        RECT 6.785000 68.065000 7.105000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 68.475000 7.105000 68.795000 ;
      LAYER met4 ;
        RECT 6.785000 68.475000 7.105000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 68.885000 7.105000 69.205000 ;
      LAYER met4 ;
        RECT 6.785000 68.885000 7.105000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 69.295000 7.105000 69.615000 ;
      LAYER met4 ;
        RECT 6.785000 69.295000 7.105000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 69.705000 7.105000 70.025000 ;
      LAYER met4 ;
        RECT 6.785000 69.705000 7.105000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 70.115000 7.105000 70.435000 ;
      LAYER met4 ;
        RECT 6.785000 70.115000 7.105000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 70.525000 7.105000 70.845000 ;
      LAYER met4 ;
        RECT 6.785000 70.525000 7.105000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 70.935000 7.105000 71.255000 ;
      LAYER met4 ;
        RECT 6.785000 70.935000 7.105000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 71.345000 7.105000 71.665000 ;
      LAYER met4 ;
        RECT 6.785000 71.345000 7.105000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 71.755000 7.105000 72.075000 ;
      LAYER met4 ;
        RECT 6.785000 71.755000 7.105000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 72.165000 7.105000 72.485000 ;
      LAYER met4 ;
        RECT 6.785000 72.165000 7.105000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 72.575000 7.105000 72.895000 ;
      LAYER met4 ;
        RECT 6.785000 72.575000 7.105000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 72.985000 7.105000 73.305000 ;
      LAYER met4 ;
        RECT 6.785000 72.985000 7.105000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 73.390000 7.105000 73.710000 ;
      LAYER met4 ;
        RECT 6.785000 73.390000 7.105000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 73.795000 7.105000 74.115000 ;
      LAYER met4 ;
        RECT 6.785000 73.795000 7.105000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 74.200000 7.105000 74.520000 ;
      LAYER met4 ;
        RECT 6.785000 74.200000 7.105000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 74.605000 7.105000 74.925000 ;
      LAYER met4 ;
        RECT 6.785000 74.605000 7.105000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 75.010000 7.105000 75.330000 ;
      LAYER met4 ;
        RECT 6.785000 75.010000 7.105000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 75.415000 7.105000 75.735000 ;
      LAYER met4 ;
        RECT 6.785000 75.415000 7.105000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 75.820000 7.105000 76.140000 ;
      LAYER met4 ;
        RECT 6.785000 75.820000 7.105000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 76.225000 7.105000 76.545000 ;
      LAYER met4 ;
        RECT 6.785000 76.225000 7.105000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 76.630000 7.105000 76.950000 ;
      LAYER met4 ;
        RECT 6.785000 76.630000 7.105000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 77.035000 7.105000 77.355000 ;
      LAYER met4 ;
        RECT 6.785000 77.035000 7.105000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 77.440000 7.105000 77.760000 ;
      LAYER met4 ;
        RECT 6.785000 77.440000 7.105000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 77.845000 7.105000 78.165000 ;
      LAYER met4 ;
        RECT 6.785000 77.845000 7.105000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 78.250000 7.105000 78.570000 ;
      LAYER met4 ;
        RECT 6.785000 78.250000 7.105000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 78.655000 7.105000 78.975000 ;
      LAYER met4 ;
        RECT 6.785000 78.655000 7.105000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 79.060000 7.105000 79.380000 ;
      LAYER met4 ;
        RECT 6.785000 79.060000 7.105000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 79.465000 7.105000 79.785000 ;
      LAYER met4 ;
        RECT 6.785000 79.465000 7.105000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 79.870000 7.105000 80.190000 ;
      LAYER met4 ;
        RECT 6.785000 79.870000 7.105000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 80.275000 7.105000 80.595000 ;
      LAYER met4 ;
        RECT 6.785000 80.275000 7.105000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 80.680000 7.105000 81.000000 ;
      LAYER met4 ;
        RECT 6.785000 80.680000 7.105000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 81.085000 7.105000 81.405000 ;
      LAYER met4 ;
        RECT 6.785000 81.085000 7.105000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 81.490000 7.105000 81.810000 ;
      LAYER met4 ;
        RECT 6.785000 81.490000 7.105000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 81.895000 7.105000 82.215000 ;
      LAYER met4 ;
        RECT 6.785000 81.895000 7.105000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785000 82.300000 7.105000 82.620000 ;
      LAYER met4 ;
        RECT 6.785000 82.300000 7.105000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 82.795000 7.145000 83.115000 ;
      LAYER met4 ;
        RECT 6.825000 82.795000 7.145000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 83.205000 7.145000 83.525000 ;
      LAYER met4 ;
        RECT 6.825000 83.205000 7.145000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 83.615000 7.145000 83.935000 ;
      LAYER met4 ;
        RECT 6.825000 83.615000 7.145000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 84.025000 7.145000 84.345000 ;
      LAYER met4 ;
        RECT 6.825000 84.025000 7.145000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 84.435000 7.145000 84.755000 ;
      LAYER met4 ;
        RECT 6.825000 84.435000 7.145000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 84.845000 7.145000 85.165000 ;
      LAYER met4 ;
        RECT 6.825000 84.845000 7.145000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 85.255000 7.145000 85.575000 ;
      LAYER met4 ;
        RECT 6.825000 85.255000 7.145000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 85.665000 7.145000 85.985000 ;
      LAYER met4 ;
        RECT 6.825000 85.665000 7.145000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 86.075000 7.145000 86.395000 ;
      LAYER met4 ;
        RECT 6.825000 86.075000 7.145000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 86.485000 7.145000 86.805000 ;
      LAYER met4 ;
        RECT 6.825000 86.485000 7.145000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 86.895000 7.145000 87.215000 ;
      LAYER met4 ;
        RECT 6.825000 86.895000 7.145000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 87.305000 7.145000 87.625000 ;
      LAYER met4 ;
        RECT 6.825000 87.305000 7.145000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 87.715000 7.145000 88.035000 ;
      LAYER met4 ;
        RECT 6.825000 87.715000 7.145000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 88.125000 7.145000 88.445000 ;
      LAYER met4 ;
        RECT 6.825000 88.125000 7.145000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 88.535000 7.145000 88.855000 ;
      LAYER met4 ;
        RECT 6.825000 88.535000 7.145000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 88.945000 7.145000 89.265000 ;
      LAYER met4 ;
        RECT 6.825000 88.945000 7.145000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 89.355000 7.145000 89.675000 ;
      LAYER met4 ;
        RECT 6.825000 89.355000 7.145000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 89.765000 7.145000 90.085000 ;
      LAYER met4 ;
        RECT 6.825000 89.765000 7.145000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 90.175000 7.145000 90.495000 ;
      LAYER met4 ;
        RECT 6.825000 90.175000 7.145000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 90.585000 7.145000 90.905000 ;
      LAYER met4 ;
        RECT 6.825000 90.585000 7.145000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 90.995000 7.145000 91.315000 ;
      LAYER met4 ;
        RECT 6.825000 90.995000 7.145000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 91.405000 7.145000 91.725000 ;
      LAYER met4 ;
        RECT 6.825000 91.405000 7.145000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 91.815000 7.145000 92.135000 ;
      LAYER met4 ;
        RECT 6.825000 91.815000 7.145000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 92.225000 7.145000 92.545000 ;
      LAYER met4 ;
        RECT 6.825000 92.225000 7.145000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825000 92.635000 7.145000 92.955000 ;
      LAYER met4 ;
        RECT 6.825000 92.635000 7.145000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.100000 17.800000 60.420000 18.120000 ;
      LAYER met4 ;
        RECT 60.100000 17.800000 60.420000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.100000 18.230000 60.420000 18.550000 ;
      LAYER met4 ;
        RECT 60.100000 18.230000 60.420000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.100000 18.660000 60.420000 18.980000 ;
      LAYER met4 ;
        RECT 60.100000 18.660000 60.420000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.100000 19.090000 60.420000 19.410000 ;
      LAYER met4 ;
        RECT 60.100000 19.090000 60.420000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.100000 19.520000 60.420000 19.840000 ;
      LAYER met4 ;
        RECT 60.100000 19.520000 60.420000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.100000 19.950000 60.420000 20.270000 ;
      LAYER met4 ;
        RECT 60.100000 19.950000 60.420000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.100000 20.380000 60.420000 20.700000 ;
      LAYER met4 ;
        RECT 60.100000 20.380000 60.420000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.100000 20.810000 60.420000 21.130000 ;
      LAYER met4 ;
        RECT 60.100000 20.810000 60.420000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.100000 21.240000 60.420000 21.560000 ;
      LAYER met4 ;
        RECT 60.100000 21.240000 60.420000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.100000 21.670000 60.420000 21.990000 ;
      LAYER met4 ;
        RECT 60.100000 21.670000 60.420000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.100000 22.100000 60.420000 22.420000 ;
      LAYER met4 ;
        RECT 60.100000 22.100000 60.420000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120000 82.995000 60.440000 83.315000 ;
      LAYER met4 ;
        RECT 60.120000 82.995000 60.440000 83.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120000 83.395000 60.440000 83.715000 ;
      LAYER met4 ;
        RECT 60.120000 83.395000 60.440000 83.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120000 83.795000 60.440000 84.115000 ;
      LAYER met4 ;
        RECT 60.120000 83.795000 60.440000 84.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120000 84.195000 60.440000 84.515000 ;
      LAYER met4 ;
        RECT 60.120000 84.195000 60.440000 84.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120000 84.595000 60.440000 84.915000 ;
      LAYER met4 ;
        RECT 60.120000 84.595000 60.440000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120000 84.995000 60.440000 85.315000 ;
      LAYER met4 ;
        RECT 60.120000 84.995000 60.440000 85.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120000 85.395000 60.440000 85.715000 ;
      LAYER met4 ;
        RECT 60.120000 85.395000 60.440000 85.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120000 85.795000 60.440000 86.115000 ;
      LAYER met4 ;
        RECT 60.120000 85.795000 60.440000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120000 86.195000 60.440000 86.515000 ;
      LAYER met4 ;
        RECT 60.120000 86.195000 60.440000 86.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120000 86.600000 60.440000 86.920000 ;
      LAYER met4 ;
        RECT 60.120000 86.600000 60.440000 86.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120000 87.005000 60.440000 87.325000 ;
      LAYER met4 ;
        RECT 60.120000 87.005000 60.440000 87.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120000 87.410000 60.440000 87.730000 ;
      LAYER met4 ;
        RECT 60.120000 87.410000 60.440000 87.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120000 87.815000 60.440000 88.135000 ;
      LAYER met4 ;
        RECT 60.120000 87.815000 60.440000 88.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 68.065000 60.470000 68.385000 ;
      LAYER met4 ;
        RECT 60.150000 68.065000 60.470000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 68.475000 60.470000 68.795000 ;
      LAYER met4 ;
        RECT 60.150000 68.475000 60.470000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 68.885000 60.470000 69.205000 ;
      LAYER met4 ;
        RECT 60.150000 68.885000 60.470000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 69.295000 60.470000 69.615000 ;
      LAYER met4 ;
        RECT 60.150000 69.295000 60.470000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 69.705000 60.470000 70.025000 ;
      LAYER met4 ;
        RECT 60.150000 69.705000 60.470000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 70.115000 60.470000 70.435000 ;
      LAYER met4 ;
        RECT 60.150000 70.115000 60.470000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 70.525000 60.470000 70.845000 ;
      LAYER met4 ;
        RECT 60.150000 70.525000 60.470000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 70.935000 60.470000 71.255000 ;
      LAYER met4 ;
        RECT 60.150000 70.935000 60.470000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 71.345000 60.470000 71.665000 ;
      LAYER met4 ;
        RECT 60.150000 71.345000 60.470000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 71.755000 60.470000 72.075000 ;
      LAYER met4 ;
        RECT 60.150000 71.755000 60.470000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 72.165000 60.470000 72.485000 ;
      LAYER met4 ;
        RECT 60.150000 72.165000 60.470000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 72.575000 60.470000 72.895000 ;
      LAYER met4 ;
        RECT 60.150000 72.575000 60.470000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 72.985000 60.470000 73.305000 ;
      LAYER met4 ;
        RECT 60.150000 72.985000 60.470000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 73.390000 60.470000 73.710000 ;
      LAYER met4 ;
        RECT 60.150000 73.390000 60.470000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 73.795000 60.470000 74.115000 ;
      LAYER met4 ;
        RECT 60.150000 73.795000 60.470000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 74.200000 60.470000 74.520000 ;
      LAYER met4 ;
        RECT 60.150000 74.200000 60.470000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 74.605000 60.470000 74.925000 ;
      LAYER met4 ;
        RECT 60.150000 74.605000 60.470000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 75.010000 60.470000 75.330000 ;
      LAYER met4 ;
        RECT 60.150000 75.010000 60.470000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 75.415000 60.470000 75.735000 ;
      LAYER met4 ;
        RECT 60.150000 75.415000 60.470000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 75.820000 60.470000 76.140000 ;
      LAYER met4 ;
        RECT 60.150000 75.820000 60.470000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 76.225000 60.470000 76.545000 ;
      LAYER met4 ;
        RECT 60.150000 76.225000 60.470000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 76.630000 60.470000 76.950000 ;
      LAYER met4 ;
        RECT 60.150000 76.630000 60.470000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 77.035000 60.470000 77.355000 ;
      LAYER met4 ;
        RECT 60.150000 77.035000 60.470000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 77.440000 60.470000 77.760000 ;
      LAYER met4 ;
        RECT 60.150000 77.440000 60.470000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 77.845000 60.470000 78.165000 ;
      LAYER met4 ;
        RECT 60.150000 77.845000 60.470000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 78.250000 60.470000 78.570000 ;
      LAYER met4 ;
        RECT 60.150000 78.250000 60.470000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 78.655000 60.470000 78.975000 ;
      LAYER met4 ;
        RECT 60.150000 78.655000 60.470000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 79.060000 60.470000 79.380000 ;
      LAYER met4 ;
        RECT 60.150000 79.060000 60.470000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 79.465000 60.470000 79.785000 ;
      LAYER met4 ;
        RECT 60.150000 79.465000 60.470000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 79.870000 60.470000 80.190000 ;
      LAYER met4 ;
        RECT 60.150000 79.870000 60.470000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 80.275000 60.470000 80.595000 ;
      LAYER met4 ;
        RECT 60.150000 80.275000 60.470000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 80.680000 60.470000 81.000000 ;
      LAYER met4 ;
        RECT 60.150000 80.680000 60.470000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 81.085000 60.470000 81.405000 ;
      LAYER met4 ;
        RECT 60.150000 81.085000 60.470000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 81.490000 60.470000 81.810000 ;
      LAYER met4 ;
        RECT 60.150000 81.490000 60.470000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 81.895000 60.470000 82.215000 ;
      LAYER met4 ;
        RECT 60.150000 81.895000 60.470000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.150000 82.300000 60.470000 82.620000 ;
      LAYER met4 ;
        RECT 60.150000 82.300000 60.470000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.245000 88.350000 60.565000 88.670000 ;
      LAYER met4 ;
        RECT 60.245000 88.350000 60.565000 88.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.245000 88.775000 60.565000 89.095000 ;
      LAYER met4 ;
        RECT 60.245000 88.775000 60.565000 89.095000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.245000 89.205000 60.565000 89.525000 ;
      LAYER met4 ;
        RECT 60.245000 89.205000 60.565000 89.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.245000 89.635000 60.565000 89.955000 ;
      LAYER met4 ;
        RECT 60.245000 89.635000 60.565000 89.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.245000 90.065000 60.565000 90.385000 ;
      LAYER met4 ;
        RECT 60.245000 90.065000 60.565000 90.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.245000 90.495000 60.565000 90.815000 ;
      LAYER met4 ;
        RECT 60.245000 90.495000 60.565000 90.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 17.800000 60.825000 18.120000 ;
      LAYER met4 ;
        RECT 60.505000 17.800000 60.825000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 18.230000 60.825000 18.550000 ;
      LAYER met4 ;
        RECT 60.505000 18.230000 60.825000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 18.660000 60.825000 18.980000 ;
      LAYER met4 ;
        RECT 60.505000 18.660000 60.825000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 19.090000 60.825000 19.410000 ;
      LAYER met4 ;
        RECT 60.505000 19.090000 60.825000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 19.520000 60.825000 19.840000 ;
      LAYER met4 ;
        RECT 60.505000 19.520000 60.825000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 19.950000 60.825000 20.270000 ;
      LAYER met4 ;
        RECT 60.505000 19.950000 60.825000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 20.380000 60.825000 20.700000 ;
      LAYER met4 ;
        RECT 60.505000 20.380000 60.825000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 20.810000 60.825000 21.130000 ;
      LAYER met4 ;
        RECT 60.505000 20.810000 60.825000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 21.240000 60.825000 21.560000 ;
      LAYER met4 ;
        RECT 60.505000 21.240000 60.825000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 21.670000 60.825000 21.990000 ;
      LAYER met4 ;
        RECT 60.505000 21.670000 60.825000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 22.100000 60.825000 22.420000 ;
      LAYER met4 ;
        RECT 60.505000 22.100000 60.825000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530000 82.995000 60.850000 83.315000 ;
      LAYER met4 ;
        RECT 60.530000 82.995000 60.850000 83.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530000 83.395000 60.850000 83.715000 ;
      LAYER met4 ;
        RECT 60.530000 83.395000 60.850000 83.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530000 83.795000 60.850000 84.115000 ;
      LAYER met4 ;
        RECT 60.530000 83.795000 60.850000 84.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530000 84.195000 60.850000 84.515000 ;
      LAYER met4 ;
        RECT 60.530000 84.195000 60.850000 84.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530000 84.595000 60.850000 84.915000 ;
      LAYER met4 ;
        RECT 60.530000 84.595000 60.850000 84.915000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530000 84.995000 60.850000 85.315000 ;
      LAYER met4 ;
        RECT 60.530000 84.995000 60.850000 85.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530000 85.395000 60.850000 85.715000 ;
      LAYER met4 ;
        RECT 60.530000 85.395000 60.850000 85.715000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530000 85.795000 60.850000 86.115000 ;
      LAYER met4 ;
        RECT 60.530000 85.795000 60.850000 86.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530000 86.195000 60.850000 86.515000 ;
      LAYER met4 ;
        RECT 60.530000 86.195000 60.850000 86.515000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530000 86.600000 60.850000 86.920000 ;
      LAYER met4 ;
        RECT 60.530000 86.600000 60.850000 86.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530000 87.005000 60.850000 87.325000 ;
      LAYER met4 ;
        RECT 60.530000 87.005000 60.850000 87.325000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530000 87.410000 60.850000 87.730000 ;
      LAYER met4 ;
        RECT 60.530000 87.410000 60.850000 87.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530000 87.815000 60.850000 88.135000 ;
      LAYER met4 ;
        RECT 60.530000 87.815000 60.850000 88.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 68.065000 60.870000 68.385000 ;
      LAYER met4 ;
        RECT 60.550000 68.065000 60.870000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 68.475000 60.870000 68.795000 ;
      LAYER met4 ;
        RECT 60.550000 68.475000 60.870000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 68.885000 60.870000 69.205000 ;
      LAYER met4 ;
        RECT 60.550000 68.885000 60.870000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 69.295000 60.870000 69.615000 ;
      LAYER met4 ;
        RECT 60.550000 69.295000 60.870000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 69.705000 60.870000 70.025000 ;
      LAYER met4 ;
        RECT 60.550000 69.705000 60.870000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 70.115000 60.870000 70.435000 ;
      LAYER met4 ;
        RECT 60.550000 70.115000 60.870000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 70.525000 60.870000 70.845000 ;
      LAYER met4 ;
        RECT 60.550000 70.525000 60.870000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 70.935000 60.870000 71.255000 ;
      LAYER met4 ;
        RECT 60.550000 70.935000 60.870000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 71.345000 60.870000 71.665000 ;
      LAYER met4 ;
        RECT 60.550000 71.345000 60.870000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 71.755000 60.870000 72.075000 ;
      LAYER met4 ;
        RECT 60.550000 71.755000 60.870000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 72.165000 60.870000 72.485000 ;
      LAYER met4 ;
        RECT 60.550000 72.165000 60.870000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 72.575000 60.870000 72.895000 ;
      LAYER met4 ;
        RECT 60.550000 72.575000 60.870000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 72.985000 60.870000 73.305000 ;
      LAYER met4 ;
        RECT 60.550000 72.985000 60.870000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 73.390000 60.870000 73.710000 ;
      LAYER met4 ;
        RECT 60.550000 73.390000 60.870000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 73.795000 60.870000 74.115000 ;
      LAYER met4 ;
        RECT 60.550000 73.795000 60.870000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 74.200000 60.870000 74.520000 ;
      LAYER met4 ;
        RECT 60.550000 74.200000 60.870000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 74.605000 60.870000 74.925000 ;
      LAYER met4 ;
        RECT 60.550000 74.605000 60.870000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 75.010000 60.870000 75.330000 ;
      LAYER met4 ;
        RECT 60.550000 75.010000 60.870000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 75.415000 60.870000 75.735000 ;
      LAYER met4 ;
        RECT 60.550000 75.415000 60.870000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 75.820000 60.870000 76.140000 ;
      LAYER met4 ;
        RECT 60.550000 75.820000 60.870000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 76.225000 60.870000 76.545000 ;
      LAYER met4 ;
        RECT 60.550000 76.225000 60.870000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 76.630000 60.870000 76.950000 ;
      LAYER met4 ;
        RECT 60.550000 76.630000 60.870000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 77.035000 60.870000 77.355000 ;
      LAYER met4 ;
        RECT 60.550000 77.035000 60.870000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 77.440000 60.870000 77.760000 ;
      LAYER met4 ;
        RECT 60.550000 77.440000 60.870000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 77.845000 60.870000 78.165000 ;
      LAYER met4 ;
        RECT 60.550000 77.845000 60.870000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 78.250000 60.870000 78.570000 ;
      LAYER met4 ;
        RECT 60.550000 78.250000 60.870000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 78.655000 60.870000 78.975000 ;
      LAYER met4 ;
        RECT 60.550000 78.655000 60.870000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 79.060000 60.870000 79.380000 ;
      LAYER met4 ;
        RECT 60.550000 79.060000 60.870000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 79.465000 60.870000 79.785000 ;
      LAYER met4 ;
        RECT 60.550000 79.465000 60.870000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 79.870000 60.870000 80.190000 ;
      LAYER met4 ;
        RECT 60.550000 79.870000 60.870000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 80.275000 60.870000 80.595000 ;
      LAYER met4 ;
        RECT 60.550000 80.275000 60.870000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 80.680000 60.870000 81.000000 ;
      LAYER met4 ;
        RECT 60.550000 80.680000 60.870000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 81.085000 60.870000 81.405000 ;
      LAYER met4 ;
        RECT 60.550000 81.085000 60.870000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 81.490000 60.870000 81.810000 ;
      LAYER met4 ;
        RECT 60.550000 81.490000 60.870000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 81.895000 60.870000 82.215000 ;
      LAYER met4 ;
        RECT 60.550000 81.895000 60.870000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550000 82.300000 60.870000 82.620000 ;
      LAYER met4 ;
        RECT 60.550000 82.300000 60.870000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.655000 88.350000 60.975000 88.670000 ;
      LAYER met4 ;
        RECT 60.655000 88.350000 60.975000 88.670000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.655000 88.775000 60.975000 89.095000 ;
      LAYER met4 ;
        RECT 60.655000 88.775000 60.975000 89.095000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.655000 89.205000 60.975000 89.525000 ;
      LAYER met4 ;
        RECT 60.655000 89.205000 60.975000 89.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.655000 89.635000 60.975000 89.955000 ;
      LAYER met4 ;
        RECT 60.655000 89.635000 60.975000 89.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.655000 90.065000 60.975000 90.385000 ;
      LAYER met4 ;
        RECT 60.655000 90.065000 60.975000 90.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.655000 90.495000 60.975000 90.815000 ;
      LAYER met4 ;
        RECT 60.655000 90.495000 60.975000 90.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.675000 90.955000 60.995000 91.275000 ;
      LAYER met4 ;
        RECT 60.675000 90.955000 60.995000 91.275000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.675000 91.385000 60.995000 91.705000 ;
      LAYER met4 ;
        RECT 60.675000 91.385000 60.995000 91.705000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.910000 17.800000 61.230000 18.120000 ;
      LAYER met4 ;
        RECT 60.910000 17.800000 61.230000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.910000 18.230000 61.230000 18.550000 ;
      LAYER met4 ;
        RECT 60.910000 18.230000 61.230000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.910000 18.660000 61.230000 18.980000 ;
      LAYER met4 ;
        RECT 60.910000 18.660000 61.230000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.910000 19.090000 61.230000 19.410000 ;
      LAYER met4 ;
        RECT 60.910000 19.090000 61.230000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.910000 19.520000 61.230000 19.840000 ;
      LAYER met4 ;
        RECT 60.910000 19.520000 61.230000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.910000 19.950000 61.230000 20.270000 ;
      LAYER met4 ;
        RECT 60.910000 19.950000 61.230000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.910000 20.380000 61.230000 20.700000 ;
      LAYER met4 ;
        RECT 60.910000 20.380000 61.230000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.910000 20.810000 61.230000 21.130000 ;
      LAYER met4 ;
        RECT 60.910000 20.810000 61.230000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.910000 21.240000 61.230000 21.560000 ;
      LAYER met4 ;
        RECT 60.910000 21.240000 61.230000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.910000 21.670000 61.230000 21.990000 ;
      LAYER met4 ;
        RECT 60.910000 21.670000 61.230000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.910000 22.100000 61.230000 22.420000 ;
      LAYER met4 ;
        RECT 60.910000 22.100000 61.230000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 68.065000 61.270000 68.385000 ;
      LAYER met4 ;
        RECT 60.950000 68.065000 61.270000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 68.475000 61.270000 68.795000 ;
      LAYER met4 ;
        RECT 60.950000 68.475000 61.270000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 68.885000 61.270000 69.205000 ;
      LAYER met4 ;
        RECT 60.950000 68.885000 61.270000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 69.295000 61.270000 69.615000 ;
      LAYER met4 ;
        RECT 60.950000 69.295000 61.270000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 69.705000 61.270000 70.025000 ;
      LAYER met4 ;
        RECT 60.950000 69.705000 61.270000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 70.115000 61.270000 70.435000 ;
      LAYER met4 ;
        RECT 60.950000 70.115000 61.270000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 70.525000 61.270000 70.845000 ;
      LAYER met4 ;
        RECT 60.950000 70.525000 61.270000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 70.935000 61.270000 71.255000 ;
      LAYER met4 ;
        RECT 60.950000 70.935000 61.270000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 71.345000 61.270000 71.665000 ;
      LAYER met4 ;
        RECT 60.950000 71.345000 61.270000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 71.755000 61.270000 72.075000 ;
      LAYER met4 ;
        RECT 60.950000 71.755000 61.270000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 72.165000 61.270000 72.485000 ;
      LAYER met4 ;
        RECT 60.950000 72.165000 61.270000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 72.575000 61.270000 72.895000 ;
      LAYER met4 ;
        RECT 60.950000 72.575000 61.270000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 72.985000 61.270000 73.305000 ;
      LAYER met4 ;
        RECT 60.950000 72.985000 61.270000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 73.390000 61.270000 73.710000 ;
      LAYER met4 ;
        RECT 60.950000 73.390000 61.270000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 73.795000 61.270000 74.115000 ;
      LAYER met4 ;
        RECT 60.950000 73.795000 61.270000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 74.200000 61.270000 74.520000 ;
      LAYER met4 ;
        RECT 60.950000 74.200000 61.270000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 74.605000 61.270000 74.925000 ;
      LAYER met4 ;
        RECT 60.950000 74.605000 61.270000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 75.010000 61.270000 75.330000 ;
      LAYER met4 ;
        RECT 60.950000 75.010000 61.270000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 75.415000 61.270000 75.735000 ;
      LAYER met4 ;
        RECT 60.950000 75.415000 61.270000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 75.820000 61.270000 76.140000 ;
      LAYER met4 ;
        RECT 60.950000 75.820000 61.270000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 76.225000 61.270000 76.545000 ;
      LAYER met4 ;
        RECT 60.950000 76.225000 61.270000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 76.630000 61.270000 76.950000 ;
      LAYER met4 ;
        RECT 60.950000 76.630000 61.270000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 77.035000 61.270000 77.355000 ;
      LAYER met4 ;
        RECT 60.950000 77.035000 61.270000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 77.440000 61.270000 77.760000 ;
      LAYER met4 ;
        RECT 60.950000 77.440000 61.270000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 77.845000 61.270000 78.165000 ;
      LAYER met4 ;
        RECT 60.950000 77.845000 61.270000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 78.250000 61.270000 78.570000 ;
      LAYER met4 ;
        RECT 60.950000 78.250000 61.270000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 78.655000 61.270000 78.975000 ;
      LAYER met4 ;
        RECT 60.950000 78.655000 61.270000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 79.060000 61.270000 79.380000 ;
      LAYER met4 ;
        RECT 60.950000 79.060000 61.270000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 79.465000 61.270000 79.785000 ;
      LAYER met4 ;
        RECT 60.950000 79.465000 61.270000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 79.870000 61.270000 80.190000 ;
      LAYER met4 ;
        RECT 60.950000 79.870000 61.270000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 80.275000 61.270000 80.595000 ;
      LAYER met4 ;
        RECT 60.950000 80.275000 61.270000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 80.680000 61.270000 81.000000 ;
      LAYER met4 ;
        RECT 60.950000 80.680000 61.270000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 81.085000 61.270000 81.405000 ;
      LAYER met4 ;
        RECT 60.950000 81.085000 61.270000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 81.490000 61.270000 81.810000 ;
      LAYER met4 ;
        RECT 60.950000 81.490000 61.270000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 81.895000 61.270000 82.215000 ;
      LAYER met4 ;
        RECT 60.950000 81.895000 61.270000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 82.300000 61.270000 82.620000 ;
      LAYER met4 ;
        RECT 60.950000 82.300000 61.270000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 82.795000 61.475000 83.115000 ;
      LAYER met4 ;
        RECT 61.155000 82.795000 61.475000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 83.205000 61.475000 83.525000 ;
      LAYER met4 ;
        RECT 61.155000 83.205000 61.475000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 83.615000 61.475000 83.935000 ;
      LAYER met4 ;
        RECT 61.155000 83.615000 61.475000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 84.025000 61.475000 84.345000 ;
      LAYER met4 ;
        RECT 61.155000 84.025000 61.475000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 84.435000 61.475000 84.755000 ;
      LAYER met4 ;
        RECT 61.155000 84.435000 61.475000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 84.845000 61.475000 85.165000 ;
      LAYER met4 ;
        RECT 61.155000 84.845000 61.475000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 85.255000 61.475000 85.575000 ;
      LAYER met4 ;
        RECT 61.155000 85.255000 61.475000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 85.665000 61.475000 85.985000 ;
      LAYER met4 ;
        RECT 61.155000 85.665000 61.475000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 86.075000 61.475000 86.395000 ;
      LAYER met4 ;
        RECT 61.155000 86.075000 61.475000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 86.485000 61.475000 86.805000 ;
      LAYER met4 ;
        RECT 61.155000 86.485000 61.475000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 86.895000 61.475000 87.215000 ;
      LAYER met4 ;
        RECT 61.155000 86.895000 61.475000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 87.305000 61.475000 87.625000 ;
      LAYER met4 ;
        RECT 61.155000 87.305000 61.475000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 87.715000 61.475000 88.035000 ;
      LAYER met4 ;
        RECT 61.155000 87.715000 61.475000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 88.125000 61.475000 88.445000 ;
      LAYER met4 ;
        RECT 61.155000 88.125000 61.475000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 88.535000 61.475000 88.855000 ;
      LAYER met4 ;
        RECT 61.155000 88.535000 61.475000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 88.945000 61.475000 89.265000 ;
      LAYER met4 ;
        RECT 61.155000 88.945000 61.475000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 89.355000 61.475000 89.675000 ;
      LAYER met4 ;
        RECT 61.155000 89.355000 61.475000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 89.765000 61.475000 90.085000 ;
      LAYER met4 ;
        RECT 61.155000 89.765000 61.475000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 90.175000 61.475000 90.495000 ;
      LAYER met4 ;
        RECT 61.155000 90.175000 61.475000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 90.585000 61.475000 90.905000 ;
      LAYER met4 ;
        RECT 61.155000 90.585000 61.475000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 90.995000 61.475000 91.315000 ;
      LAYER met4 ;
        RECT 61.155000 90.995000 61.475000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 91.405000 61.475000 91.725000 ;
      LAYER met4 ;
        RECT 61.155000 91.405000 61.475000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 91.815000 61.475000 92.135000 ;
      LAYER met4 ;
        RECT 61.155000 91.815000 61.475000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 92.225000 61.475000 92.545000 ;
      LAYER met4 ;
        RECT 61.155000 92.225000 61.475000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155000 92.635000 61.475000 92.955000 ;
      LAYER met4 ;
        RECT 61.155000 92.635000 61.475000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.315000 17.800000 61.635000 18.120000 ;
      LAYER met4 ;
        RECT 61.315000 17.800000 61.635000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.315000 18.230000 61.635000 18.550000 ;
      LAYER met4 ;
        RECT 61.315000 18.230000 61.635000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.315000 18.660000 61.635000 18.980000 ;
      LAYER met4 ;
        RECT 61.315000 18.660000 61.635000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.315000 19.090000 61.635000 19.410000 ;
      LAYER met4 ;
        RECT 61.315000 19.090000 61.635000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.315000 19.520000 61.635000 19.840000 ;
      LAYER met4 ;
        RECT 61.315000 19.520000 61.635000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.315000 19.950000 61.635000 20.270000 ;
      LAYER met4 ;
        RECT 61.315000 19.950000 61.635000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.315000 20.380000 61.635000 20.700000 ;
      LAYER met4 ;
        RECT 61.315000 20.380000 61.635000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.315000 20.810000 61.635000 21.130000 ;
      LAYER met4 ;
        RECT 61.315000 20.810000 61.635000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.315000 21.240000 61.635000 21.560000 ;
      LAYER met4 ;
        RECT 61.315000 21.240000 61.635000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.315000 21.670000 61.635000 21.990000 ;
      LAYER met4 ;
        RECT 61.315000 21.670000 61.635000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.315000 22.100000 61.635000 22.420000 ;
      LAYER met4 ;
        RECT 61.315000 22.100000 61.635000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 68.065000 61.670000 68.385000 ;
      LAYER met4 ;
        RECT 61.350000 68.065000 61.670000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 68.475000 61.670000 68.795000 ;
      LAYER met4 ;
        RECT 61.350000 68.475000 61.670000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 68.885000 61.670000 69.205000 ;
      LAYER met4 ;
        RECT 61.350000 68.885000 61.670000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 69.295000 61.670000 69.615000 ;
      LAYER met4 ;
        RECT 61.350000 69.295000 61.670000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 69.705000 61.670000 70.025000 ;
      LAYER met4 ;
        RECT 61.350000 69.705000 61.670000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 70.115000 61.670000 70.435000 ;
      LAYER met4 ;
        RECT 61.350000 70.115000 61.670000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 70.525000 61.670000 70.845000 ;
      LAYER met4 ;
        RECT 61.350000 70.525000 61.670000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 70.935000 61.670000 71.255000 ;
      LAYER met4 ;
        RECT 61.350000 70.935000 61.670000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 71.345000 61.670000 71.665000 ;
      LAYER met4 ;
        RECT 61.350000 71.345000 61.670000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 71.755000 61.670000 72.075000 ;
      LAYER met4 ;
        RECT 61.350000 71.755000 61.670000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 72.165000 61.670000 72.485000 ;
      LAYER met4 ;
        RECT 61.350000 72.165000 61.670000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 72.575000 61.670000 72.895000 ;
      LAYER met4 ;
        RECT 61.350000 72.575000 61.670000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 72.985000 61.670000 73.305000 ;
      LAYER met4 ;
        RECT 61.350000 72.985000 61.670000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 73.390000 61.670000 73.710000 ;
      LAYER met4 ;
        RECT 61.350000 73.390000 61.670000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 73.795000 61.670000 74.115000 ;
      LAYER met4 ;
        RECT 61.350000 73.795000 61.670000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 74.200000 61.670000 74.520000 ;
      LAYER met4 ;
        RECT 61.350000 74.200000 61.670000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 74.605000 61.670000 74.925000 ;
      LAYER met4 ;
        RECT 61.350000 74.605000 61.670000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 75.010000 61.670000 75.330000 ;
      LAYER met4 ;
        RECT 61.350000 75.010000 61.670000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 75.415000 61.670000 75.735000 ;
      LAYER met4 ;
        RECT 61.350000 75.415000 61.670000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 75.820000 61.670000 76.140000 ;
      LAYER met4 ;
        RECT 61.350000 75.820000 61.670000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 76.225000 61.670000 76.545000 ;
      LAYER met4 ;
        RECT 61.350000 76.225000 61.670000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 76.630000 61.670000 76.950000 ;
      LAYER met4 ;
        RECT 61.350000 76.630000 61.670000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 77.035000 61.670000 77.355000 ;
      LAYER met4 ;
        RECT 61.350000 77.035000 61.670000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 77.440000 61.670000 77.760000 ;
      LAYER met4 ;
        RECT 61.350000 77.440000 61.670000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 77.845000 61.670000 78.165000 ;
      LAYER met4 ;
        RECT 61.350000 77.845000 61.670000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 78.250000 61.670000 78.570000 ;
      LAYER met4 ;
        RECT 61.350000 78.250000 61.670000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 78.655000 61.670000 78.975000 ;
      LAYER met4 ;
        RECT 61.350000 78.655000 61.670000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 79.060000 61.670000 79.380000 ;
      LAYER met4 ;
        RECT 61.350000 79.060000 61.670000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 79.465000 61.670000 79.785000 ;
      LAYER met4 ;
        RECT 61.350000 79.465000 61.670000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 79.870000 61.670000 80.190000 ;
      LAYER met4 ;
        RECT 61.350000 79.870000 61.670000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 80.275000 61.670000 80.595000 ;
      LAYER met4 ;
        RECT 61.350000 80.275000 61.670000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 80.680000 61.670000 81.000000 ;
      LAYER met4 ;
        RECT 61.350000 80.680000 61.670000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 81.085000 61.670000 81.405000 ;
      LAYER met4 ;
        RECT 61.350000 81.085000 61.670000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 81.490000 61.670000 81.810000 ;
      LAYER met4 ;
        RECT 61.350000 81.490000 61.670000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 81.895000 61.670000 82.215000 ;
      LAYER met4 ;
        RECT 61.350000 81.895000 61.670000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.350000 82.300000 61.670000 82.620000 ;
      LAYER met4 ;
        RECT 61.350000 82.300000 61.670000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 82.795000 61.880000 83.115000 ;
      LAYER met4 ;
        RECT 61.560000 82.795000 61.880000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 83.205000 61.880000 83.525000 ;
      LAYER met4 ;
        RECT 61.560000 83.205000 61.880000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 83.615000 61.880000 83.935000 ;
      LAYER met4 ;
        RECT 61.560000 83.615000 61.880000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 84.025000 61.880000 84.345000 ;
      LAYER met4 ;
        RECT 61.560000 84.025000 61.880000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 84.435000 61.880000 84.755000 ;
      LAYER met4 ;
        RECT 61.560000 84.435000 61.880000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 84.845000 61.880000 85.165000 ;
      LAYER met4 ;
        RECT 61.560000 84.845000 61.880000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 85.255000 61.880000 85.575000 ;
      LAYER met4 ;
        RECT 61.560000 85.255000 61.880000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 85.665000 61.880000 85.985000 ;
      LAYER met4 ;
        RECT 61.560000 85.665000 61.880000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 86.075000 61.880000 86.395000 ;
      LAYER met4 ;
        RECT 61.560000 86.075000 61.880000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 86.485000 61.880000 86.805000 ;
      LAYER met4 ;
        RECT 61.560000 86.485000 61.880000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 86.895000 61.880000 87.215000 ;
      LAYER met4 ;
        RECT 61.560000 86.895000 61.880000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 87.305000 61.880000 87.625000 ;
      LAYER met4 ;
        RECT 61.560000 87.305000 61.880000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 87.715000 61.880000 88.035000 ;
      LAYER met4 ;
        RECT 61.560000 87.715000 61.880000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 88.125000 61.880000 88.445000 ;
      LAYER met4 ;
        RECT 61.560000 88.125000 61.880000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 88.535000 61.880000 88.855000 ;
      LAYER met4 ;
        RECT 61.560000 88.535000 61.880000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 88.945000 61.880000 89.265000 ;
      LAYER met4 ;
        RECT 61.560000 88.945000 61.880000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 89.355000 61.880000 89.675000 ;
      LAYER met4 ;
        RECT 61.560000 89.355000 61.880000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 89.765000 61.880000 90.085000 ;
      LAYER met4 ;
        RECT 61.560000 89.765000 61.880000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 90.175000 61.880000 90.495000 ;
      LAYER met4 ;
        RECT 61.560000 90.175000 61.880000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 90.585000 61.880000 90.905000 ;
      LAYER met4 ;
        RECT 61.560000 90.585000 61.880000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 90.995000 61.880000 91.315000 ;
      LAYER met4 ;
        RECT 61.560000 90.995000 61.880000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 91.405000 61.880000 91.725000 ;
      LAYER met4 ;
        RECT 61.560000 91.405000 61.880000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 91.815000 61.880000 92.135000 ;
      LAYER met4 ;
        RECT 61.560000 91.815000 61.880000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 92.225000 61.880000 92.545000 ;
      LAYER met4 ;
        RECT 61.560000 92.225000 61.880000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560000 92.635000 61.880000 92.955000 ;
      LAYER met4 ;
        RECT 61.560000 92.635000 61.880000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.720000 17.800000 62.040000 18.120000 ;
      LAYER met4 ;
        RECT 61.720000 17.800000 62.040000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.720000 18.230000 62.040000 18.550000 ;
      LAYER met4 ;
        RECT 61.720000 18.230000 62.040000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.720000 18.660000 62.040000 18.980000 ;
      LAYER met4 ;
        RECT 61.720000 18.660000 62.040000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.720000 19.090000 62.040000 19.410000 ;
      LAYER met4 ;
        RECT 61.720000 19.090000 62.040000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.720000 19.520000 62.040000 19.840000 ;
      LAYER met4 ;
        RECT 61.720000 19.520000 62.040000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.720000 19.950000 62.040000 20.270000 ;
      LAYER met4 ;
        RECT 61.720000 19.950000 62.040000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.720000 20.380000 62.040000 20.700000 ;
      LAYER met4 ;
        RECT 61.720000 20.380000 62.040000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.720000 20.810000 62.040000 21.130000 ;
      LAYER met4 ;
        RECT 61.720000 20.810000 62.040000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.720000 21.240000 62.040000 21.560000 ;
      LAYER met4 ;
        RECT 61.720000 21.240000 62.040000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.720000 21.670000 62.040000 21.990000 ;
      LAYER met4 ;
        RECT 61.720000 21.670000 62.040000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.720000 22.100000 62.040000 22.420000 ;
      LAYER met4 ;
        RECT 61.720000 22.100000 62.040000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 68.065000 62.070000 68.385000 ;
      LAYER met4 ;
        RECT 61.750000 68.065000 62.070000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 68.475000 62.070000 68.795000 ;
      LAYER met4 ;
        RECT 61.750000 68.475000 62.070000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 68.885000 62.070000 69.205000 ;
      LAYER met4 ;
        RECT 61.750000 68.885000 62.070000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 69.295000 62.070000 69.615000 ;
      LAYER met4 ;
        RECT 61.750000 69.295000 62.070000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 69.705000 62.070000 70.025000 ;
      LAYER met4 ;
        RECT 61.750000 69.705000 62.070000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 70.115000 62.070000 70.435000 ;
      LAYER met4 ;
        RECT 61.750000 70.115000 62.070000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 70.525000 62.070000 70.845000 ;
      LAYER met4 ;
        RECT 61.750000 70.525000 62.070000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 70.935000 62.070000 71.255000 ;
      LAYER met4 ;
        RECT 61.750000 70.935000 62.070000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 71.345000 62.070000 71.665000 ;
      LAYER met4 ;
        RECT 61.750000 71.345000 62.070000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 71.755000 62.070000 72.075000 ;
      LAYER met4 ;
        RECT 61.750000 71.755000 62.070000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 72.165000 62.070000 72.485000 ;
      LAYER met4 ;
        RECT 61.750000 72.165000 62.070000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 72.575000 62.070000 72.895000 ;
      LAYER met4 ;
        RECT 61.750000 72.575000 62.070000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 72.985000 62.070000 73.305000 ;
      LAYER met4 ;
        RECT 61.750000 72.985000 62.070000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 73.390000 62.070000 73.710000 ;
      LAYER met4 ;
        RECT 61.750000 73.390000 62.070000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 73.795000 62.070000 74.115000 ;
      LAYER met4 ;
        RECT 61.750000 73.795000 62.070000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 74.200000 62.070000 74.520000 ;
      LAYER met4 ;
        RECT 61.750000 74.200000 62.070000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 74.605000 62.070000 74.925000 ;
      LAYER met4 ;
        RECT 61.750000 74.605000 62.070000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 75.010000 62.070000 75.330000 ;
      LAYER met4 ;
        RECT 61.750000 75.010000 62.070000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 75.415000 62.070000 75.735000 ;
      LAYER met4 ;
        RECT 61.750000 75.415000 62.070000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 75.820000 62.070000 76.140000 ;
      LAYER met4 ;
        RECT 61.750000 75.820000 62.070000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 76.225000 62.070000 76.545000 ;
      LAYER met4 ;
        RECT 61.750000 76.225000 62.070000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 76.630000 62.070000 76.950000 ;
      LAYER met4 ;
        RECT 61.750000 76.630000 62.070000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 77.035000 62.070000 77.355000 ;
      LAYER met4 ;
        RECT 61.750000 77.035000 62.070000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 77.440000 62.070000 77.760000 ;
      LAYER met4 ;
        RECT 61.750000 77.440000 62.070000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 77.845000 62.070000 78.165000 ;
      LAYER met4 ;
        RECT 61.750000 77.845000 62.070000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 78.250000 62.070000 78.570000 ;
      LAYER met4 ;
        RECT 61.750000 78.250000 62.070000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 78.655000 62.070000 78.975000 ;
      LAYER met4 ;
        RECT 61.750000 78.655000 62.070000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 79.060000 62.070000 79.380000 ;
      LAYER met4 ;
        RECT 61.750000 79.060000 62.070000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 79.465000 62.070000 79.785000 ;
      LAYER met4 ;
        RECT 61.750000 79.465000 62.070000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 79.870000 62.070000 80.190000 ;
      LAYER met4 ;
        RECT 61.750000 79.870000 62.070000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 80.275000 62.070000 80.595000 ;
      LAYER met4 ;
        RECT 61.750000 80.275000 62.070000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 80.680000 62.070000 81.000000 ;
      LAYER met4 ;
        RECT 61.750000 80.680000 62.070000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 81.085000 62.070000 81.405000 ;
      LAYER met4 ;
        RECT 61.750000 81.085000 62.070000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 81.490000 62.070000 81.810000 ;
      LAYER met4 ;
        RECT 61.750000 81.490000 62.070000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 81.895000 62.070000 82.215000 ;
      LAYER met4 ;
        RECT 61.750000 81.895000 62.070000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 82.300000 62.070000 82.620000 ;
      LAYER met4 ;
        RECT 61.750000 82.300000 62.070000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 82.795000 62.285000 83.115000 ;
      LAYER met4 ;
        RECT 61.965000 82.795000 62.285000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 83.205000 62.285000 83.525000 ;
      LAYER met4 ;
        RECT 61.965000 83.205000 62.285000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 83.615000 62.285000 83.935000 ;
      LAYER met4 ;
        RECT 61.965000 83.615000 62.285000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 84.025000 62.285000 84.345000 ;
      LAYER met4 ;
        RECT 61.965000 84.025000 62.285000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 84.435000 62.285000 84.755000 ;
      LAYER met4 ;
        RECT 61.965000 84.435000 62.285000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 84.845000 62.285000 85.165000 ;
      LAYER met4 ;
        RECT 61.965000 84.845000 62.285000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 85.255000 62.285000 85.575000 ;
      LAYER met4 ;
        RECT 61.965000 85.255000 62.285000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 85.665000 62.285000 85.985000 ;
      LAYER met4 ;
        RECT 61.965000 85.665000 62.285000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 86.075000 62.285000 86.395000 ;
      LAYER met4 ;
        RECT 61.965000 86.075000 62.285000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 86.485000 62.285000 86.805000 ;
      LAYER met4 ;
        RECT 61.965000 86.485000 62.285000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 86.895000 62.285000 87.215000 ;
      LAYER met4 ;
        RECT 61.965000 86.895000 62.285000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 87.305000 62.285000 87.625000 ;
      LAYER met4 ;
        RECT 61.965000 87.305000 62.285000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 87.715000 62.285000 88.035000 ;
      LAYER met4 ;
        RECT 61.965000 87.715000 62.285000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 88.125000 62.285000 88.445000 ;
      LAYER met4 ;
        RECT 61.965000 88.125000 62.285000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 88.535000 62.285000 88.855000 ;
      LAYER met4 ;
        RECT 61.965000 88.535000 62.285000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 88.945000 62.285000 89.265000 ;
      LAYER met4 ;
        RECT 61.965000 88.945000 62.285000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 89.355000 62.285000 89.675000 ;
      LAYER met4 ;
        RECT 61.965000 89.355000 62.285000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 89.765000 62.285000 90.085000 ;
      LAYER met4 ;
        RECT 61.965000 89.765000 62.285000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 90.175000 62.285000 90.495000 ;
      LAYER met4 ;
        RECT 61.965000 90.175000 62.285000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 90.585000 62.285000 90.905000 ;
      LAYER met4 ;
        RECT 61.965000 90.585000 62.285000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 90.995000 62.285000 91.315000 ;
      LAYER met4 ;
        RECT 61.965000 90.995000 62.285000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 91.405000 62.285000 91.725000 ;
      LAYER met4 ;
        RECT 61.965000 91.405000 62.285000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 91.815000 62.285000 92.135000 ;
      LAYER met4 ;
        RECT 61.965000 91.815000 62.285000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 92.225000 62.285000 92.545000 ;
      LAYER met4 ;
        RECT 61.965000 92.225000 62.285000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965000 92.635000 62.285000 92.955000 ;
      LAYER met4 ;
        RECT 61.965000 92.635000 62.285000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.125000 17.800000 62.445000 18.120000 ;
      LAYER met4 ;
        RECT 62.125000 17.800000 62.445000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.125000 18.230000 62.445000 18.550000 ;
      LAYER met4 ;
        RECT 62.125000 18.230000 62.445000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.125000 18.660000 62.445000 18.980000 ;
      LAYER met4 ;
        RECT 62.125000 18.660000 62.445000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.125000 19.090000 62.445000 19.410000 ;
      LAYER met4 ;
        RECT 62.125000 19.090000 62.445000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.125000 19.520000 62.445000 19.840000 ;
      LAYER met4 ;
        RECT 62.125000 19.520000 62.445000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.125000 19.950000 62.445000 20.270000 ;
      LAYER met4 ;
        RECT 62.125000 19.950000 62.445000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.125000 20.380000 62.445000 20.700000 ;
      LAYER met4 ;
        RECT 62.125000 20.380000 62.445000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.125000 20.810000 62.445000 21.130000 ;
      LAYER met4 ;
        RECT 62.125000 20.810000 62.445000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.125000 21.240000 62.445000 21.560000 ;
      LAYER met4 ;
        RECT 62.125000 21.240000 62.445000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.125000 21.670000 62.445000 21.990000 ;
      LAYER met4 ;
        RECT 62.125000 21.670000 62.445000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.125000 22.100000 62.445000 22.420000 ;
      LAYER met4 ;
        RECT 62.125000 22.100000 62.445000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 68.065000 62.470000 68.385000 ;
      LAYER met4 ;
        RECT 62.150000 68.065000 62.470000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 68.475000 62.470000 68.795000 ;
      LAYER met4 ;
        RECT 62.150000 68.475000 62.470000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 68.885000 62.470000 69.205000 ;
      LAYER met4 ;
        RECT 62.150000 68.885000 62.470000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 69.295000 62.470000 69.615000 ;
      LAYER met4 ;
        RECT 62.150000 69.295000 62.470000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 69.705000 62.470000 70.025000 ;
      LAYER met4 ;
        RECT 62.150000 69.705000 62.470000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 70.115000 62.470000 70.435000 ;
      LAYER met4 ;
        RECT 62.150000 70.115000 62.470000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 70.525000 62.470000 70.845000 ;
      LAYER met4 ;
        RECT 62.150000 70.525000 62.470000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 70.935000 62.470000 71.255000 ;
      LAYER met4 ;
        RECT 62.150000 70.935000 62.470000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 71.345000 62.470000 71.665000 ;
      LAYER met4 ;
        RECT 62.150000 71.345000 62.470000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 71.755000 62.470000 72.075000 ;
      LAYER met4 ;
        RECT 62.150000 71.755000 62.470000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 72.165000 62.470000 72.485000 ;
      LAYER met4 ;
        RECT 62.150000 72.165000 62.470000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 72.575000 62.470000 72.895000 ;
      LAYER met4 ;
        RECT 62.150000 72.575000 62.470000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 72.985000 62.470000 73.305000 ;
      LAYER met4 ;
        RECT 62.150000 72.985000 62.470000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 73.390000 62.470000 73.710000 ;
      LAYER met4 ;
        RECT 62.150000 73.390000 62.470000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 73.795000 62.470000 74.115000 ;
      LAYER met4 ;
        RECT 62.150000 73.795000 62.470000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 74.200000 62.470000 74.520000 ;
      LAYER met4 ;
        RECT 62.150000 74.200000 62.470000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 74.605000 62.470000 74.925000 ;
      LAYER met4 ;
        RECT 62.150000 74.605000 62.470000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 75.010000 62.470000 75.330000 ;
      LAYER met4 ;
        RECT 62.150000 75.010000 62.470000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 75.415000 62.470000 75.735000 ;
      LAYER met4 ;
        RECT 62.150000 75.415000 62.470000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 75.820000 62.470000 76.140000 ;
      LAYER met4 ;
        RECT 62.150000 75.820000 62.470000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 76.225000 62.470000 76.545000 ;
      LAYER met4 ;
        RECT 62.150000 76.225000 62.470000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 76.630000 62.470000 76.950000 ;
      LAYER met4 ;
        RECT 62.150000 76.630000 62.470000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 77.035000 62.470000 77.355000 ;
      LAYER met4 ;
        RECT 62.150000 77.035000 62.470000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 77.440000 62.470000 77.760000 ;
      LAYER met4 ;
        RECT 62.150000 77.440000 62.470000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 77.845000 62.470000 78.165000 ;
      LAYER met4 ;
        RECT 62.150000 77.845000 62.470000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 78.250000 62.470000 78.570000 ;
      LAYER met4 ;
        RECT 62.150000 78.250000 62.470000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 78.655000 62.470000 78.975000 ;
      LAYER met4 ;
        RECT 62.150000 78.655000 62.470000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 79.060000 62.470000 79.380000 ;
      LAYER met4 ;
        RECT 62.150000 79.060000 62.470000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 79.465000 62.470000 79.785000 ;
      LAYER met4 ;
        RECT 62.150000 79.465000 62.470000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 79.870000 62.470000 80.190000 ;
      LAYER met4 ;
        RECT 62.150000 79.870000 62.470000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 80.275000 62.470000 80.595000 ;
      LAYER met4 ;
        RECT 62.150000 80.275000 62.470000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 80.680000 62.470000 81.000000 ;
      LAYER met4 ;
        RECT 62.150000 80.680000 62.470000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 81.085000 62.470000 81.405000 ;
      LAYER met4 ;
        RECT 62.150000 81.085000 62.470000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 81.490000 62.470000 81.810000 ;
      LAYER met4 ;
        RECT 62.150000 81.490000 62.470000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 81.895000 62.470000 82.215000 ;
      LAYER met4 ;
        RECT 62.150000 81.895000 62.470000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.150000 82.300000 62.470000 82.620000 ;
      LAYER met4 ;
        RECT 62.150000 82.300000 62.470000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 82.795000 62.690000 83.115000 ;
      LAYER met4 ;
        RECT 62.370000 82.795000 62.690000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 83.205000 62.690000 83.525000 ;
      LAYER met4 ;
        RECT 62.370000 83.205000 62.690000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 83.615000 62.690000 83.935000 ;
      LAYER met4 ;
        RECT 62.370000 83.615000 62.690000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 84.025000 62.690000 84.345000 ;
      LAYER met4 ;
        RECT 62.370000 84.025000 62.690000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 84.435000 62.690000 84.755000 ;
      LAYER met4 ;
        RECT 62.370000 84.435000 62.690000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 84.845000 62.690000 85.165000 ;
      LAYER met4 ;
        RECT 62.370000 84.845000 62.690000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 85.255000 62.690000 85.575000 ;
      LAYER met4 ;
        RECT 62.370000 85.255000 62.690000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 85.665000 62.690000 85.985000 ;
      LAYER met4 ;
        RECT 62.370000 85.665000 62.690000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 86.075000 62.690000 86.395000 ;
      LAYER met4 ;
        RECT 62.370000 86.075000 62.690000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 86.485000 62.690000 86.805000 ;
      LAYER met4 ;
        RECT 62.370000 86.485000 62.690000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 86.895000 62.690000 87.215000 ;
      LAYER met4 ;
        RECT 62.370000 86.895000 62.690000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 87.305000 62.690000 87.625000 ;
      LAYER met4 ;
        RECT 62.370000 87.305000 62.690000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 87.715000 62.690000 88.035000 ;
      LAYER met4 ;
        RECT 62.370000 87.715000 62.690000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 88.125000 62.690000 88.445000 ;
      LAYER met4 ;
        RECT 62.370000 88.125000 62.690000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 88.535000 62.690000 88.855000 ;
      LAYER met4 ;
        RECT 62.370000 88.535000 62.690000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 88.945000 62.690000 89.265000 ;
      LAYER met4 ;
        RECT 62.370000 88.945000 62.690000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 89.355000 62.690000 89.675000 ;
      LAYER met4 ;
        RECT 62.370000 89.355000 62.690000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 89.765000 62.690000 90.085000 ;
      LAYER met4 ;
        RECT 62.370000 89.765000 62.690000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 90.175000 62.690000 90.495000 ;
      LAYER met4 ;
        RECT 62.370000 90.175000 62.690000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 90.585000 62.690000 90.905000 ;
      LAYER met4 ;
        RECT 62.370000 90.585000 62.690000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 90.995000 62.690000 91.315000 ;
      LAYER met4 ;
        RECT 62.370000 90.995000 62.690000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 91.405000 62.690000 91.725000 ;
      LAYER met4 ;
        RECT 62.370000 91.405000 62.690000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 91.815000 62.690000 92.135000 ;
      LAYER met4 ;
        RECT 62.370000 91.815000 62.690000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 92.225000 62.690000 92.545000 ;
      LAYER met4 ;
        RECT 62.370000 92.225000 62.690000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370000 92.635000 62.690000 92.955000 ;
      LAYER met4 ;
        RECT 62.370000 92.635000 62.690000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.530000 17.800000 62.850000 18.120000 ;
      LAYER met4 ;
        RECT 62.530000 17.800000 62.850000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.530000 18.230000 62.850000 18.550000 ;
      LAYER met4 ;
        RECT 62.530000 18.230000 62.850000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.530000 18.660000 62.850000 18.980000 ;
      LAYER met4 ;
        RECT 62.530000 18.660000 62.850000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.530000 19.090000 62.850000 19.410000 ;
      LAYER met4 ;
        RECT 62.530000 19.090000 62.850000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.530000 19.520000 62.850000 19.840000 ;
      LAYER met4 ;
        RECT 62.530000 19.520000 62.850000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.530000 19.950000 62.850000 20.270000 ;
      LAYER met4 ;
        RECT 62.530000 19.950000 62.850000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.530000 20.380000 62.850000 20.700000 ;
      LAYER met4 ;
        RECT 62.530000 20.380000 62.850000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.530000 20.810000 62.850000 21.130000 ;
      LAYER met4 ;
        RECT 62.530000 20.810000 62.850000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.530000 21.240000 62.850000 21.560000 ;
      LAYER met4 ;
        RECT 62.530000 21.240000 62.850000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.530000 21.670000 62.850000 21.990000 ;
      LAYER met4 ;
        RECT 62.530000 21.670000 62.850000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.530000 22.100000 62.850000 22.420000 ;
      LAYER met4 ;
        RECT 62.530000 22.100000 62.850000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 68.065000 62.870000 68.385000 ;
      LAYER met4 ;
        RECT 62.550000 68.065000 62.870000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 68.475000 62.870000 68.795000 ;
      LAYER met4 ;
        RECT 62.550000 68.475000 62.870000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 68.885000 62.870000 69.205000 ;
      LAYER met4 ;
        RECT 62.550000 68.885000 62.870000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 69.295000 62.870000 69.615000 ;
      LAYER met4 ;
        RECT 62.550000 69.295000 62.870000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 69.705000 62.870000 70.025000 ;
      LAYER met4 ;
        RECT 62.550000 69.705000 62.870000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 70.115000 62.870000 70.435000 ;
      LAYER met4 ;
        RECT 62.550000 70.115000 62.870000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 70.525000 62.870000 70.845000 ;
      LAYER met4 ;
        RECT 62.550000 70.525000 62.870000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 70.935000 62.870000 71.255000 ;
      LAYER met4 ;
        RECT 62.550000 70.935000 62.870000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 71.345000 62.870000 71.665000 ;
      LAYER met4 ;
        RECT 62.550000 71.345000 62.870000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 71.755000 62.870000 72.075000 ;
      LAYER met4 ;
        RECT 62.550000 71.755000 62.870000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 72.165000 62.870000 72.485000 ;
      LAYER met4 ;
        RECT 62.550000 72.165000 62.870000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 72.575000 62.870000 72.895000 ;
      LAYER met4 ;
        RECT 62.550000 72.575000 62.870000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 72.985000 62.870000 73.305000 ;
      LAYER met4 ;
        RECT 62.550000 72.985000 62.870000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 73.390000 62.870000 73.710000 ;
      LAYER met4 ;
        RECT 62.550000 73.390000 62.870000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 73.795000 62.870000 74.115000 ;
      LAYER met4 ;
        RECT 62.550000 73.795000 62.870000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 74.200000 62.870000 74.520000 ;
      LAYER met4 ;
        RECT 62.550000 74.200000 62.870000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 74.605000 62.870000 74.925000 ;
      LAYER met4 ;
        RECT 62.550000 74.605000 62.870000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 75.010000 62.870000 75.330000 ;
      LAYER met4 ;
        RECT 62.550000 75.010000 62.870000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 75.415000 62.870000 75.735000 ;
      LAYER met4 ;
        RECT 62.550000 75.415000 62.870000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 75.820000 62.870000 76.140000 ;
      LAYER met4 ;
        RECT 62.550000 75.820000 62.870000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 76.225000 62.870000 76.545000 ;
      LAYER met4 ;
        RECT 62.550000 76.225000 62.870000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 76.630000 62.870000 76.950000 ;
      LAYER met4 ;
        RECT 62.550000 76.630000 62.870000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 77.035000 62.870000 77.355000 ;
      LAYER met4 ;
        RECT 62.550000 77.035000 62.870000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 77.440000 62.870000 77.760000 ;
      LAYER met4 ;
        RECT 62.550000 77.440000 62.870000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 77.845000 62.870000 78.165000 ;
      LAYER met4 ;
        RECT 62.550000 77.845000 62.870000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 78.250000 62.870000 78.570000 ;
      LAYER met4 ;
        RECT 62.550000 78.250000 62.870000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 78.655000 62.870000 78.975000 ;
      LAYER met4 ;
        RECT 62.550000 78.655000 62.870000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 79.060000 62.870000 79.380000 ;
      LAYER met4 ;
        RECT 62.550000 79.060000 62.870000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 79.465000 62.870000 79.785000 ;
      LAYER met4 ;
        RECT 62.550000 79.465000 62.870000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 79.870000 62.870000 80.190000 ;
      LAYER met4 ;
        RECT 62.550000 79.870000 62.870000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 80.275000 62.870000 80.595000 ;
      LAYER met4 ;
        RECT 62.550000 80.275000 62.870000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 80.680000 62.870000 81.000000 ;
      LAYER met4 ;
        RECT 62.550000 80.680000 62.870000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 81.085000 62.870000 81.405000 ;
      LAYER met4 ;
        RECT 62.550000 81.085000 62.870000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 81.490000 62.870000 81.810000 ;
      LAYER met4 ;
        RECT 62.550000 81.490000 62.870000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 81.895000 62.870000 82.215000 ;
      LAYER met4 ;
        RECT 62.550000 81.895000 62.870000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550000 82.300000 62.870000 82.620000 ;
      LAYER met4 ;
        RECT 62.550000 82.300000 62.870000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 82.795000 63.100000 83.115000 ;
      LAYER met4 ;
        RECT 62.780000 82.795000 63.100000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 83.205000 63.100000 83.525000 ;
      LAYER met4 ;
        RECT 62.780000 83.205000 63.100000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 83.615000 63.100000 83.935000 ;
      LAYER met4 ;
        RECT 62.780000 83.615000 63.100000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 84.025000 63.100000 84.345000 ;
      LAYER met4 ;
        RECT 62.780000 84.025000 63.100000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 84.435000 63.100000 84.755000 ;
      LAYER met4 ;
        RECT 62.780000 84.435000 63.100000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 84.845000 63.100000 85.165000 ;
      LAYER met4 ;
        RECT 62.780000 84.845000 63.100000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 85.255000 63.100000 85.575000 ;
      LAYER met4 ;
        RECT 62.780000 85.255000 63.100000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 85.665000 63.100000 85.985000 ;
      LAYER met4 ;
        RECT 62.780000 85.665000 63.100000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 86.075000 63.100000 86.395000 ;
      LAYER met4 ;
        RECT 62.780000 86.075000 63.100000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 86.485000 63.100000 86.805000 ;
      LAYER met4 ;
        RECT 62.780000 86.485000 63.100000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 86.895000 63.100000 87.215000 ;
      LAYER met4 ;
        RECT 62.780000 86.895000 63.100000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 87.305000 63.100000 87.625000 ;
      LAYER met4 ;
        RECT 62.780000 87.305000 63.100000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 87.715000 63.100000 88.035000 ;
      LAYER met4 ;
        RECT 62.780000 87.715000 63.100000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 88.125000 63.100000 88.445000 ;
      LAYER met4 ;
        RECT 62.780000 88.125000 63.100000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 88.535000 63.100000 88.855000 ;
      LAYER met4 ;
        RECT 62.780000 88.535000 63.100000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 88.945000 63.100000 89.265000 ;
      LAYER met4 ;
        RECT 62.780000 88.945000 63.100000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 89.355000 63.100000 89.675000 ;
      LAYER met4 ;
        RECT 62.780000 89.355000 63.100000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 89.765000 63.100000 90.085000 ;
      LAYER met4 ;
        RECT 62.780000 89.765000 63.100000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 90.175000 63.100000 90.495000 ;
      LAYER met4 ;
        RECT 62.780000 90.175000 63.100000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 90.585000 63.100000 90.905000 ;
      LAYER met4 ;
        RECT 62.780000 90.585000 63.100000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 90.995000 63.100000 91.315000 ;
      LAYER met4 ;
        RECT 62.780000 90.995000 63.100000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 91.405000 63.100000 91.725000 ;
      LAYER met4 ;
        RECT 62.780000 91.405000 63.100000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 91.815000 63.100000 92.135000 ;
      LAYER met4 ;
        RECT 62.780000 91.815000 63.100000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 92.225000 63.100000 92.545000 ;
      LAYER met4 ;
        RECT 62.780000 92.225000 63.100000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780000 92.635000 63.100000 92.955000 ;
      LAYER met4 ;
        RECT 62.780000 92.635000 63.100000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.935000 17.800000 63.255000 18.120000 ;
      LAYER met4 ;
        RECT 62.935000 17.800000 63.255000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.935000 18.230000 63.255000 18.550000 ;
      LAYER met4 ;
        RECT 62.935000 18.230000 63.255000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.935000 18.660000 63.255000 18.980000 ;
      LAYER met4 ;
        RECT 62.935000 18.660000 63.255000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.935000 19.090000 63.255000 19.410000 ;
      LAYER met4 ;
        RECT 62.935000 19.090000 63.255000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.935000 19.520000 63.255000 19.840000 ;
      LAYER met4 ;
        RECT 62.935000 19.520000 63.255000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.935000 19.950000 63.255000 20.270000 ;
      LAYER met4 ;
        RECT 62.935000 19.950000 63.255000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.935000 20.380000 63.255000 20.700000 ;
      LAYER met4 ;
        RECT 62.935000 20.380000 63.255000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.935000 20.810000 63.255000 21.130000 ;
      LAYER met4 ;
        RECT 62.935000 20.810000 63.255000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.935000 21.240000 63.255000 21.560000 ;
      LAYER met4 ;
        RECT 62.935000 21.240000 63.255000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.935000 21.670000 63.255000 21.990000 ;
      LAYER met4 ;
        RECT 62.935000 21.670000 63.255000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.935000 22.100000 63.255000 22.420000 ;
      LAYER met4 ;
        RECT 62.935000 22.100000 63.255000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 68.065000 63.270000 68.385000 ;
      LAYER met4 ;
        RECT 62.950000 68.065000 63.270000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 68.475000 63.270000 68.795000 ;
      LAYER met4 ;
        RECT 62.950000 68.475000 63.270000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 68.885000 63.270000 69.205000 ;
      LAYER met4 ;
        RECT 62.950000 68.885000 63.270000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 69.295000 63.270000 69.615000 ;
      LAYER met4 ;
        RECT 62.950000 69.295000 63.270000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 69.705000 63.270000 70.025000 ;
      LAYER met4 ;
        RECT 62.950000 69.705000 63.270000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 70.115000 63.270000 70.435000 ;
      LAYER met4 ;
        RECT 62.950000 70.115000 63.270000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 70.525000 63.270000 70.845000 ;
      LAYER met4 ;
        RECT 62.950000 70.525000 63.270000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 70.935000 63.270000 71.255000 ;
      LAYER met4 ;
        RECT 62.950000 70.935000 63.270000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 71.345000 63.270000 71.665000 ;
      LAYER met4 ;
        RECT 62.950000 71.345000 63.270000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 71.755000 63.270000 72.075000 ;
      LAYER met4 ;
        RECT 62.950000 71.755000 63.270000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 72.165000 63.270000 72.485000 ;
      LAYER met4 ;
        RECT 62.950000 72.165000 63.270000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 72.575000 63.270000 72.895000 ;
      LAYER met4 ;
        RECT 62.950000 72.575000 63.270000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 72.985000 63.270000 73.305000 ;
      LAYER met4 ;
        RECT 62.950000 72.985000 63.270000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 73.390000 63.270000 73.710000 ;
      LAYER met4 ;
        RECT 62.950000 73.390000 63.270000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 73.795000 63.270000 74.115000 ;
      LAYER met4 ;
        RECT 62.950000 73.795000 63.270000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 74.200000 63.270000 74.520000 ;
      LAYER met4 ;
        RECT 62.950000 74.200000 63.270000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 74.605000 63.270000 74.925000 ;
      LAYER met4 ;
        RECT 62.950000 74.605000 63.270000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 75.010000 63.270000 75.330000 ;
      LAYER met4 ;
        RECT 62.950000 75.010000 63.270000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 75.415000 63.270000 75.735000 ;
      LAYER met4 ;
        RECT 62.950000 75.415000 63.270000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 75.820000 63.270000 76.140000 ;
      LAYER met4 ;
        RECT 62.950000 75.820000 63.270000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 76.225000 63.270000 76.545000 ;
      LAYER met4 ;
        RECT 62.950000 76.225000 63.270000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 76.630000 63.270000 76.950000 ;
      LAYER met4 ;
        RECT 62.950000 76.630000 63.270000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 77.035000 63.270000 77.355000 ;
      LAYER met4 ;
        RECT 62.950000 77.035000 63.270000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 77.440000 63.270000 77.760000 ;
      LAYER met4 ;
        RECT 62.950000 77.440000 63.270000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 77.845000 63.270000 78.165000 ;
      LAYER met4 ;
        RECT 62.950000 77.845000 63.270000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 78.250000 63.270000 78.570000 ;
      LAYER met4 ;
        RECT 62.950000 78.250000 63.270000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 78.655000 63.270000 78.975000 ;
      LAYER met4 ;
        RECT 62.950000 78.655000 63.270000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 79.060000 63.270000 79.380000 ;
      LAYER met4 ;
        RECT 62.950000 79.060000 63.270000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 79.465000 63.270000 79.785000 ;
      LAYER met4 ;
        RECT 62.950000 79.465000 63.270000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 79.870000 63.270000 80.190000 ;
      LAYER met4 ;
        RECT 62.950000 79.870000 63.270000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 80.275000 63.270000 80.595000 ;
      LAYER met4 ;
        RECT 62.950000 80.275000 63.270000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 80.680000 63.270000 81.000000 ;
      LAYER met4 ;
        RECT 62.950000 80.680000 63.270000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 81.085000 63.270000 81.405000 ;
      LAYER met4 ;
        RECT 62.950000 81.085000 63.270000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 81.490000 63.270000 81.810000 ;
      LAYER met4 ;
        RECT 62.950000 81.490000 63.270000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 81.895000 63.270000 82.215000 ;
      LAYER met4 ;
        RECT 62.950000 81.895000 63.270000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.950000 82.300000 63.270000 82.620000 ;
      LAYER met4 ;
        RECT 62.950000 82.300000 63.270000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 82.795000 63.510000 83.115000 ;
      LAYER met4 ;
        RECT 63.190000 82.795000 63.510000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 83.205000 63.510000 83.525000 ;
      LAYER met4 ;
        RECT 63.190000 83.205000 63.510000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 83.615000 63.510000 83.935000 ;
      LAYER met4 ;
        RECT 63.190000 83.615000 63.510000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 84.025000 63.510000 84.345000 ;
      LAYER met4 ;
        RECT 63.190000 84.025000 63.510000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 84.435000 63.510000 84.755000 ;
      LAYER met4 ;
        RECT 63.190000 84.435000 63.510000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 84.845000 63.510000 85.165000 ;
      LAYER met4 ;
        RECT 63.190000 84.845000 63.510000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 85.255000 63.510000 85.575000 ;
      LAYER met4 ;
        RECT 63.190000 85.255000 63.510000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 85.665000 63.510000 85.985000 ;
      LAYER met4 ;
        RECT 63.190000 85.665000 63.510000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 86.075000 63.510000 86.395000 ;
      LAYER met4 ;
        RECT 63.190000 86.075000 63.510000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 86.485000 63.510000 86.805000 ;
      LAYER met4 ;
        RECT 63.190000 86.485000 63.510000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 86.895000 63.510000 87.215000 ;
      LAYER met4 ;
        RECT 63.190000 86.895000 63.510000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 87.305000 63.510000 87.625000 ;
      LAYER met4 ;
        RECT 63.190000 87.305000 63.510000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 87.715000 63.510000 88.035000 ;
      LAYER met4 ;
        RECT 63.190000 87.715000 63.510000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 88.125000 63.510000 88.445000 ;
      LAYER met4 ;
        RECT 63.190000 88.125000 63.510000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 88.535000 63.510000 88.855000 ;
      LAYER met4 ;
        RECT 63.190000 88.535000 63.510000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 88.945000 63.510000 89.265000 ;
      LAYER met4 ;
        RECT 63.190000 88.945000 63.510000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 89.355000 63.510000 89.675000 ;
      LAYER met4 ;
        RECT 63.190000 89.355000 63.510000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 89.765000 63.510000 90.085000 ;
      LAYER met4 ;
        RECT 63.190000 89.765000 63.510000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 90.175000 63.510000 90.495000 ;
      LAYER met4 ;
        RECT 63.190000 90.175000 63.510000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 90.585000 63.510000 90.905000 ;
      LAYER met4 ;
        RECT 63.190000 90.585000 63.510000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 90.995000 63.510000 91.315000 ;
      LAYER met4 ;
        RECT 63.190000 90.995000 63.510000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 91.405000 63.510000 91.725000 ;
      LAYER met4 ;
        RECT 63.190000 91.405000 63.510000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 91.815000 63.510000 92.135000 ;
      LAYER met4 ;
        RECT 63.190000 91.815000 63.510000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 92.225000 63.510000 92.545000 ;
      LAYER met4 ;
        RECT 63.190000 92.225000 63.510000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190000 92.635000 63.510000 92.955000 ;
      LAYER met4 ;
        RECT 63.190000 92.635000 63.510000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.340000 17.800000 63.660000 18.120000 ;
      LAYER met4 ;
        RECT 63.340000 17.800000 63.660000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.340000 18.230000 63.660000 18.550000 ;
      LAYER met4 ;
        RECT 63.340000 18.230000 63.660000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.340000 18.660000 63.660000 18.980000 ;
      LAYER met4 ;
        RECT 63.340000 18.660000 63.660000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.340000 19.090000 63.660000 19.410000 ;
      LAYER met4 ;
        RECT 63.340000 19.090000 63.660000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.340000 19.520000 63.660000 19.840000 ;
      LAYER met4 ;
        RECT 63.340000 19.520000 63.660000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.340000 19.950000 63.660000 20.270000 ;
      LAYER met4 ;
        RECT 63.340000 19.950000 63.660000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.340000 20.380000 63.660000 20.700000 ;
      LAYER met4 ;
        RECT 63.340000 20.380000 63.660000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.340000 20.810000 63.660000 21.130000 ;
      LAYER met4 ;
        RECT 63.340000 20.810000 63.660000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.340000 21.240000 63.660000 21.560000 ;
      LAYER met4 ;
        RECT 63.340000 21.240000 63.660000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.340000 21.670000 63.660000 21.990000 ;
      LAYER met4 ;
        RECT 63.340000 21.670000 63.660000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.340000 22.100000 63.660000 22.420000 ;
      LAYER met4 ;
        RECT 63.340000 22.100000 63.660000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 68.065000 63.670000 68.385000 ;
      LAYER met4 ;
        RECT 63.350000 68.065000 63.670000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 68.475000 63.670000 68.795000 ;
      LAYER met4 ;
        RECT 63.350000 68.475000 63.670000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 68.885000 63.670000 69.205000 ;
      LAYER met4 ;
        RECT 63.350000 68.885000 63.670000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 69.295000 63.670000 69.615000 ;
      LAYER met4 ;
        RECT 63.350000 69.295000 63.670000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 69.705000 63.670000 70.025000 ;
      LAYER met4 ;
        RECT 63.350000 69.705000 63.670000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 70.115000 63.670000 70.435000 ;
      LAYER met4 ;
        RECT 63.350000 70.115000 63.670000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 70.525000 63.670000 70.845000 ;
      LAYER met4 ;
        RECT 63.350000 70.525000 63.670000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 70.935000 63.670000 71.255000 ;
      LAYER met4 ;
        RECT 63.350000 70.935000 63.670000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 71.345000 63.670000 71.665000 ;
      LAYER met4 ;
        RECT 63.350000 71.345000 63.670000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 71.755000 63.670000 72.075000 ;
      LAYER met4 ;
        RECT 63.350000 71.755000 63.670000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 72.165000 63.670000 72.485000 ;
      LAYER met4 ;
        RECT 63.350000 72.165000 63.670000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 72.575000 63.670000 72.895000 ;
      LAYER met4 ;
        RECT 63.350000 72.575000 63.670000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 72.985000 63.670000 73.305000 ;
      LAYER met4 ;
        RECT 63.350000 72.985000 63.670000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 73.390000 63.670000 73.710000 ;
      LAYER met4 ;
        RECT 63.350000 73.390000 63.670000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 73.795000 63.670000 74.115000 ;
      LAYER met4 ;
        RECT 63.350000 73.795000 63.670000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 74.200000 63.670000 74.520000 ;
      LAYER met4 ;
        RECT 63.350000 74.200000 63.670000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 74.605000 63.670000 74.925000 ;
      LAYER met4 ;
        RECT 63.350000 74.605000 63.670000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 75.010000 63.670000 75.330000 ;
      LAYER met4 ;
        RECT 63.350000 75.010000 63.670000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 75.415000 63.670000 75.735000 ;
      LAYER met4 ;
        RECT 63.350000 75.415000 63.670000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 75.820000 63.670000 76.140000 ;
      LAYER met4 ;
        RECT 63.350000 75.820000 63.670000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 76.225000 63.670000 76.545000 ;
      LAYER met4 ;
        RECT 63.350000 76.225000 63.670000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 76.630000 63.670000 76.950000 ;
      LAYER met4 ;
        RECT 63.350000 76.630000 63.670000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 77.035000 63.670000 77.355000 ;
      LAYER met4 ;
        RECT 63.350000 77.035000 63.670000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 77.440000 63.670000 77.760000 ;
      LAYER met4 ;
        RECT 63.350000 77.440000 63.670000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 77.845000 63.670000 78.165000 ;
      LAYER met4 ;
        RECT 63.350000 77.845000 63.670000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 78.250000 63.670000 78.570000 ;
      LAYER met4 ;
        RECT 63.350000 78.250000 63.670000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 78.655000 63.670000 78.975000 ;
      LAYER met4 ;
        RECT 63.350000 78.655000 63.670000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 79.060000 63.670000 79.380000 ;
      LAYER met4 ;
        RECT 63.350000 79.060000 63.670000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 79.465000 63.670000 79.785000 ;
      LAYER met4 ;
        RECT 63.350000 79.465000 63.670000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 79.870000 63.670000 80.190000 ;
      LAYER met4 ;
        RECT 63.350000 79.870000 63.670000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 80.275000 63.670000 80.595000 ;
      LAYER met4 ;
        RECT 63.350000 80.275000 63.670000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 80.680000 63.670000 81.000000 ;
      LAYER met4 ;
        RECT 63.350000 80.680000 63.670000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 81.085000 63.670000 81.405000 ;
      LAYER met4 ;
        RECT 63.350000 81.085000 63.670000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 81.490000 63.670000 81.810000 ;
      LAYER met4 ;
        RECT 63.350000 81.490000 63.670000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 81.895000 63.670000 82.215000 ;
      LAYER met4 ;
        RECT 63.350000 81.895000 63.670000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.350000 82.300000 63.670000 82.620000 ;
      LAYER met4 ;
        RECT 63.350000 82.300000 63.670000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 82.795000 63.920000 83.115000 ;
      LAYER met4 ;
        RECT 63.600000 82.795000 63.920000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 83.205000 63.920000 83.525000 ;
      LAYER met4 ;
        RECT 63.600000 83.205000 63.920000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 83.615000 63.920000 83.935000 ;
      LAYER met4 ;
        RECT 63.600000 83.615000 63.920000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 84.025000 63.920000 84.345000 ;
      LAYER met4 ;
        RECT 63.600000 84.025000 63.920000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 84.435000 63.920000 84.755000 ;
      LAYER met4 ;
        RECT 63.600000 84.435000 63.920000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 84.845000 63.920000 85.165000 ;
      LAYER met4 ;
        RECT 63.600000 84.845000 63.920000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 85.255000 63.920000 85.575000 ;
      LAYER met4 ;
        RECT 63.600000 85.255000 63.920000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 85.665000 63.920000 85.985000 ;
      LAYER met4 ;
        RECT 63.600000 85.665000 63.920000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 86.075000 63.920000 86.395000 ;
      LAYER met4 ;
        RECT 63.600000 86.075000 63.920000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 86.485000 63.920000 86.805000 ;
      LAYER met4 ;
        RECT 63.600000 86.485000 63.920000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 86.895000 63.920000 87.215000 ;
      LAYER met4 ;
        RECT 63.600000 86.895000 63.920000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 87.305000 63.920000 87.625000 ;
      LAYER met4 ;
        RECT 63.600000 87.305000 63.920000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 87.715000 63.920000 88.035000 ;
      LAYER met4 ;
        RECT 63.600000 87.715000 63.920000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 88.125000 63.920000 88.445000 ;
      LAYER met4 ;
        RECT 63.600000 88.125000 63.920000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 88.535000 63.920000 88.855000 ;
      LAYER met4 ;
        RECT 63.600000 88.535000 63.920000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 88.945000 63.920000 89.265000 ;
      LAYER met4 ;
        RECT 63.600000 88.945000 63.920000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 89.355000 63.920000 89.675000 ;
      LAYER met4 ;
        RECT 63.600000 89.355000 63.920000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 89.765000 63.920000 90.085000 ;
      LAYER met4 ;
        RECT 63.600000 89.765000 63.920000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 90.175000 63.920000 90.495000 ;
      LAYER met4 ;
        RECT 63.600000 90.175000 63.920000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 90.585000 63.920000 90.905000 ;
      LAYER met4 ;
        RECT 63.600000 90.585000 63.920000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 90.995000 63.920000 91.315000 ;
      LAYER met4 ;
        RECT 63.600000 90.995000 63.920000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 91.405000 63.920000 91.725000 ;
      LAYER met4 ;
        RECT 63.600000 91.405000 63.920000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 91.815000 63.920000 92.135000 ;
      LAYER met4 ;
        RECT 63.600000 91.815000 63.920000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 92.225000 63.920000 92.545000 ;
      LAYER met4 ;
        RECT 63.600000 92.225000 63.920000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600000 92.635000 63.920000 92.955000 ;
      LAYER met4 ;
        RECT 63.600000 92.635000 63.920000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.745000 17.800000 64.065000 18.120000 ;
      LAYER met4 ;
        RECT 63.745000 17.800000 64.065000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.745000 18.230000 64.065000 18.550000 ;
      LAYER met4 ;
        RECT 63.745000 18.230000 64.065000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.745000 18.660000 64.065000 18.980000 ;
      LAYER met4 ;
        RECT 63.745000 18.660000 64.065000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.745000 19.090000 64.065000 19.410000 ;
      LAYER met4 ;
        RECT 63.745000 19.090000 64.065000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.745000 19.520000 64.065000 19.840000 ;
      LAYER met4 ;
        RECT 63.745000 19.520000 64.065000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.745000 19.950000 64.065000 20.270000 ;
      LAYER met4 ;
        RECT 63.745000 19.950000 64.065000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.745000 20.380000 64.065000 20.700000 ;
      LAYER met4 ;
        RECT 63.745000 20.380000 64.065000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.745000 20.810000 64.065000 21.130000 ;
      LAYER met4 ;
        RECT 63.745000 20.810000 64.065000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.745000 21.240000 64.065000 21.560000 ;
      LAYER met4 ;
        RECT 63.745000 21.240000 64.065000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.745000 21.670000 64.065000 21.990000 ;
      LAYER met4 ;
        RECT 63.745000 21.670000 64.065000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.745000 22.100000 64.065000 22.420000 ;
      LAYER met4 ;
        RECT 63.745000 22.100000 64.065000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 68.065000 64.070000 68.385000 ;
      LAYER met4 ;
        RECT 63.750000 68.065000 64.070000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 68.475000 64.070000 68.795000 ;
      LAYER met4 ;
        RECT 63.750000 68.475000 64.070000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 68.885000 64.070000 69.205000 ;
      LAYER met4 ;
        RECT 63.750000 68.885000 64.070000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 69.295000 64.070000 69.615000 ;
      LAYER met4 ;
        RECT 63.750000 69.295000 64.070000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 69.705000 64.070000 70.025000 ;
      LAYER met4 ;
        RECT 63.750000 69.705000 64.070000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 70.115000 64.070000 70.435000 ;
      LAYER met4 ;
        RECT 63.750000 70.115000 64.070000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 70.525000 64.070000 70.845000 ;
      LAYER met4 ;
        RECT 63.750000 70.525000 64.070000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 70.935000 64.070000 71.255000 ;
      LAYER met4 ;
        RECT 63.750000 70.935000 64.070000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 71.345000 64.070000 71.665000 ;
      LAYER met4 ;
        RECT 63.750000 71.345000 64.070000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 71.755000 64.070000 72.075000 ;
      LAYER met4 ;
        RECT 63.750000 71.755000 64.070000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 72.165000 64.070000 72.485000 ;
      LAYER met4 ;
        RECT 63.750000 72.165000 64.070000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 72.575000 64.070000 72.895000 ;
      LAYER met4 ;
        RECT 63.750000 72.575000 64.070000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 72.985000 64.070000 73.305000 ;
      LAYER met4 ;
        RECT 63.750000 72.985000 64.070000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 73.390000 64.070000 73.710000 ;
      LAYER met4 ;
        RECT 63.750000 73.390000 64.070000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 73.795000 64.070000 74.115000 ;
      LAYER met4 ;
        RECT 63.750000 73.795000 64.070000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 74.200000 64.070000 74.520000 ;
      LAYER met4 ;
        RECT 63.750000 74.200000 64.070000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 74.605000 64.070000 74.925000 ;
      LAYER met4 ;
        RECT 63.750000 74.605000 64.070000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 75.010000 64.070000 75.330000 ;
      LAYER met4 ;
        RECT 63.750000 75.010000 64.070000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 75.415000 64.070000 75.735000 ;
      LAYER met4 ;
        RECT 63.750000 75.415000 64.070000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 75.820000 64.070000 76.140000 ;
      LAYER met4 ;
        RECT 63.750000 75.820000 64.070000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 76.225000 64.070000 76.545000 ;
      LAYER met4 ;
        RECT 63.750000 76.225000 64.070000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 76.630000 64.070000 76.950000 ;
      LAYER met4 ;
        RECT 63.750000 76.630000 64.070000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 77.035000 64.070000 77.355000 ;
      LAYER met4 ;
        RECT 63.750000 77.035000 64.070000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 77.440000 64.070000 77.760000 ;
      LAYER met4 ;
        RECT 63.750000 77.440000 64.070000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 77.845000 64.070000 78.165000 ;
      LAYER met4 ;
        RECT 63.750000 77.845000 64.070000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 78.250000 64.070000 78.570000 ;
      LAYER met4 ;
        RECT 63.750000 78.250000 64.070000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 78.655000 64.070000 78.975000 ;
      LAYER met4 ;
        RECT 63.750000 78.655000 64.070000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 79.060000 64.070000 79.380000 ;
      LAYER met4 ;
        RECT 63.750000 79.060000 64.070000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 79.465000 64.070000 79.785000 ;
      LAYER met4 ;
        RECT 63.750000 79.465000 64.070000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 79.870000 64.070000 80.190000 ;
      LAYER met4 ;
        RECT 63.750000 79.870000 64.070000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 80.275000 64.070000 80.595000 ;
      LAYER met4 ;
        RECT 63.750000 80.275000 64.070000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 80.680000 64.070000 81.000000 ;
      LAYER met4 ;
        RECT 63.750000 80.680000 64.070000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 81.085000 64.070000 81.405000 ;
      LAYER met4 ;
        RECT 63.750000 81.085000 64.070000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 81.490000 64.070000 81.810000 ;
      LAYER met4 ;
        RECT 63.750000 81.490000 64.070000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 81.895000 64.070000 82.215000 ;
      LAYER met4 ;
        RECT 63.750000 81.895000 64.070000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.750000 82.300000 64.070000 82.620000 ;
      LAYER met4 ;
        RECT 63.750000 82.300000 64.070000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 82.795000 64.330000 83.115000 ;
      LAYER met4 ;
        RECT 64.010000 82.795000 64.330000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 83.205000 64.330000 83.525000 ;
      LAYER met4 ;
        RECT 64.010000 83.205000 64.330000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 83.615000 64.330000 83.935000 ;
      LAYER met4 ;
        RECT 64.010000 83.615000 64.330000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 84.025000 64.330000 84.345000 ;
      LAYER met4 ;
        RECT 64.010000 84.025000 64.330000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 84.435000 64.330000 84.755000 ;
      LAYER met4 ;
        RECT 64.010000 84.435000 64.330000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 84.845000 64.330000 85.165000 ;
      LAYER met4 ;
        RECT 64.010000 84.845000 64.330000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 85.255000 64.330000 85.575000 ;
      LAYER met4 ;
        RECT 64.010000 85.255000 64.330000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 85.665000 64.330000 85.985000 ;
      LAYER met4 ;
        RECT 64.010000 85.665000 64.330000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 86.075000 64.330000 86.395000 ;
      LAYER met4 ;
        RECT 64.010000 86.075000 64.330000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 86.485000 64.330000 86.805000 ;
      LAYER met4 ;
        RECT 64.010000 86.485000 64.330000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 86.895000 64.330000 87.215000 ;
      LAYER met4 ;
        RECT 64.010000 86.895000 64.330000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 87.305000 64.330000 87.625000 ;
      LAYER met4 ;
        RECT 64.010000 87.305000 64.330000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 87.715000 64.330000 88.035000 ;
      LAYER met4 ;
        RECT 64.010000 87.715000 64.330000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 88.125000 64.330000 88.445000 ;
      LAYER met4 ;
        RECT 64.010000 88.125000 64.330000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 88.535000 64.330000 88.855000 ;
      LAYER met4 ;
        RECT 64.010000 88.535000 64.330000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 88.945000 64.330000 89.265000 ;
      LAYER met4 ;
        RECT 64.010000 88.945000 64.330000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 89.355000 64.330000 89.675000 ;
      LAYER met4 ;
        RECT 64.010000 89.355000 64.330000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 89.765000 64.330000 90.085000 ;
      LAYER met4 ;
        RECT 64.010000 89.765000 64.330000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 90.175000 64.330000 90.495000 ;
      LAYER met4 ;
        RECT 64.010000 90.175000 64.330000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 90.585000 64.330000 90.905000 ;
      LAYER met4 ;
        RECT 64.010000 90.585000 64.330000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 90.995000 64.330000 91.315000 ;
      LAYER met4 ;
        RECT 64.010000 90.995000 64.330000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 91.405000 64.330000 91.725000 ;
      LAYER met4 ;
        RECT 64.010000 91.405000 64.330000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 91.815000 64.330000 92.135000 ;
      LAYER met4 ;
        RECT 64.010000 91.815000 64.330000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 92.225000 64.330000 92.545000 ;
      LAYER met4 ;
        RECT 64.010000 92.225000 64.330000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010000 92.635000 64.330000 92.955000 ;
      LAYER met4 ;
        RECT 64.010000 92.635000 64.330000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 17.800000 64.470000 18.120000 ;
      LAYER met4 ;
        RECT 64.150000 17.800000 64.470000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 18.230000 64.470000 18.550000 ;
      LAYER met4 ;
        RECT 64.150000 18.230000 64.470000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 18.660000 64.470000 18.980000 ;
      LAYER met4 ;
        RECT 64.150000 18.660000 64.470000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 19.090000 64.470000 19.410000 ;
      LAYER met4 ;
        RECT 64.150000 19.090000 64.470000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 19.520000 64.470000 19.840000 ;
      LAYER met4 ;
        RECT 64.150000 19.520000 64.470000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 19.950000 64.470000 20.270000 ;
      LAYER met4 ;
        RECT 64.150000 19.950000 64.470000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 20.380000 64.470000 20.700000 ;
      LAYER met4 ;
        RECT 64.150000 20.380000 64.470000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 20.810000 64.470000 21.130000 ;
      LAYER met4 ;
        RECT 64.150000 20.810000 64.470000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 21.240000 64.470000 21.560000 ;
      LAYER met4 ;
        RECT 64.150000 21.240000 64.470000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 21.670000 64.470000 21.990000 ;
      LAYER met4 ;
        RECT 64.150000 21.670000 64.470000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 22.100000 64.470000 22.420000 ;
      LAYER met4 ;
        RECT 64.150000 22.100000 64.470000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 68.065000 64.470000 68.385000 ;
      LAYER met4 ;
        RECT 64.150000 68.065000 64.470000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 68.475000 64.470000 68.795000 ;
      LAYER met4 ;
        RECT 64.150000 68.475000 64.470000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 68.885000 64.470000 69.205000 ;
      LAYER met4 ;
        RECT 64.150000 68.885000 64.470000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 69.295000 64.470000 69.615000 ;
      LAYER met4 ;
        RECT 64.150000 69.295000 64.470000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 69.705000 64.470000 70.025000 ;
      LAYER met4 ;
        RECT 64.150000 69.705000 64.470000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 70.115000 64.470000 70.435000 ;
      LAYER met4 ;
        RECT 64.150000 70.115000 64.470000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 70.525000 64.470000 70.845000 ;
      LAYER met4 ;
        RECT 64.150000 70.525000 64.470000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 70.935000 64.470000 71.255000 ;
      LAYER met4 ;
        RECT 64.150000 70.935000 64.470000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 71.345000 64.470000 71.665000 ;
      LAYER met4 ;
        RECT 64.150000 71.345000 64.470000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 71.755000 64.470000 72.075000 ;
      LAYER met4 ;
        RECT 64.150000 71.755000 64.470000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 72.165000 64.470000 72.485000 ;
      LAYER met4 ;
        RECT 64.150000 72.165000 64.470000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 72.575000 64.470000 72.895000 ;
      LAYER met4 ;
        RECT 64.150000 72.575000 64.470000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 72.985000 64.470000 73.305000 ;
      LAYER met4 ;
        RECT 64.150000 72.985000 64.470000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 73.390000 64.470000 73.710000 ;
      LAYER met4 ;
        RECT 64.150000 73.390000 64.470000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 73.795000 64.470000 74.115000 ;
      LAYER met4 ;
        RECT 64.150000 73.795000 64.470000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 74.200000 64.470000 74.520000 ;
      LAYER met4 ;
        RECT 64.150000 74.200000 64.470000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 74.605000 64.470000 74.925000 ;
      LAYER met4 ;
        RECT 64.150000 74.605000 64.470000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 75.010000 64.470000 75.330000 ;
      LAYER met4 ;
        RECT 64.150000 75.010000 64.470000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 75.415000 64.470000 75.735000 ;
      LAYER met4 ;
        RECT 64.150000 75.415000 64.470000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 75.820000 64.470000 76.140000 ;
      LAYER met4 ;
        RECT 64.150000 75.820000 64.470000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 76.225000 64.470000 76.545000 ;
      LAYER met4 ;
        RECT 64.150000 76.225000 64.470000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 76.630000 64.470000 76.950000 ;
      LAYER met4 ;
        RECT 64.150000 76.630000 64.470000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 77.035000 64.470000 77.355000 ;
      LAYER met4 ;
        RECT 64.150000 77.035000 64.470000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 77.440000 64.470000 77.760000 ;
      LAYER met4 ;
        RECT 64.150000 77.440000 64.470000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 77.845000 64.470000 78.165000 ;
      LAYER met4 ;
        RECT 64.150000 77.845000 64.470000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 78.250000 64.470000 78.570000 ;
      LAYER met4 ;
        RECT 64.150000 78.250000 64.470000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 78.655000 64.470000 78.975000 ;
      LAYER met4 ;
        RECT 64.150000 78.655000 64.470000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 79.060000 64.470000 79.380000 ;
      LAYER met4 ;
        RECT 64.150000 79.060000 64.470000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 79.465000 64.470000 79.785000 ;
      LAYER met4 ;
        RECT 64.150000 79.465000 64.470000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 79.870000 64.470000 80.190000 ;
      LAYER met4 ;
        RECT 64.150000 79.870000 64.470000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 80.275000 64.470000 80.595000 ;
      LAYER met4 ;
        RECT 64.150000 80.275000 64.470000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 80.680000 64.470000 81.000000 ;
      LAYER met4 ;
        RECT 64.150000 80.680000 64.470000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 81.085000 64.470000 81.405000 ;
      LAYER met4 ;
        RECT 64.150000 81.085000 64.470000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 81.490000 64.470000 81.810000 ;
      LAYER met4 ;
        RECT 64.150000 81.490000 64.470000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 81.895000 64.470000 82.215000 ;
      LAYER met4 ;
        RECT 64.150000 81.895000 64.470000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 82.300000 64.470000 82.620000 ;
      LAYER met4 ;
        RECT 64.150000 82.300000 64.470000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 82.795000 64.740000 83.115000 ;
      LAYER met4 ;
        RECT 64.420000 82.795000 64.740000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 83.205000 64.740000 83.525000 ;
      LAYER met4 ;
        RECT 64.420000 83.205000 64.740000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 83.615000 64.740000 83.935000 ;
      LAYER met4 ;
        RECT 64.420000 83.615000 64.740000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 84.025000 64.740000 84.345000 ;
      LAYER met4 ;
        RECT 64.420000 84.025000 64.740000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 84.435000 64.740000 84.755000 ;
      LAYER met4 ;
        RECT 64.420000 84.435000 64.740000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 84.845000 64.740000 85.165000 ;
      LAYER met4 ;
        RECT 64.420000 84.845000 64.740000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 85.255000 64.740000 85.575000 ;
      LAYER met4 ;
        RECT 64.420000 85.255000 64.740000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 85.665000 64.740000 85.985000 ;
      LAYER met4 ;
        RECT 64.420000 85.665000 64.740000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 86.075000 64.740000 86.395000 ;
      LAYER met4 ;
        RECT 64.420000 86.075000 64.740000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 86.485000 64.740000 86.805000 ;
      LAYER met4 ;
        RECT 64.420000 86.485000 64.740000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 86.895000 64.740000 87.215000 ;
      LAYER met4 ;
        RECT 64.420000 86.895000 64.740000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 87.305000 64.740000 87.625000 ;
      LAYER met4 ;
        RECT 64.420000 87.305000 64.740000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 87.715000 64.740000 88.035000 ;
      LAYER met4 ;
        RECT 64.420000 87.715000 64.740000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 88.125000 64.740000 88.445000 ;
      LAYER met4 ;
        RECT 64.420000 88.125000 64.740000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 88.535000 64.740000 88.855000 ;
      LAYER met4 ;
        RECT 64.420000 88.535000 64.740000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 88.945000 64.740000 89.265000 ;
      LAYER met4 ;
        RECT 64.420000 88.945000 64.740000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 89.355000 64.740000 89.675000 ;
      LAYER met4 ;
        RECT 64.420000 89.355000 64.740000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 89.765000 64.740000 90.085000 ;
      LAYER met4 ;
        RECT 64.420000 89.765000 64.740000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 90.175000 64.740000 90.495000 ;
      LAYER met4 ;
        RECT 64.420000 90.175000 64.740000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 90.585000 64.740000 90.905000 ;
      LAYER met4 ;
        RECT 64.420000 90.585000 64.740000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 90.995000 64.740000 91.315000 ;
      LAYER met4 ;
        RECT 64.420000 90.995000 64.740000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 91.405000 64.740000 91.725000 ;
      LAYER met4 ;
        RECT 64.420000 91.405000 64.740000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 91.815000 64.740000 92.135000 ;
      LAYER met4 ;
        RECT 64.420000 91.815000 64.740000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 92.225000 64.740000 92.545000 ;
      LAYER met4 ;
        RECT 64.420000 92.225000 64.740000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420000 92.635000 64.740000 92.955000 ;
      LAYER met4 ;
        RECT 64.420000 92.635000 64.740000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 68.065000 64.870000 68.385000 ;
      LAYER met4 ;
        RECT 64.550000 68.065000 64.870000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 68.475000 64.870000 68.795000 ;
      LAYER met4 ;
        RECT 64.550000 68.475000 64.870000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 68.885000 64.870000 69.205000 ;
      LAYER met4 ;
        RECT 64.550000 68.885000 64.870000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 69.295000 64.870000 69.615000 ;
      LAYER met4 ;
        RECT 64.550000 69.295000 64.870000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 69.705000 64.870000 70.025000 ;
      LAYER met4 ;
        RECT 64.550000 69.705000 64.870000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 70.115000 64.870000 70.435000 ;
      LAYER met4 ;
        RECT 64.550000 70.115000 64.870000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 70.525000 64.870000 70.845000 ;
      LAYER met4 ;
        RECT 64.550000 70.525000 64.870000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 70.935000 64.870000 71.255000 ;
      LAYER met4 ;
        RECT 64.550000 70.935000 64.870000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 71.345000 64.870000 71.665000 ;
      LAYER met4 ;
        RECT 64.550000 71.345000 64.870000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 71.755000 64.870000 72.075000 ;
      LAYER met4 ;
        RECT 64.550000 71.755000 64.870000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 72.165000 64.870000 72.485000 ;
      LAYER met4 ;
        RECT 64.550000 72.165000 64.870000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 72.575000 64.870000 72.895000 ;
      LAYER met4 ;
        RECT 64.550000 72.575000 64.870000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 72.985000 64.870000 73.305000 ;
      LAYER met4 ;
        RECT 64.550000 72.985000 64.870000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 73.390000 64.870000 73.710000 ;
      LAYER met4 ;
        RECT 64.550000 73.390000 64.870000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 73.795000 64.870000 74.115000 ;
      LAYER met4 ;
        RECT 64.550000 73.795000 64.870000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 74.200000 64.870000 74.520000 ;
      LAYER met4 ;
        RECT 64.550000 74.200000 64.870000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 74.605000 64.870000 74.925000 ;
      LAYER met4 ;
        RECT 64.550000 74.605000 64.870000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 75.010000 64.870000 75.330000 ;
      LAYER met4 ;
        RECT 64.550000 75.010000 64.870000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 75.415000 64.870000 75.735000 ;
      LAYER met4 ;
        RECT 64.550000 75.415000 64.870000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 75.820000 64.870000 76.140000 ;
      LAYER met4 ;
        RECT 64.550000 75.820000 64.870000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 76.225000 64.870000 76.545000 ;
      LAYER met4 ;
        RECT 64.550000 76.225000 64.870000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 76.630000 64.870000 76.950000 ;
      LAYER met4 ;
        RECT 64.550000 76.630000 64.870000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 77.035000 64.870000 77.355000 ;
      LAYER met4 ;
        RECT 64.550000 77.035000 64.870000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 77.440000 64.870000 77.760000 ;
      LAYER met4 ;
        RECT 64.550000 77.440000 64.870000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 77.845000 64.870000 78.165000 ;
      LAYER met4 ;
        RECT 64.550000 77.845000 64.870000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 78.250000 64.870000 78.570000 ;
      LAYER met4 ;
        RECT 64.550000 78.250000 64.870000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 78.655000 64.870000 78.975000 ;
      LAYER met4 ;
        RECT 64.550000 78.655000 64.870000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 79.060000 64.870000 79.380000 ;
      LAYER met4 ;
        RECT 64.550000 79.060000 64.870000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 79.465000 64.870000 79.785000 ;
      LAYER met4 ;
        RECT 64.550000 79.465000 64.870000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 79.870000 64.870000 80.190000 ;
      LAYER met4 ;
        RECT 64.550000 79.870000 64.870000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 80.275000 64.870000 80.595000 ;
      LAYER met4 ;
        RECT 64.550000 80.275000 64.870000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 80.680000 64.870000 81.000000 ;
      LAYER met4 ;
        RECT 64.550000 80.680000 64.870000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 81.085000 64.870000 81.405000 ;
      LAYER met4 ;
        RECT 64.550000 81.085000 64.870000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 81.490000 64.870000 81.810000 ;
      LAYER met4 ;
        RECT 64.550000 81.490000 64.870000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 81.895000 64.870000 82.215000 ;
      LAYER met4 ;
        RECT 64.550000 81.895000 64.870000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.550000 82.300000 64.870000 82.620000 ;
      LAYER met4 ;
        RECT 64.550000 82.300000 64.870000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.555000 17.800000 64.875000 18.120000 ;
      LAYER met4 ;
        RECT 64.555000 17.800000 64.875000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.555000 18.230000 64.875000 18.550000 ;
      LAYER met4 ;
        RECT 64.555000 18.230000 64.875000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.555000 18.660000 64.875000 18.980000 ;
      LAYER met4 ;
        RECT 64.555000 18.660000 64.875000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.555000 19.090000 64.875000 19.410000 ;
      LAYER met4 ;
        RECT 64.555000 19.090000 64.875000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.555000 19.520000 64.875000 19.840000 ;
      LAYER met4 ;
        RECT 64.555000 19.520000 64.875000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.555000 19.950000 64.875000 20.270000 ;
      LAYER met4 ;
        RECT 64.555000 19.950000 64.875000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.555000 20.380000 64.875000 20.700000 ;
      LAYER met4 ;
        RECT 64.555000 20.380000 64.875000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.555000 20.810000 64.875000 21.130000 ;
      LAYER met4 ;
        RECT 64.555000 20.810000 64.875000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.555000 21.240000 64.875000 21.560000 ;
      LAYER met4 ;
        RECT 64.555000 21.240000 64.875000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.555000 21.670000 64.875000 21.990000 ;
      LAYER met4 ;
        RECT 64.555000 21.670000 64.875000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.555000 22.100000 64.875000 22.420000 ;
      LAYER met4 ;
        RECT 64.555000 22.100000 64.875000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 82.795000 65.150000 83.115000 ;
      LAYER met4 ;
        RECT 64.830000 82.795000 65.150000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 83.205000 65.150000 83.525000 ;
      LAYER met4 ;
        RECT 64.830000 83.205000 65.150000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 83.615000 65.150000 83.935000 ;
      LAYER met4 ;
        RECT 64.830000 83.615000 65.150000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 84.025000 65.150000 84.345000 ;
      LAYER met4 ;
        RECT 64.830000 84.025000 65.150000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 84.435000 65.150000 84.755000 ;
      LAYER met4 ;
        RECT 64.830000 84.435000 65.150000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 84.845000 65.150000 85.165000 ;
      LAYER met4 ;
        RECT 64.830000 84.845000 65.150000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 85.255000 65.150000 85.575000 ;
      LAYER met4 ;
        RECT 64.830000 85.255000 65.150000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 85.665000 65.150000 85.985000 ;
      LAYER met4 ;
        RECT 64.830000 85.665000 65.150000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 86.075000 65.150000 86.395000 ;
      LAYER met4 ;
        RECT 64.830000 86.075000 65.150000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 86.485000 65.150000 86.805000 ;
      LAYER met4 ;
        RECT 64.830000 86.485000 65.150000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 86.895000 65.150000 87.215000 ;
      LAYER met4 ;
        RECT 64.830000 86.895000 65.150000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 87.305000 65.150000 87.625000 ;
      LAYER met4 ;
        RECT 64.830000 87.305000 65.150000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 87.715000 65.150000 88.035000 ;
      LAYER met4 ;
        RECT 64.830000 87.715000 65.150000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 88.125000 65.150000 88.445000 ;
      LAYER met4 ;
        RECT 64.830000 88.125000 65.150000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 88.535000 65.150000 88.855000 ;
      LAYER met4 ;
        RECT 64.830000 88.535000 65.150000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 88.945000 65.150000 89.265000 ;
      LAYER met4 ;
        RECT 64.830000 88.945000 65.150000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 89.355000 65.150000 89.675000 ;
      LAYER met4 ;
        RECT 64.830000 89.355000 65.150000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 89.765000 65.150000 90.085000 ;
      LAYER met4 ;
        RECT 64.830000 89.765000 65.150000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 90.175000 65.150000 90.495000 ;
      LAYER met4 ;
        RECT 64.830000 90.175000 65.150000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 90.585000 65.150000 90.905000 ;
      LAYER met4 ;
        RECT 64.830000 90.585000 65.150000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 90.995000 65.150000 91.315000 ;
      LAYER met4 ;
        RECT 64.830000 90.995000 65.150000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 91.405000 65.150000 91.725000 ;
      LAYER met4 ;
        RECT 64.830000 91.405000 65.150000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 91.815000 65.150000 92.135000 ;
      LAYER met4 ;
        RECT 64.830000 91.815000 65.150000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 92.225000 65.150000 92.545000 ;
      LAYER met4 ;
        RECT 64.830000 92.225000 65.150000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830000 92.635000 65.150000 92.955000 ;
      LAYER met4 ;
        RECT 64.830000 92.635000 65.150000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 68.065000 65.270000 68.385000 ;
      LAYER met4 ;
        RECT 64.950000 68.065000 65.270000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 68.475000 65.270000 68.795000 ;
      LAYER met4 ;
        RECT 64.950000 68.475000 65.270000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 68.885000 65.270000 69.205000 ;
      LAYER met4 ;
        RECT 64.950000 68.885000 65.270000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 69.295000 65.270000 69.615000 ;
      LAYER met4 ;
        RECT 64.950000 69.295000 65.270000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 69.705000 65.270000 70.025000 ;
      LAYER met4 ;
        RECT 64.950000 69.705000 65.270000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 70.115000 65.270000 70.435000 ;
      LAYER met4 ;
        RECT 64.950000 70.115000 65.270000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 70.525000 65.270000 70.845000 ;
      LAYER met4 ;
        RECT 64.950000 70.525000 65.270000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 70.935000 65.270000 71.255000 ;
      LAYER met4 ;
        RECT 64.950000 70.935000 65.270000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 71.345000 65.270000 71.665000 ;
      LAYER met4 ;
        RECT 64.950000 71.345000 65.270000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 71.755000 65.270000 72.075000 ;
      LAYER met4 ;
        RECT 64.950000 71.755000 65.270000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 72.165000 65.270000 72.485000 ;
      LAYER met4 ;
        RECT 64.950000 72.165000 65.270000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 72.575000 65.270000 72.895000 ;
      LAYER met4 ;
        RECT 64.950000 72.575000 65.270000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 72.985000 65.270000 73.305000 ;
      LAYER met4 ;
        RECT 64.950000 72.985000 65.270000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 73.390000 65.270000 73.710000 ;
      LAYER met4 ;
        RECT 64.950000 73.390000 65.270000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 73.795000 65.270000 74.115000 ;
      LAYER met4 ;
        RECT 64.950000 73.795000 65.270000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 74.200000 65.270000 74.520000 ;
      LAYER met4 ;
        RECT 64.950000 74.200000 65.270000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 74.605000 65.270000 74.925000 ;
      LAYER met4 ;
        RECT 64.950000 74.605000 65.270000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 75.010000 65.270000 75.330000 ;
      LAYER met4 ;
        RECT 64.950000 75.010000 65.270000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 75.415000 65.270000 75.735000 ;
      LAYER met4 ;
        RECT 64.950000 75.415000 65.270000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 75.820000 65.270000 76.140000 ;
      LAYER met4 ;
        RECT 64.950000 75.820000 65.270000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 76.225000 65.270000 76.545000 ;
      LAYER met4 ;
        RECT 64.950000 76.225000 65.270000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 76.630000 65.270000 76.950000 ;
      LAYER met4 ;
        RECT 64.950000 76.630000 65.270000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 77.035000 65.270000 77.355000 ;
      LAYER met4 ;
        RECT 64.950000 77.035000 65.270000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 77.440000 65.270000 77.760000 ;
      LAYER met4 ;
        RECT 64.950000 77.440000 65.270000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 77.845000 65.270000 78.165000 ;
      LAYER met4 ;
        RECT 64.950000 77.845000 65.270000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 78.250000 65.270000 78.570000 ;
      LAYER met4 ;
        RECT 64.950000 78.250000 65.270000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 78.655000 65.270000 78.975000 ;
      LAYER met4 ;
        RECT 64.950000 78.655000 65.270000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 79.060000 65.270000 79.380000 ;
      LAYER met4 ;
        RECT 64.950000 79.060000 65.270000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 79.465000 65.270000 79.785000 ;
      LAYER met4 ;
        RECT 64.950000 79.465000 65.270000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 79.870000 65.270000 80.190000 ;
      LAYER met4 ;
        RECT 64.950000 79.870000 65.270000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 80.275000 65.270000 80.595000 ;
      LAYER met4 ;
        RECT 64.950000 80.275000 65.270000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 80.680000 65.270000 81.000000 ;
      LAYER met4 ;
        RECT 64.950000 80.680000 65.270000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 81.085000 65.270000 81.405000 ;
      LAYER met4 ;
        RECT 64.950000 81.085000 65.270000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 81.490000 65.270000 81.810000 ;
      LAYER met4 ;
        RECT 64.950000 81.490000 65.270000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 81.895000 65.270000 82.215000 ;
      LAYER met4 ;
        RECT 64.950000 81.895000 65.270000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.950000 82.300000 65.270000 82.620000 ;
      LAYER met4 ;
        RECT 64.950000 82.300000 65.270000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.960000 17.800000 65.280000 18.120000 ;
      LAYER met4 ;
        RECT 64.960000 17.800000 65.280000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.960000 18.230000 65.280000 18.550000 ;
      LAYER met4 ;
        RECT 64.960000 18.230000 65.280000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.960000 18.660000 65.280000 18.980000 ;
      LAYER met4 ;
        RECT 64.960000 18.660000 65.280000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.960000 19.090000 65.280000 19.410000 ;
      LAYER met4 ;
        RECT 64.960000 19.090000 65.280000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.960000 19.520000 65.280000 19.840000 ;
      LAYER met4 ;
        RECT 64.960000 19.520000 65.280000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.960000 19.950000 65.280000 20.270000 ;
      LAYER met4 ;
        RECT 64.960000 19.950000 65.280000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.960000 20.380000 65.280000 20.700000 ;
      LAYER met4 ;
        RECT 64.960000 20.380000 65.280000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.960000 20.810000 65.280000 21.130000 ;
      LAYER met4 ;
        RECT 64.960000 20.810000 65.280000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.960000 21.240000 65.280000 21.560000 ;
      LAYER met4 ;
        RECT 64.960000 21.240000 65.280000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.960000 21.670000 65.280000 21.990000 ;
      LAYER met4 ;
        RECT 64.960000 21.670000 65.280000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.960000 22.100000 65.280000 22.420000 ;
      LAYER met4 ;
        RECT 64.960000 22.100000 65.280000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 82.795000 65.560000 83.115000 ;
      LAYER met4 ;
        RECT 65.240000 82.795000 65.560000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 83.205000 65.560000 83.525000 ;
      LAYER met4 ;
        RECT 65.240000 83.205000 65.560000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 83.615000 65.560000 83.935000 ;
      LAYER met4 ;
        RECT 65.240000 83.615000 65.560000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 84.025000 65.560000 84.345000 ;
      LAYER met4 ;
        RECT 65.240000 84.025000 65.560000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 84.435000 65.560000 84.755000 ;
      LAYER met4 ;
        RECT 65.240000 84.435000 65.560000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 84.845000 65.560000 85.165000 ;
      LAYER met4 ;
        RECT 65.240000 84.845000 65.560000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 85.255000 65.560000 85.575000 ;
      LAYER met4 ;
        RECT 65.240000 85.255000 65.560000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 85.665000 65.560000 85.985000 ;
      LAYER met4 ;
        RECT 65.240000 85.665000 65.560000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 86.075000 65.560000 86.395000 ;
      LAYER met4 ;
        RECT 65.240000 86.075000 65.560000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 86.485000 65.560000 86.805000 ;
      LAYER met4 ;
        RECT 65.240000 86.485000 65.560000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 86.895000 65.560000 87.215000 ;
      LAYER met4 ;
        RECT 65.240000 86.895000 65.560000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 87.305000 65.560000 87.625000 ;
      LAYER met4 ;
        RECT 65.240000 87.305000 65.560000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 87.715000 65.560000 88.035000 ;
      LAYER met4 ;
        RECT 65.240000 87.715000 65.560000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 88.125000 65.560000 88.445000 ;
      LAYER met4 ;
        RECT 65.240000 88.125000 65.560000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 88.535000 65.560000 88.855000 ;
      LAYER met4 ;
        RECT 65.240000 88.535000 65.560000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 88.945000 65.560000 89.265000 ;
      LAYER met4 ;
        RECT 65.240000 88.945000 65.560000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 89.355000 65.560000 89.675000 ;
      LAYER met4 ;
        RECT 65.240000 89.355000 65.560000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 89.765000 65.560000 90.085000 ;
      LAYER met4 ;
        RECT 65.240000 89.765000 65.560000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 90.175000 65.560000 90.495000 ;
      LAYER met4 ;
        RECT 65.240000 90.175000 65.560000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 90.585000 65.560000 90.905000 ;
      LAYER met4 ;
        RECT 65.240000 90.585000 65.560000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 90.995000 65.560000 91.315000 ;
      LAYER met4 ;
        RECT 65.240000 90.995000 65.560000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 91.405000 65.560000 91.725000 ;
      LAYER met4 ;
        RECT 65.240000 91.405000 65.560000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 91.815000 65.560000 92.135000 ;
      LAYER met4 ;
        RECT 65.240000 91.815000 65.560000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 92.225000 65.560000 92.545000 ;
      LAYER met4 ;
        RECT 65.240000 92.225000 65.560000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240000 92.635000 65.560000 92.955000 ;
      LAYER met4 ;
        RECT 65.240000 92.635000 65.560000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 68.065000 65.670000 68.385000 ;
      LAYER met4 ;
        RECT 65.350000 68.065000 65.670000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 68.475000 65.670000 68.795000 ;
      LAYER met4 ;
        RECT 65.350000 68.475000 65.670000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 68.885000 65.670000 69.205000 ;
      LAYER met4 ;
        RECT 65.350000 68.885000 65.670000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 69.295000 65.670000 69.615000 ;
      LAYER met4 ;
        RECT 65.350000 69.295000 65.670000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 69.705000 65.670000 70.025000 ;
      LAYER met4 ;
        RECT 65.350000 69.705000 65.670000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 70.115000 65.670000 70.435000 ;
      LAYER met4 ;
        RECT 65.350000 70.115000 65.670000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 70.525000 65.670000 70.845000 ;
      LAYER met4 ;
        RECT 65.350000 70.525000 65.670000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 70.935000 65.670000 71.255000 ;
      LAYER met4 ;
        RECT 65.350000 70.935000 65.670000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 71.345000 65.670000 71.665000 ;
      LAYER met4 ;
        RECT 65.350000 71.345000 65.670000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 71.755000 65.670000 72.075000 ;
      LAYER met4 ;
        RECT 65.350000 71.755000 65.670000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 72.165000 65.670000 72.485000 ;
      LAYER met4 ;
        RECT 65.350000 72.165000 65.670000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 72.575000 65.670000 72.895000 ;
      LAYER met4 ;
        RECT 65.350000 72.575000 65.670000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 72.985000 65.670000 73.305000 ;
      LAYER met4 ;
        RECT 65.350000 72.985000 65.670000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 73.390000 65.670000 73.710000 ;
      LAYER met4 ;
        RECT 65.350000 73.390000 65.670000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 73.795000 65.670000 74.115000 ;
      LAYER met4 ;
        RECT 65.350000 73.795000 65.670000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 74.200000 65.670000 74.520000 ;
      LAYER met4 ;
        RECT 65.350000 74.200000 65.670000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 74.605000 65.670000 74.925000 ;
      LAYER met4 ;
        RECT 65.350000 74.605000 65.670000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 75.010000 65.670000 75.330000 ;
      LAYER met4 ;
        RECT 65.350000 75.010000 65.670000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 75.415000 65.670000 75.735000 ;
      LAYER met4 ;
        RECT 65.350000 75.415000 65.670000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 75.820000 65.670000 76.140000 ;
      LAYER met4 ;
        RECT 65.350000 75.820000 65.670000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 76.225000 65.670000 76.545000 ;
      LAYER met4 ;
        RECT 65.350000 76.225000 65.670000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 76.630000 65.670000 76.950000 ;
      LAYER met4 ;
        RECT 65.350000 76.630000 65.670000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 77.035000 65.670000 77.355000 ;
      LAYER met4 ;
        RECT 65.350000 77.035000 65.670000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 77.440000 65.670000 77.760000 ;
      LAYER met4 ;
        RECT 65.350000 77.440000 65.670000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 77.845000 65.670000 78.165000 ;
      LAYER met4 ;
        RECT 65.350000 77.845000 65.670000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 78.250000 65.670000 78.570000 ;
      LAYER met4 ;
        RECT 65.350000 78.250000 65.670000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 78.655000 65.670000 78.975000 ;
      LAYER met4 ;
        RECT 65.350000 78.655000 65.670000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 79.060000 65.670000 79.380000 ;
      LAYER met4 ;
        RECT 65.350000 79.060000 65.670000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 79.465000 65.670000 79.785000 ;
      LAYER met4 ;
        RECT 65.350000 79.465000 65.670000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 79.870000 65.670000 80.190000 ;
      LAYER met4 ;
        RECT 65.350000 79.870000 65.670000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 80.275000 65.670000 80.595000 ;
      LAYER met4 ;
        RECT 65.350000 80.275000 65.670000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 80.680000 65.670000 81.000000 ;
      LAYER met4 ;
        RECT 65.350000 80.680000 65.670000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 81.085000 65.670000 81.405000 ;
      LAYER met4 ;
        RECT 65.350000 81.085000 65.670000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 81.490000 65.670000 81.810000 ;
      LAYER met4 ;
        RECT 65.350000 81.490000 65.670000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 81.895000 65.670000 82.215000 ;
      LAYER met4 ;
        RECT 65.350000 81.895000 65.670000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.350000 82.300000 65.670000 82.620000 ;
      LAYER met4 ;
        RECT 65.350000 82.300000 65.670000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.365000 17.800000 65.685000 18.120000 ;
      LAYER met4 ;
        RECT 65.365000 17.800000 65.685000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.365000 18.230000 65.685000 18.550000 ;
      LAYER met4 ;
        RECT 65.365000 18.230000 65.685000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.365000 18.660000 65.685000 18.980000 ;
      LAYER met4 ;
        RECT 65.365000 18.660000 65.685000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.365000 19.090000 65.685000 19.410000 ;
      LAYER met4 ;
        RECT 65.365000 19.090000 65.685000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.365000 19.520000 65.685000 19.840000 ;
      LAYER met4 ;
        RECT 65.365000 19.520000 65.685000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.365000 19.950000 65.685000 20.270000 ;
      LAYER met4 ;
        RECT 65.365000 19.950000 65.685000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.365000 20.380000 65.685000 20.700000 ;
      LAYER met4 ;
        RECT 65.365000 20.380000 65.685000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.365000 20.810000 65.685000 21.130000 ;
      LAYER met4 ;
        RECT 65.365000 20.810000 65.685000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.365000 21.240000 65.685000 21.560000 ;
      LAYER met4 ;
        RECT 65.365000 21.240000 65.685000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.365000 21.670000 65.685000 21.990000 ;
      LAYER met4 ;
        RECT 65.365000 21.670000 65.685000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.365000 22.100000 65.685000 22.420000 ;
      LAYER met4 ;
        RECT 65.365000 22.100000 65.685000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 82.795000 65.970000 83.115000 ;
      LAYER met4 ;
        RECT 65.650000 82.795000 65.970000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 83.205000 65.970000 83.525000 ;
      LAYER met4 ;
        RECT 65.650000 83.205000 65.970000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 83.615000 65.970000 83.935000 ;
      LAYER met4 ;
        RECT 65.650000 83.615000 65.970000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 84.025000 65.970000 84.345000 ;
      LAYER met4 ;
        RECT 65.650000 84.025000 65.970000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 84.435000 65.970000 84.755000 ;
      LAYER met4 ;
        RECT 65.650000 84.435000 65.970000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 84.845000 65.970000 85.165000 ;
      LAYER met4 ;
        RECT 65.650000 84.845000 65.970000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 85.255000 65.970000 85.575000 ;
      LAYER met4 ;
        RECT 65.650000 85.255000 65.970000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 85.665000 65.970000 85.985000 ;
      LAYER met4 ;
        RECT 65.650000 85.665000 65.970000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 86.075000 65.970000 86.395000 ;
      LAYER met4 ;
        RECT 65.650000 86.075000 65.970000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 86.485000 65.970000 86.805000 ;
      LAYER met4 ;
        RECT 65.650000 86.485000 65.970000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 86.895000 65.970000 87.215000 ;
      LAYER met4 ;
        RECT 65.650000 86.895000 65.970000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 87.305000 65.970000 87.625000 ;
      LAYER met4 ;
        RECT 65.650000 87.305000 65.970000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 87.715000 65.970000 88.035000 ;
      LAYER met4 ;
        RECT 65.650000 87.715000 65.970000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 88.125000 65.970000 88.445000 ;
      LAYER met4 ;
        RECT 65.650000 88.125000 65.970000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 88.535000 65.970000 88.855000 ;
      LAYER met4 ;
        RECT 65.650000 88.535000 65.970000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 88.945000 65.970000 89.265000 ;
      LAYER met4 ;
        RECT 65.650000 88.945000 65.970000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 89.355000 65.970000 89.675000 ;
      LAYER met4 ;
        RECT 65.650000 89.355000 65.970000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 89.765000 65.970000 90.085000 ;
      LAYER met4 ;
        RECT 65.650000 89.765000 65.970000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 90.175000 65.970000 90.495000 ;
      LAYER met4 ;
        RECT 65.650000 90.175000 65.970000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 90.585000 65.970000 90.905000 ;
      LAYER met4 ;
        RECT 65.650000 90.585000 65.970000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 90.995000 65.970000 91.315000 ;
      LAYER met4 ;
        RECT 65.650000 90.995000 65.970000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 91.405000 65.970000 91.725000 ;
      LAYER met4 ;
        RECT 65.650000 91.405000 65.970000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 91.815000 65.970000 92.135000 ;
      LAYER met4 ;
        RECT 65.650000 91.815000 65.970000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 92.225000 65.970000 92.545000 ;
      LAYER met4 ;
        RECT 65.650000 92.225000 65.970000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650000 92.635000 65.970000 92.955000 ;
      LAYER met4 ;
        RECT 65.650000 92.635000 65.970000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 68.065000 66.070000 68.385000 ;
      LAYER met4 ;
        RECT 65.750000 68.065000 66.070000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 68.475000 66.070000 68.795000 ;
      LAYER met4 ;
        RECT 65.750000 68.475000 66.070000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 68.885000 66.070000 69.205000 ;
      LAYER met4 ;
        RECT 65.750000 68.885000 66.070000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 69.295000 66.070000 69.615000 ;
      LAYER met4 ;
        RECT 65.750000 69.295000 66.070000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 69.705000 66.070000 70.025000 ;
      LAYER met4 ;
        RECT 65.750000 69.705000 66.070000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 70.115000 66.070000 70.435000 ;
      LAYER met4 ;
        RECT 65.750000 70.115000 66.070000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 70.525000 66.070000 70.845000 ;
      LAYER met4 ;
        RECT 65.750000 70.525000 66.070000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 70.935000 66.070000 71.255000 ;
      LAYER met4 ;
        RECT 65.750000 70.935000 66.070000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 71.345000 66.070000 71.665000 ;
      LAYER met4 ;
        RECT 65.750000 71.345000 66.070000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 71.755000 66.070000 72.075000 ;
      LAYER met4 ;
        RECT 65.750000 71.755000 66.070000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 72.165000 66.070000 72.485000 ;
      LAYER met4 ;
        RECT 65.750000 72.165000 66.070000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 72.575000 66.070000 72.895000 ;
      LAYER met4 ;
        RECT 65.750000 72.575000 66.070000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 72.985000 66.070000 73.305000 ;
      LAYER met4 ;
        RECT 65.750000 72.985000 66.070000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 73.390000 66.070000 73.710000 ;
      LAYER met4 ;
        RECT 65.750000 73.390000 66.070000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 73.795000 66.070000 74.115000 ;
      LAYER met4 ;
        RECT 65.750000 73.795000 66.070000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 74.200000 66.070000 74.520000 ;
      LAYER met4 ;
        RECT 65.750000 74.200000 66.070000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 74.605000 66.070000 74.925000 ;
      LAYER met4 ;
        RECT 65.750000 74.605000 66.070000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 75.010000 66.070000 75.330000 ;
      LAYER met4 ;
        RECT 65.750000 75.010000 66.070000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 75.415000 66.070000 75.735000 ;
      LAYER met4 ;
        RECT 65.750000 75.415000 66.070000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 75.820000 66.070000 76.140000 ;
      LAYER met4 ;
        RECT 65.750000 75.820000 66.070000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 76.225000 66.070000 76.545000 ;
      LAYER met4 ;
        RECT 65.750000 76.225000 66.070000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 76.630000 66.070000 76.950000 ;
      LAYER met4 ;
        RECT 65.750000 76.630000 66.070000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 77.035000 66.070000 77.355000 ;
      LAYER met4 ;
        RECT 65.750000 77.035000 66.070000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 77.440000 66.070000 77.760000 ;
      LAYER met4 ;
        RECT 65.750000 77.440000 66.070000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 77.845000 66.070000 78.165000 ;
      LAYER met4 ;
        RECT 65.750000 77.845000 66.070000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 78.250000 66.070000 78.570000 ;
      LAYER met4 ;
        RECT 65.750000 78.250000 66.070000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 78.655000 66.070000 78.975000 ;
      LAYER met4 ;
        RECT 65.750000 78.655000 66.070000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 79.060000 66.070000 79.380000 ;
      LAYER met4 ;
        RECT 65.750000 79.060000 66.070000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 79.465000 66.070000 79.785000 ;
      LAYER met4 ;
        RECT 65.750000 79.465000 66.070000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 79.870000 66.070000 80.190000 ;
      LAYER met4 ;
        RECT 65.750000 79.870000 66.070000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 80.275000 66.070000 80.595000 ;
      LAYER met4 ;
        RECT 65.750000 80.275000 66.070000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 80.680000 66.070000 81.000000 ;
      LAYER met4 ;
        RECT 65.750000 80.680000 66.070000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 81.085000 66.070000 81.405000 ;
      LAYER met4 ;
        RECT 65.750000 81.085000 66.070000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 81.490000 66.070000 81.810000 ;
      LAYER met4 ;
        RECT 65.750000 81.490000 66.070000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 81.895000 66.070000 82.215000 ;
      LAYER met4 ;
        RECT 65.750000 81.895000 66.070000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.750000 82.300000 66.070000 82.620000 ;
      LAYER met4 ;
        RECT 65.750000 82.300000 66.070000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 17.800000 66.090000 18.120000 ;
      LAYER met4 ;
        RECT 65.770000 17.800000 66.090000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 18.230000 66.090000 18.550000 ;
      LAYER met4 ;
        RECT 65.770000 18.230000 66.090000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 18.660000 66.090000 18.980000 ;
      LAYER met4 ;
        RECT 65.770000 18.660000 66.090000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 19.090000 66.090000 19.410000 ;
      LAYER met4 ;
        RECT 65.770000 19.090000 66.090000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 19.520000 66.090000 19.840000 ;
      LAYER met4 ;
        RECT 65.770000 19.520000 66.090000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 19.950000 66.090000 20.270000 ;
      LAYER met4 ;
        RECT 65.770000 19.950000 66.090000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 20.380000 66.090000 20.700000 ;
      LAYER met4 ;
        RECT 65.770000 20.380000 66.090000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 20.810000 66.090000 21.130000 ;
      LAYER met4 ;
        RECT 65.770000 20.810000 66.090000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 21.240000 66.090000 21.560000 ;
      LAYER met4 ;
        RECT 65.770000 21.240000 66.090000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 21.670000 66.090000 21.990000 ;
      LAYER met4 ;
        RECT 65.770000 21.670000 66.090000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 22.100000 66.090000 22.420000 ;
      LAYER met4 ;
        RECT 65.770000 22.100000 66.090000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 82.795000 66.380000 83.115000 ;
      LAYER met4 ;
        RECT 66.060000 82.795000 66.380000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 83.205000 66.380000 83.525000 ;
      LAYER met4 ;
        RECT 66.060000 83.205000 66.380000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 83.615000 66.380000 83.935000 ;
      LAYER met4 ;
        RECT 66.060000 83.615000 66.380000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 84.025000 66.380000 84.345000 ;
      LAYER met4 ;
        RECT 66.060000 84.025000 66.380000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 84.435000 66.380000 84.755000 ;
      LAYER met4 ;
        RECT 66.060000 84.435000 66.380000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 84.845000 66.380000 85.165000 ;
      LAYER met4 ;
        RECT 66.060000 84.845000 66.380000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 85.255000 66.380000 85.575000 ;
      LAYER met4 ;
        RECT 66.060000 85.255000 66.380000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 85.665000 66.380000 85.985000 ;
      LAYER met4 ;
        RECT 66.060000 85.665000 66.380000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 86.075000 66.380000 86.395000 ;
      LAYER met4 ;
        RECT 66.060000 86.075000 66.380000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 86.485000 66.380000 86.805000 ;
      LAYER met4 ;
        RECT 66.060000 86.485000 66.380000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 86.895000 66.380000 87.215000 ;
      LAYER met4 ;
        RECT 66.060000 86.895000 66.380000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 87.305000 66.380000 87.625000 ;
      LAYER met4 ;
        RECT 66.060000 87.305000 66.380000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 87.715000 66.380000 88.035000 ;
      LAYER met4 ;
        RECT 66.060000 87.715000 66.380000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 88.125000 66.380000 88.445000 ;
      LAYER met4 ;
        RECT 66.060000 88.125000 66.380000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 88.535000 66.380000 88.855000 ;
      LAYER met4 ;
        RECT 66.060000 88.535000 66.380000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 88.945000 66.380000 89.265000 ;
      LAYER met4 ;
        RECT 66.060000 88.945000 66.380000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 89.355000 66.380000 89.675000 ;
      LAYER met4 ;
        RECT 66.060000 89.355000 66.380000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 89.765000 66.380000 90.085000 ;
      LAYER met4 ;
        RECT 66.060000 89.765000 66.380000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 90.175000 66.380000 90.495000 ;
      LAYER met4 ;
        RECT 66.060000 90.175000 66.380000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 90.585000 66.380000 90.905000 ;
      LAYER met4 ;
        RECT 66.060000 90.585000 66.380000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 90.995000 66.380000 91.315000 ;
      LAYER met4 ;
        RECT 66.060000 90.995000 66.380000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 91.405000 66.380000 91.725000 ;
      LAYER met4 ;
        RECT 66.060000 91.405000 66.380000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 91.815000 66.380000 92.135000 ;
      LAYER met4 ;
        RECT 66.060000 91.815000 66.380000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 92.225000 66.380000 92.545000 ;
      LAYER met4 ;
        RECT 66.060000 92.225000 66.380000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060000 92.635000 66.380000 92.955000 ;
      LAYER met4 ;
        RECT 66.060000 92.635000 66.380000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 68.065000 66.470000 68.385000 ;
      LAYER met4 ;
        RECT 66.150000 68.065000 66.470000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 68.475000 66.470000 68.795000 ;
      LAYER met4 ;
        RECT 66.150000 68.475000 66.470000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 68.885000 66.470000 69.205000 ;
      LAYER met4 ;
        RECT 66.150000 68.885000 66.470000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 69.295000 66.470000 69.615000 ;
      LAYER met4 ;
        RECT 66.150000 69.295000 66.470000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 69.705000 66.470000 70.025000 ;
      LAYER met4 ;
        RECT 66.150000 69.705000 66.470000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 70.115000 66.470000 70.435000 ;
      LAYER met4 ;
        RECT 66.150000 70.115000 66.470000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 70.525000 66.470000 70.845000 ;
      LAYER met4 ;
        RECT 66.150000 70.525000 66.470000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 70.935000 66.470000 71.255000 ;
      LAYER met4 ;
        RECT 66.150000 70.935000 66.470000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 71.345000 66.470000 71.665000 ;
      LAYER met4 ;
        RECT 66.150000 71.345000 66.470000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 71.755000 66.470000 72.075000 ;
      LAYER met4 ;
        RECT 66.150000 71.755000 66.470000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 72.165000 66.470000 72.485000 ;
      LAYER met4 ;
        RECT 66.150000 72.165000 66.470000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 72.575000 66.470000 72.895000 ;
      LAYER met4 ;
        RECT 66.150000 72.575000 66.470000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 72.985000 66.470000 73.305000 ;
      LAYER met4 ;
        RECT 66.150000 72.985000 66.470000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 73.390000 66.470000 73.710000 ;
      LAYER met4 ;
        RECT 66.150000 73.390000 66.470000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 73.795000 66.470000 74.115000 ;
      LAYER met4 ;
        RECT 66.150000 73.795000 66.470000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 74.200000 66.470000 74.520000 ;
      LAYER met4 ;
        RECT 66.150000 74.200000 66.470000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 74.605000 66.470000 74.925000 ;
      LAYER met4 ;
        RECT 66.150000 74.605000 66.470000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 75.010000 66.470000 75.330000 ;
      LAYER met4 ;
        RECT 66.150000 75.010000 66.470000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 75.415000 66.470000 75.735000 ;
      LAYER met4 ;
        RECT 66.150000 75.415000 66.470000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 75.820000 66.470000 76.140000 ;
      LAYER met4 ;
        RECT 66.150000 75.820000 66.470000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 76.225000 66.470000 76.545000 ;
      LAYER met4 ;
        RECT 66.150000 76.225000 66.470000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 76.630000 66.470000 76.950000 ;
      LAYER met4 ;
        RECT 66.150000 76.630000 66.470000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 77.035000 66.470000 77.355000 ;
      LAYER met4 ;
        RECT 66.150000 77.035000 66.470000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 77.440000 66.470000 77.760000 ;
      LAYER met4 ;
        RECT 66.150000 77.440000 66.470000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 77.845000 66.470000 78.165000 ;
      LAYER met4 ;
        RECT 66.150000 77.845000 66.470000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 78.250000 66.470000 78.570000 ;
      LAYER met4 ;
        RECT 66.150000 78.250000 66.470000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 78.655000 66.470000 78.975000 ;
      LAYER met4 ;
        RECT 66.150000 78.655000 66.470000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 79.060000 66.470000 79.380000 ;
      LAYER met4 ;
        RECT 66.150000 79.060000 66.470000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 79.465000 66.470000 79.785000 ;
      LAYER met4 ;
        RECT 66.150000 79.465000 66.470000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 79.870000 66.470000 80.190000 ;
      LAYER met4 ;
        RECT 66.150000 79.870000 66.470000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 80.275000 66.470000 80.595000 ;
      LAYER met4 ;
        RECT 66.150000 80.275000 66.470000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 80.680000 66.470000 81.000000 ;
      LAYER met4 ;
        RECT 66.150000 80.680000 66.470000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 81.085000 66.470000 81.405000 ;
      LAYER met4 ;
        RECT 66.150000 81.085000 66.470000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 81.490000 66.470000 81.810000 ;
      LAYER met4 ;
        RECT 66.150000 81.490000 66.470000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 81.895000 66.470000 82.215000 ;
      LAYER met4 ;
        RECT 66.150000 81.895000 66.470000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.150000 82.300000 66.470000 82.620000 ;
      LAYER met4 ;
        RECT 66.150000 82.300000 66.470000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.175000 17.800000 66.495000 18.120000 ;
      LAYER met4 ;
        RECT 66.175000 17.800000 66.495000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.175000 18.230000 66.495000 18.550000 ;
      LAYER met4 ;
        RECT 66.175000 18.230000 66.495000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.175000 18.660000 66.495000 18.980000 ;
      LAYER met4 ;
        RECT 66.175000 18.660000 66.495000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.175000 19.090000 66.495000 19.410000 ;
      LAYER met4 ;
        RECT 66.175000 19.090000 66.495000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.175000 19.520000 66.495000 19.840000 ;
      LAYER met4 ;
        RECT 66.175000 19.520000 66.495000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.175000 19.950000 66.495000 20.270000 ;
      LAYER met4 ;
        RECT 66.175000 19.950000 66.495000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.175000 20.380000 66.495000 20.700000 ;
      LAYER met4 ;
        RECT 66.175000 20.380000 66.495000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.175000 20.810000 66.495000 21.130000 ;
      LAYER met4 ;
        RECT 66.175000 20.810000 66.495000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.175000 21.240000 66.495000 21.560000 ;
      LAYER met4 ;
        RECT 66.175000 21.240000 66.495000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.175000 21.670000 66.495000 21.990000 ;
      LAYER met4 ;
        RECT 66.175000 21.670000 66.495000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.175000 22.100000 66.495000 22.420000 ;
      LAYER met4 ;
        RECT 66.175000 22.100000 66.495000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 82.795000 66.790000 83.115000 ;
      LAYER met4 ;
        RECT 66.470000 82.795000 66.790000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 83.205000 66.790000 83.525000 ;
      LAYER met4 ;
        RECT 66.470000 83.205000 66.790000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 83.615000 66.790000 83.935000 ;
      LAYER met4 ;
        RECT 66.470000 83.615000 66.790000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 84.025000 66.790000 84.345000 ;
      LAYER met4 ;
        RECT 66.470000 84.025000 66.790000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 84.435000 66.790000 84.755000 ;
      LAYER met4 ;
        RECT 66.470000 84.435000 66.790000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 84.845000 66.790000 85.165000 ;
      LAYER met4 ;
        RECT 66.470000 84.845000 66.790000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 85.255000 66.790000 85.575000 ;
      LAYER met4 ;
        RECT 66.470000 85.255000 66.790000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 85.665000 66.790000 85.985000 ;
      LAYER met4 ;
        RECT 66.470000 85.665000 66.790000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 86.075000 66.790000 86.395000 ;
      LAYER met4 ;
        RECT 66.470000 86.075000 66.790000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 86.485000 66.790000 86.805000 ;
      LAYER met4 ;
        RECT 66.470000 86.485000 66.790000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 86.895000 66.790000 87.215000 ;
      LAYER met4 ;
        RECT 66.470000 86.895000 66.790000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 87.305000 66.790000 87.625000 ;
      LAYER met4 ;
        RECT 66.470000 87.305000 66.790000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 87.715000 66.790000 88.035000 ;
      LAYER met4 ;
        RECT 66.470000 87.715000 66.790000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 88.125000 66.790000 88.445000 ;
      LAYER met4 ;
        RECT 66.470000 88.125000 66.790000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 88.535000 66.790000 88.855000 ;
      LAYER met4 ;
        RECT 66.470000 88.535000 66.790000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 88.945000 66.790000 89.265000 ;
      LAYER met4 ;
        RECT 66.470000 88.945000 66.790000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 89.355000 66.790000 89.675000 ;
      LAYER met4 ;
        RECT 66.470000 89.355000 66.790000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 89.765000 66.790000 90.085000 ;
      LAYER met4 ;
        RECT 66.470000 89.765000 66.790000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 90.175000 66.790000 90.495000 ;
      LAYER met4 ;
        RECT 66.470000 90.175000 66.790000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 90.585000 66.790000 90.905000 ;
      LAYER met4 ;
        RECT 66.470000 90.585000 66.790000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 90.995000 66.790000 91.315000 ;
      LAYER met4 ;
        RECT 66.470000 90.995000 66.790000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 91.405000 66.790000 91.725000 ;
      LAYER met4 ;
        RECT 66.470000 91.405000 66.790000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 91.815000 66.790000 92.135000 ;
      LAYER met4 ;
        RECT 66.470000 91.815000 66.790000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 92.225000 66.790000 92.545000 ;
      LAYER met4 ;
        RECT 66.470000 92.225000 66.790000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470000 92.635000 66.790000 92.955000 ;
      LAYER met4 ;
        RECT 66.470000 92.635000 66.790000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 68.065000 66.870000 68.385000 ;
      LAYER met4 ;
        RECT 66.550000 68.065000 66.870000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 68.475000 66.870000 68.795000 ;
      LAYER met4 ;
        RECT 66.550000 68.475000 66.870000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 68.885000 66.870000 69.205000 ;
      LAYER met4 ;
        RECT 66.550000 68.885000 66.870000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 69.295000 66.870000 69.615000 ;
      LAYER met4 ;
        RECT 66.550000 69.295000 66.870000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 69.705000 66.870000 70.025000 ;
      LAYER met4 ;
        RECT 66.550000 69.705000 66.870000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 70.115000 66.870000 70.435000 ;
      LAYER met4 ;
        RECT 66.550000 70.115000 66.870000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 70.525000 66.870000 70.845000 ;
      LAYER met4 ;
        RECT 66.550000 70.525000 66.870000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 70.935000 66.870000 71.255000 ;
      LAYER met4 ;
        RECT 66.550000 70.935000 66.870000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 71.345000 66.870000 71.665000 ;
      LAYER met4 ;
        RECT 66.550000 71.345000 66.870000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 71.755000 66.870000 72.075000 ;
      LAYER met4 ;
        RECT 66.550000 71.755000 66.870000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 72.165000 66.870000 72.485000 ;
      LAYER met4 ;
        RECT 66.550000 72.165000 66.870000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 72.575000 66.870000 72.895000 ;
      LAYER met4 ;
        RECT 66.550000 72.575000 66.870000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 72.985000 66.870000 73.305000 ;
      LAYER met4 ;
        RECT 66.550000 72.985000 66.870000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 73.390000 66.870000 73.710000 ;
      LAYER met4 ;
        RECT 66.550000 73.390000 66.870000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 73.795000 66.870000 74.115000 ;
      LAYER met4 ;
        RECT 66.550000 73.795000 66.870000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 74.200000 66.870000 74.520000 ;
      LAYER met4 ;
        RECT 66.550000 74.200000 66.870000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 74.605000 66.870000 74.925000 ;
      LAYER met4 ;
        RECT 66.550000 74.605000 66.870000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 75.010000 66.870000 75.330000 ;
      LAYER met4 ;
        RECT 66.550000 75.010000 66.870000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 75.415000 66.870000 75.735000 ;
      LAYER met4 ;
        RECT 66.550000 75.415000 66.870000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 75.820000 66.870000 76.140000 ;
      LAYER met4 ;
        RECT 66.550000 75.820000 66.870000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 76.225000 66.870000 76.545000 ;
      LAYER met4 ;
        RECT 66.550000 76.225000 66.870000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 76.630000 66.870000 76.950000 ;
      LAYER met4 ;
        RECT 66.550000 76.630000 66.870000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 77.035000 66.870000 77.355000 ;
      LAYER met4 ;
        RECT 66.550000 77.035000 66.870000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 77.440000 66.870000 77.760000 ;
      LAYER met4 ;
        RECT 66.550000 77.440000 66.870000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 77.845000 66.870000 78.165000 ;
      LAYER met4 ;
        RECT 66.550000 77.845000 66.870000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 78.250000 66.870000 78.570000 ;
      LAYER met4 ;
        RECT 66.550000 78.250000 66.870000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 78.655000 66.870000 78.975000 ;
      LAYER met4 ;
        RECT 66.550000 78.655000 66.870000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 79.060000 66.870000 79.380000 ;
      LAYER met4 ;
        RECT 66.550000 79.060000 66.870000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 79.465000 66.870000 79.785000 ;
      LAYER met4 ;
        RECT 66.550000 79.465000 66.870000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 79.870000 66.870000 80.190000 ;
      LAYER met4 ;
        RECT 66.550000 79.870000 66.870000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 80.275000 66.870000 80.595000 ;
      LAYER met4 ;
        RECT 66.550000 80.275000 66.870000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 80.680000 66.870000 81.000000 ;
      LAYER met4 ;
        RECT 66.550000 80.680000 66.870000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 81.085000 66.870000 81.405000 ;
      LAYER met4 ;
        RECT 66.550000 81.085000 66.870000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 81.490000 66.870000 81.810000 ;
      LAYER met4 ;
        RECT 66.550000 81.490000 66.870000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 81.895000 66.870000 82.215000 ;
      LAYER met4 ;
        RECT 66.550000 81.895000 66.870000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.550000 82.300000 66.870000 82.620000 ;
      LAYER met4 ;
        RECT 66.550000 82.300000 66.870000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.580000 17.800000 66.900000 18.120000 ;
      LAYER met4 ;
        RECT 66.580000 17.800000 66.900000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.580000 18.230000 66.900000 18.550000 ;
      LAYER met4 ;
        RECT 66.580000 18.230000 66.900000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.580000 18.660000 66.900000 18.980000 ;
      LAYER met4 ;
        RECT 66.580000 18.660000 66.900000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.580000 19.090000 66.900000 19.410000 ;
      LAYER met4 ;
        RECT 66.580000 19.090000 66.900000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.580000 19.520000 66.900000 19.840000 ;
      LAYER met4 ;
        RECT 66.580000 19.520000 66.900000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.580000 19.950000 66.900000 20.270000 ;
      LAYER met4 ;
        RECT 66.580000 19.950000 66.900000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.580000 20.380000 66.900000 20.700000 ;
      LAYER met4 ;
        RECT 66.580000 20.380000 66.900000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.580000 20.810000 66.900000 21.130000 ;
      LAYER met4 ;
        RECT 66.580000 20.810000 66.900000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.580000 21.240000 66.900000 21.560000 ;
      LAYER met4 ;
        RECT 66.580000 21.240000 66.900000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.580000 21.670000 66.900000 21.990000 ;
      LAYER met4 ;
        RECT 66.580000 21.670000 66.900000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.580000 22.100000 66.900000 22.420000 ;
      LAYER met4 ;
        RECT 66.580000 22.100000 66.900000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 82.795000 67.200000 83.115000 ;
      LAYER met4 ;
        RECT 66.880000 82.795000 67.200000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 83.205000 67.200000 83.525000 ;
      LAYER met4 ;
        RECT 66.880000 83.205000 67.200000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 83.615000 67.200000 83.935000 ;
      LAYER met4 ;
        RECT 66.880000 83.615000 67.200000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 84.025000 67.200000 84.345000 ;
      LAYER met4 ;
        RECT 66.880000 84.025000 67.200000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 84.435000 67.200000 84.755000 ;
      LAYER met4 ;
        RECT 66.880000 84.435000 67.200000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 84.845000 67.200000 85.165000 ;
      LAYER met4 ;
        RECT 66.880000 84.845000 67.200000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 85.255000 67.200000 85.575000 ;
      LAYER met4 ;
        RECT 66.880000 85.255000 67.200000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 85.665000 67.200000 85.985000 ;
      LAYER met4 ;
        RECT 66.880000 85.665000 67.200000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 86.075000 67.200000 86.395000 ;
      LAYER met4 ;
        RECT 66.880000 86.075000 67.200000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 86.485000 67.200000 86.805000 ;
      LAYER met4 ;
        RECT 66.880000 86.485000 67.200000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 86.895000 67.200000 87.215000 ;
      LAYER met4 ;
        RECT 66.880000 86.895000 67.200000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 87.305000 67.200000 87.625000 ;
      LAYER met4 ;
        RECT 66.880000 87.305000 67.200000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 87.715000 67.200000 88.035000 ;
      LAYER met4 ;
        RECT 66.880000 87.715000 67.200000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 88.125000 67.200000 88.445000 ;
      LAYER met4 ;
        RECT 66.880000 88.125000 67.200000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 88.535000 67.200000 88.855000 ;
      LAYER met4 ;
        RECT 66.880000 88.535000 67.200000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 88.945000 67.200000 89.265000 ;
      LAYER met4 ;
        RECT 66.880000 88.945000 67.200000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 89.355000 67.200000 89.675000 ;
      LAYER met4 ;
        RECT 66.880000 89.355000 67.200000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 89.765000 67.200000 90.085000 ;
      LAYER met4 ;
        RECT 66.880000 89.765000 67.200000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 90.175000 67.200000 90.495000 ;
      LAYER met4 ;
        RECT 66.880000 90.175000 67.200000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 90.585000 67.200000 90.905000 ;
      LAYER met4 ;
        RECT 66.880000 90.585000 67.200000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 90.995000 67.200000 91.315000 ;
      LAYER met4 ;
        RECT 66.880000 90.995000 67.200000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 91.405000 67.200000 91.725000 ;
      LAYER met4 ;
        RECT 66.880000 91.405000 67.200000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 91.815000 67.200000 92.135000 ;
      LAYER met4 ;
        RECT 66.880000 91.815000 67.200000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 92.225000 67.200000 92.545000 ;
      LAYER met4 ;
        RECT 66.880000 92.225000 67.200000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880000 92.635000 67.200000 92.955000 ;
      LAYER met4 ;
        RECT 66.880000 92.635000 67.200000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 68.065000 67.270000 68.385000 ;
      LAYER met4 ;
        RECT 66.950000 68.065000 67.270000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 68.475000 67.270000 68.795000 ;
      LAYER met4 ;
        RECT 66.950000 68.475000 67.270000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 68.885000 67.270000 69.205000 ;
      LAYER met4 ;
        RECT 66.950000 68.885000 67.270000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 69.295000 67.270000 69.615000 ;
      LAYER met4 ;
        RECT 66.950000 69.295000 67.270000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 69.705000 67.270000 70.025000 ;
      LAYER met4 ;
        RECT 66.950000 69.705000 67.270000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 70.115000 67.270000 70.435000 ;
      LAYER met4 ;
        RECT 66.950000 70.115000 67.270000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 70.525000 67.270000 70.845000 ;
      LAYER met4 ;
        RECT 66.950000 70.525000 67.270000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 70.935000 67.270000 71.255000 ;
      LAYER met4 ;
        RECT 66.950000 70.935000 67.270000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 71.345000 67.270000 71.665000 ;
      LAYER met4 ;
        RECT 66.950000 71.345000 67.270000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 71.755000 67.270000 72.075000 ;
      LAYER met4 ;
        RECT 66.950000 71.755000 67.270000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 72.165000 67.270000 72.485000 ;
      LAYER met4 ;
        RECT 66.950000 72.165000 67.270000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 72.575000 67.270000 72.895000 ;
      LAYER met4 ;
        RECT 66.950000 72.575000 67.270000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 72.985000 67.270000 73.305000 ;
      LAYER met4 ;
        RECT 66.950000 72.985000 67.270000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 73.390000 67.270000 73.710000 ;
      LAYER met4 ;
        RECT 66.950000 73.390000 67.270000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 73.795000 67.270000 74.115000 ;
      LAYER met4 ;
        RECT 66.950000 73.795000 67.270000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 74.200000 67.270000 74.520000 ;
      LAYER met4 ;
        RECT 66.950000 74.200000 67.270000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 74.605000 67.270000 74.925000 ;
      LAYER met4 ;
        RECT 66.950000 74.605000 67.270000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 75.010000 67.270000 75.330000 ;
      LAYER met4 ;
        RECT 66.950000 75.010000 67.270000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 75.415000 67.270000 75.735000 ;
      LAYER met4 ;
        RECT 66.950000 75.415000 67.270000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 75.820000 67.270000 76.140000 ;
      LAYER met4 ;
        RECT 66.950000 75.820000 67.270000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 76.225000 67.270000 76.545000 ;
      LAYER met4 ;
        RECT 66.950000 76.225000 67.270000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 76.630000 67.270000 76.950000 ;
      LAYER met4 ;
        RECT 66.950000 76.630000 67.270000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 77.035000 67.270000 77.355000 ;
      LAYER met4 ;
        RECT 66.950000 77.035000 67.270000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 77.440000 67.270000 77.760000 ;
      LAYER met4 ;
        RECT 66.950000 77.440000 67.270000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 77.845000 67.270000 78.165000 ;
      LAYER met4 ;
        RECT 66.950000 77.845000 67.270000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 78.250000 67.270000 78.570000 ;
      LAYER met4 ;
        RECT 66.950000 78.250000 67.270000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 78.655000 67.270000 78.975000 ;
      LAYER met4 ;
        RECT 66.950000 78.655000 67.270000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 79.060000 67.270000 79.380000 ;
      LAYER met4 ;
        RECT 66.950000 79.060000 67.270000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 79.465000 67.270000 79.785000 ;
      LAYER met4 ;
        RECT 66.950000 79.465000 67.270000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 79.870000 67.270000 80.190000 ;
      LAYER met4 ;
        RECT 66.950000 79.870000 67.270000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 80.275000 67.270000 80.595000 ;
      LAYER met4 ;
        RECT 66.950000 80.275000 67.270000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 80.680000 67.270000 81.000000 ;
      LAYER met4 ;
        RECT 66.950000 80.680000 67.270000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 81.085000 67.270000 81.405000 ;
      LAYER met4 ;
        RECT 66.950000 81.085000 67.270000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 81.490000 67.270000 81.810000 ;
      LAYER met4 ;
        RECT 66.950000 81.490000 67.270000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 81.895000 67.270000 82.215000 ;
      LAYER met4 ;
        RECT 66.950000 81.895000 67.270000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.950000 82.300000 67.270000 82.620000 ;
      LAYER met4 ;
        RECT 66.950000 82.300000 67.270000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.985000 17.800000 67.305000 18.120000 ;
      LAYER met4 ;
        RECT 66.985000 17.800000 67.305000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.985000 18.230000 67.305000 18.550000 ;
      LAYER met4 ;
        RECT 66.985000 18.230000 67.305000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.985000 18.660000 67.305000 18.980000 ;
      LAYER met4 ;
        RECT 66.985000 18.660000 67.305000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.985000 19.090000 67.305000 19.410000 ;
      LAYER met4 ;
        RECT 66.985000 19.090000 67.305000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.985000 19.520000 67.305000 19.840000 ;
      LAYER met4 ;
        RECT 66.985000 19.520000 67.305000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.985000 19.950000 67.305000 20.270000 ;
      LAYER met4 ;
        RECT 66.985000 19.950000 67.305000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.985000 20.380000 67.305000 20.700000 ;
      LAYER met4 ;
        RECT 66.985000 20.380000 67.305000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.985000 20.810000 67.305000 21.130000 ;
      LAYER met4 ;
        RECT 66.985000 20.810000 67.305000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.985000 21.240000 67.305000 21.560000 ;
      LAYER met4 ;
        RECT 66.985000 21.240000 67.305000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.985000 21.670000 67.305000 21.990000 ;
      LAYER met4 ;
        RECT 66.985000 21.670000 67.305000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.985000 22.100000 67.305000 22.420000 ;
      LAYER met4 ;
        RECT 66.985000 22.100000 67.305000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 82.795000 67.610000 83.115000 ;
      LAYER met4 ;
        RECT 67.290000 82.795000 67.610000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 83.205000 67.610000 83.525000 ;
      LAYER met4 ;
        RECT 67.290000 83.205000 67.610000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 83.615000 67.610000 83.935000 ;
      LAYER met4 ;
        RECT 67.290000 83.615000 67.610000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 84.025000 67.610000 84.345000 ;
      LAYER met4 ;
        RECT 67.290000 84.025000 67.610000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 84.435000 67.610000 84.755000 ;
      LAYER met4 ;
        RECT 67.290000 84.435000 67.610000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 84.845000 67.610000 85.165000 ;
      LAYER met4 ;
        RECT 67.290000 84.845000 67.610000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 85.255000 67.610000 85.575000 ;
      LAYER met4 ;
        RECT 67.290000 85.255000 67.610000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 85.665000 67.610000 85.985000 ;
      LAYER met4 ;
        RECT 67.290000 85.665000 67.610000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 86.075000 67.610000 86.395000 ;
      LAYER met4 ;
        RECT 67.290000 86.075000 67.610000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 86.485000 67.610000 86.805000 ;
      LAYER met4 ;
        RECT 67.290000 86.485000 67.610000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 86.895000 67.610000 87.215000 ;
      LAYER met4 ;
        RECT 67.290000 86.895000 67.610000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 87.305000 67.610000 87.625000 ;
      LAYER met4 ;
        RECT 67.290000 87.305000 67.610000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 87.715000 67.610000 88.035000 ;
      LAYER met4 ;
        RECT 67.290000 87.715000 67.610000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 88.125000 67.610000 88.445000 ;
      LAYER met4 ;
        RECT 67.290000 88.125000 67.610000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 88.535000 67.610000 88.855000 ;
      LAYER met4 ;
        RECT 67.290000 88.535000 67.610000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 88.945000 67.610000 89.265000 ;
      LAYER met4 ;
        RECT 67.290000 88.945000 67.610000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 89.355000 67.610000 89.675000 ;
      LAYER met4 ;
        RECT 67.290000 89.355000 67.610000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 89.765000 67.610000 90.085000 ;
      LAYER met4 ;
        RECT 67.290000 89.765000 67.610000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 90.175000 67.610000 90.495000 ;
      LAYER met4 ;
        RECT 67.290000 90.175000 67.610000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 90.585000 67.610000 90.905000 ;
      LAYER met4 ;
        RECT 67.290000 90.585000 67.610000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 90.995000 67.610000 91.315000 ;
      LAYER met4 ;
        RECT 67.290000 90.995000 67.610000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 91.405000 67.610000 91.725000 ;
      LAYER met4 ;
        RECT 67.290000 91.405000 67.610000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 91.815000 67.610000 92.135000 ;
      LAYER met4 ;
        RECT 67.290000 91.815000 67.610000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 92.225000 67.610000 92.545000 ;
      LAYER met4 ;
        RECT 67.290000 92.225000 67.610000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290000 92.635000 67.610000 92.955000 ;
      LAYER met4 ;
        RECT 67.290000 92.635000 67.610000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 68.065000 67.670000 68.385000 ;
      LAYER met4 ;
        RECT 67.350000 68.065000 67.670000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 68.475000 67.670000 68.795000 ;
      LAYER met4 ;
        RECT 67.350000 68.475000 67.670000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 68.885000 67.670000 69.205000 ;
      LAYER met4 ;
        RECT 67.350000 68.885000 67.670000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 69.295000 67.670000 69.615000 ;
      LAYER met4 ;
        RECT 67.350000 69.295000 67.670000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 69.705000 67.670000 70.025000 ;
      LAYER met4 ;
        RECT 67.350000 69.705000 67.670000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 70.115000 67.670000 70.435000 ;
      LAYER met4 ;
        RECT 67.350000 70.115000 67.670000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 70.525000 67.670000 70.845000 ;
      LAYER met4 ;
        RECT 67.350000 70.525000 67.670000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 70.935000 67.670000 71.255000 ;
      LAYER met4 ;
        RECT 67.350000 70.935000 67.670000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 71.345000 67.670000 71.665000 ;
      LAYER met4 ;
        RECT 67.350000 71.345000 67.670000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 71.755000 67.670000 72.075000 ;
      LAYER met4 ;
        RECT 67.350000 71.755000 67.670000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 72.165000 67.670000 72.485000 ;
      LAYER met4 ;
        RECT 67.350000 72.165000 67.670000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 72.575000 67.670000 72.895000 ;
      LAYER met4 ;
        RECT 67.350000 72.575000 67.670000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 72.985000 67.670000 73.305000 ;
      LAYER met4 ;
        RECT 67.350000 72.985000 67.670000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 73.390000 67.670000 73.710000 ;
      LAYER met4 ;
        RECT 67.350000 73.390000 67.670000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 73.795000 67.670000 74.115000 ;
      LAYER met4 ;
        RECT 67.350000 73.795000 67.670000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 74.200000 67.670000 74.520000 ;
      LAYER met4 ;
        RECT 67.350000 74.200000 67.670000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 74.605000 67.670000 74.925000 ;
      LAYER met4 ;
        RECT 67.350000 74.605000 67.670000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 75.010000 67.670000 75.330000 ;
      LAYER met4 ;
        RECT 67.350000 75.010000 67.670000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 75.415000 67.670000 75.735000 ;
      LAYER met4 ;
        RECT 67.350000 75.415000 67.670000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 75.820000 67.670000 76.140000 ;
      LAYER met4 ;
        RECT 67.350000 75.820000 67.670000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 76.225000 67.670000 76.545000 ;
      LAYER met4 ;
        RECT 67.350000 76.225000 67.670000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 76.630000 67.670000 76.950000 ;
      LAYER met4 ;
        RECT 67.350000 76.630000 67.670000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 77.035000 67.670000 77.355000 ;
      LAYER met4 ;
        RECT 67.350000 77.035000 67.670000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 77.440000 67.670000 77.760000 ;
      LAYER met4 ;
        RECT 67.350000 77.440000 67.670000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 77.845000 67.670000 78.165000 ;
      LAYER met4 ;
        RECT 67.350000 77.845000 67.670000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 78.250000 67.670000 78.570000 ;
      LAYER met4 ;
        RECT 67.350000 78.250000 67.670000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 78.655000 67.670000 78.975000 ;
      LAYER met4 ;
        RECT 67.350000 78.655000 67.670000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 79.060000 67.670000 79.380000 ;
      LAYER met4 ;
        RECT 67.350000 79.060000 67.670000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 79.465000 67.670000 79.785000 ;
      LAYER met4 ;
        RECT 67.350000 79.465000 67.670000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 79.870000 67.670000 80.190000 ;
      LAYER met4 ;
        RECT 67.350000 79.870000 67.670000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 80.275000 67.670000 80.595000 ;
      LAYER met4 ;
        RECT 67.350000 80.275000 67.670000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 80.680000 67.670000 81.000000 ;
      LAYER met4 ;
        RECT 67.350000 80.680000 67.670000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 81.085000 67.670000 81.405000 ;
      LAYER met4 ;
        RECT 67.350000 81.085000 67.670000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 81.490000 67.670000 81.810000 ;
      LAYER met4 ;
        RECT 67.350000 81.490000 67.670000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 81.895000 67.670000 82.215000 ;
      LAYER met4 ;
        RECT 67.350000 81.895000 67.670000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350000 82.300000 67.670000 82.620000 ;
      LAYER met4 ;
        RECT 67.350000 82.300000 67.670000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 17.800000 67.710000 18.120000 ;
      LAYER met4 ;
        RECT 67.390000 17.800000 67.710000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 18.230000 67.710000 18.550000 ;
      LAYER met4 ;
        RECT 67.390000 18.230000 67.710000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 18.660000 67.710000 18.980000 ;
      LAYER met4 ;
        RECT 67.390000 18.660000 67.710000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 19.090000 67.710000 19.410000 ;
      LAYER met4 ;
        RECT 67.390000 19.090000 67.710000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 19.520000 67.710000 19.840000 ;
      LAYER met4 ;
        RECT 67.390000 19.520000 67.710000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 19.950000 67.710000 20.270000 ;
      LAYER met4 ;
        RECT 67.390000 19.950000 67.710000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 20.380000 67.710000 20.700000 ;
      LAYER met4 ;
        RECT 67.390000 20.380000 67.710000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 20.810000 67.710000 21.130000 ;
      LAYER met4 ;
        RECT 67.390000 20.810000 67.710000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 21.240000 67.710000 21.560000 ;
      LAYER met4 ;
        RECT 67.390000 21.240000 67.710000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 21.670000 67.710000 21.990000 ;
      LAYER met4 ;
        RECT 67.390000 21.670000 67.710000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 22.100000 67.710000 22.420000 ;
      LAYER met4 ;
        RECT 67.390000 22.100000 67.710000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 82.795000 68.020000 83.115000 ;
      LAYER met4 ;
        RECT 67.700000 82.795000 68.020000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 83.205000 68.020000 83.525000 ;
      LAYER met4 ;
        RECT 67.700000 83.205000 68.020000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 83.615000 68.020000 83.935000 ;
      LAYER met4 ;
        RECT 67.700000 83.615000 68.020000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 84.025000 68.020000 84.345000 ;
      LAYER met4 ;
        RECT 67.700000 84.025000 68.020000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 84.435000 68.020000 84.755000 ;
      LAYER met4 ;
        RECT 67.700000 84.435000 68.020000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 84.845000 68.020000 85.165000 ;
      LAYER met4 ;
        RECT 67.700000 84.845000 68.020000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 85.255000 68.020000 85.575000 ;
      LAYER met4 ;
        RECT 67.700000 85.255000 68.020000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 85.665000 68.020000 85.985000 ;
      LAYER met4 ;
        RECT 67.700000 85.665000 68.020000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 86.075000 68.020000 86.395000 ;
      LAYER met4 ;
        RECT 67.700000 86.075000 68.020000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 86.485000 68.020000 86.805000 ;
      LAYER met4 ;
        RECT 67.700000 86.485000 68.020000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 86.895000 68.020000 87.215000 ;
      LAYER met4 ;
        RECT 67.700000 86.895000 68.020000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 87.305000 68.020000 87.625000 ;
      LAYER met4 ;
        RECT 67.700000 87.305000 68.020000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 87.715000 68.020000 88.035000 ;
      LAYER met4 ;
        RECT 67.700000 87.715000 68.020000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 88.125000 68.020000 88.445000 ;
      LAYER met4 ;
        RECT 67.700000 88.125000 68.020000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 88.535000 68.020000 88.855000 ;
      LAYER met4 ;
        RECT 67.700000 88.535000 68.020000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 88.945000 68.020000 89.265000 ;
      LAYER met4 ;
        RECT 67.700000 88.945000 68.020000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 89.355000 68.020000 89.675000 ;
      LAYER met4 ;
        RECT 67.700000 89.355000 68.020000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 89.765000 68.020000 90.085000 ;
      LAYER met4 ;
        RECT 67.700000 89.765000 68.020000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 90.175000 68.020000 90.495000 ;
      LAYER met4 ;
        RECT 67.700000 90.175000 68.020000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 90.585000 68.020000 90.905000 ;
      LAYER met4 ;
        RECT 67.700000 90.585000 68.020000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 90.995000 68.020000 91.315000 ;
      LAYER met4 ;
        RECT 67.700000 90.995000 68.020000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 91.405000 68.020000 91.725000 ;
      LAYER met4 ;
        RECT 67.700000 91.405000 68.020000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 91.815000 68.020000 92.135000 ;
      LAYER met4 ;
        RECT 67.700000 91.815000 68.020000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 92.225000 68.020000 92.545000 ;
      LAYER met4 ;
        RECT 67.700000 92.225000 68.020000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700000 92.635000 68.020000 92.955000 ;
      LAYER met4 ;
        RECT 67.700000 92.635000 68.020000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 68.065000 68.070000 68.385000 ;
      LAYER met4 ;
        RECT 67.750000 68.065000 68.070000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 68.475000 68.070000 68.795000 ;
      LAYER met4 ;
        RECT 67.750000 68.475000 68.070000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 68.885000 68.070000 69.205000 ;
      LAYER met4 ;
        RECT 67.750000 68.885000 68.070000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 69.295000 68.070000 69.615000 ;
      LAYER met4 ;
        RECT 67.750000 69.295000 68.070000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 69.705000 68.070000 70.025000 ;
      LAYER met4 ;
        RECT 67.750000 69.705000 68.070000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 70.115000 68.070000 70.435000 ;
      LAYER met4 ;
        RECT 67.750000 70.115000 68.070000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 70.525000 68.070000 70.845000 ;
      LAYER met4 ;
        RECT 67.750000 70.525000 68.070000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 70.935000 68.070000 71.255000 ;
      LAYER met4 ;
        RECT 67.750000 70.935000 68.070000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 71.345000 68.070000 71.665000 ;
      LAYER met4 ;
        RECT 67.750000 71.345000 68.070000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 71.755000 68.070000 72.075000 ;
      LAYER met4 ;
        RECT 67.750000 71.755000 68.070000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 72.165000 68.070000 72.485000 ;
      LAYER met4 ;
        RECT 67.750000 72.165000 68.070000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 72.575000 68.070000 72.895000 ;
      LAYER met4 ;
        RECT 67.750000 72.575000 68.070000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 72.985000 68.070000 73.305000 ;
      LAYER met4 ;
        RECT 67.750000 72.985000 68.070000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 73.390000 68.070000 73.710000 ;
      LAYER met4 ;
        RECT 67.750000 73.390000 68.070000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 73.795000 68.070000 74.115000 ;
      LAYER met4 ;
        RECT 67.750000 73.795000 68.070000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 74.200000 68.070000 74.520000 ;
      LAYER met4 ;
        RECT 67.750000 74.200000 68.070000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 74.605000 68.070000 74.925000 ;
      LAYER met4 ;
        RECT 67.750000 74.605000 68.070000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 75.010000 68.070000 75.330000 ;
      LAYER met4 ;
        RECT 67.750000 75.010000 68.070000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 75.415000 68.070000 75.735000 ;
      LAYER met4 ;
        RECT 67.750000 75.415000 68.070000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 75.820000 68.070000 76.140000 ;
      LAYER met4 ;
        RECT 67.750000 75.820000 68.070000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 76.225000 68.070000 76.545000 ;
      LAYER met4 ;
        RECT 67.750000 76.225000 68.070000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 76.630000 68.070000 76.950000 ;
      LAYER met4 ;
        RECT 67.750000 76.630000 68.070000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 77.035000 68.070000 77.355000 ;
      LAYER met4 ;
        RECT 67.750000 77.035000 68.070000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 77.440000 68.070000 77.760000 ;
      LAYER met4 ;
        RECT 67.750000 77.440000 68.070000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 77.845000 68.070000 78.165000 ;
      LAYER met4 ;
        RECT 67.750000 77.845000 68.070000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 78.250000 68.070000 78.570000 ;
      LAYER met4 ;
        RECT 67.750000 78.250000 68.070000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 78.655000 68.070000 78.975000 ;
      LAYER met4 ;
        RECT 67.750000 78.655000 68.070000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 79.060000 68.070000 79.380000 ;
      LAYER met4 ;
        RECT 67.750000 79.060000 68.070000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 79.465000 68.070000 79.785000 ;
      LAYER met4 ;
        RECT 67.750000 79.465000 68.070000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 79.870000 68.070000 80.190000 ;
      LAYER met4 ;
        RECT 67.750000 79.870000 68.070000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 80.275000 68.070000 80.595000 ;
      LAYER met4 ;
        RECT 67.750000 80.275000 68.070000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 80.680000 68.070000 81.000000 ;
      LAYER met4 ;
        RECT 67.750000 80.680000 68.070000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 81.085000 68.070000 81.405000 ;
      LAYER met4 ;
        RECT 67.750000 81.085000 68.070000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 81.490000 68.070000 81.810000 ;
      LAYER met4 ;
        RECT 67.750000 81.490000 68.070000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 81.895000 68.070000 82.215000 ;
      LAYER met4 ;
        RECT 67.750000 81.895000 68.070000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.750000 82.300000 68.070000 82.620000 ;
      LAYER met4 ;
        RECT 67.750000 82.300000 68.070000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.795000 17.800000 68.115000 18.120000 ;
      LAYER met4 ;
        RECT 67.795000 17.800000 68.115000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.795000 18.230000 68.115000 18.550000 ;
      LAYER met4 ;
        RECT 67.795000 18.230000 68.115000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.795000 18.660000 68.115000 18.980000 ;
      LAYER met4 ;
        RECT 67.795000 18.660000 68.115000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.795000 19.090000 68.115000 19.410000 ;
      LAYER met4 ;
        RECT 67.795000 19.090000 68.115000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.795000 19.520000 68.115000 19.840000 ;
      LAYER met4 ;
        RECT 67.795000 19.520000 68.115000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.795000 19.950000 68.115000 20.270000 ;
      LAYER met4 ;
        RECT 67.795000 19.950000 68.115000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.795000 20.380000 68.115000 20.700000 ;
      LAYER met4 ;
        RECT 67.795000 20.380000 68.115000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.795000 20.810000 68.115000 21.130000 ;
      LAYER met4 ;
        RECT 67.795000 20.810000 68.115000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.795000 21.240000 68.115000 21.560000 ;
      LAYER met4 ;
        RECT 67.795000 21.240000 68.115000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.795000 21.670000 68.115000 21.990000 ;
      LAYER met4 ;
        RECT 67.795000 21.670000 68.115000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.795000 22.100000 68.115000 22.420000 ;
      LAYER met4 ;
        RECT 67.795000 22.100000 68.115000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 82.795000 68.430000 83.115000 ;
      LAYER met4 ;
        RECT 68.110000 82.795000 68.430000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 83.205000 68.430000 83.525000 ;
      LAYER met4 ;
        RECT 68.110000 83.205000 68.430000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 83.615000 68.430000 83.935000 ;
      LAYER met4 ;
        RECT 68.110000 83.615000 68.430000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 84.025000 68.430000 84.345000 ;
      LAYER met4 ;
        RECT 68.110000 84.025000 68.430000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 84.435000 68.430000 84.755000 ;
      LAYER met4 ;
        RECT 68.110000 84.435000 68.430000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 84.845000 68.430000 85.165000 ;
      LAYER met4 ;
        RECT 68.110000 84.845000 68.430000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 85.255000 68.430000 85.575000 ;
      LAYER met4 ;
        RECT 68.110000 85.255000 68.430000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 85.665000 68.430000 85.985000 ;
      LAYER met4 ;
        RECT 68.110000 85.665000 68.430000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 86.075000 68.430000 86.395000 ;
      LAYER met4 ;
        RECT 68.110000 86.075000 68.430000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 86.485000 68.430000 86.805000 ;
      LAYER met4 ;
        RECT 68.110000 86.485000 68.430000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 86.895000 68.430000 87.215000 ;
      LAYER met4 ;
        RECT 68.110000 86.895000 68.430000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 87.305000 68.430000 87.625000 ;
      LAYER met4 ;
        RECT 68.110000 87.305000 68.430000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 87.715000 68.430000 88.035000 ;
      LAYER met4 ;
        RECT 68.110000 87.715000 68.430000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 88.125000 68.430000 88.445000 ;
      LAYER met4 ;
        RECT 68.110000 88.125000 68.430000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 88.535000 68.430000 88.855000 ;
      LAYER met4 ;
        RECT 68.110000 88.535000 68.430000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 88.945000 68.430000 89.265000 ;
      LAYER met4 ;
        RECT 68.110000 88.945000 68.430000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 89.355000 68.430000 89.675000 ;
      LAYER met4 ;
        RECT 68.110000 89.355000 68.430000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 89.765000 68.430000 90.085000 ;
      LAYER met4 ;
        RECT 68.110000 89.765000 68.430000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 90.175000 68.430000 90.495000 ;
      LAYER met4 ;
        RECT 68.110000 90.175000 68.430000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 90.585000 68.430000 90.905000 ;
      LAYER met4 ;
        RECT 68.110000 90.585000 68.430000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 90.995000 68.430000 91.315000 ;
      LAYER met4 ;
        RECT 68.110000 90.995000 68.430000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 91.405000 68.430000 91.725000 ;
      LAYER met4 ;
        RECT 68.110000 91.405000 68.430000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 91.815000 68.430000 92.135000 ;
      LAYER met4 ;
        RECT 68.110000 91.815000 68.430000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 92.225000 68.430000 92.545000 ;
      LAYER met4 ;
        RECT 68.110000 92.225000 68.430000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110000 92.635000 68.430000 92.955000 ;
      LAYER met4 ;
        RECT 68.110000 92.635000 68.430000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 68.065000 68.470000 68.385000 ;
      LAYER met4 ;
        RECT 68.150000 68.065000 68.470000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 68.475000 68.470000 68.795000 ;
      LAYER met4 ;
        RECT 68.150000 68.475000 68.470000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 68.885000 68.470000 69.205000 ;
      LAYER met4 ;
        RECT 68.150000 68.885000 68.470000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 69.295000 68.470000 69.615000 ;
      LAYER met4 ;
        RECT 68.150000 69.295000 68.470000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 69.705000 68.470000 70.025000 ;
      LAYER met4 ;
        RECT 68.150000 69.705000 68.470000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 70.115000 68.470000 70.435000 ;
      LAYER met4 ;
        RECT 68.150000 70.115000 68.470000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 70.525000 68.470000 70.845000 ;
      LAYER met4 ;
        RECT 68.150000 70.525000 68.470000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 70.935000 68.470000 71.255000 ;
      LAYER met4 ;
        RECT 68.150000 70.935000 68.470000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 71.345000 68.470000 71.665000 ;
      LAYER met4 ;
        RECT 68.150000 71.345000 68.470000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 71.755000 68.470000 72.075000 ;
      LAYER met4 ;
        RECT 68.150000 71.755000 68.470000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 72.165000 68.470000 72.485000 ;
      LAYER met4 ;
        RECT 68.150000 72.165000 68.470000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 72.575000 68.470000 72.895000 ;
      LAYER met4 ;
        RECT 68.150000 72.575000 68.470000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 72.985000 68.470000 73.305000 ;
      LAYER met4 ;
        RECT 68.150000 72.985000 68.470000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 73.390000 68.470000 73.710000 ;
      LAYER met4 ;
        RECT 68.150000 73.390000 68.470000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 73.795000 68.470000 74.115000 ;
      LAYER met4 ;
        RECT 68.150000 73.795000 68.470000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 74.200000 68.470000 74.520000 ;
      LAYER met4 ;
        RECT 68.150000 74.200000 68.470000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 74.605000 68.470000 74.925000 ;
      LAYER met4 ;
        RECT 68.150000 74.605000 68.470000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 75.010000 68.470000 75.330000 ;
      LAYER met4 ;
        RECT 68.150000 75.010000 68.470000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 75.415000 68.470000 75.735000 ;
      LAYER met4 ;
        RECT 68.150000 75.415000 68.470000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 75.820000 68.470000 76.140000 ;
      LAYER met4 ;
        RECT 68.150000 75.820000 68.470000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 76.225000 68.470000 76.545000 ;
      LAYER met4 ;
        RECT 68.150000 76.225000 68.470000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 76.630000 68.470000 76.950000 ;
      LAYER met4 ;
        RECT 68.150000 76.630000 68.470000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 77.035000 68.470000 77.355000 ;
      LAYER met4 ;
        RECT 68.150000 77.035000 68.470000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 77.440000 68.470000 77.760000 ;
      LAYER met4 ;
        RECT 68.150000 77.440000 68.470000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 77.845000 68.470000 78.165000 ;
      LAYER met4 ;
        RECT 68.150000 77.845000 68.470000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 78.250000 68.470000 78.570000 ;
      LAYER met4 ;
        RECT 68.150000 78.250000 68.470000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 78.655000 68.470000 78.975000 ;
      LAYER met4 ;
        RECT 68.150000 78.655000 68.470000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 79.060000 68.470000 79.380000 ;
      LAYER met4 ;
        RECT 68.150000 79.060000 68.470000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 79.465000 68.470000 79.785000 ;
      LAYER met4 ;
        RECT 68.150000 79.465000 68.470000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 79.870000 68.470000 80.190000 ;
      LAYER met4 ;
        RECT 68.150000 79.870000 68.470000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 80.275000 68.470000 80.595000 ;
      LAYER met4 ;
        RECT 68.150000 80.275000 68.470000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 80.680000 68.470000 81.000000 ;
      LAYER met4 ;
        RECT 68.150000 80.680000 68.470000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 81.085000 68.470000 81.405000 ;
      LAYER met4 ;
        RECT 68.150000 81.085000 68.470000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 81.490000 68.470000 81.810000 ;
      LAYER met4 ;
        RECT 68.150000 81.490000 68.470000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 81.895000 68.470000 82.215000 ;
      LAYER met4 ;
        RECT 68.150000 81.895000 68.470000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.150000 82.300000 68.470000 82.620000 ;
      LAYER met4 ;
        RECT 68.150000 82.300000 68.470000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.200000 17.800000 68.520000 18.120000 ;
      LAYER met4 ;
        RECT 68.200000 17.800000 68.520000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.200000 18.230000 68.520000 18.550000 ;
      LAYER met4 ;
        RECT 68.200000 18.230000 68.520000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.200000 18.660000 68.520000 18.980000 ;
      LAYER met4 ;
        RECT 68.200000 18.660000 68.520000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.200000 19.090000 68.520000 19.410000 ;
      LAYER met4 ;
        RECT 68.200000 19.090000 68.520000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.200000 19.520000 68.520000 19.840000 ;
      LAYER met4 ;
        RECT 68.200000 19.520000 68.520000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.200000 19.950000 68.520000 20.270000 ;
      LAYER met4 ;
        RECT 68.200000 19.950000 68.520000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.200000 20.380000 68.520000 20.700000 ;
      LAYER met4 ;
        RECT 68.200000 20.380000 68.520000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.200000 20.810000 68.520000 21.130000 ;
      LAYER met4 ;
        RECT 68.200000 20.810000 68.520000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.200000 21.240000 68.520000 21.560000 ;
      LAYER met4 ;
        RECT 68.200000 21.240000 68.520000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.200000 21.670000 68.520000 21.990000 ;
      LAYER met4 ;
        RECT 68.200000 21.670000 68.520000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.200000 22.100000 68.520000 22.420000 ;
      LAYER met4 ;
        RECT 68.200000 22.100000 68.520000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 82.795000 68.840000 83.115000 ;
      LAYER met4 ;
        RECT 68.520000 82.795000 68.840000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 83.205000 68.840000 83.525000 ;
      LAYER met4 ;
        RECT 68.520000 83.205000 68.840000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 83.615000 68.840000 83.935000 ;
      LAYER met4 ;
        RECT 68.520000 83.615000 68.840000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 84.025000 68.840000 84.345000 ;
      LAYER met4 ;
        RECT 68.520000 84.025000 68.840000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 84.435000 68.840000 84.755000 ;
      LAYER met4 ;
        RECT 68.520000 84.435000 68.840000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 84.845000 68.840000 85.165000 ;
      LAYER met4 ;
        RECT 68.520000 84.845000 68.840000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 85.255000 68.840000 85.575000 ;
      LAYER met4 ;
        RECT 68.520000 85.255000 68.840000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 85.665000 68.840000 85.985000 ;
      LAYER met4 ;
        RECT 68.520000 85.665000 68.840000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 86.075000 68.840000 86.395000 ;
      LAYER met4 ;
        RECT 68.520000 86.075000 68.840000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 86.485000 68.840000 86.805000 ;
      LAYER met4 ;
        RECT 68.520000 86.485000 68.840000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 86.895000 68.840000 87.215000 ;
      LAYER met4 ;
        RECT 68.520000 86.895000 68.840000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 87.305000 68.840000 87.625000 ;
      LAYER met4 ;
        RECT 68.520000 87.305000 68.840000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 87.715000 68.840000 88.035000 ;
      LAYER met4 ;
        RECT 68.520000 87.715000 68.840000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 88.125000 68.840000 88.445000 ;
      LAYER met4 ;
        RECT 68.520000 88.125000 68.840000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 88.535000 68.840000 88.855000 ;
      LAYER met4 ;
        RECT 68.520000 88.535000 68.840000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 88.945000 68.840000 89.265000 ;
      LAYER met4 ;
        RECT 68.520000 88.945000 68.840000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 89.355000 68.840000 89.675000 ;
      LAYER met4 ;
        RECT 68.520000 89.355000 68.840000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 89.765000 68.840000 90.085000 ;
      LAYER met4 ;
        RECT 68.520000 89.765000 68.840000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 90.175000 68.840000 90.495000 ;
      LAYER met4 ;
        RECT 68.520000 90.175000 68.840000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 90.585000 68.840000 90.905000 ;
      LAYER met4 ;
        RECT 68.520000 90.585000 68.840000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 90.995000 68.840000 91.315000 ;
      LAYER met4 ;
        RECT 68.520000 90.995000 68.840000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 91.405000 68.840000 91.725000 ;
      LAYER met4 ;
        RECT 68.520000 91.405000 68.840000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 91.815000 68.840000 92.135000 ;
      LAYER met4 ;
        RECT 68.520000 91.815000 68.840000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 92.225000 68.840000 92.545000 ;
      LAYER met4 ;
        RECT 68.520000 92.225000 68.840000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520000 92.635000 68.840000 92.955000 ;
      LAYER met4 ;
        RECT 68.520000 92.635000 68.840000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 68.065000 68.870000 68.385000 ;
      LAYER met4 ;
        RECT 68.550000 68.065000 68.870000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 68.475000 68.870000 68.795000 ;
      LAYER met4 ;
        RECT 68.550000 68.475000 68.870000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 68.885000 68.870000 69.205000 ;
      LAYER met4 ;
        RECT 68.550000 68.885000 68.870000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 69.295000 68.870000 69.615000 ;
      LAYER met4 ;
        RECT 68.550000 69.295000 68.870000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 69.705000 68.870000 70.025000 ;
      LAYER met4 ;
        RECT 68.550000 69.705000 68.870000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 70.115000 68.870000 70.435000 ;
      LAYER met4 ;
        RECT 68.550000 70.115000 68.870000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 70.525000 68.870000 70.845000 ;
      LAYER met4 ;
        RECT 68.550000 70.525000 68.870000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 70.935000 68.870000 71.255000 ;
      LAYER met4 ;
        RECT 68.550000 70.935000 68.870000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 71.345000 68.870000 71.665000 ;
      LAYER met4 ;
        RECT 68.550000 71.345000 68.870000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 71.755000 68.870000 72.075000 ;
      LAYER met4 ;
        RECT 68.550000 71.755000 68.870000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 72.165000 68.870000 72.485000 ;
      LAYER met4 ;
        RECT 68.550000 72.165000 68.870000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 72.575000 68.870000 72.895000 ;
      LAYER met4 ;
        RECT 68.550000 72.575000 68.870000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 72.985000 68.870000 73.305000 ;
      LAYER met4 ;
        RECT 68.550000 72.985000 68.870000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 73.390000 68.870000 73.710000 ;
      LAYER met4 ;
        RECT 68.550000 73.390000 68.870000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 73.795000 68.870000 74.115000 ;
      LAYER met4 ;
        RECT 68.550000 73.795000 68.870000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 74.200000 68.870000 74.520000 ;
      LAYER met4 ;
        RECT 68.550000 74.200000 68.870000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 74.605000 68.870000 74.925000 ;
      LAYER met4 ;
        RECT 68.550000 74.605000 68.870000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 75.010000 68.870000 75.330000 ;
      LAYER met4 ;
        RECT 68.550000 75.010000 68.870000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 75.415000 68.870000 75.735000 ;
      LAYER met4 ;
        RECT 68.550000 75.415000 68.870000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 75.820000 68.870000 76.140000 ;
      LAYER met4 ;
        RECT 68.550000 75.820000 68.870000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 76.225000 68.870000 76.545000 ;
      LAYER met4 ;
        RECT 68.550000 76.225000 68.870000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 76.630000 68.870000 76.950000 ;
      LAYER met4 ;
        RECT 68.550000 76.630000 68.870000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 77.035000 68.870000 77.355000 ;
      LAYER met4 ;
        RECT 68.550000 77.035000 68.870000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 77.440000 68.870000 77.760000 ;
      LAYER met4 ;
        RECT 68.550000 77.440000 68.870000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 77.845000 68.870000 78.165000 ;
      LAYER met4 ;
        RECT 68.550000 77.845000 68.870000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 78.250000 68.870000 78.570000 ;
      LAYER met4 ;
        RECT 68.550000 78.250000 68.870000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 78.655000 68.870000 78.975000 ;
      LAYER met4 ;
        RECT 68.550000 78.655000 68.870000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 79.060000 68.870000 79.380000 ;
      LAYER met4 ;
        RECT 68.550000 79.060000 68.870000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 79.465000 68.870000 79.785000 ;
      LAYER met4 ;
        RECT 68.550000 79.465000 68.870000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 79.870000 68.870000 80.190000 ;
      LAYER met4 ;
        RECT 68.550000 79.870000 68.870000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 80.275000 68.870000 80.595000 ;
      LAYER met4 ;
        RECT 68.550000 80.275000 68.870000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 80.680000 68.870000 81.000000 ;
      LAYER met4 ;
        RECT 68.550000 80.680000 68.870000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 81.085000 68.870000 81.405000 ;
      LAYER met4 ;
        RECT 68.550000 81.085000 68.870000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 81.490000 68.870000 81.810000 ;
      LAYER met4 ;
        RECT 68.550000 81.490000 68.870000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 81.895000 68.870000 82.215000 ;
      LAYER met4 ;
        RECT 68.550000 81.895000 68.870000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.550000 82.300000 68.870000 82.620000 ;
      LAYER met4 ;
        RECT 68.550000 82.300000 68.870000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.605000 17.800000 68.925000 18.120000 ;
      LAYER met4 ;
        RECT 68.605000 17.800000 68.925000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.605000 18.230000 68.925000 18.550000 ;
      LAYER met4 ;
        RECT 68.605000 18.230000 68.925000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.605000 18.660000 68.925000 18.980000 ;
      LAYER met4 ;
        RECT 68.605000 18.660000 68.925000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.605000 19.090000 68.925000 19.410000 ;
      LAYER met4 ;
        RECT 68.605000 19.090000 68.925000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.605000 19.520000 68.925000 19.840000 ;
      LAYER met4 ;
        RECT 68.605000 19.520000 68.925000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.605000 19.950000 68.925000 20.270000 ;
      LAYER met4 ;
        RECT 68.605000 19.950000 68.925000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.605000 20.380000 68.925000 20.700000 ;
      LAYER met4 ;
        RECT 68.605000 20.380000 68.925000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.605000 20.810000 68.925000 21.130000 ;
      LAYER met4 ;
        RECT 68.605000 20.810000 68.925000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.605000 21.240000 68.925000 21.560000 ;
      LAYER met4 ;
        RECT 68.605000 21.240000 68.925000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.605000 21.670000 68.925000 21.990000 ;
      LAYER met4 ;
        RECT 68.605000 21.670000 68.925000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.605000 22.100000 68.925000 22.420000 ;
      LAYER met4 ;
        RECT 68.605000 22.100000 68.925000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 82.795000 69.250000 83.115000 ;
      LAYER met4 ;
        RECT 68.930000 82.795000 69.250000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 83.205000 69.250000 83.525000 ;
      LAYER met4 ;
        RECT 68.930000 83.205000 69.250000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 83.615000 69.250000 83.935000 ;
      LAYER met4 ;
        RECT 68.930000 83.615000 69.250000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 84.025000 69.250000 84.345000 ;
      LAYER met4 ;
        RECT 68.930000 84.025000 69.250000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 84.435000 69.250000 84.755000 ;
      LAYER met4 ;
        RECT 68.930000 84.435000 69.250000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 84.845000 69.250000 85.165000 ;
      LAYER met4 ;
        RECT 68.930000 84.845000 69.250000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 85.255000 69.250000 85.575000 ;
      LAYER met4 ;
        RECT 68.930000 85.255000 69.250000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 85.665000 69.250000 85.985000 ;
      LAYER met4 ;
        RECT 68.930000 85.665000 69.250000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 86.075000 69.250000 86.395000 ;
      LAYER met4 ;
        RECT 68.930000 86.075000 69.250000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 86.485000 69.250000 86.805000 ;
      LAYER met4 ;
        RECT 68.930000 86.485000 69.250000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 86.895000 69.250000 87.215000 ;
      LAYER met4 ;
        RECT 68.930000 86.895000 69.250000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 87.305000 69.250000 87.625000 ;
      LAYER met4 ;
        RECT 68.930000 87.305000 69.250000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 87.715000 69.250000 88.035000 ;
      LAYER met4 ;
        RECT 68.930000 87.715000 69.250000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 88.125000 69.250000 88.445000 ;
      LAYER met4 ;
        RECT 68.930000 88.125000 69.250000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 88.535000 69.250000 88.855000 ;
      LAYER met4 ;
        RECT 68.930000 88.535000 69.250000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 88.945000 69.250000 89.265000 ;
      LAYER met4 ;
        RECT 68.930000 88.945000 69.250000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 89.355000 69.250000 89.675000 ;
      LAYER met4 ;
        RECT 68.930000 89.355000 69.250000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 89.765000 69.250000 90.085000 ;
      LAYER met4 ;
        RECT 68.930000 89.765000 69.250000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 90.175000 69.250000 90.495000 ;
      LAYER met4 ;
        RECT 68.930000 90.175000 69.250000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 90.585000 69.250000 90.905000 ;
      LAYER met4 ;
        RECT 68.930000 90.585000 69.250000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 90.995000 69.250000 91.315000 ;
      LAYER met4 ;
        RECT 68.930000 90.995000 69.250000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 91.405000 69.250000 91.725000 ;
      LAYER met4 ;
        RECT 68.930000 91.405000 69.250000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 91.815000 69.250000 92.135000 ;
      LAYER met4 ;
        RECT 68.930000 91.815000 69.250000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 92.225000 69.250000 92.545000 ;
      LAYER met4 ;
        RECT 68.930000 92.225000 69.250000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930000 92.635000 69.250000 92.955000 ;
      LAYER met4 ;
        RECT 68.930000 92.635000 69.250000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 68.065000 69.270000 68.385000 ;
      LAYER met4 ;
        RECT 68.950000 68.065000 69.270000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 68.475000 69.270000 68.795000 ;
      LAYER met4 ;
        RECT 68.950000 68.475000 69.270000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 68.885000 69.270000 69.205000 ;
      LAYER met4 ;
        RECT 68.950000 68.885000 69.270000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 69.295000 69.270000 69.615000 ;
      LAYER met4 ;
        RECT 68.950000 69.295000 69.270000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 69.705000 69.270000 70.025000 ;
      LAYER met4 ;
        RECT 68.950000 69.705000 69.270000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 70.115000 69.270000 70.435000 ;
      LAYER met4 ;
        RECT 68.950000 70.115000 69.270000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 70.525000 69.270000 70.845000 ;
      LAYER met4 ;
        RECT 68.950000 70.525000 69.270000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 70.935000 69.270000 71.255000 ;
      LAYER met4 ;
        RECT 68.950000 70.935000 69.270000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 71.345000 69.270000 71.665000 ;
      LAYER met4 ;
        RECT 68.950000 71.345000 69.270000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 71.755000 69.270000 72.075000 ;
      LAYER met4 ;
        RECT 68.950000 71.755000 69.270000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 72.165000 69.270000 72.485000 ;
      LAYER met4 ;
        RECT 68.950000 72.165000 69.270000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 72.575000 69.270000 72.895000 ;
      LAYER met4 ;
        RECT 68.950000 72.575000 69.270000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 72.985000 69.270000 73.305000 ;
      LAYER met4 ;
        RECT 68.950000 72.985000 69.270000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 73.390000 69.270000 73.710000 ;
      LAYER met4 ;
        RECT 68.950000 73.390000 69.270000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 73.795000 69.270000 74.115000 ;
      LAYER met4 ;
        RECT 68.950000 73.795000 69.270000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 74.200000 69.270000 74.520000 ;
      LAYER met4 ;
        RECT 68.950000 74.200000 69.270000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 74.605000 69.270000 74.925000 ;
      LAYER met4 ;
        RECT 68.950000 74.605000 69.270000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 75.010000 69.270000 75.330000 ;
      LAYER met4 ;
        RECT 68.950000 75.010000 69.270000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 75.415000 69.270000 75.735000 ;
      LAYER met4 ;
        RECT 68.950000 75.415000 69.270000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 75.820000 69.270000 76.140000 ;
      LAYER met4 ;
        RECT 68.950000 75.820000 69.270000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 76.225000 69.270000 76.545000 ;
      LAYER met4 ;
        RECT 68.950000 76.225000 69.270000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 76.630000 69.270000 76.950000 ;
      LAYER met4 ;
        RECT 68.950000 76.630000 69.270000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 77.035000 69.270000 77.355000 ;
      LAYER met4 ;
        RECT 68.950000 77.035000 69.270000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 77.440000 69.270000 77.760000 ;
      LAYER met4 ;
        RECT 68.950000 77.440000 69.270000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 77.845000 69.270000 78.165000 ;
      LAYER met4 ;
        RECT 68.950000 77.845000 69.270000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 78.250000 69.270000 78.570000 ;
      LAYER met4 ;
        RECT 68.950000 78.250000 69.270000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 78.655000 69.270000 78.975000 ;
      LAYER met4 ;
        RECT 68.950000 78.655000 69.270000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 79.060000 69.270000 79.380000 ;
      LAYER met4 ;
        RECT 68.950000 79.060000 69.270000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 79.465000 69.270000 79.785000 ;
      LAYER met4 ;
        RECT 68.950000 79.465000 69.270000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 79.870000 69.270000 80.190000 ;
      LAYER met4 ;
        RECT 68.950000 79.870000 69.270000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 80.275000 69.270000 80.595000 ;
      LAYER met4 ;
        RECT 68.950000 80.275000 69.270000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 80.680000 69.270000 81.000000 ;
      LAYER met4 ;
        RECT 68.950000 80.680000 69.270000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 81.085000 69.270000 81.405000 ;
      LAYER met4 ;
        RECT 68.950000 81.085000 69.270000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 81.490000 69.270000 81.810000 ;
      LAYER met4 ;
        RECT 68.950000 81.490000 69.270000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 81.895000 69.270000 82.215000 ;
      LAYER met4 ;
        RECT 68.950000 81.895000 69.270000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.950000 82.300000 69.270000 82.620000 ;
      LAYER met4 ;
        RECT 68.950000 82.300000 69.270000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010000 17.800000 69.330000 18.120000 ;
      LAYER met4 ;
        RECT 69.010000 17.800000 69.330000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010000 18.230000 69.330000 18.550000 ;
      LAYER met4 ;
        RECT 69.010000 18.230000 69.330000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010000 18.660000 69.330000 18.980000 ;
      LAYER met4 ;
        RECT 69.010000 18.660000 69.330000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010000 19.090000 69.330000 19.410000 ;
      LAYER met4 ;
        RECT 69.010000 19.090000 69.330000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010000 19.520000 69.330000 19.840000 ;
      LAYER met4 ;
        RECT 69.010000 19.520000 69.330000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010000 19.950000 69.330000 20.270000 ;
      LAYER met4 ;
        RECT 69.010000 19.950000 69.330000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010000 20.380000 69.330000 20.700000 ;
      LAYER met4 ;
        RECT 69.010000 20.380000 69.330000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010000 20.810000 69.330000 21.130000 ;
      LAYER met4 ;
        RECT 69.010000 20.810000 69.330000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010000 21.240000 69.330000 21.560000 ;
      LAYER met4 ;
        RECT 69.010000 21.240000 69.330000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010000 21.670000 69.330000 21.990000 ;
      LAYER met4 ;
        RECT 69.010000 21.670000 69.330000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010000 22.100000 69.330000 22.420000 ;
      LAYER met4 ;
        RECT 69.010000 22.100000 69.330000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 82.795000 69.660000 83.115000 ;
      LAYER met4 ;
        RECT 69.340000 82.795000 69.660000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 83.205000 69.660000 83.525000 ;
      LAYER met4 ;
        RECT 69.340000 83.205000 69.660000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 83.615000 69.660000 83.935000 ;
      LAYER met4 ;
        RECT 69.340000 83.615000 69.660000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 84.025000 69.660000 84.345000 ;
      LAYER met4 ;
        RECT 69.340000 84.025000 69.660000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 84.435000 69.660000 84.755000 ;
      LAYER met4 ;
        RECT 69.340000 84.435000 69.660000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 84.845000 69.660000 85.165000 ;
      LAYER met4 ;
        RECT 69.340000 84.845000 69.660000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 85.255000 69.660000 85.575000 ;
      LAYER met4 ;
        RECT 69.340000 85.255000 69.660000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 85.665000 69.660000 85.985000 ;
      LAYER met4 ;
        RECT 69.340000 85.665000 69.660000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 86.075000 69.660000 86.395000 ;
      LAYER met4 ;
        RECT 69.340000 86.075000 69.660000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 86.485000 69.660000 86.805000 ;
      LAYER met4 ;
        RECT 69.340000 86.485000 69.660000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 86.895000 69.660000 87.215000 ;
      LAYER met4 ;
        RECT 69.340000 86.895000 69.660000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 87.305000 69.660000 87.625000 ;
      LAYER met4 ;
        RECT 69.340000 87.305000 69.660000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 87.715000 69.660000 88.035000 ;
      LAYER met4 ;
        RECT 69.340000 87.715000 69.660000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 88.125000 69.660000 88.445000 ;
      LAYER met4 ;
        RECT 69.340000 88.125000 69.660000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 88.535000 69.660000 88.855000 ;
      LAYER met4 ;
        RECT 69.340000 88.535000 69.660000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 88.945000 69.660000 89.265000 ;
      LAYER met4 ;
        RECT 69.340000 88.945000 69.660000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 89.355000 69.660000 89.675000 ;
      LAYER met4 ;
        RECT 69.340000 89.355000 69.660000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 89.765000 69.660000 90.085000 ;
      LAYER met4 ;
        RECT 69.340000 89.765000 69.660000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 90.175000 69.660000 90.495000 ;
      LAYER met4 ;
        RECT 69.340000 90.175000 69.660000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 90.585000 69.660000 90.905000 ;
      LAYER met4 ;
        RECT 69.340000 90.585000 69.660000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 90.995000 69.660000 91.315000 ;
      LAYER met4 ;
        RECT 69.340000 90.995000 69.660000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 91.405000 69.660000 91.725000 ;
      LAYER met4 ;
        RECT 69.340000 91.405000 69.660000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 91.815000 69.660000 92.135000 ;
      LAYER met4 ;
        RECT 69.340000 91.815000 69.660000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 92.225000 69.660000 92.545000 ;
      LAYER met4 ;
        RECT 69.340000 92.225000 69.660000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340000 92.635000 69.660000 92.955000 ;
      LAYER met4 ;
        RECT 69.340000 92.635000 69.660000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 68.065000 69.670000 68.385000 ;
      LAYER met4 ;
        RECT 69.350000 68.065000 69.670000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 68.475000 69.670000 68.795000 ;
      LAYER met4 ;
        RECT 69.350000 68.475000 69.670000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 68.885000 69.670000 69.205000 ;
      LAYER met4 ;
        RECT 69.350000 68.885000 69.670000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 69.295000 69.670000 69.615000 ;
      LAYER met4 ;
        RECT 69.350000 69.295000 69.670000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 69.705000 69.670000 70.025000 ;
      LAYER met4 ;
        RECT 69.350000 69.705000 69.670000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 70.115000 69.670000 70.435000 ;
      LAYER met4 ;
        RECT 69.350000 70.115000 69.670000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 70.525000 69.670000 70.845000 ;
      LAYER met4 ;
        RECT 69.350000 70.525000 69.670000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 70.935000 69.670000 71.255000 ;
      LAYER met4 ;
        RECT 69.350000 70.935000 69.670000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 71.345000 69.670000 71.665000 ;
      LAYER met4 ;
        RECT 69.350000 71.345000 69.670000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 71.755000 69.670000 72.075000 ;
      LAYER met4 ;
        RECT 69.350000 71.755000 69.670000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 72.165000 69.670000 72.485000 ;
      LAYER met4 ;
        RECT 69.350000 72.165000 69.670000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 72.575000 69.670000 72.895000 ;
      LAYER met4 ;
        RECT 69.350000 72.575000 69.670000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 72.985000 69.670000 73.305000 ;
      LAYER met4 ;
        RECT 69.350000 72.985000 69.670000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 73.390000 69.670000 73.710000 ;
      LAYER met4 ;
        RECT 69.350000 73.390000 69.670000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 73.795000 69.670000 74.115000 ;
      LAYER met4 ;
        RECT 69.350000 73.795000 69.670000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 74.200000 69.670000 74.520000 ;
      LAYER met4 ;
        RECT 69.350000 74.200000 69.670000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 74.605000 69.670000 74.925000 ;
      LAYER met4 ;
        RECT 69.350000 74.605000 69.670000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 75.010000 69.670000 75.330000 ;
      LAYER met4 ;
        RECT 69.350000 75.010000 69.670000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 75.415000 69.670000 75.735000 ;
      LAYER met4 ;
        RECT 69.350000 75.415000 69.670000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 75.820000 69.670000 76.140000 ;
      LAYER met4 ;
        RECT 69.350000 75.820000 69.670000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 76.225000 69.670000 76.545000 ;
      LAYER met4 ;
        RECT 69.350000 76.225000 69.670000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 76.630000 69.670000 76.950000 ;
      LAYER met4 ;
        RECT 69.350000 76.630000 69.670000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 77.035000 69.670000 77.355000 ;
      LAYER met4 ;
        RECT 69.350000 77.035000 69.670000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 77.440000 69.670000 77.760000 ;
      LAYER met4 ;
        RECT 69.350000 77.440000 69.670000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 77.845000 69.670000 78.165000 ;
      LAYER met4 ;
        RECT 69.350000 77.845000 69.670000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 78.250000 69.670000 78.570000 ;
      LAYER met4 ;
        RECT 69.350000 78.250000 69.670000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 78.655000 69.670000 78.975000 ;
      LAYER met4 ;
        RECT 69.350000 78.655000 69.670000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 79.060000 69.670000 79.380000 ;
      LAYER met4 ;
        RECT 69.350000 79.060000 69.670000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 79.465000 69.670000 79.785000 ;
      LAYER met4 ;
        RECT 69.350000 79.465000 69.670000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 79.870000 69.670000 80.190000 ;
      LAYER met4 ;
        RECT 69.350000 79.870000 69.670000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 80.275000 69.670000 80.595000 ;
      LAYER met4 ;
        RECT 69.350000 80.275000 69.670000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 80.680000 69.670000 81.000000 ;
      LAYER met4 ;
        RECT 69.350000 80.680000 69.670000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 81.085000 69.670000 81.405000 ;
      LAYER met4 ;
        RECT 69.350000 81.085000 69.670000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 81.490000 69.670000 81.810000 ;
      LAYER met4 ;
        RECT 69.350000 81.490000 69.670000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 81.895000 69.670000 82.215000 ;
      LAYER met4 ;
        RECT 69.350000 81.895000 69.670000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.350000 82.300000 69.670000 82.620000 ;
      LAYER met4 ;
        RECT 69.350000 82.300000 69.670000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.415000 17.800000 69.735000 18.120000 ;
      LAYER met4 ;
        RECT 69.415000 17.800000 69.735000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.415000 18.230000 69.735000 18.550000 ;
      LAYER met4 ;
        RECT 69.415000 18.230000 69.735000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.415000 18.660000 69.735000 18.980000 ;
      LAYER met4 ;
        RECT 69.415000 18.660000 69.735000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.415000 19.090000 69.735000 19.410000 ;
      LAYER met4 ;
        RECT 69.415000 19.090000 69.735000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.415000 19.520000 69.735000 19.840000 ;
      LAYER met4 ;
        RECT 69.415000 19.520000 69.735000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.415000 19.950000 69.735000 20.270000 ;
      LAYER met4 ;
        RECT 69.415000 19.950000 69.735000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.415000 20.380000 69.735000 20.700000 ;
      LAYER met4 ;
        RECT 69.415000 20.380000 69.735000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.415000 20.810000 69.735000 21.130000 ;
      LAYER met4 ;
        RECT 69.415000 20.810000 69.735000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.415000 21.240000 69.735000 21.560000 ;
      LAYER met4 ;
        RECT 69.415000 21.240000 69.735000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.415000 21.670000 69.735000 21.990000 ;
      LAYER met4 ;
        RECT 69.415000 21.670000 69.735000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.415000 22.100000 69.735000 22.420000 ;
      LAYER met4 ;
        RECT 69.415000 22.100000 69.735000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 68.065000 70.070000 68.385000 ;
      LAYER met4 ;
        RECT 69.750000 68.065000 70.070000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 68.475000 70.070000 68.795000 ;
      LAYER met4 ;
        RECT 69.750000 68.475000 70.070000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 68.885000 70.070000 69.205000 ;
      LAYER met4 ;
        RECT 69.750000 68.885000 70.070000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 69.295000 70.070000 69.615000 ;
      LAYER met4 ;
        RECT 69.750000 69.295000 70.070000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 69.705000 70.070000 70.025000 ;
      LAYER met4 ;
        RECT 69.750000 69.705000 70.070000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 70.115000 70.070000 70.435000 ;
      LAYER met4 ;
        RECT 69.750000 70.115000 70.070000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 70.525000 70.070000 70.845000 ;
      LAYER met4 ;
        RECT 69.750000 70.525000 70.070000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 70.935000 70.070000 71.255000 ;
      LAYER met4 ;
        RECT 69.750000 70.935000 70.070000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 71.345000 70.070000 71.665000 ;
      LAYER met4 ;
        RECT 69.750000 71.345000 70.070000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 71.755000 70.070000 72.075000 ;
      LAYER met4 ;
        RECT 69.750000 71.755000 70.070000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 72.165000 70.070000 72.485000 ;
      LAYER met4 ;
        RECT 69.750000 72.165000 70.070000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 72.575000 70.070000 72.895000 ;
      LAYER met4 ;
        RECT 69.750000 72.575000 70.070000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 72.985000 70.070000 73.305000 ;
      LAYER met4 ;
        RECT 69.750000 72.985000 70.070000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 73.390000 70.070000 73.710000 ;
      LAYER met4 ;
        RECT 69.750000 73.390000 70.070000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 73.795000 70.070000 74.115000 ;
      LAYER met4 ;
        RECT 69.750000 73.795000 70.070000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 74.200000 70.070000 74.520000 ;
      LAYER met4 ;
        RECT 69.750000 74.200000 70.070000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 74.605000 70.070000 74.925000 ;
      LAYER met4 ;
        RECT 69.750000 74.605000 70.070000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 75.010000 70.070000 75.330000 ;
      LAYER met4 ;
        RECT 69.750000 75.010000 70.070000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 75.415000 70.070000 75.735000 ;
      LAYER met4 ;
        RECT 69.750000 75.415000 70.070000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 75.820000 70.070000 76.140000 ;
      LAYER met4 ;
        RECT 69.750000 75.820000 70.070000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 76.225000 70.070000 76.545000 ;
      LAYER met4 ;
        RECT 69.750000 76.225000 70.070000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 76.630000 70.070000 76.950000 ;
      LAYER met4 ;
        RECT 69.750000 76.630000 70.070000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 77.035000 70.070000 77.355000 ;
      LAYER met4 ;
        RECT 69.750000 77.035000 70.070000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 77.440000 70.070000 77.760000 ;
      LAYER met4 ;
        RECT 69.750000 77.440000 70.070000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 77.845000 70.070000 78.165000 ;
      LAYER met4 ;
        RECT 69.750000 77.845000 70.070000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 78.250000 70.070000 78.570000 ;
      LAYER met4 ;
        RECT 69.750000 78.250000 70.070000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 78.655000 70.070000 78.975000 ;
      LAYER met4 ;
        RECT 69.750000 78.655000 70.070000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 79.060000 70.070000 79.380000 ;
      LAYER met4 ;
        RECT 69.750000 79.060000 70.070000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 79.465000 70.070000 79.785000 ;
      LAYER met4 ;
        RECT 69.750000 79.465000 70.070000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 79.870000 70.070000 80.190000 ;
      LAYER met4 ;
        RECT 69.750000 79.870000 70.070000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 80.275000 70.070000 80.595000 ;
      LAYER met4 ;
        RECT 69.750000 80.275000 70.070000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 80.680000 70.070000 81.000000 ;
      LAYER met4 ;
        RECT 69.750000 80.680000 70.070000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 81.085000 70.070000 81.405000 ;
      LAYER met4 ;
        RECT 69.750000 81.085000 70.070000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 81.490000 70.070000 81.810000 ;
      LAYER met4 ;
        RECT 69.750000 81.490000 70.070000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 81.895000 70.070000 82.215000 ;
      LAYER met4 ;
        RECT 69.750000 81.895000 70.070000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 82.300000 70.070000 82.620000 ;
      LAYER met4 ;
        RECT 69.750000 82.300000 70.070000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 82.795000 70.070000 83.115000 ;
      LAYER met4 ;
        RECT 69.750000 82.795000 70.070000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 83.205000 70.070000 83.525000 ;
      LAYER met4 ;
        RECT 69.750000 83.205000 70.070000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 83.615000 70.070000 83.935000 ;
      LAYER met4 ;
        RECT 69.750000 83.615000 70.070000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 84.025000 70.070000 84.345000 ;
      LAYER met4 ;
        RECT 69.750000 84.025000 70.070000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 84.435000 70.070000 84.755000 ;
      LAYER met4 ;
        RECT 69.750000 84.435000 70.070000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 84.845000 70.070000 85.165000 ;
      LAYER met4 ;
        RECT 69.750000 84.845000 70.070000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 85.255000 70.070000 85.575000 ;
      LAYER met4 ;
        RECT 69.750000 85.255000 70.070000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 85.665000 70.070000 85.985000 ;
      LAYER met4 ;
        RECT 69.750000 85.665000 70.070000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 86.075000 70.070000 86.395000 ;
      LAYER met4 ;
        RECT 69.750000 86.075000 70.070000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 86.485000 70.070000 86.805000 ;
      LAYER met4 ;
        RECT 69.750000 86.485000 70.070000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 86.895000 70.070000 87.215000 ;
      LAYER met4 ;
        RECT 69.750000 86.895000 70.070000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 87.305000 70.070000 87.625000 ;
      LAYER met4 ;
        RECT 69.750000 87.305000 70.070000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 87.715000 70.070000 88.035000 ;
      LAYER met4 ;
        RECT 69.750000 87.715000 70.070000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 88.125000 70.070000 88.445000 ;
      LAYER met4 ;
        RECT 69.750000 88.125000 70.070000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 88.535000 70.070000 88.855000 ;
      LAYER met4 ;
        RECT 69.750000 88.535000 70.070000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 88.945000 70.070000 89.265000 ;
      LAYER met4 ;
        RECT 69.750000 88.945000 70.070000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 89.355000 70.070000 89.675000 ;
      LAYER met4 ;
        RECT 69.750000 89.355000 70.070000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 89.765000 70.070000 90.085000 ;
      LAYER met4 ;
        RECT 69.750000 89.765000 70.070000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 90.175000 70.070000 90.495000 ;
      LAYER met4 ;
        RECT 69.750000 90.175000 70.070000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 90.585000 70.070000 90.905000 ;
      LAYER met4 ;
        RECT 69.750000 90.585000 70.070000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 90.995000 70.070000 91.315000 ;
      LAYER met4 ;
        RECT 69.750000 90.995000 70.070000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 91.405000 70.070000 91.725000 ;
      LAYER met4 ;
        RECT 69.750000 91.405000 70.070000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 91.815000 70.070000 92.135000 ;
      LAYER met4 ;
        RECT 69.750000 91.815000 70.070000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 92.225000 70.070000 92.545000 ;
      LAYER met4 ;
        RECT 69.750000 92.225000 70.070000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750000 92.635000 70.070000 92.955000 ;
      LAYER met4 ;
        RECT 69.750000 92.635000 70.070000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.820000 17.800000 70.140000 18.120000 ;
      LAYER met4 ;
        RECT 69.820000 17.800000 70.140000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.820000 18.230000 70.140000 18.550000 ;
      LAYER met4 ;
        RECT 69.820000 18.230000 70.140000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.820000 18.660000 70.140000 18.980000 ;
      LAYER met4 ;
        RECT 69.820000 18.660000 70.140000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.820000 19.090000 70.140000 19.410000 ;
      LAYER met4 ;
        RECT 69.820000 19.090000 70.140000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.820000 19.520000 70.140000 19.840000 ;
      LAYER met4 ;
        RECT 69.820000 19.520000 70.140000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.820000 19.950000 70.140000 20.270000 ;
      LAYER met4 ;
        RECT 69.820000 19.950000 70.140000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.820000 20.380000 70.140000 20.700000 ;
      LAYER met4 ;
        RECT 69.820000 20.380000 70.140000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.820000 20.810000 70.140000 21.130000 ;
      LAYER met4 ;
        RECT 69.820000 20.810000 70.140000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.820000 21.240000 70.140000 21.560000 ;
      LAYER met4 ;
        RECT 69.820000 21.240000 70.140000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.820000 21.670000 70.140000 21.990000 ;
      LAYER met4 ;
        RECT 69.820000 21.670000 70.140000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.820000 22.100000 70.140000 22.420000 ;
      LAYER met4 ;
        RECT 69.820000 22.100000 70.140000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110000 17.800000 7.430000 18.120000 ;
      LAYER met4 ;
        RECT 7.110000 17.800000 7.430000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110000 18.230000 7.430000 18.550000 ;
      LAYER met4 ;
        RECT 7.110000 18.230000 7.430000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110000 18.660000 7.430000 18.980000 ;
      LAYER met4 ;
        RECT 7.110000 18.660000 7.430000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110000 19.090000 7.430000 19.410000 ;
      LAYER met4 ;
        RECT 7.110000 19.090000 7.430000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110000 19.520000 7.430000 19.840000 ;
      LAYER met4 ;
        RECT 7.110000 19.520000 7.430000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110000 19.950000 7.430000 20.270000 ;
      LAYER met4 ;
        RECT 7.110000 19.950000 7.430000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110000 20.380000 7.430000 20.700000 ;
      LAYER met4 ;
        RECT 7.110000 20.380000 7.430000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110000 20.810000 7.430000 21.130000 ;
      LAYER met4 ;
        RECT 7.110000 20.810000 7.430000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110000 21.240000 7.430000 21.560000 ;
      LAYER met4 ;
        RECT 7.110000 21.240000 7.430000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110000 21.670000 7.430000 21.990000 ;
      LAYER met4 ;
        RECT 7.110000 21.670000 7.430000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110000 22.100000 7.430000 22.420000 ;
      LAYER met4 ;
        RECT 7.110000 22.100000 7.430000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 68.065000 7.505000 68.385000 ;
      LAYER met4 ;
        RECT 7.185000 68.065000 7.505000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 68.475000 7.505000 68.795000 ;
      LAYER met4 ;
        RECT 7.185000 68.475000 7.505000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 68.885000 7.505000 69.205000 ;
      LAYER met4 ;
        RECT 7.185000 68.885000 7.505000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 69.295000 7.505000 69.615000 ;
      LAYER met4 ;
        RECT 7.185000 69.295000 7.505000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 69.705000 7.505000 70.025000 ;
      LAYER met4 ;
        RECT 7.185000 69.705000 7.505000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 70.115000 7.505000 70.435000 ;
      LAYER met4 ;
        RECT 7.185000 70.115000 7.505000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 70.525000 7.505000 70.845000 ;
      LAYER met4 ;
        RECT 7.185000 70.525000 7.505000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 70.935000 7.505000 71.255000 ;
      LAYER met4 ;
        RECT 7.185000 70.935000 7.505000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 71.345000 7.505000 71.665000 ;
      LAYER met4 ;
        RECT 7.185000 71.345000 7.505000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 71.755000 7.505000 72.075000 ;
      LAYER met4 ;
        RECT 7.185000 71.755000 7.505000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 72.165000 7.505000 72.485000 ;
      LAYER met4 ;
        RECT 7.185000 72.165000 7.505000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 72.575000 7.505000 72.895000 ;
      LAYER met4 ;
        RECT 7.185000 72.575000 7.505000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 72.985000 7.505000 73.305000 ;
      LAYER met4 ;
        RECT 7.185000 72.985000 7.505000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 73.390000 7.505000 73.710000 ;
      LAYER met4 ;
        RECT 7.185000 73.390000 7.505000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 73.795000 7.505000 74.115000 ;
      LAYER met4 ;
        RECT 7.185000 73.795000 7.505000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 74.200000 7.505000 74.520000 ;
      LAYER met4 ;
        RECT 7.185000 74.200000 7.505000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 74.605000 7.505000 74.925000 ;
      LAYER met4 ;
        RECT 7.185000 74.605000 7.505000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 75.010000 7.505000 75.330000 ;
      LAYER met4 ;
        RECT 7.185000 75.010000 7.505000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 75.415000 7.505000 75.735000 ;
      LAYER met4 ;
        RECT 7.185000 75.415000 7.505000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 75.820000 7.505000 76.140000 ;
      LAYER met4 ;
        RECT 7.185000 75.820000 7.505000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 76.225000 7.505000 76.545000 ;
      LAYER met4 ;
        RECT 7.185000 76.225000 7.505000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 76.630000 7.505000 76.950000 ;
      LAYER met4 ;
        RECT 7.185000 76.630000 7.505000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 77.035000 7.505000 77.355000 ;
      LAYER met4 ;
        RECT 7.185000 77.035000 7.505000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 77.440000 7.505000 77.760000 ;
      LAYER met4 ;
        RECT 7.185000 77.440000 7.505000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 77.845000 7.505000 78.165000 ;
      LAYER met4 ;
        RECT 7.185000 77.845000 7.505000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 78.250000 7.505000 78.570000 ;
      LAYER met4 ;
        RECT 7.185000 78.250000 7.505000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 78.655000 7.505000 78.975000 ;
      LAYER met4 ;
        RECT 7.185000 78.655000 7.505000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 79.060000 7.505000 79.380000 ;
      LAYER met4 ;
        RECT 7.185000 79.060000 7.505000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 79.465000 7.505000 79.785000 ;
      LAYER met4 ;
        RECT 7.185000 79.465000 7.505000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 79.870000 7.505000 80.190000 ;
      LAYER met4 ;
        RECT 7.185000 79.870000 7.505000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 80.275000 7.505000 80.595000 ;
      LAYER met4 ;
        RECT 7.185000 80.275000 7.505000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 80.680000 7.505000 81.000000 ;
      LAYER met4 ;
        RECT 7.185000 80.680000 7.505000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 81.085000 7.505000 81.405000 ;
      LAYER met4 ;
        RECT 7.185000 81.085000 7.505000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 81.490000 7.505000 81.810000 ;
      LAYER met4 ;
        RECT 7.185000 81.490000 7.505000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 81.895000 7.505000 82.215000 ;
      LAYER met4 ;
        RECT 7.185000 81.895000 7.505000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185000 82.300000 7.505000 82.620000 ;
      LAYER met4 ;
        RECT 7.185000 82.300000 7.505000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 82.795000 7.555000 83.115000 ;
      LAYER met4 ;
        RECT 7.235000 82.795000 7.555000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 83.205000 7.555000 83.525000 ;
      LAYER met4 ;
        RECT 7.235000 83.205000 7.555000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 83.615000 7.555000 83.935000 ;
      LAYER met4 ;
        RECT 7.235000 83.615000 7.555000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 84.025000 7.555000 84.345000 ;
      LAYER met4 ;
        RECT 7.235000 84.025000 7.555000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 84.435000 7.555000 84.755000 ;
      LAYER met4 ;
        RECT 7.235000 84.435000 7.555000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 84.845000 7.555000 85.165000 ;
      LAYER met4 ;
        RECT 7.235000 84.845000 7.555000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 85.255000 7.555000 85.575000 ;
      LAYER met4 ;
        RECT 7.235000 85.255000 7.555000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 85.665000 7.555000 85.985000 ;
      LAYER met4 ;
        RECT 7.235000 85.665000 7.555000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 86.075000 7.555000 86.395000 ;
      LAYER met4 ;
        RECT 7.235000 86.075000 7.555000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 86.485000 7.555000 86.805000 ;
      LAYER met4 ;
        RECT 7.235000 86.485000 7.555000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 86.895000 7.555000 87.215000 ;
      LAYER met4 ;
        RECT 7.235000 86.895000 7.555000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 87.305000 7.555000 87.625000 ;
      LAYER met4 ;
        RECT 7.235000 87.305000 7.555000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 87.715000 7.555000 88.035000 ;
      LAYER met4 ;
        RECT 7.235000 87.715000 7.555000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 88.125000 7.555000 88.445000 ;
      LAYER met4 ;
        RECT 7.235000 88.125000 7.555000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 88.535000 7.555000 88.855000 ;
      LAYER met4 ;
        RECT 7.235000 88.535000 7.555000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 88.945000 7.555000 89.265000 ;
      LAYER met4 ;
        RECT 7.235000 88.945000 7.555000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 89.355000 7.555000 89.675000 ;
      LAYER met4 ;
        RECT 7.235000 89.355000 7.555000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 89.765000 7.555000 90.085000 ;
      LAYER met4 ;
        RECT 7.235000 89.765000 7.555000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 90.175000 7.555000 90.495000 ;
      LAYER met4 ;
        RECT 7.235000 90.175000 7.555000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 90.585000 7.555000 90.905000 ;
      LAYER met4 ;
        RECT 7.235000 90.585000 7.555000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 90.995000 7.555000 91.315000 ;
      LAYER met4 ;
        RECT 7.235000 90.995000 7.555000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 91.405000 7.555000 91.725000 ;
      LAYER met4 ;
        RECT 7.235000 91.405000 7.555000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 91.815000 7.555000 92.135000 ;
      LAYER met4 ;
        RECT 7.235000 91.815000 7.555000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 92.225000 7.555000 92.545000 ;
      LAYER met4 ;
        RECT 7.235000 92.225000 7.555000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235000 92.635000 7.555000 92.955000 ;
      LAYER met4 ;
        RECT 7.235000 92.635000 7.555000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515000 17.800000 7.835000 18.120000 ;
      LAYER met4 ;
        RECT 7.515000 17.800000 7.835000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515000 18.230000 7.835000 18.550000 ;
      LAYER met4 ;
        RECT 7.515000 18.230000 7.835000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515000 18.660000 7.835000 18.980000 ;
      LAYER met4 ;
        RECT 7.515000 18.660000 7.835000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515000 19.090000 7.835000 19.410000 ;
      LAYER met4 ;
        RECT 7.515000 19.090000 7.835000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515000 19.520000 7.835000 19.840000 ;
      LAYER met4 ;
        RECT 7.515000 19.520000 7.835000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515000 19.950000 7.835000 20.270000 ;
      LAYER met4 ;
        RECT 7.515000 19.950000 7.835000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515000 20.380000 7.835000 20.700000 ;
      LAYER met4 ;
        RECT 7.515000 20.380000 7.835000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515000 20.810000 7.835000 21.130000 ;
      LAYER met4 ;
        RECT 7.515000 20.810000 7.835000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515000 21.240000 7.835000 21.560000 ;
      LAYER met4 ;
        RECT 7.515000 21.240000 7.835000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515000 21.670000 7.835000 21.990000 ;
      LAYER met4 ;
        RECT 7.515000 21.670000 7.835000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515000 22.100000 7.835000 22.420000 ;
      LAYER met4 ;
        RECT 7.515000 22.100000 7.835000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 68.065000 7.905000 68.385000 ;
      LAYER met4 ;
        RECT 7.585000 68.065000 7.905000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 68.475000 7.905000 68.795000 ;
      LAYER met4 ;
        RECT 7.585000 68.475000 7.905000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 68.885000 7.905000 69.205000 ;
      LAYER met4 ;
        RECT 7.585000 68.885000 7.905000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 69.295000 7.905000 69.615000 ;
      LAYER met4 ;
        RECT 7.585000 69.295000 7.905000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 69.705000 7.905000 70.025000 ;
      LAYER met4 ;
        RECT 7.585000 69.705000 7.905000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 70.115000 7.905000 70.435000 ;
      LAYER met4 ;
        RECT 7.585000 70.115000 7.905000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 70.525000 7.905000 70.845000 ;
      LAYER met4 ;
        RECT 7.585000 70.525000 7.905000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 70.935000 7.905000 71.255000 ;
      LAYER met4 ;
        RECT 7.585000 70.935000 7.905000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 71.345000 7.905000 71.665000 ;
      LAYER met4 ;
        RECT 7.585000 71.345000 7.905000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 71.755000 7.905000 72.075000 ;
      LAYER met4 ;
        RECT 7.585000 71.755000 7.905000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 72.165000 7.905000 72.485000 ;
      LAYER met4 ;
        RECT 7.585000 72.165000 7.905000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 72.575000 7.905000 72.895000 ;
      LAYER met4 ;
        RECT 7.585000 72.575000 7.905000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 72.985000 7.905000 73.305000 ;
      LAYER met4 ;
        RECT 7.585000 72.985000 7.905000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 73.390000 7.905000 73.710000 ;
      LAYER met4 ;
        RECT 7.585000 73.390000 7.905000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 73.795000 7.905000 74.115000 ;
      LAYER met4 ;
        RECT 7.585000 73.795000 7.905000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 74.200000 7.905000 74.520000 ;
      LAYER met4 ;
        RECT 7.585000 74.200000 7.905000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 74.605000 7.905000 74.925000 ;
      LAYER met4 ;
        RECT 7.585000 74.605000 7.905000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 75.010000 7.905000 75.330000 ;
      LAYER met4 ;
        RECT 7.585000 75.010000 7.905000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 75.415000 7.905000 75.735000 ;
      LAYER met4 ;
        RECT 7.585000 75.415000 7.905000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 75.820000 7.905000 76.140000 ;
      LAYER met4 ;
        RECT 7.585000 75.820000 7.905000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 76.225000 7.905000 76.545000 ;
      LAYER met4 ;
        RECT 7.585000 76.225000 7.905000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 76.630000 7.905000 76.950000 ;
      LAYER met4 ;
        RECT 7.585000 76.630000 7.905000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 77.035000 7.905000 77.355000 ;
      LAYER met4 ;
        RECT 7.585000 77.035000 7.905000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 77.440000 7.905000 77.760000 ;
      LAYER met4 ;
        RECT 7.585000 77.440000 7.905000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 77.845000 7.905000 78.165000 ;
      LAYER met4 ;
        RECT 7.585000 77.845000 7.905000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 78.250000 7.905000 78.570000 ;
      LAYER met4 ;
        RECT 7.585000 78.250000 7.905000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 78.655000 7.905000 78.975000 ;
      LAYER met4 ;
        RECT 7.585000 78.655000 7.905000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 79.060000 7.905000 79.380000 ;
      LAYER met4 ;
        RECT 7.585000 79.060000 7.905000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 79.465000 7.905000 79.785000 ;
      LAYER met4 ;
        RECT 7.585000 79.465000 7.905000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 79.870000 7.905000 80.190000 ;
      LAYER met4 ;
        RECT 7.585000 79.870000 7.905000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 80.275000 7.905000 80.595000 ;
      LAYER met4 ;
        RECT 7.585000 80.275000 7.905000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 80.680000 7.905000 81.000000 ;
      LAYER met4 ;
        RECT 7.585000 80.680000 7.905000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 81.085000 7.905000 81.405000 ;
      LAYER met4 ;
        RECT 7.585000 81.085000 7.905000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 81.490000 7.905000 81.810000 ;
      LAYER met4 ;
        RECT 7.585000 81.490000 7.905000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 81.895000 7.905000 82.215000 ;
      LAYER met4 ;
        RECT 7.585000 81.895000 7.905000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585000 82.300000 7.905000 82.620000 ;
      LAYER met4 ;
        RECT 7.585000 82.300000 7.905000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 82.795000 7.965000 83.115000 ;
      LAYER met4 ;
        RECT 7.645000 82.795000 7.965000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 83.205000 7.965000 83.525000 ;
      LAYER met4 ;
        RECT 7.645000 83.205000 7.965000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 83.615000 7.965000 83.935000 ;
      LAYER met4 ;
        RECT 7.645000 83.615000 7.965000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 84.025000 7.965000 84.345000 ;
      LAYER met4 ;
        RECT 7.645000 84.025000 7.965000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 84.435000 7.965000 84.755000 ;
      LAYER met4 ;
        RECT 7.645000 84.435000 7.965000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 84.845000 7.965000 85.165000 ;
      LAYER met4 ;
        RECT 7.645000 84.845000 7.965000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 85.255000 7.965000 85.575000 ;
      LAYER met4 ;
        RECT 7.645000 85.255000 7.965000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 85.665000 7.965000 85.985000 ;
      LAYER met4 ;
        RECT 7.645000 85.665000 7.965000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 86.075000 7.965000 86.395000 ;
      LAYER met4 ;
        RECT 7.645000 86.075000 7.965000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 86.485000 7.965000 86.805000 ;
      LAYER met4 ;
        RECT 7.645000 86.485000 7.965000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 86.895000 7.965000 87.215000 ;
      LAYER met4 ;
        RECT 7.645000 86.895000 7.965000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 87.305000 7.965000 87.625000 ;
      LAYER met4 ;
        RECT 7.645000 87.305000 7.965000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 87.715000 7.965000 88.035000 ;
      LAYER met4 ;
        RECT 7.645000 87.715000 7.965000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 88.125000 7.965000 88.445000 ;
      LAYER met4 ;
        RECT 7.645000 88.125000 7.965000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 88.535000 7.965000 88.855000 ;
      LAYER met4 ;
        RECT 7.645000 88.535000 7.965000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 88.945000 7.965000 89.265000 ;
      LAYER met4 ;
        RECT 7.645000 88.945000 7.965000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 89.355000 7.965000 89.675000 ;
      LAYER met4 ;
        RECT 7.645000 89.355000 7.965000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 89.765000 7.965000 90.085000 ;
      LAYER met4 ;
        RECT 7.645000 89.765000 7.965000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 90.175000 7.965000 90.495000 ;
      LAYER met4 ;
        RECT 7.645000 90.175000 7.965000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 90.585000 7.965000 90.905000 ;
      LAYER met4 ;
        RECT 7.645000 90.585000 7.965000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 90.995000 7.965000 91.315000 ;
      LAYER met4 ;
        RECT 7.645000 90.995000 7.965000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 91.405000 7.965000 91.725000 ;
      LAYER met4 ;
        RECT 7.645000 91.405000 7.965000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 91.815000 7.965000 92.135000 ;
      LAYER met4 ;
        RECT 7.645000 91.815000 7.965000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 92.225000 7.965000 92.545000 ;
      LAYER met4 ;
        RECT 7.645000 92.225000 7.965000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645000 92.635000 7.965000 92.955000 ;
      LAYER met4 ;
        RECT 7.645000 92.635000 7.965000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920000 17.800000 8.240000 18.120000 ;
      LAYER met4 ;
        RECT 7.920000 17.800000 8.240000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920000 18.230000 8.240000 18.550000 ;
      LAYER met4 ;
        RECT 7.920000 18.230000 8.240000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920000 18.660000 8.240000 18.980000 ;
      LAYER met4 ;
        RECT 7.920000 18.660000 8.240000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920000 19.090000 8.240000 19.410000 ;
      LAYER met4 ;
        RECT 7.920000 19.090000 8.240000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920000 19.520000 8.240000 19.840000 ;
      LAYER met4 ;
        RECT 7.920000 19.520000 8.240000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920000 19.950000 8.240000 20.270000 ;
      LAYER met4 ;
        RECT 7.920000 19.950000 8.240000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920000 20.380000 8.240000 20.700000 ;
      LAYER met4 ;
        RECT 7.920000 20.380000 8.240000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920000 20.810000 8.240000 21.130000 ;
      LAYER met4 ;
        RECT 7.920000 20.810000 8.240000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920000 21.240000 8.240000 21.560000 ;
      LAYER met4 ;
        RECT 7.920000 21.240000 8.240000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920000 21.670000 8.240000 21.990000 ;
      LAYER met4 ;
        RECT 7.920000 21.670000 8.240000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920000 22.100000 8.240000 22.420000 ;
      LAYER met4 ;
        RECT 7.920000 22.100000 8.240000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 68.065000 8.305000 68.385000 ;
      LAYER met4 ;
        RECT 7.985000 68.065000 8.305000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 68.475000 8.305000 68.795000 ;
      LAYER met4 ;
        RECT 7.985000 68.475000 8.305000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 68.885000 8.305000 69.205000 ;
      LAYER met4 ;
        RECT 7.985000 68.885000 8.305000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 69.295000 8.305000 69.615000 ;
      LAYER met4 ;
        RECT 7.985000 69.295000 8.305000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 69.705000 8.305000 70.025000 ;
      LAYER met4 ;
        RECT 7.985000 69.705000 8.305000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 70.115000 8.305000 70.435000 ;
      LAYER met4 ;
        RECT 7.985000 70.115000 8.305000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 70.525000 8.305000 70.845000 ;
      LAYER met4 ;
        RECT 7.985000 70.525000 8.305000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 70.935000 8.305000 71.255000 ;
      LAYER met4 ;
        RECT 7.985000 70.935000 8.305000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 71.345000 8.305000 71.665000 ;
      LAYER met4 ;
        RECT 7.985000 71.345000 8.305000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 71.755000 8.305000 72.075000 ;
      LAYER met4 ;
        RECT 7.985000 71.755000 8.305000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 72.165000 8.305000 72.485000 ;
      LAYER met4 ;
        RECT 7.985000 72.165000 8.305000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 72.575000 8.305000 72.895000 ;
      LAYER met4 ;
        RECT 7.985000 72.575000 8.305000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 72.985000 8.305000 73.305000 ;
      LAYER met4 ;
        RECT 7.985000 72.985000 8.305000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 73.390000 8.305000 73.710000 ;
      LAYER met4 ;
        RECT 7.985000 73.390000 8.305000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 73.795000 8.305000 74.115000 ;
      LAYER met4 ;
        RECT 7.985000 73.795000 8.305000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 74.200000 8.305000 74.520000 ;
      LAYER met4 ;
        RECT 7.985000 74.200000 8.305000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 74.605000 8.305000 74.925000 ;
      LAYER met4 ;
        RECT 7.985000 74.605000 8.305000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 75.010000 8.305000 75.330000 ;
      LAYER met4 ;
        RECT 7.985000 75.010000 8.305000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 75.415000 8.305000 75.735000 ;
      LAYER met4 ;
        RECT 7.985000 75.415000 8.305000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 75.820000 8.305000 76.140000 ;
      LAYER met4 ;
        RECT 7.985000 75.820000 8.305000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 76.225000 8.305000 76.545000 ;
      LAYER met4 ;
        RECT 7.985000 76.225000 8.305000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 76.630000 8.305000 76.950000 ;
      LAYER met4 ;
        RECT 7.985000 76.630000 8.305000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 77.035000 8.305000 77.355000 ;
      LAYER met4 ;
        RECT 7.985000 77.035000 8.305000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 77.440000 8.305000 77.760000 ;
      LAYER met4 ;
        RECT 7.985000 77.440000 8.305000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 77.845000 8.305000 78.165000 ;
      LAYER met4 ;
        RECT 7.985000 77.845000 8.305000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 78.250000 8.305000 78.570000 ;
      LAYER met4 ;
        RECT 7.985000 78.250000 8.305000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 78.655000 8.305000 78.975000 ;
      LAYER met4 ;
        RECT 7.985000 78.655000 8.305000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 79.060000 8.305000 79.380000 ;
      LAYER met4 ;
        RECT 7.985000 79.060000 8.305000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 79.465000 8.305000 79.785000 ;
      LAYER met4 ;
        RECT 7.985000 79.465000 8.305000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 79.870000 8.305000 80.190000 ;
      LAYER met4 ;
        RECT 7.985000 79.870000 8.305000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 80.275000 8.305000 80.595000 ;
      LAYER met4 ;
        RECT 7.985000 80.275000 8.305000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 80.680000 8.305000 81.000000 ;
      LAYER met4 ;
        RECT 7.985000 80.680000 8.305000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 81.085000 8.305000 81.405000 ;
      LAYER met4 ;
        RECT 7.985000 81.085000 8.305000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 81.490000 8.305000 81.810000 ;
      LAYER met4 ;
        RECT 7.985000 81.490000 8.305000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 81.895000 8.305000 82.215000 ;
      LAYER met4 ;
        RECT 7.985000 81.895000 8.305000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985000 82.300000 8.305000 82.620000 ;
      LAYER met4 ;
        RECT 7.985000 82.300000 8.305000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 68.065000 70.470000 68.385000 ;
      LAYER met4 ;
        RECT 70.150000 68.065000 70.470000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 68.475000 70.470000 68.795000 ;
      LAYER met4 ;
        RECT 70.150000 68.475000 70.470000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 68.885000 70.470000 69.205000 ;
      LAYER met4 ;
        RECT 70.150000 68.885000 70.470000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 69.295000 70.470000 69.615000 ;
      LAYER met4 ;
        RECT 70.150000 69.295000 70.470000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 69.705000 70.470000 70.025000 ;
      LAYER met4 ;
        RECT 70.150000 69.705000 70.470000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 70.115000 70.470000 70.435000 ;
      LAYER met4 ;
        RECT 70.150000 70.115000 70.470000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 70.525000 70.470000 70.845000 ;
      LAYER met4 ;
        RECT 70.150000 70.525000 70.470000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 70.935000 70.470000 71.255000 ;
      LAYER met4 ;
        RECT 70.150000 70.935000 70.470000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 71.345000 70.470000 71.665000 ;
      LAYER met4 ;
        RECT 70.150000 71.345000 70.470000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 71.755000 70.470000 72.075000 ;
      LAYER met4 ;
        RECT 70.150000 71.755000 70.470000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 72.165000 70.470000 72.485000 ;
      LAYER met4 ;
        RECT 70.150000 72.165000 70.470000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 72.575000 70.470000 72.895000 ;
      LAYER met4 ;
        RECT 70.150000 72.575000 70.470000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 72.985000 70.470000 73.305000 ;
      LAYER met4 ;
        RECT 70.150000 72.985000 70.470000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 73.390000 70.470000 73.710000 ;
      LAYER met4 ;
        RECT 70.150000 73.390000 70.470000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 73.795000 70.470000 74.115000 ;
      LAYER met4 ;
        RECT 70.150000 73.795000 70.470000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 74.200000 70.470000 74.520000 ;
      LAYER met4 ;
        RECT 70.150000 74.200000 70.470000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 74.605000 70.470000 74.925000 ;
      LAYER met4 ;
        RECT 70.150000 74.605000 70.470000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 75.010000 70.470000 75.330000 ;
      LAYER met4 ;
        RECT 70.150000 75.010000 70.470000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 75.415000 70.470000 75.735000 ;
      LAYER met4 ;
        RECT 70.150000 75.415000 70.470000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 75.820000 70.470000 76.140000 ;
      LAYER met4 ;
        RECT 70.150000 75.820000 70.470000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 76.225000 70.470000 76.545000 ;
      LAYER met4 ;
        RECT 70.150000 76.225000 70.470000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 76.630000 70.470000 76.950000 ;
      LAYER met4 ;
        RECT 70.150000 76.630000 70.470000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 77.035000 70.470000 77.355000 ;
      LAYER met4 ;
        RECT 70.150000 77.035000 70.470000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 77.440000 70.470000 77.760000 ;
      LAYER met4 ;
        RECT 70.150000 77.440000 70.470000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 77.845000 70.470000 78.165000 ;
      LAYER met4 ;
        RECT 70.150000 77.845000 70.470000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 78.250000 70.470000 78.570000 ;
      LAYER met4 ;
        RECT 70.150000 78.250000 70.470000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 78.655000 70.470000 78.975000 ;
      LAYER met4 ;
        RECT 70.150000 78.655000 70.470000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 79.060000 70.470000 79.380000 ;
      LAYER met4 ;
        RECT 70.150000 79.060000 70.470000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 79.465000 70.470000 79.785000 ;
      LAYER met4 ;
        RECT 70.150000 79.465000 70.470000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 79.870000 70.470000 80.190000 ;
      LAYER met4 ;
        RECT 70.150000 79.870000 70.470000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 80.275000 70.470000 80.595000 ;
      LAYER met4 ;
        RECT 70.150000 80.275000 70.470000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 80.680000 70.470000 81.000000 ;
      LAYER met4 ;
        RECT 70.150000 80.680000 70.470000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 81.085000 70.470000 81.405000 ;
      LAYER met4 ;
        RECT 70.150000 81.085000 70.470000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 81.490000 70.470000 81.810000 ;
      LAYER met4 ;
        RECT 70.150000 81.490000 70.470000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 81.895000 70.470000 82.215000 ;
      LAYER met4 ;
        RECT 70.150000 81.895000 70.470000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.150000 82.300000 70.470000 82.620000 ;
      LAYER met4 ;
        RECT 70.150000 82.300000 70.470000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 82.795000 70.480000 83.115000 ;
      LAYER met4 ;
        RECT 70.160000 82.795000 70.480000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 83.205000 70.480000 83.525000 ;
      LAYER met4 ;
        RECT 70.160000 83.205000 70.480000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 83.615000 70.480000 83.935000 ;
      LAYER met4 ;
        RECT 70.160000 83.615000 70.480000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 84.025000 70.480000 84.345000 ;
      LAYER met4 ;
        RECT 70.160000 84.025000 70.480000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 84.435000 70.480000 84.755000 ;
      LAYER met4 ;
        RECT 70.160000 84.435000 70.480000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 84.845000 70.480000 85.165000 ;
      LAYER met4 ;
        RECT 70.160000 84.845000 70.480000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 85.255000 70.480000 85.575000 ;
      LAYER met4 ;
        RECT 70.160000 85.255000 70.480000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 85.665000 70.480000 85.985000 ;
      LAYER met4 ;
        RECT 70.160000 85.665000 70.480000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 86.075000 70.480000 86.395000 ;
      LAYER met4 ;
        RECT 70.160000 86.075000 70.480000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 86.485000 70.480000 86.805000 ;
      LAYER met4 ;
        RECT 70.160000 86.485000 70.480000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 86.895000 70.480000 87.215000 ;
      LAYER met4 ;
        RECT 70.160000 86.895000 70.480000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 87.305000 70.480000 87.625000 ;
      LAYER met4 ;
        RECT 70.160000 87.305000 70.480000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 87.715000 70.480000 88.035000 ;
      LAYER met4 ;
        RECT 70.160000 87.715000 70.480000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 88.125000 70.480000 88.445000 ;
      LAYER met4 ;
        RECT 70.160000 88.125000 70.480000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 88.535000 70.480000 88.855000 ;
      LAYER met4 ;
        RECT 70.160000 88.535000 70.480000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 88.945000 70.480000 89.265000 ;
      LAYER met4 ;
        RECT 70.160000 88.945000 70.480000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 89.355000 70.480000 89.675000 ;
      LAYER met4 ;
        RECT 70.160000 89.355000 70.480000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 89.765000 70.480000 90.085000 ;
      LAYER met4 ;
        RECT 70.160000 89.765000 70.480000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 90.175000 70.480000 90.495000 ;
      LAYER met4 ;
        RECT 70.160000 90.175000 70.480000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 90.585000 70.480000 90.905000 ;
      LAYER met4 ;
        RECT 70.160000 90.585000 70.480000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 90.995000 70.480000 91.315000 ;
      LAYER met4 ;
        RECT 70.160000 90.995000 70.480000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 91.405000 70.480000 91.725000 ;
      LAYER met4 ;
        RECT 70.160000 91.405000 70.480000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 91.815000 70.480000 92.135000 ;
      LAYER met4 ;
        RECT 70.160000 91.815000 70.480000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 92.225000 70.480000 92.545000 ;
      LAYER met4 ;
        RECT 70.160000 92.225000 70.480000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160000 92.635000 70.480000 92.955000 ;
      LAYER met4 ;
        RECT 70.160000 92.635000 70.480000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.225000 17.800000 70.545000 18.120000 ;
      LAYER met4 ;
        RECT 70.225000 17.800000 70.545000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.225000 18.230000 70.545000 18.550000 ;
      LAYER met4 ;
        RECT 70.225000 18.230000 70.545000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.225000 18.660000 70.545000 18.980000 ;
      LAYER met4 ;
        RECT 70.225000 18.660000 70.545000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.225000 19.090000 70.545000 19.410000 ;
      LAYER met4 ;
        RECT 70.225000 19.090000 70.545000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.225000 19.520000 70.545000 19.840000 ;
      LAYER met4 ;
        RECT 70.225000 19.520000 70.545000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.225000 19.950000 70.545000 20.270000 ;
      LAYER met4 ;
        RECT 70.225000 19.950000 70.545000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.225000 20.380000 70.545000 20.700000 ;
      LAYER met4 ;
        RECT 70.225000 20.380000 70.545000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.225000 20.810000 70.545000 21.130000 ;
      LAYER met4 ;
        RECT 70.225000 20.810000 70.545000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.225000 21.240000 70.545000 21.560000 ;
      LAYER met4 ;
        RECT 70.225000 21.240000 70.545000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.225000 21.670000 70.545000 21.990000 ;
      LAYER met4 ;
        RECT 70.225000 21.670000 70.545000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.225000 22.100000 70.545000 22.420000 ;
      LAYER met4 ;
        RECT 70.225000 22.100000 70.545000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 68.065000 70.870000 68.385000 ;
      LAYER met4 ;
        RECT 70.550000 68.065000 70.870000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 68.475000 70.870000 68.795000 ;
      LAYER met4 ;
        RECT 70.550000 68.475000 70.870000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 68.885000 70.870000 69.205000 ;
      LAYER met4 ;
        RECT 70.550000 68.885000 70.870000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 69.295000 70.870000 69.615000 ;
      LAYER met4 ;
        RECT 70.550000 69.295000 70.870000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 69.705000 70.870000 70.025000 ;
      LAYER met4 ;
        RECT 70.550000 69.705000 70.870000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 70.115000 70.870000 70.435000 ;
      LAYER met4 ;
        RECT 70.550000 70.115000 70.870000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 70.525000 70.870000 70.845000 ;
      LAYER met4 ;
        RECT 70.550000 70.525000 70.870000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 70.935000 70.870000 71.255000 ;
      LAYER met4 ;
        RECT 70.550000 70.935000 70.870000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 71.345000 70.870000 71.665000 ;
      LAYER met4 ;
        RECT 70.550000 71.345000 70.870000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 71.755000 70.870000 72.075000 ;
      LAYER met4 ;
        RECT 70.550000 71.755000 70.870000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 72.165000 70.870000 72.485000 ;
      LAYER met4 ;
        RECT 70.550000 72.165000 70.870000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 72.575000 70.870000 72.895000 ;
      LAYER met4 ;
        RECT 70.550000 72.575000 70.870000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 72.985000 70.870000 73.305000 ;
      LAYER met4 ;
        RECT 70.550000 72.985000 70.870000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 73.390000 70.870000 73.710000 ;
      LAYER met4 ;
        RECT 70.550000 73.390000 70.870000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 73.795000 70.870000 74.115000 ;
      LAYER met4 ;
        RECT 70.550000 73.795000 70.870000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 74.200000 70.870000 74.520000 ;
      LAYER met4 ;
        RECT 70.550000 74.200000 70.870000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 74.605000 70.870000 74.925000 ;
      LAYER met4 ;
        RECT 70.550000 74.605000 70.870000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 75.010000 70.870000 75.330000 ;
      LAYER met4 ;
        RECT 70.550000 75.010000 70.870000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 75.415000 70.870000 75.735000 ;
      LAYER met4 ;
        RECT 70.550000 75.415000 70.870000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 75.820000 70.870000 76.140000 ;
      LAYER met4 ;
        RECT 70.550000 75.820000 70.870000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 76.225000 70.870000 76.545000 ;
      LAYER met4 ;
        RECT 70.550000 76.225000 70.870000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 76.630000 70.870000 76.950000 ;
      LAYER met4 ;
        RECT 70.550000 76.630000 70.870000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 77.035000 70.870000 77.355000 ;
      LAYER met4 ;
        RECT 70.550000 77.035000 70.870000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 77.440000 70.870000 77.760000 ;
      LAYER met4 ;
        RECT 70.550000 77.440000 70.870000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 77.845000 70.870000 78.165000 ;
      LAYER met4 ;
        RECT 70.550000 77.845000 70.870000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 78.250000 70.870000 78.570000 ;
      LAYER met4 ;
        RECT 70.550000 78.250000 70.870000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 78.655000 70.870000 78.975000 ;
      LAYER met4 ;
        RECT 70.550000 78.655000 70.870000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 79.060000 70.870000 79.380000 ;
      LAYER met4 ;
        RECT 70.550000 79.060000 70.870000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 79.465000 70.870000 79.785000 ;
      LAYER met4 ;
        RECT 70.550000 79.465000 70.870000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 79.870000 70.870000 80.190000 ;
      LAYER met4 ;
        RECT 70.550000 79.870000 70.870000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 80.275000 70.870000 80.595000 ;
      LAYER met4 ;
        RECT 70.550000 80.275000 70.870000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 80.680000 70.870000 81.000000 ;
      LAYER met4 ;
        RECT 70.550000 80.680000 70.870000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 81.085000 70.870000 81.405000 ;
      LAYER met4 ;
        RECT 70.550000 81.085000 70.870000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 81.490000 70.870000 81.810000 ;
      LAYER met4 ;
        RECT 70.550000 81.490000 70.870000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 81.895000 70.870000 82.215000 ;
      LAYER met4 ;
        RECT 70.550000 81.895000 70.870000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.550000 82.300000 70.870000 82.620000 ;
      LAYER met4 ;
        RECT 70.550000 82.300000 70.870000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 82.795000 70.890000 83.115000 ;
      LAYER met4 ;
        RECT 70.570000 82.795000 70.890000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 83.205000 70.890000 83.525000 ;
      LAYER met4 ;
        RECT 70.570000 83.205000 70.890000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 83.615000 70.890000 83.935000 ;
      LAYER met4 ;
        RECT 70.570000 83.615000 70.890000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 84.025000 70.890000 84.345000 ;
      LAYER met4 ;
        RECT 70.570000 84.025000 70.890000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 84.435000 70.890000 84.755000 ;
      LAYER met4 ;
        RECT 70.570000 84.435000 70.890000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 84.845000 70.890000 85.165000 ;
      LAYER met4 ;
        RECT 70.570000 84.845000 70.890000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 85.255000 70.890000 85.575000 ;
      LAYER met4 ;
        RECT 70.570000 85.255000 70.890000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 85.665000 70.890000 85.985000 ;
      LAYER met4 ;
        RECT 70.570000 85.665000 70.890000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 86.075000 70.890000 86.395000 ;
      LAYER met4 ;
        RECT 70.570000 86.075000 70.890000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 86.485000 70.890000 86.805000 ;
      LAYER met4 ;
        RECT 70.570000 86.485000 70.890000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 86.895000 70.890000 87.215000 ;
      LAYER met4 ;
        RECT 70.570000 86.895000 70.890000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 87.305000 70.890000 87.625000 ;
      LAYER met4 ;
        RECT 70.570000 87.305000 70.890000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 87.715000 70.890000 88.035000 ;
      LAYER met4 ;
        RECT 70.570000 87.715000 70.890000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 88.125000 70.890000 88.445000 ;
      LAYER met4 ;
        RECT 70.570000 88.125000 70.890000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 88.535000 70.890000 88.855000 ;
      LAYER met4 ;
        RECT 70.570000 88.535000 70.890000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 88.945000 70.890000 89.265000 ;
      LAYER met4 ;
        RECT 70.570000 88.945000 70.890000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 89.355000 70.890000 89.675000 ;
      LAYER met4 ;
        RECT 70.570000 89.355000 70.890000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 89.765000 70.890000 90.085000 ;
      LAYER met4 ;
        RECT 70.570000 89.765000 70.890000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 90.175000 70.890000 90.495000 ;
      LAYER met4 ;
        RECT 70.570000 90.175000 70.890000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 90.585000 70.890000 90.905000 ;
      LAYER met4 ;
        RECT 70.570000 90.585000 70.890000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 90.995000 70.890000 91.315000 ;
      LAYER met4 ;
        RECT 70.570000 90.995000 70.890000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 91.405000 70.890000 91.725000 ;
      LAYER met4 ;
        RECT 70.570000 91.405000 70.890000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 91.815000 70.890000 92.135000 ;
      LAYER met4 ;
        RECT 70.570000 91.815000 70.890000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 92.225000 70.890000 92.545000 ;
      LAYER met4 ;
        RECT 70.570000 92.225000 70.890000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570000 92.635000 70.890000 92.955000 ;
      LAYER met4 ;
        RECT 70.570000 92.635000 70.890000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630000 17.800000 70.950000 18.120000 ;
      LAYER met4 ;
        RECT 70.630000 17.800000 70.950000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630000 18.230000 70.950000 18.550000 ;
      LAYER met4 ;
        RECT 70.630000 18.230000 70.950000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630000 18.660000 70.950000 18.980000 ;
      LAYER met4 ;
        RECT 70.630000 18.660000 70.950000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630000 19.090000 70.950000 19.410000 ;
      LAYER met4 ;
        RECT 70.630000 19.090000 70.950000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630000 19.520000 70.950000 19.840000 ;
      LAYER met4 ;
        RECT 70.630000 19.520000 70.950000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630000 19.950000 70.950000 20.270000 ;
      LAYER met4 ;
        RECT 70.630000 19.950000 70.950000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630000 20.380000 70.950000 20.700000 ;
      LAYER met4 ;
        RECT 70.630000 20.380000 70.950000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630000 20.810000 70.950000 21.130000 ;
      LAYER met4 ;
        RECT 70.630000 20.810000 70.950000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630000 21.240000 70.950000 21.560000 ;
      LAYER met4 ;
        RECT 70.630000 21.240000 70.950000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630000 21.670000 70.950000 21.990000 ;
      LAYER met4 ;
        RECT 70.630000 21.670000 70.950000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630000 22.100000 70.950000 22.420000 ;
      LAYER met4 ;
        RECT 70.630000 22.100000 70.950000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 68.065000 71.270000 68.385000 ;
      LAYER met4 ;
        RECT 70.950000 68.065000 71.270000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 68.475000 71.270000 68.795000 ;
      LAYER met4 ;
        RECT 70.950000 68.475000 71.270000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 68.885000 71.270000 69.205000 ;
      LAYER met4 ;
        RECT 70.950000 68.885000 71.270000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 69.295000 71.270000 69.615000 ;
      LAYER met4 ;
        RECT 70.950000 69.295000 71.270000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 69.705000 71.270000 70.025000 ;
      LAYER met4 ;
        RECT 70.950000 69.705000 71.270000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 70.115000 71.270000 70.435000 ;
      LAYER met4 ;
        RECT 70.950000 70.115000 71.270000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 70.525000 71.270000 70.845000 ;
      LAYER met4 ;
        RECT 70.950000 70.525000 71.270000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 70.935000 71.270000 71.255000 ;
      LAYER met4 ;
        RECT 70.950000 70.935000 71.270000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 71.345000 71.270000 71.665000 ;
      LAYER met4 ;
        RECT 70.950000 71.345000 71.270000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 71.755000 71.270000 72.075000 ;
      LAYER met4 ;
        RECT 70.950000 71.755000 71.270000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 72.165000 71.270000 72.485000 ;
      LAYER met4 ;
        RECT 70.950000 72.165000 71.270000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 72.575000 71.270000 72.895000 ;
      LAYER met4 ;
        RECT 70.950000 72.575000 71.270000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 72.985000 71.270000 73.305000 ;
      LAYER met4 ;
        RECT 70.950000 72.985000 71.270000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 73.390000 71.270000 73.710000 ;
      LAYER met4 ;
        RECT 70.950000 73.390000 71.270000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 73.795000 71.270000 74.115000 ;
      LAYER met4 ;
        RECT 70.950000 73.795000 71.270000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 74.200000 71.270000 74.520000 ;
      LAYER met4 ;
        RECT 70.950000 74.200000 71.270000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 74.605000 71.270000 74.925000 ;
      LAYER met4 ;
        RECT 70.950000 74.605000 71.270000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 75.010000 71.270000 75.330000 ;
      LAYER met4 ;
        RECT 70.950000 75.010000 71.270000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 75.415000 71.270000 75.735000 ;
      LAYER met4 ;
        RECT 70.950000 75.415000 71.270000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 75.820000 71.270000 76.140000 ;
      LAYER met4 ;
        RECT 70.950000 75.820000 71.270000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 76.225000 71.270000 76.545000 ;
      LAYER met4 ;
        RECT 70.950000 76.225000 71.270000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 76.630000 71.270000 76.950000 ;
      LAYER met4 ;
        RECT 70.950000 76.630000 71.270000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 77.035000 71.270000 77.355000 ;
      LAYER met4 ;
        RECT 70.950000 77.035000 71.270000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 77.440000 71.270000 77.760000 ;
      LAYER met4 ;
        RECT 70.950000 77.440000 71.270000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 77.845000 71.270000 78.165000 ;
      LAYER met4 ;
        RECT 70.950000 77.845000 71.270000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 78.250000 71.270000 78.570000 ;
      LAYER met4 ;
        RECT 70.950000 78.250000 71.270000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 78.655000 71.270000 78.975000 ;
      LAYER met4 ;
        RECT 70.950000 78.655000 71.270000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 79.060000 71.270000 79.380000 ;
      LAYER met4 ;
        RECT 70.950000 79.060000 71.270000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 79.465000 71.270000 79.785000 ;
      LAYER met4 ;
        RECT 70.950000 79.465000 71.270000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 79.870000 71.270000 80.190000 ;
      LAYER met4 ;
        RECT 70.950000 79.870000 71.270000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 80.275000 71.270000 80.595000 ;
      LAYER met4 ;
        RECT 70.950000 80.275000 71.270000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 80.680000 71.270000 81.000000 ;
      LAYER met4 ;
        RECT 70.950000 80.680000 71.270000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 81.085000 71.270000 81.405000 ;
      LAYER met4 ;
        RECT 70.950000 81.085000 71.270000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 81.490000 71.270000 81.810000 ;
      LAYER met4 ;
        RECT 70.950000 81.490000 71.270000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 81.895000 71.270000 82.215000 ;
      LAYER met4 ;
        RECT 70.950000 81.895000 71.270000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.950000 82.300000 71.270000 82.620000 ;
      LAYER met4 ;
        RECT 70.950000 82.300000 71.270000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 82.795000 71.300000 83.115000 ;
      LAYER met4 ;
        RECT 70.980000 82.795000 71.300000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 83.205000 71.300000 83.525000 ;
      LAYER met4 ;
        RECT 70.980000 83.205000 71.300000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 83.615000 71.300000 83.935000 ;
      LAYER met4 ;
        RECT 70.980000 83.615000 71.300000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 84.025000 71.300000 84.345000 ;
      LAYER met4 ;
        RECT 70.980000 84.025000 71.300000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 84.435000 71.300000 84.755000 ;
      LAYER met4 ;
        RECT 70.980000 84.435000 71.300000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 84.845000 71.300000 85.165000 ;
      LAYER met4 ;
        RECT 70.980000 84.845000 71.300000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 85.255000 71.300000 85.575000 ;
      LAYER met4 ;
        RECT 70.980000 85.255000 71.300000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 85.665000 71.300000 85.985000 ;
      LAYER met4 ;
        RECT 70.980000 85.665000 71.300000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 86.075000 71.300000 86.395000 ;
      LAYER met4 ;
        RECT 70.980000 86.075000 71.300000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 86.485000 71.300000 86.805000 ;
      LAYER met4 ;
        RECT 70.980000 86.485000 71.300000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 86.895000 71.300000 87.215000 ;
      LAYER met4 ;
        RECT 70.980000 86.895000 71.300000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 87.305000 71.300000 87.625000 ;
      LAYER met4 ;
        RECT 70.980000 87.305000 71.300000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 87.715000 71.300000 88.035000 ;
      LAYER met4 ;
        RECT 70.980000 87.715000 71.300000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 88.125000 71.300000 88.445000 ;
      LAYER met4 ;
        RECT 70.980000 88.125000 71.300000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 88.535000 71.300000 88.855000 ;
      LAYER met4 ;
        RECT 70.980000 88.535000 71.300000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 88.945000 71.300000 89.265000 ;
      LAYER met4 ;
        RECT 70.980000 88.945000 71.300000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 89.355000 71.300000 89.675000 ;
      LAYER met4 ;
        RECT 70.980000 89.355000 71.300000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 89.765000 71.300000 90.085000 ;
      LAYER met4 ;
        RECT 70.980000 89.765000 71.300000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 90.175000 71.300000 90.495000 ;
      LAYER met4 ;
        RECT 70.980000 90.175000 71.300000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 90.585000 71.300000 90.905000 ;
      LAYER met4 ;
        RECT 70.980000 90.585000 71.300000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 90.995000 71.300000 91.315000 ;
      LAYER met4 ;
        RECT 70.980000 90.995000 71.300000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 91.405000 71.300000 91.725000 ;
      LAYER met4 ;
        RECT 70.980000 91.405000 71.300000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 91.815000 71.300000 92.135000 ;
      LAYER met4 ;
        RECT 70.980000 91.815000 71.300000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 92.225000 71.300000 92.545000 ;
      LAYER met4 ;
        RECT 70.980000 92.225000 71.300000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980000 92.635000 71.300000 92.955000 ;
      LAYER met4 ;
        RECT 70.980000 92.635000 71.300000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.035000 17.800000 71.355000 18.120000 ;
      LAYER met4 ;
        RECT 71.035000 17.800000 71.355000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.035000 18.230000 71.355000 18.550000 ;
      LAYER met4 ;
        RECT 71.035000 18.230000 71.355000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.035000 18.660000 71.355000 18.980000 ;
      LAYER met4 ;
        RECT 71.035000 18.660000 71.355000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.035000 19.090000 71.355000 19.410000 ;
      LAYER met4 ;
        RECT 71.035000 19.090000 71.355000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.035000 19.520000 71.355000 19.840000 ;
      LAYER met4 ;
        RECT 71.035000 19.520000 71.355000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.035000 19.950000 71.355000 20.270000 ;
      LAYER met4 ;
        RECT 71.035000 19.950000 71.355000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.035000 20.380000 71.355000 20.700000 ;
      LAYER met4 ;
        RECT 71.035000 20.380000 71.355000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.035000 20.810000 71.355000 21.130000 ;
      LAYER met4 ;
        RECT 71.035000 20.810000 71.355000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.035000 21.240000 71.355000 21.560000 ;
      LAYER met4 ;
        RECT 71.035000 21.240000 71.355000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.035000 21.670000 71.355000 21.990000 ;
      LAYER met4 ;
        RECT 71.035000 21.670000 71.355000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.035000 22.100000 71.355000 22.420000 ;
      LAYER met4 ;
        RECT 71.035000 22.100000 71.355000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 68.065000 71.670000 68.385000 ;
      LAYER met4 ;
        RECT 71.350000 68.065000 71.670000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 68.475000 71.670000 68.795000 ;
      LAYER met4 ;
        RECT 71.350000 68.475000 71.670000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 68.885000 71.670000 69.205000 ;
      LAYER met4 ;
        RECT 71.350000 68.885000 71.670000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 69.295000 71.670000 69.615000 ;
      LAYER met4 ;
        RECT 71.350000 69.295000 71.670000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 69.705000 71.670000 70.025000 ;
      LAYER met4 ;
        RECT 71.350000 69.705000 71.670000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 70.115000 71.670000 70.435000 ;
      LAYER met4 ;
        RECT 71.350000 70.115000 71.670000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 70.525000 71.670000 70.845000 ;
      LAYER met4 ;
        RECT 71.350000 70.525000 71.670000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 70.935000 71.670000 71.255000 ;
      LAYER met4 ;
        RECT 71.350000 70.935000 71.670000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 71.345000 71.670000 71.665000 ;
      LAYER met4 ;
        RECT 71.350000 71.345000 71.670000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 71.755000 71.670000 72.075000 ;
      LAYER met4 ;
        RECT 71.350000 71.755000 71.670000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 72.165000 71.670000 72.485000 ;
      LAYER met4 ;
        RECT 71.350000 72.165000 71.670000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 72.575000 71.670000 72.895000 ;
      LAYER met4 ;
        RECT 71.350000 72.575000 71.670000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 72.985000 71.670000 73.305000 ;
      LAYER met4 ;
        RECT 71.350000 72.985000 71.670000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 73.390000 71.670000 73.710000 ;
      LAYER met4 ;
        RECT 71.350000 73.390000 71.670000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 73.795000 71.670000 74.115000 ;
      LAYER met4 ;
        RECT 71.350000 73.795000 71.670000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 74.200000 71.670000 74.520000 ;
      LAYER met4 ;
        RECT 71.350000 74.200000 71.670000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 74.605000 71.670000 74.925000 ;
      LAYER met4 ;
        RECT 71.350000 74.605000 71.670000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 75.010000 71.670000 75.330000 ;
      LAYER met4 ;
        RECT 71.350000 75.010000 71.670000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 75.415000 71.670000 75.735000 ;
      LAYER met4 ;
        RECT 71.350000 75.415000 71.670000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 75.820000 71.670000 76.140000 ;
      LAYER met4 ;
        RECT 71.350000 75.820000 71.670000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 76.225000 71.670000 76.545000 ;
      LAYER met4 ;
        RECT 71.350000 76.225000 71.670000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 76.630000 71.670000 76.950000 ;
      LAYER met4 ;
        RECT 71.350000 76.630000 71.670000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 77.035000 71.670000 77.355000 ;
      LAYER met4 ;
        RECT 71.350000 77.035000 71.670000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 77.440000 71.670000 77.760000 ;
      LAYER met4 ;
        RECT 71.350000 77.440000 71.670000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 77.845000 71.670000 78.165000 ;
      LAYER met4 ;
        RECT 71.350000 77.845000 71.670000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 78.250000 71.670000 78.570000 ;
      LAYER met4 ;
        RECT 71.350000 78.250000 71.670000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 78.655000 71.670000 78.975000 ;
      LAYER met4 ;
        RECT 71.350000 78.655000 71.670000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 79.060000 71.670000 79.380000 ;
      LAYER met4 ;
        RECT 71.350000 79.060000 71.670000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 79.465000 71.670000 79.785000 ;
      LAYER met4 ;
        RECT 71.350000 79.465000 71.670000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 79.870000 71.670000 80.190000 ;
      LAYER met4 ;
        RECT 71.350000 79.870000 71.670000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 80.275000 71.670000 80.595000 ;
      LAYER met4 ;
        RECT 71.350000 80.275000 71.670000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 80.680000 71.670000 81.000000 ;
      LAYER met4 ;
        RECT 71.350000 80.680000 71.670000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 81.085000 71.670000 81.405000 ;
      LAYER met4 ;
        RECT 71.350000 81.085000 71.670000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 81.490000 71.670000 81.810000 ;
      LAYER met4 ;
        RECT 71.350000 81.490000 71.670000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 81.895000 71.670000 82.215000 ;
      LAYER met4 ;
        RECT 71.350000 81.895000 71.670000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.350000 82.300000 71.670000 82.620000 ;
      LAYER met4 ;
        RECT 71.350000 82.300000 71.670000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 82.795000 71.710000 83.115000 ;
      LAYER met4 ;
        RECT 71.390000 82.795000 71.710000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 83.205000 71.710000 83.525000 ;
      LAYER met4 ;
        RECT 71.390000 83.205000 71.710000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 83.615000 71.710000 83.935000 ;
      LAYER met4 ;
        RECT 71.390000 83.615000 71.710000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 84.025000 71.710000 84.345000 ;
      LAYER met4 ;
        RECT 71.390000 84.025000 71.710000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 84.435000 71.710000 84.755000 ;
      LAYER met4 ;
        RECT 71.390000 84.435000 71.710000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 84.845000 71.710000 85.165000 ;
      LAYER met4 ;
        RECT 71.390000 84.845000 71.710000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 85.255000 71.710000 85.575000 ;
      LAYER met4 ;
        RECT 71.390000 85.255000 71.710000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 85.665000 71.710000 85.985000 ;
      LAYER met4 ;
        RECT 71.390000 85.665000 71.710000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 86.075000 71.710000 86.395000 ;
      LAYER met4 ;
        RECT 71.390000 86.075000 71.710000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 86.485000 71.710000 86.805000 ;
      LAYER met4 ;
        RECT 71.390000 86.485000 71.710000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 86.895000 71.710000 87.215000 ;
      LAYER met4 ;
        RECT 71.390000 86.895000 71.710000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 87.305000 71.710000 87.625000 ;
      LAYER met4 ;
        RECT 71.390000 87.305000 71.710000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 87.715000 71.710000 88.035000 ;
      LAYER met4 ;
        RECT 71.390000 87.715000 71.710000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 88.125000 71.710000 88.445000 ;
      LAYER met4 ;
        RECT 71.390000 88.125000 71.710000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 88.535000 71.710000 88.855000 ;
      LAYER met4 ;
        RECT 71.390000 88.535000 71.710000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 88.945000 71.710000 89.265000 ;
      LAYER met4 ;
        RECT 71.390000 88.945000 71.710000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 89.355000 71.710000 89.675000 ;
      LAYER met4 ;
        RECT 71.390000 89.355000 71.710000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 89.765000 71.710000 90.085000 ;
      LAYER met4 ;
        RECT 71.390000 89.765000 71.710000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 90.175000 71.710000 90.495000 ;
      LAYER met4 ;
        RECT 71.390000 90.175000 71.710000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 90.585000 71.710000 90.905000 ;
      LAYER met4 ;
        RECT 71.390000 90.585000 71.710000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 90.995000 71.710000 91.315000 ;
      LAYER met4 ;
        RECT 71.390000 90.995000 71.710000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 91.405000 71.710000 91.725000 ;
      LAYER met4 ;
        RECT 71.390000 91.405000 71.710000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 91.815000 71.710000 92.135000 ;
      LAYER met4 ;
        RECT 71.390000 91.815000 71.710000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 92.225000 71.710000 92.545000 ;
      LAYER met4 ;
        RECT 71.390000 92.225000 71.710000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390000 92.635000 71.710000 92.955000 ;
      LAYER met4 ;
        RECT 71.390000 92.635000 71.710000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 17.800000 71.760000 18.120000 ;
      LAYER met4 ;
        RECT 71.440000 17.800000 71.760000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 18.230000 71.760000 18.550000 ;
      LAYER met4 ;
        RECT 71.440000 18.230000 71.760000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 18.660000 71.760000 18.980000 ;
      LAYER met4 ;
        RECT 71.440000 18.660000 71.760000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 19.090000 71.760000 19.410000 ;
      LAYER met4 ;
        RECT 71.440000 19.090000 71.760000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 19.520000 71.760000 19.840000 ;
      LAYER met4 ;
        RECT 71.440000 19.520000 71.760000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 19.950000 71.760000 20.270000 ;
      LAYER met4 ;
        RECT 71.440000 19.950000 71.760000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 20.380000 71.760000 20.700000 ;
      LAYER met4 ;
        RECT 71.440000 20.380000 71.760000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 20.810000 71.760000 21.130000 ;
      LAYER met4 ;
        RECT 71.440000 20.810000 71.760000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 21.240000 71.760000 21.560000 ;
      LAYER met4 ;
        RECT 71.440000 21.240000 71.760000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 21.670000 71.760000 21.990000 ;
      LAYER met4 ;
        RECT 71.440000 21.670000 71.760000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 22.100000 71.760000 22.420000 ;
      LAYER met4 ;
        RECT 71.440000 22.100000 71.760000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 68.065000 72.070000 68.385000 ;
      LAYER met4 ;
        RECT 71.750000 68.065000 72.070000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 68.475000 72.070000 68.795000 ;
      LAYER met4 ;
        RECT 71.750000 68.475000 72.070000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 68.885000 72.070000 69.205000 ;
      LAYER met4 ;
        RECT 71.750000 68.885000 72.070000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 69.295000 72.070000 69.615000 ;
      LAYER met4 ;
        RECT 71.750000 69.295000 72.070000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 69.705000 72.070000 70.025000 ;
      LAYER met4 ;
        RECT 71.750000 69.705000 72.070000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 70.115000 72.070000 70.435000 ;
      LAYER met4 ;
        RECT 71.750000 70.115000 72.070000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 70.525000 72.070000 70.845000 ;
      LAYER met4 ;
        RECT 71.750000 70.525000 72.070000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 70.935000 72.070000 71.255000 ;
      LAYER met4 ;
        RECT 71.750000 70.935000 72.070000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 71.345000 72.070000 71.665000 ;
      LAYER met4 ;
        RECT 71.750000 71.345000 72.070000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 71.755000 72.070000 72.075000 ;
      LAYER met4 ;
        RECT 71.750000 71.755000 72.070000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 72.165000 72.070000 72.485000 ;
      LAYER met4 ;
        RECT 71.750000 72.165000 72.070000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 72.575000 72.070000 72.895000 ;
      LAYER met4 ;
        RECT 71.750000 72.575000 72.070000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 72.985000 72.070000 73.305000 ;
      LAYER met4 ;
        RECT 71.750000 72.985000 72.070000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 73.390000 72.070000 73.710000 ;
      LAYER met4 ;
        RECT 71.750000 73.390000 72.070000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 73.795000 72.070000 74.115000 ;
      LAYER met4 ;
        RECT 71.750000 73.795000 72.070000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 74.200000 72.070000 74.520000 ;
      LAYER met4 ;
        RECT 71.750000 74.200000 72.070000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 74.605000 72.070000 74.925000 ;
      LAYER met4 ;
        RECT 71.750000 74.605000 72.070000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 75.010000 72.070000 75.330000 ;
      LAYER met4 ;
        RECT 71.750000 75.010000 72.070000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 75.415000 72.070000 75.735000 ;
      LAYER met4 ;
        RECT 71.750000 75.415000 72.070000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 75.820000 72.070000 76.140000 ;
      LAYER met4 ;
        RECT 71.750000 75.820000 72.070000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 76.225000 72.070000 76.545000 ;
      LAYER met4 ;
        RECT 71.750000 76.225000 72.070000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 76.630000 72.070000 76.950000 ;
      LAYER met4 ;
        RECT 71.750000 76.630000 72.070000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 77.035000 72.070000 77.355000 ;
      LAYER met4 ;
        RECT 71.750000 77.035000 72.070000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 77.440000 72.070000 77.760000 ;
      LAYER met4 ;
        RECT 71.750000 77.440000 72.070000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 77.845000 72.070000 78.165000 ;
      LAYER met4 ;
        RECT 71.750000 77.845000 72.070000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 78.250000 72.070000 78.570000 ;
      LAYER met4 ;
        RECT 71.750000 78.250000 72.070000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 78.655000 72.070000 78.975000 ;
      LAYER met4 ;
        RECT 71.750000 78.655000 72.070000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 79.060000 72.070000 79.380000 ;
      LAYER met4 ;
        RECT 71.750000 79.060000 72.070000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 79.465000 72.070000 79.785000 ;
      LAYER met4 ;
        RECT 71.750000 79.465000 72.070000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 79.870000 72.070000 80.190000 ;
      LAYER met4 ;
        RECT 71.750000 79.870000 72.070000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 80.275000 72.070000 80.595000 ;
      LAYER met4 ;
        RECT 71.750000 80.275000 72.070000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 80.680000 72.070000 81.000000 ;
      LAYER met4 ;
        RECT 71.750000 80.680000 72.070000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 81.085000 72.070000 81.405000 ;
      LAYER met4 ;
        RECT 71.750000 81.085000 72.070000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 81.490000 72.070000 81.810000 ;
      LAYER met4 ;
        RECT 71.750000 81.490000 72.070000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 81.895000 72.070000 82.215000 ;
      LAYER met4 ;
        RECT 71.750000 81.895000 72.070000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.750000 82.300000 72.070000 82.620000 ;
      LAYER met4 ;
        RECT 71.750000 82.300000 72.070000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 82.795000 72.120000 83.115000 ;
      LAYER met4 ;
        RECT 71.800000 82.795000 72.120000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 83.205000 72.120000 83.525000 ;
      LAYER met4 ;
        RECT 71.800000 83.205000 72.120000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 83.615000 72.120000 83.935000 ;
      LAYER met4 ;
        RECT 71.800000 83.615000 72.120000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 84.025000 72.120000 84.345000 ;
      LAYER met4 ;
        RECT 71.800000 84.025000 72.120000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 84.435000 72.120000 84.755000 ;
      LAYER met4 ;
        RECT 71.800000 84.435000 72.120000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 84.845000 72.120000 85.165000 ;
      LAYER met4 ;
        RECT 71.800000 84.845000 72.120000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 85.255000 72.120000 85.575000 ;
      LAYER met4 ;
        RECT 71.800000 85.255000 72.120000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 85.665000 72.120000 85.985000 ;
      LAYER met4 ;
        RECT 71.800000 85.665000 72.120000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 86.075000 72.120000 86.395000 ;
      LAYER met4 ;
        RECT 71.800000 86.075000 72.120000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 86.485000 72.120000 86.805000 ;
      LAYER met4 ;
        RECT 71.800000 86.485000 72.120000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 86.895000 72.120000 87.215000 ;
      LAYER met4 ;
        RECT 71.800000 86.895000 72.120000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 87.305000 72.120000 87.625000 ;
      LAYER met4 ;
        RECT 71.800000 87.305000 72.120000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 87.715000 72.120000 88.035000 ;
      LAYER met4 ;
        RECT 71.800000 87.715000 72.120000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 88.125000 72.120000 88.445000 ;
      LAYER met4 ;
        RECT 71.800000 88.125000 72.120000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 88.535000 72.120000 88.855000 ;
      LAYER met4 ;
        RECT 71.800000 88.535000 72.120000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 88.945000 72.120000 89.265000 ;
      LAYER met4 ;
        RECT 71.800000 88.945000 72.120000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 89.355000 72.120000 89.675000 ;
      LAYER met4 ;
        RECT 71.800000 89.355000 72.120000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 89.765000 72.120000 90.085000 ;
      LAYER met4 ;
        RECT 71.800000 89.765000 72.120000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 90.175000 72.120000 90.495000 ;
      LAYER met4 ;
        RECT 71.800000 90.175000 72.120000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 90.585000 72.120000 90.905000 ;
      LAYER met4 ;
        RECT 71.800000 90.585000 72.120000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 90.995000 72.120000 91.315000 ;
      LAYER met4 ;
        RECT 71.800000 90.995000 72.120000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 91.405000 72.120000 91.725000 ;
      LAYER met4 ;
        RECT 71.800000 91.405000 72.120000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 91.815000 72.120000 92.135000 ;
      LAYER met4 ;
        RECT 71.800000 91.815000 72.120000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 92.225000 72.120000 92.545000 ;
      LAYER met4 ;
        RECT 71.800000 92.225000 72.120000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800000 92.635000 72.120000 92.955000 ;
      LAYER met4 ;
        RECT 71.800000 92.635000 72.120000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.845000 17.800000 72.165000 18.120000 ;
      LAYER met4 ;
        RECT 71.845000 17.800000 72.165000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.845000 18.230000 72.165000 18.550000 ;
      LAYER met4 ;
        RECT 71.845000 18.230000 72.165000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.845000 18.660000 72.165000 18.980000 ;
      LAYER met4 ;
        RECT 71.845000 18.660000 72.165000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.845000 19.090000 72.165000 19.410000 ;
      LAYER met4 ;
        RECT 71.845000 19.090000 72.165000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.845000 19.520000 72.165000 19.840000 ;
      LAYER met4 ;
        RECT 71.845000 19.520000 72.165000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.845000 19.950000 72.165000 20.270000 ;
      LAYER met4 ;
        RECT 71.845000 19.950000 72.165000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.845000 20.380000 72.165000 20.700000 ;
      LAYER met4 ;
        RECT 71.845000 20.380000 72.165000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.845000 20.810000 72.165000 21.130000 ;
      LAYER met4 ;
        RECT 71.845000 20.810000 72.165000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.845000 21.240000 72.165000 21.560000 ;
      LAYER met4 ;
        RECT 71.845000 21.240000 72.165000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.845000 21.670000 72.165000 21.990000 ;
      LAYER met4 ;
        RECT 71.845000 21.670000 72.165000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.845000 22.100000 72.165000 22.420000 ;
      LAYER met4 ;
        RECT 71.845000 22.100000 72.165000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 68.065000 72.470000 68.385000 ;
      LAYER met4 ;
        RECT 72.150000 68.065000 72.470000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 68.475000 72.470000 68.795000 ;
      LAYER met4 ;
        RECT 72.150000 68.475000 72.470000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 68.885000 72.470000 69.205000 ;
      LAYER met4 ;
        RECT 72.150000 68.885000 72.470000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 69.295000 72.470000 69.615000 ;
      LAYER met4 ;
        RECT 72.150000 69.295000 72.470000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 69.705000 72.470000 70.025000 ;
      LAYER met4 ;
        RECT 72.150000 69.705000 72.470000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 70.115000 72.470000 70.435000 ;
      LAYER met4 ;
        RECT 72.150000 70.115000 72.470000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 70.525000 72.470000 70.845000 ;
      LAYER met4 ;
        RECT 72.150000 70.525000 72.470000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 70.935000 72.470000 71.255000 ;
      LAYER met4 ;
        RECT 72.150000 70.935000 72.470000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 71.345000 72.470000 71.665000 ;
      LAYER met4 ;
        RECT 72.150000 71.345000 72.470000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 71.755000 72.470000 72.075000 ;
      LAYER met4 ;
        RECT 72.150000 71.755000 72.470000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 72.165000 72.470000 72.485000 ;
      LAYER met4 ;
        RECT 72.150000 72.165000 72.470000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 72.575000 72.470000 72.895000 ;
      LAYER met4 ;
        RECT 72.150000 72.575000 72.470000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 72.985000 72.470000 73.305000 ;
      LAYER met4 ;
        RECT 72.150000 72.985000 72.470000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 73.390000 72.470000 73.710000 ;
      LAYER met4 ;
        RECT 72.150000 73.390000 72.470000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 73.795000 72.470000 74.115000 ;
      LAYER met4 ;
        RECT 72.150000 73.795000 72.470000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 74.200000 72.470000 74.520000 ;
      LAYER met4 ;
        RECT 72.150000 74.200000 72.470000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 74.605000 72.470000 74.925000 ;
      LAYER met4 ;
        RECT 72.150000 74.605000 72.470000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 75.010000 72.470000 75.330000 ;
      LAYER met4 ;
        RECT 72.150000 75.010000 72.470000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 75.415000 72.470000 75.735000 ;
      LAYER met4 ;
        RECT 72.150000 75.415000 72.470000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 75.820000 72.470000 76.140000 ;
      LAYER met4 ;
        RECT 72.150000 75.820000 72.470000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 76.225000 72.470000 76.545000 ;
      LAYER met4 ;
        RECT 72.150000 76.225000 72.470000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 76.630000 72.470000 76.950000 ;
      LAYER met4 ;
        RECT 72.150000 76.630000 72.470000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 77.035000 72.470000 77.355000 ;
      LAYER met4 ;
        RECT 72.150000 77.035000 72.470000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 77.440000 72.470000 77.760000 ;
      LAYER met4 ;
        RECT 72.150000 77.440000 72.470000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 77.845000 72.470000 78.165000 ;
      LAYER met4 ;
        RECT 72.150000 77.845000 72.470000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 78.250000 72.470000 78.570000 ;
      LAYER met4 ;
        RECT 72.150000 78.250000 72.470000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 78.655000 72.470000 78.975000 ;
      LAYER met4 ;
        RECT 72.150000 78.655000 72.470000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 79.060000 72.470000 79.380000 ;
      LAYER met4 ;
        RECT 72.150000 79.060000 72.470000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 79.465000 72.470000 79.785000 ;
      LAYER met4 ;
        RECT 72.150000 79.465000 72.470000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 79.870000 72.470000 80.190000 ;
      LAYER met4 ;
        RECT 72.150000 79.870000 72.470000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 80.275000 72.470000 80.595000 ;
      LAYER met4 ;
        RECT 72.150000 80.275000 72.470000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 80.680000 72.470000 81.000000 ;
      LAYER met4 ;
        RECT 72.150000 80.680000 72.470000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 81.085000 72.470000 81.405000 ;
      LAYER met4 ;
        RECT 72.150000 81.085000 72.470000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 81.490000 72.470000 81.810000 ;
      LAYER met4 ;
        RECT 72.150000 81.490000 72.470000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 81.895000 72.470000 82.215000 ;
      LAYER met4 ;
        RECT 72.150000 81.895000 72.470000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.150000 82.300000 72.470000 82.620000 ;
      LAYER met4 ;
        RECT 72.150000 82.300000 72.470000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 82.795000 72.530000 83.115000 ;
      LAYER met4 ;
        RECT 72.210000 82.795000 72.530000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 83.205000 72.530000 83.525000 ;
      LAYER met4 ;
        RECT 72.210000 83.205000 72.530000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 83.615000 72.530000 83.935000 ;
      LAYER met4 ;
        RECT 72.210000 83.615000 72.530000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 84.025000 72.530000 84.345000 ;
      LAYER met4 ;
        RECT 72.210000 84.025000 72.530000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 84.435000 72.530000 84.755000 ;
      LAYER met4 ;
        RECT 72.210000 84.435000 72.530000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 84.845000 72.530000 85.165000 ;
      LAYER met4 ;
        RECT 72.210000 84.845000 72.530000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 85.255000 72.530000 85.575000 ;
      LAYER met4 ;
        RECT 72.210000 85.255000 72.530000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 85.665000 72.530000 85.985000 ;
      LAYER met4 ;
        RECT 72.210000 85.665000 72.530000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 86.075000 72.530000 86.395000 ;
      LAYER met4 ;
        RECT 72.210000 86.075000 72.530000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 86.485000 72.530000 86.805000 ;
      LAYER met4 ;
        RECT 72.210000 86.485000 72.530000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 86.895000 72.530000 87.215000 ;
      LAYER met4 ;
        RECT 72.210000 86.895000 72.530000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 87.305000 72.530000 87.625000 ;
      LAYER met4 ;
        RECT 72.210000 87.305000 72.530000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 87.715000 72.530000 88.035000 ;
      LAYER met4 ;
        RECT 72.210000 87.715000 72.530000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 88.125000 72.530000 88.445000 ;
      LAYER met4 ;
        RECT 72.210000 88.125000 72.530000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 88.535000 72.530000 88.855000 ;
      LAYER met4 ;
        RECT 72.210000 88.535000 72.530000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 88.945000 72.530000 89.265000 ;
      LAYER met4 ;
        RECT 72.210000 88.945000 72.530000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 89.355000 72.530000 89.675000 ;
      LAYER met4 ;
        RECT 72.210000 89.355000 72.530000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 89.765000 72.530000 90.085000 ;
      LAYER met4 ;
        RECT 72.210000 89.765000 72.530000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 90.175000 72.530000 90.495000 ;
      LAYER met4 ;
        RECT 72.210000 90.175000 72.530000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 90.585000 72.530000 90.905000 ;
      LAYER met4 ;
        RECT 72.210000 90.585000 72.530000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 90.995000 72.530000 91.315000 ;
      LAYER met4 ;
        RECT 72.210000 90.995000 72.530000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 91.405000 72.530000 91.725000 ;
      LAYER met4 ;
        RECT 72.210000 91.405000 72.530000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 91.815000 72.530000 92.135000 ;
      LAYER met4 ;
        RECT 72.210000 91.815000 72.530000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 92.225000 72.530000 92.545000 ;
      LAYER met4 ;
        RECT 72.210000 92.225000 72.530000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210000 92.635000 72.530000 92.955000 ;
      LAYER met4 ;
        RECT 72.210000 92.635000 72.530000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.255000 17.800000 72.575000 18.120000 ;
      LAYER met4 ;
        RECT 72.255000 17.800000 72.575000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.255000 18.230000 72.575000 18.550000 ;
      LAYER met4 ;
        RECT 72.255000 18.230000 72.575000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.255000 18.660000 72.575000 18.980000 ;
      LAYER met4 ;
        RECT 72.255000 18.660000 72.575000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.255000 19.090000 72.575000 19.410000 ;
      LAYER met4 ;
        RECT 72.255000 19.090000 72.575000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.255000 19.520000 72.575000 19.840000 ;
      LAYER met4 ;
        RECT 72.255000 19.520000 72.575000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.255000 19.950000 72.575000 20.270000 ;
      LAYER met4 ;
        RECT 72.255000 19.950000 72.575000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.255000 20.380000 72.575000 20.700000 ;
      LAYER met4 ;
        RECT 72.255000 20.380000 72.575000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.255000 20.810000 72.575000 21.130000 ;
      LAYER met4 ;
        RECT 72.255000 20.810000 72.575000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.255000 21.240000 72.575000 21.560000 ;
      LAYER met4 ;
        RECT 72.255000 21.240000 72.575000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.255000 21.670000 72.575000 21.990000 ;
      LAYER met4 ;
        RECT 72.255000 21.670000 72.575000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.255000 22.100000 72.575000 22.420000 ;
      LAYER met4 ;
        RECT 72.255000 22.100000 72.575000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 68.065000 72.870000 68.385000 ;
      LAYER met4 ;
        RECT 72.550000 68.065000 72.870000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 68.475000 72.870000 68.795000 ;
      LAYER met4 ;
        RECT 72.550000 68.475000 72.870000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 68.885000 72.870000 69.205000 ;
      LAYER met4 ;
        RECT 72.550000 68.885000 72.870000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 69.295000 72.870000 69.615000 ;
      LAYER met4 ;
        RECT 72.550000 69.295000 72.870000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 69.705000 72.870000 70.025000 ;
      LAYER met4 ;
        RECT 72.550000 69.705000 72.870000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 70.115000 72.870000 70.435000 ;
      LAYER met4 ;
        RECT 72.550000 70.115000 72.870000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 70.525000 72.870000 70.845000 ;
      LAYER met4 ;
        RECT 72.550000 70.525000 72.870000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 70.935000 72.870000 71.255000 ;
      LAYER met4 ;
        RECT 72.550000 70.935000 72.870000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 71.345000 72.870000 71.665000 ;
      LAYER met4 ;
        RECT 72.550000 71.345000 72.870000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 71.755000 72.870000 72.075000 ;
      LAYER met4 ;
        RECT 72.550000 71.755000 72.870000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 72.165000 72.870000 72.485000 ;
      LAYER met4 ;
        RECT 72.550000 72.165000 72.870000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 72.575000 72.870000 72.895000 ;
      LAYER met4 ;
        RECT 72.550000 72.575000 72.870000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 72.985000 72.870000 73.305000 ;
      LAYER met4 ;
        RECT 72.550000 72.985000 72.870000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 73.390000 72.870000 73.710000 ;
      LAYER met4 ;
        RECT 72.550000 73.390000 72.870000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 73.795000 72.870000 74.115000 ;
      LAYER met4 ;
        RECT 72.550000 73.795000 72.870000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 74.200000 72.870000 74.520000 ;
      LAYER met4 ;
        RECT 72.550000 74.200000 72.870000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 74.605000 72.870000 74.925000 ;
      LAYER met4 ;
        RECT 72.550000 74.605000 72.870000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 75.010000 72.870000 75.330000 ;
      LAYER met4 ;
        RECT 72.550000 75.010000 72.870000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 75.415000 72.870000 75.735000 ;
      LAYER met4 ;
        RECT 72.550000 75.415000 72.870000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 75.820000 72.870000 76.140000 ;
      LAYER met4 ;
        RECT 72.550000 75.820000 72.870000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 76.225000 72.870000 76.545000 ;
      LAYER met4 ;
        RECT 72.550000 76.225000 72.870000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 76.630000 72.870000 76.950000 ;
      LAYER met4 ;
        RECT 72.550000 76.630000 72.870000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 77.035000 72.870000 77.355000 ;
      LAYER met4 ;
        RECT 72.550000 77.035000 72.870000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 77.440000 72.870000 77.760000 ;
      LAYER met4 ;
        RECT 72.550000 77.440000 72.870000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 77.845000 72.870000 78.165000 ;
      LAYER met4 ;
        RECT 72.550000 77.845000 72.870000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 78.250000 72.870000 78.570000 ;
      LAYER met4 ;
        RECT 72.550000 78.250000 72.870000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 78.655000 72.870000 78.975000 ;
      LAYER met4 ;
        RECT 72.550000 78.655000 72.870000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 79.060000 72.870000 79.380000 ;
      LAYER met4 ;
        RECT 72.550000 79.060000 72.870000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 79.465000 72.870000 79.785000 ;
      LAYER met4 ;
        RECT 72.550000 79.465000 72.870000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 79.870000 72.870000 80.190000 ;
      LAYER met4 ;
        RECT 72.550000 79.870000 72.870000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 80.275000 72.870000 80.595000 ;
      LAYER met4 ;
        RECT 72.550000 80.275000 72.870000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 80.680000 72.870000 81.000000 ;
      LAYER met4 ;
        RECT 72.550000 80.680000 72.870000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 81.085000 72.870000 81.405000 ;
      LAYER met4 ;
        RECT 72.550000 81.085000 72.870000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 81.490000 72.870000 81.810000 ;
      LAYER met4 ;
        RECT 72.550000 81.490000 72.870000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 81.895000 72.870000 82.215000 ;
      LAYER met4 ;
        RECT 72.550000 81.895000 72.870000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.550000 82.300000 72.870000 82.620000 ;
      LAYER met4 ;
        RECT 72.550000 82.300000 72.870000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 82.795000 72.940000 83.115000 ;
      LAYER met4 ;
        RECT 72.620000 82.795000 72.940000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 83.205000 72.940000 83.525000 ;
      LAYER met4 ;
        RECT 72.620000 83.205000 72.940000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 83.615000 72.940000 83.935000 ;
      LAYER met4 ;
        RECT 72.620000 83.615000 72.940000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 84.025000 72.940000 84.345000 ;
      LAYER met4 ;
        RECT 72.620000 84.025000 72.940000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 84.435000 72.940000 84.755000 ;
      LAYER met4 ;
        RECT 72.620000 84.435000 72.940000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 84.845000 72.940000 85.165000 ;
      LAYER met4 ;
        RECT 72.620000 84.845000 72.940000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 85.255000 72.940000 85.575000 ;
      LAYER met4 ;
        RECT 72.620000 85.255000 72.940000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 85.665000 72.940000 85.985000 ;
      LAYER met4 ;
        RECT 72.620000 85.665000 72.940000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 86.075000 72.940000 86.395000 ;
      LAYER met4 ;
        RECT 72.620000 86.075000 72.940000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 86.485000 72.940000 86.805000 ;
      LAYER met4 ;
        RECT 72.620000 86.485000 72.940000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 86.895000 72.940000 87.215000 ;
      LAYER met4 ;
        RECT 72.620000 86.895000 72.940000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 87.305000 72.940000 87.625000 ;
      LAYER met4 ;
        RECT 72.620000 87.305000 72.940000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 87.715000 72.940000 88.035000 ;
      LAYER met4 ;
        RECT 72.620000 87.715000 72.940000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 88.125000 72.940000 88.445000 ;
      LAYER met4 ;
        RECT 72.620000 88.125000 72.940000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 88.535000 72.940000 88.855000 ;
      LAYER met4 ;
        RECT 72.620000 88.535000 72.940000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 88.945000 72.940000 89.265000 ;
      LAYER met4 ;
        RECT 72.620000 88.945000 72.940000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 89.355000 72.940000 89.675000 ;
      LAYER met4 ;
        RECT 72.620000 89.355000 72.940000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 89.765000 72.940000 90.085000 ;
      LAYER met4 ;
        RECT 72.620000 89.765000 72.940000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 90.175000 72.940000 90.495000 ;
      LAYER met4 ;
        RECT 72.620000 90.175000 72.940000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 90.585000 72.940000 90.905000 ;
      LAYER met4 ;
        RECT 72.620000 90.585000 72.940000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 90.995000 72.940000 91.315000 ;
      LAYER met4 ;
        RECT 72.620000 90.995000 72.940000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 91.405000 72.940000 91.725000 ;
      LAYER met4 ;
        RECT 72.620000 91.405000 72.940000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 91.815000 72.940000 92.135000 ;
      LAYER met4 ;
        RECT 72.620000 91.815000 72.940000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 92.225000 72.940000 92.545000 ;
      LAYER met4 ;
        RECT 72.620000 92.225000 72.940000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620000 92.635000 72.940000 92.955000 ;
      LAYER met4 ;
        RECT 72.620000 92.635000 72.940000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.665000 17.800000 72.985000 18.120000 ;
      LAYER met4 ;
        RECT 72.665000 17.800000 72.985000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.665000 18.230000 72.985000 18.550000 ;
      LAYER met4 ;
        RECT 72.665000 18.230000 72.985000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.665000 18.660000 72.985000 18.980000 ;
      LAYER met4 ;
        RECT 72.665000 18.660000 72.985000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.665000 19.090000 72.985000 19.410000 ;
      LAYER met4 ;
        RECT 72.665000 19.090000 72.985000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.665000 19.520000 72.985000 19.840000 ;
      LAYER met4 ;
        RECT 72.665000 19.520000 72.985000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.665000 19.950000 72.985000 20.270000 ;
      LAYER met4 ;
        RECT 72.665000 19.950000 72.985000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.665000 20.380000 72.985000 20.700000 ;
      LAYER met4 ;
        RECT 72.665000 20.380000 72.985000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.665000 20.810000 72.985000 21.130000 ;
      LAYER met4 ;
        RECT 72.665000 20.810000 72.985000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.665000 21.240000 72.985000 21.560000 ;
      LAYER met4 ;
        RECT 72.665000 21.240000 72.985000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.665000 21.670000 72.985000 21.990000 ;
      LAYER met4 ;
        RECT 72.665000 21.670000 72.985000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.665000 22.100000 72.985000 22.420000 ;
      LAYER met4 ;
        RECT 72.665000 22.100000 72.985000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 68.065000 73.270000 68.385000 ;
      LAYER met4 ;
        RECT 72.950000 68.065000 73.270000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 68.475000 73.270000 68.795000 ;
      LAYER met4 ;
        RECT 72.950000 68.475000 73.270000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 68.885000 73.270000 69.205000 ;
      LAYER met4 ;
        RECT 72.950000 68.885000 73.270000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 69.295000 73.270000 69.615000 ;
      LAYER met4 ;
        RECT 72.950000 69.295000 73.270000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 69.705000 73.270000 70.025000 ;
      LAYER met4 ;
        RECT 72.950000 69.705000 73.270000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 70.115000 73.270000 70.435000 ;
      LAYER met4 ;
        RECT 72.950000 70.115000 73.270000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 70.525000 73.270000 70.845000 ;
      LAYER met4 ;
        RECT 72.950000 70.525000 73.270000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 70.935000 73.270000 71.255000 ;
      LAYER met4 ;
        RECT 72.950000 70.935000 73.270000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 71.345000 73.270000 71.665000 ;
      LAYER met4 ;
        RECT 72.950000 71.345000 73.270000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 71.755000 73.270000 72.075000 ;
      LAYER met4 ;
        RECT 72.950000 71.755000 73.270000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 72.165000 73.270000 72.485000 ;
      LAYER met4 ;
        RECT 72.950000 72.165000 73.270000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 72.575000 73.270000 72.895000 ;
      LAYER met4 ;
        RECT 72.950000 72.575000 73.270000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 72.985000 73.270000 73.305000 ;
      LAYER met4 ;
        RECT 72.950000 72.985000 73.270000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 73.390000 73.270000 73.710000 ;
      LAYER met4 ;
        RECT 72.950000 73.390000 73.270000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 73.795000 73.270000 74.115000 ;
      LAYER met4 ;
        RECT 72.950000 73.795000 73.270000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 74.200000 73.270000 74.520000 ;
      LAYER met4 ;
        RECT 72.950000 74.200000 73.270000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 74.605000 73.270000 74.925000 ;
      LAYER met4 ;
        RECT 72.950000 74.605000 73.270000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 75.010000 73.270000 75.330000 ;
      LAYER met4 ;
        RECT 72.950000 75.010000 73.270000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 75.415000 73.270000 75.735000 ;
      LAYER met4 ;
        RECT 72.950000 75.415000 73.270000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 75.820000 73.270000 76.140000 ;
      LAYER met4 ;
        RECT 72.950000 75.820000 73.270000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 76.225000 73.270000 76.545000 ;
      LAYER met4 ;
        RECT 72.950000 76.225000 73.270000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 76.630000 73.270000 76.950000 ;
      LAYER met4 ;
        RECT 72.950000 76.630000 73.270000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 77.035000 73.270000 77.355000 ;
      LAYER met4 ;
        RECT 72.950000 77.035000 73.270000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 77.440000 73.270000 77.760000 ;
      LAYER met4 ;
        RECT 72.950000 77.440000 73.270000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 77.845000 73.270000 78.165000 ;
      LAYER met4 ;
        RECT 72.950000 77.845000 73.270000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 78.250000 73.270000 78.570000 ;
      LAYER met4 ;
        RECT 72.950000 78.250000 73.270000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 78.655000 73.270000 78.975000 ;
      LAYER met4 ;
        RECT 72.950000 78.655000 73.270000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 79.060000 73.270000 79.380000 ;
      LAYER met4 ;
        RECT 72.950000 79.060000 73.270000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 79.465000 73.270000 79.785000 ;
      LAYER met4 ;
        RECT 72.950000 79.465000 73.270000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 79.870000 73.270000 80.190000 ;
      LAYER met4 ;
        RECT 72.950000 79.870000 73.270000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 80.275000 73.270000 80.595000 ;
      LAYER met4 ;
        RECT 72.950000 80.275000 73.270000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 80.680000 73.270000 81.000000 ;
      LAYER met4 ;
        RECT 72.950000 80.680000 73.270000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 81.085000 73.270000 81.405000 ;
      LAYER met4 ;
        RECT 72.950000 81.085000 73.270000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 81.490000 73.270000 81.810000 ;
      LAYER met4 ;
        RECT 72.950000 81.490000 73.270000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 81.895000 73.270000 82.215000 ;
      LAYER met4 ;
        RECT 72.950000 81.895000 73.270000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.950000 82.300000 73.270000 82.620000 ;
      LAYER met4 ;
        RECT 72.950000 82.300000 73.270000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 82.795000 73.350000 83.115000 ;
      LAYER met4 ;
        RECT 73.030000 82.795000 73.350000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 83.205000 73.350000 83.525000 ;
      LAYER met4 ;
        RECT 73.030000 83.205000 73.350000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 83.615000 73.350000 83.935000 ;
      LAYER met4 ;
        RECT 73.030000 83.615000 73.350000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 84.025000 73.350000 84.345000 ;
      LAYER met4 ;
        RECT 73.030000 84.025000 73.350000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 84.435000 73.350000 84.755000 ;
      LAYER met4 ;
        RECT 73.030000 84.435000 73.350000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 84.845000 73.350000 85.165000 ;
      LAYER met4 ;
        RECT 73.030000 84.845000 73.350000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 85.255000 73.350000 85.575000 ;
      LAYER met4 ;
        RECT 73.030000 85.255000 73.350000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 85.665000 73.350000 85.985000 ;
      LAYER met4 ;
        RECT 73.030000 85.665000 73.350000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 86.075000 73.350000 86.395000 ;
      LAYER met4 ;
        RECT 73.030000 86.075000 73.350000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 86.485000 73.350000 86.805000 ;
      LAYER met4 ;
        RECT 73.030000 86.485000 73.350000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 86.895000 73.350000 87.215000 ;
      LAYER met4 ;
        RECT 73.030000 86.895000 73.350000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 87.305000 73.350000 87.625000 ;
      LAYER met4 ;
        RECT 73.030000 87.305000 73.350000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 87.715000 73.350000 88.035000 ;
      LAYER met4 ;
        RECT 73.030000 87.715000 73.350000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 88.125000 73.350000 88.445000 ;
      LAYER met4 ;
        RECT 73.030000 88.125000 73.350000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 88.535000 73.350000 88.855000 ;
      LAYER met4 ;
        RECT 73.030000 88.535000 73.350000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 88.945000 73.350000 89.265000 ;
      LAYER met4 ;
        RECT 73.030000 88.945000 73.350000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 89.355000 73.350000 89.675000 ;
      LAYER met4 ;
        RECT 73.030000 89.355000 73.350000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 89.765000 73.350000 90.085000 ;
      LAYER met4 ;
        RECT 73.030000 89.765000 73.350000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 90.175000 73.350000 90.495000 ;
      LAYER met4 ;
        RECT 73.030000 90.175000 73.350000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 90.585000 73.350000 90.905000 ;
      LAYER met4 ;
        RECT 73.030000 90.585000 73.350000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 90.995000 73.350000 91.315000 ;
      LAYER met4 ;
        RECT 73.030000 90.995000 73.350000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 91.405000 73.350000 91.725000 ;
      LAYER met4 ;
        RECT 73.030000 91.405000 73.350000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 91.815000 73.350000 92.135000 ;
      LAYER met4 ;
        RECT 73.030000 91.815000 73.350000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 92.225000 73.350000 92.545000 ;
      LAYER met4 ;
        RECT 73.030000 92.225000 73.350000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030000 92.635000 73.350000 92.955000 ;
      LAYER met4 ;
        RECT 73.030000 92.635000 73.350000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.075000 17.800000 73.395000 18.120000 ;
      LAYER met4 ;
        RECT 73.075000 17.800000 73.395000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.075000 18.230000 73.395000 18.550000 ;
      LAYER met4 ;
        RECT 73.075000 18.230000 73.395000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.075000 18.660000 73.395000 18.980000 ;
      LAYER met4 ;
        RECT 73.075000 18.660000 73.395000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.075000 19.090000 73.395000 19.410000 ;
      LAYER met4 ;
        RECT 73.075000 19.090000 73.395000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.075000 19.520000 73.395000 19.840000 ;
      LAYER met4 ;
        RECT 73.075000 19.520000 73.395000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.075000 19.950000 73.395000 20.270000 ;
      LAYER met4 ;
        RECT 73.075000 19.950000 73.395000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.075000 20.380000 73.395000 20.700000 ;
      LAYER met4 ;
        RECT 73.075000 20.380000 73.395000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.075000 20.810000 73.395000 21.130000 ;
      LAYER met4 ;
        RECT 73.075000 20.810000 73.395000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.075000 21.240000 73.395000 21.560000 ;
      LAYER met4 ;
        RECT 73.075000 21.240000 73.395000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.075000 21.670000 73.395000 21.990000 ;
      LAYER met4 ;
        RECT 73.075000 21.670000 73.395000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.075000 22.100000 73.395000 22.420000 ;
      LAYER met4 ;
        RECT 73.075000 22.100000 73.395000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 68.065000 73.670000 68.385000 ;
      LAYER met4 ;
        RECT 73.350000 68.065000 73.670000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 68.475000 73.670000 68.795000 ;
      LAYER met4 ;
        RECT 73.350000 68.475000 73.670000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 68.885000 73.670000 69.205000 ;
      LAYER met4 ;
        RECT 73.350000 68.885000 73.670000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 69.295000 73.670000 69.615000 ;
      LAYER met4 ;
        RECT 73.350000 69.295000 73.670000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 69.705000 73.670000 70.025000 ;
      LAYER met4 ;
        RECT 73.350000 69.705000 73.670000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 70.115000 73.670000 70.435000 ;
      LAYER met4 ;
        RECT 73.350000 70.115000 73.670000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 70.525000 73.670000 70.845000 ;
      LAYER met4 ;
        RECT 73.350000 70.525000 73.670000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 70.935000 73.670000 71.255000 ;
      LAYER met4 ;
        RECT 73.350000 70.935000 73.670000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 71.345000 73.670000 71.665000 ;
      LAYER met4 ;
        RECT 73.350000 71.345000 73.670000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 71.755000 73.670000 72.075000 ;
      LAYER met4 ;
        RECT 73.350000 71.755000 73.670000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 72.165000 73.670000 72.485000 ;
      LAYER met4 ;
        RECT 73.350000 72.165000 73.670000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 72.575000 73.670000 72.895000 ;
      LAYER met4 ;
        RECT 73.350000 72.575000 73.670000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 72.985000 73.670000 73.305000 ;
      LAYER met4 ;
        RECT 73.350000 72.985000 73.670000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 73.390000 73.670000 73.710000 ;
      LAYER met4 ;
        RECT 73.350000 73.390000 73.670000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 73.795000 73.670000 74.115000 ;
      LAYER met4 ;
        RECT 73.350000 73.795000 73.670000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 74.200000 73.670000 74.520000 ;
      LAYER met4 ;
        RECT 73.350000 74.200000 73.670000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 74.605000 73.670000 74.925000 ;
      LAYER met4 ;
        RECT 73.350000 74.605000 73.670000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 75.010000 73.670000 75.330000 ;
      LAYER met4 ;
        RECT 73.350000 75.010000 73.670000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 75.415000 73.670000 75.735000 ;
      LAYER met4 ;
        RECT 73.350000 75.415000 73.670000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 75.820000 73.670000 76.140000 ;
      LAYER met4 ;
        RECT 73.350000 75.820000 73.670000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 76.225000 73.670000 76.545000 ;
      LAYER met4 ;
        RECT 73.350000 76.225000 73.670000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 76.630000 73.670000 76.950000 ;
      LAYER met4 ;
        RECT 73.350000 76.630000 73.670000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 77.035000 73.670000 77.355000 ;
      LAYER met4 ;
        RECT 73.350000 77.035000 73.670000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 77.440000 73.670000 77.760000 ;
      LAYER met4 ;
        RECT 73.350000 77.440000 73.670000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 77.845000 73.670000 78.165000 ;
      LAYER met4 ;
        RECT 73.350000 77.845000 73.670000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 78.250000 73.670000 78.570000 ;
      LAYER met4 ;
        RECT 73.350000 78.250000 73.670000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 78.655000 73.670000 78.975000 ;
      LAYER met4 ;
        RECT 73.350000 78.655000 73.670000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 79.060000 73.670000 79.380000 ;
      LAYER met4 ;
        RECT 73.350000 79.060000 73.670000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 79.465000 73.670000 79.785000 ;
      LAYER met4 ;
        RECT 73.350000 79.465000 73.670000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 79.870000 73.670000 80.190000 ;
      LAYER met4 ;
        RECT 73.350000 79.870000 73.670000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 80.275000 73.670000 80.595000 ;
      LAYER met4 ;
        RECT 73.350000 80.275000 73.670000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 80.680000 73.670000 81.000000 ;
      LAYER met4 ;
        RECT 73.350000 80.680000 73.670000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 81.085000 73.670000 81.405000 ;
      LAYER met4 ;
        RECT 73.350000 81.085000 73.670000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 81.490000 73.670000 81.810000 ;
      LAYER met4 ;
        RECT 73.350000 81.490000 73.670000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 81.895000 73.670000 82.215000 ;
      LAYER met4 ;
        RECT 73.350000 81.895000 73.670000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.350000 82.300000 73.670000 82.620000 ;
      LAYER met4 ;
        RECT 73.350000 82.300000 73.670000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 82.795000 73.760000 83.115000 ;
      LAYER met4 ;
        RECT 73.440000 82.795000 73.760000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 83.205000 73.760000 83.525000 ;
      LAYER met4 ;
        RECT 73.440000 83.205000 73.760000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 83.615000 73.760000 83.935000 ;
      LAYER met4 ;
        RECT 73.440000 83.615000 73.760000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 84.025000 73.760000 84.345000 ;
      LAYER met4 ;
        RECT 73.440000 84.025000 73.760000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 84.435000 73.760000 84.755000 ;
      LAYER met4 ;
        RECT 73.440000 84.435000 73.760000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 84.845000 73.760000 85.165000 ;
      LAYER met4 ;
        RECT 73.440000 84.845000 73.760000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 85.255000 73.760000 85.575000 ;
      LAYER met4 ;
        RECT 73.440000 85.255000 73.760000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 85.665000 73.760000 85.985000 ;
      LAYER met4 ;
        RECT 73.440000 85.665000 73.760000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 86.075000 73.760000 86.395000 ;
      LAYER met4 ;
        RECT 73.440000 86.075000 73.760000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 86.485000 73.760000 86.805000 ;
      LAYER met4 ;
        RECT 73.440000 86.485000 73.760000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 86.895000 73.760000 87.215000 ;
      LAYER met4 ;
        RECT 73.440000 86.895000 73.760000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 87.305000 73.760000 87.625000 ;
      LAYER met4 ;
        RECT 73.440000 87.305000 73.760000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 87.715000 73.760000 88.035000 ;
      LAYER met4 ;
        RECT 73.440000 87.715000 73.760000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 88.125000 73.760000 88.445000 ;
      LAYER met4 ;
        RECT 73.440000 88.125000 73.760000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 88.535000 73.760000 88.855000 ;
      LAYER met4 ;
        RECT 73.440000 88.535000 73.760000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 88.945000 73.760000 89.265000 ;
      LAYER met4 ;
        RECT 73.440000 88.945000 73.760000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 89.355000 73.760000 89.675000 ;
      LAYER met4 ;
        RECT 73.440000 89.355000 73.760000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 89.765000 73.760000 90.085000 ;
      LAYER met4 ;
        RECT 73.440000 89.765000 73.760000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 90.175000 73.760000 90.495000 ;
      LAYER met4 ;
        RECT 73.440000 90.175000 73.760000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 90.585000 73.760000 90.905000 ;
      LAYER met4 ;
        RECT 73.440000 90.585000 73.760000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 90.995000 73.760000 91.315000 ;
      LAYER met4 ;
        RECT 73.440000 90.995000 73.760000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 91.405000 73.760000 91.725000 ;
      LAYER met4 ;
        RECT 73.440000 91.405000 73.760000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 91.815000 73.760000 92.135000 ;
      LAYER met4 ;
        RECT 73.440000 91.815000 73.760000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 92.225000 73.760000 92.545000 ;
      LAYER met4 ;
        RECT 73.440000 92.225000 73.760000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440000 92.635000 73.760000 92.955000 ;
      LAYER met4 ;
        RECT 73.440000 92.635000 73.760000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.485000 17.800000 73.805000 18.120000 ;
      LAYER met4 ;
        RECT 73.485000 17.800000 73.805000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.485000 18.230000 73.805000 18.550000 ;
      LAYER met4 ;
        RECT 73.485000 18.230000 73.805000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.485000 18.660000 73.805000 18.980000 ;
      LAYER met4 ;
        RECT 73.485000 18.660000 73.805000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.485000 19.090000 73.805000 19.410000 ;
      LAYER met4 ;
        RECT 73.485000 19.090000 73.805000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.485000 19.520000 73.805000 19.840000 ;
      LAYER met4 ;
        RECT 73.485000 19.520000 73.805000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.485000 19.950000 73.805000 20.270000 ;
      LAYER met4 ;
        RECT 73.485000 19.950000 73.805000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.485000 20.380000 73.805000 20.700000 ;
      LAYER met4 ;
        RECT 73.485000 20.380000 73.805000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.485000 20.810000 73.805000 21.130000 ;
      LAYER met4 ;
        RECT 73.485000 20.810000 73.805000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.485000 21.240000 73.805000 21.560000 ;
      LAYER met4 ;
        RECT 73.485000 21.240000 73.805000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.485000 21.670000 73.805000 21.990000 ;
      LAYER met4 ;
        RECT 73.485000 21.670000 73.805000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.485000 22.100000 73.805000 22.420000 ;
      LAYER met4 ;
        RECT 73.485000 22.100000 73.805000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 68.065000 74.070000 68.385000 ;
      LAYER met4 ;
        RECT 73.750000 68.065000 74.070000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 68.475000 74.070000 68.795000 ;
      LAYER met4 ;
        RECT 73.750000 68.475000 74.070000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 68.885000 74.070000 69.205000 ;
      LAYER met4 ;
        RECT 73.750000 68.885000 74.070000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 69.295000 74.070000 69.615000 ;
      LAYER met4 ;
        RECT 73.750000 69.295000 74.070000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 69.705000 74.070000 70.025000 ;
      LAYER met4 ;
        RECT 73.750000 69.705000 74.070000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 70.115000 74.070000 70.435000 ;
      LAYER met4 ;
        RECT 73.750000 70.115000 74.070000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 70.525000 74.070000 70.845000 ;
      LAYER met4 ;
        RECT 73.750000 70.525000 74.070000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 70.935000 74.070000 71.255000 ;
      LAYER met4 ;
        RECT 73.750000 70.935000 74.070000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 71.345000 74.070000 71.665000 ;
      LAYER met4 ;
        RECT 73.750000 71.345000 74.070000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 71.755000 74.070000 72.075000 ;
      LAYER met4 ;
        RECT 73.750000 71.755000 74.070000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 72.165000 74.070000 72.485000 ;
      LAYER met4 ;
        RECT 73.750000 72.165000 74.070000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 72.575000 74.070000 72.895000 ;
      LAYER met4 ;
        RECT 73.750000 72.575000 74.070000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 72.985000 74.070000 73.305000 ;
      LAYER met4 ;
        RECT 73.750000 72.985000 74.070000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 73.390000 74.070000 73.710000 ;
      LAYER met4 ;
        RECT 73.750000 73.390000 74.070000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 73.795000 74.070000 74.115000 ;
      LAYER met4 ;
        RECT 73.750000 73.795000 74.070000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 74.200000 74.070000 74.520000 ;
      LAYER met4 ;
        RECT 73.750000 74.200000 74.070000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 74.605000 74.070000 74.925000 ;
      LAYER met4 ;
        RECT 73.750000 74.605000 74.070000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 75.010000 74.070000 75.330000 ;
      LAYER met4 ;
        RECT 73.750000 75.010000 74.070000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 75.415000 74.070000 75.735000 ;
      LAYER met4 ;
        RECT 73.750000 75.415000 74.070000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 75.820000 74.070000 76.140000 ;
      LAYER met4 ;
        RECT 73.750000 75.820000 74.070000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 76.225000 74.070000 76.545000 ;
      LAYER met4 ;
        RECT 73.750000 76.225000 74.070000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 76.630000 74.070000 76.950000 ;
      LAYER met4 ;
        RECT 73.750000 76.630000 74.070000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 77.035000 74.070000 77.355000 ;
      LAYER met4 ;
        RECT 73.750000 77.035000 74.070000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 77.440000 74.070000 77.760000 ;
      LAYER met4 ;
        RECT 73.750000 77.440000 74.070000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 77.845000 74.070000 78.165000 ;
      LAYER met4 ;
        RECT 73.750000 77.845000 74.070000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 78.250000 74.070000 78.570000 ;
      LAYER met4 ;
        RECT 73.750000 78.250000 74.070000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 78.655000 74.070000 78.975000 ;
      LAYER met4 ;
        RECT 73.750000 78.655000 74.070000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 79.060000 74.070000 79.380000 ;
      LAYER met4 ;
        RECT 73.750000 79.060000 74.070000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 79.465000 74.070000 79.785000 ;
      LAYER met4 ;
        RECT 73.750000 79.465000 74.070000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 79.870000 74.070000 80.190000 ;
      LAYER met4 ;
        RECT 73.750000 79.870000 74.070000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 80.275000 74.070000 80.595000 ;
      LAYER met4 ;
        RECT 73.750000 80.275000 74.070000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 80.680000 74.070000 81.000000 ;
      LAYER met4 ;
        RECT 73.750000 80.680000 74.070000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 81.085000 74.070000 81.405000 ;
      LAYER met4 ;
        RECT 73.750000 81.085000 74.070000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 81.490000 74.070000 81.810000 ;
      LAYER met4 ;
        RECT 73.750000 81.490000 74.070000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 81.895000 74.070000 82.215000 ;
      LAYER met4 ;
        RECT 73.750000 81.895000 74.070000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.750000 82.300000 74.070000 82.620000 ;
      LAYER met4 ;
        RECT 73.750000 82.300000 74.070000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 82.795000 74.170000 83.115000 ;
      LAYER met4 ;
        RECT 73.850000 82.795000 74.170000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 83.205000 74.170000 83.525000 ;
      LAYER met4 ;
        RECT 73.850000 83.205000 74.170000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 83.615000 74.170000 83.935000 ;
      LAYER met4 ;
        RECT 73.850000 83.615000 74.170000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 84.025000 74.170000 84.345000 ;
      LAYER met4 ;
        RECT 73.850000 84.025000 74.170000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 84.435000 74.170000 84.755000 ;
      LAYER met4 ;
        RECT 73.850000 84.435000 74.170000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 84.845000 74.170000 85.165000 ;
      LAYER met4 ;
        RECT 73.850000 84.845000 74.170000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 85.255000 74.170000 85.575000 ;
      LAYER met4 ;
        RECT 73.850000 85.255000 74.170000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 85.665000 74.170000 85.985000 ;
      LAYER met4 ;
        RECT 73.850000 85.665000 74.170000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 86.075000 74.170000 86.395000 ;
      LAYER met4 ;
        RECT 73.850000 86.075000 74.170000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 86.485000 74.170000 86.805000 ;
      LAYER met4 ;
        RECT 73.850000 86.485000 74.170000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 86.895000 74.170000 87.215000 ;
      LAYER met4 ;
        RECT 73.850000 86.895000 74.170000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 87.305000 74.170000 87.625000 ;
      LAYER met4 ;
        RECT 73.850000 87.305000 74.170000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 87.715000 74.170000 88.035000 ;
      LAYER met4 ;
        RECT 73.850000 87.715000 74.170000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 88.125000 74.170000 88.445000 ;
      LAYER met4 ;
        RECT 73.850000 88.125000 74.170000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 88.535000 74.170000 88.855000 ;
      LAYER met4 ;
        RECT 73.850000 88.535000 74.170000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 88.945000 74.170000 89.265000 ;
      LAYER met4 ;
        RECT 73.850000 88.945000 74.170000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 89.355000 74.170000 89.675000 ;
      LAYER met4 ;
        RECT 73.850000 89.355000 74.170000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 89.765000 74.170000 90.085000 ;
      LAYER met4 ;
        RECT 73.850000 89.765000 74.170000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 90.175000 74.170000 90.495000 ;
      LAYER met4 ;
        RECT 73.850000 90.175000 74.170000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 90.585000 74.170000 90.905000 ;
      LAYER met4 ;
        RECT 73.850000 90.585000 74.170000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 90.995000 74.170000 91.315000 ;
      LAYER met4 ;
        RECT 73.850000 90.995000 74.170000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 91.405000 74.170000 91.725000 ;
      LAYER met4 ;
        RECT 73.850000 91.405000 74.170000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 91.815000 74.170000 92.135000 ;
      LAYER met4 ;
        RECT 73.850000 91.815000 74.170000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 92.225000 74.170000 92.545000 ;
      LAYER met4 ;
        RECT 73.850000 92.225000 74.170000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850000 92.635000 74.170000 92.955000 ;
      LAYER met4 ;
        RECT 73.850000 92.635000 74.170000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.895000 17.800000 74.215000 18.120000 ;
      LAYER met4 ;
        RECT 73.895000 17.800000 74.215000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.895000 18.230000 74.215000 18.550000 ;
      LAYER met4 ;
        RECT 73.895000 18.230000 74.215000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.895000 18.660000 74.215000 18.980000 ;
      LAYER met4 ;
        RECT 73.895000 18.660000 74.215000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.895000 19.090000 74.215000 19.410000 ;
      LAYER met4 ;
        RECT 73.895000 19.090000 74.215000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.895000 19.520000 74.215000 19.840000 ;
      LAYER met4 ;
        RECT 73.895000 19.520000 74.215000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.895000 19.950000 74.215000 20.270000 ;
      LAYER met4 ;
        RECT 73.895000 19.950000 74.215000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.895000 20.380000 74.215000 20.700000 ;
      LAYER met4 ;
        RECT 73.895000 20.380000 74.215000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.895000 20.810000 74.215000 21.130000 ;
      LAYER met4 ;
        RECT 73.895000 20.810000 74.215000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.895000 21.240000 74.215000 21.560000 ;
      LAYER met4 ;
        RECT 73.895000 21.240000 74.215000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.895000 21.670000 74.215000 21.990000 ;
      LAYER met4 ;
        RECT 73.895000 21.670000 74.215000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.895000 22.100000 74.215000 22.420000 ;
      LAYER met4 ;
        RECT 73.895000 22.100000 74.215000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 68.065000 74.470000 68.385000 ;
      LAYER met4 ;
        RECT 74.150000 68.065000 74.470000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 68.475000 74.470000 68.795000 ;
      LAYER met4 ;
        RECT 74.150000 68.475000 74.470000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 68.885000 74.470000 69.205000 ;
      LAYER met4 ;
        RECT 74.150000 68.885000 74.470000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 69.295000 74.470000 69.615000 ;
      LAYER met4 ;
        RECT 74.150000 69.295000 74.470000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 69.705000 74.470000 70.025000 ;
      LAYER met4 ;
        RECT 74.150000 69.705000 74.470000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 70.115000 74.470000 70.435000 ;
      LAYER met4 ;
        RECT 74.150000 70.115000 74.470000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 70.525000 74.470000 70.845000 ;
      LAYER met4 ;
        RECT 74.150000 70.525000 74.470000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 70.935000 74.470000 71.255000 ;
      LAYER met4 ;
        RECT 74.150000 70.935000 74.470000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 71.345000 74.470000 71.665000 ;
      LAYER met4 ;
        RECT 74.150000 71.345000 74.470000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 71.755000 74.470000 72.075000 ;
      LAYER met4 ;
        RECT 74.150000 71.755000 74.470000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 72.165000 74.470000 72.485000 ;
      LAYER met4 ;
        RECT 74.150000 72.165000 74.470000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 72.575000 74.470000 72.895000 ;
      LAYER met4 ;
        RECT 74.150000 72.575000 74.470000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 72.985000 74.470000 73.305000 ;
      LAYER met4 ;
        RECT 74.150000 72.985000 74.470000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 73.390000 74.470000 73.710000 ;
      LAYER met4 ;
        RECT 74.150000 73.390000 74.470000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 73.795000 74.470000 74.115000 ;
      LAYER met4 ;
        RECT 74.150000 73.795000 74.470000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 74.200000 74.470000 74.520000 ;
      LAYER met4 ;
        RECT 74.150000 74.200000 74.470000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 74.605000 74.470000 74.925000 ;
      LAYER met4 ;
        RECT 74.150000 74.605000 74.470000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 75.010000 74.470000 75.330000 ;
      LAYER met4 ;
        RECT 74.150000 75.010000 74.470000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 75.415000 74.470000 75.735000 ;
      LAYER met4 ;
        RECT 74.150000 75.415000 74.470000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 75.820000 74.470000 76.140000 ;
      LAYER met4 ;
        RECT 74.150000 75.820000 74.470000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 76.225000 74.470000 76.545000 ;
      LAYER met4 ;
        RECT 74.150000 76.225000 74.470000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 76.630000 74.470000 76.950000 ;
      LAYER met4 ;
        RECT 74.150000 76.630000 74.470000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 77.035000 74.470000 77.355000 ;
      LAYER met4 ;
        RECT 74.150000 77.035000 74.470000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 77.440000 74.470000 77.760000 ;
      LAYER met4 ;
        RECT 74.150000 77.440000 74.470000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 77.845000 74.470000 78.165000 ;
      LAYER met4 ;
        RECT 74.150000 77.845000 74.470000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 78.250000 74.470000 78.570000 ;
      LAYER met4 ;
        RECT 74.150000 78.250000 74.470000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 78.655000 74.470000 78.975000 ;
      LAYER met4 ;
        RECT 74.150000 78.655000 74.470000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 79.060000 74.470000 79.380000 ;
      LAYER met4 ;
        RECT 74.150000 79.060000 74.470000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 79.465000 74.470000 79.785000 ;
      LAYER met4 ;
        RECT 74.150000 79.465000 74.470000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 79.870000 74.470000 80.190000 ;
      LAYER met4 ;
        RECT 74.150000 79.870000 74.470000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 80.275000 74.470000 80.595000 ;
      LAYER met4 ;
        RECT 74.150000 80.275000 74.470000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 80.680000 74.470000 81.000000 ;
      LAYER met4 ;
        RECT 74.150000 80.680000 74.470000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 81.085000 74.470000 81.405000 ;
      LAYER met4 ;
        RECT 74.150000 81.085000 74.470000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 81.490000 74.470000 81.810000 ;
      LAYER met4 ;
        RECT 74.150000 81.490000 74.470000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 81.895000 74.470000 82.215000 ;
      LAYER met4 ;
        RECT 74.150000 81.895000 74.470000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.150000 82.300000 74.470000 82.620000 ;
      LAYER met4 ;
        RECT 74.150000 82.300000 74.470000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 82.795000 74.580000 83.115000 ;
      LAYER met4 ;
        RECT 74.260000 82.795000 74.580000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 83.205000 74.580000 83.525000 ;
      LAYER met4 ;
        RECT 74.260000 83.205000 74.580000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 83.615000 74.580000 83.935000 ;
      LAYER met4 ;
        RECT 74.260000 83.615000 74.580000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 84.025000 74.580000 84.345000 ;
      LAYER met4 ;
        RECT 74.260000 84.025000 74.580000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 84.435000 74.580000 84.755000 ;
      LAYER met4 ;
        RECT 74.260000 84.435000 74.580000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 84.845000 74.580000 85.165000 ;
      LAYER met4 ;
        RECT 74.260000 84.845000 74.580000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 85.255000 74.580000 85.575000 ;
      LAYER met4 ;
        RECT 74.260000 85.255000 74.580000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 85.665000 74.580000 85.985000 ;
      LAYER met4 ;
        RECT 74.260000 85.665000 74.580000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 86.075000 74.580000 86.395000 ;
      LAYER met4 ;
        RECT 74.260000 86.075000 74.580000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 86.485000 74.580000 86.805000 ;
      LAYER met4 ;
        RECT 74.260000 86.485000 74.580000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 86.895000 74.580000 87.215000 ;
      LAYER met4 ;
        RECT 74.260000 86.895000 74.580000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 87.305000 74.580000 87.625000 ;
      LAYER met4 ;
        RECT 74.260000 87.305000 74.580000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 87.715000 74.580000 88.035000 ;
      LAYER met4 ;
        RECT 74.260000 87.715000 74.580000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 88.125000 74.580000 88.445000 ;
      LAYER met4 ;
        RECT 74.260000 88.125000 74.580000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 88.535000 74.580000 88.855000 ;
      LAYER met4 ;
        RECT 74.260000 88.535000 74.580000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 88.945000 74.580000 89.265000 ;
      LAYER met4 ;
        RECT 74.260000 88.945000 74.580000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 89.355000 74.580000 89.675000 ;
      LAYER met4 ;
        RECT 74.260000 89.355000 74.580000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 89.765000 74.580000 90.085000 ;
      LAYER met4 ;
        RECT 74.260000 89.765000 74.580000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 90.175000 74.580000 90.495000 ;
      LAYER met4 ;
        RECT 74.260000 90.175000 74.580000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 90.585000 74.580000 90.905000 ;
      LAYER met4 ;
        RECT 74.260000 90.585000 74.580000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 90.995000 74.580000 91.315000 ;
      LAYER met4 ;
        RECT 74.260000 90.995000 74.580000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 91.405000 74.580000 91.725000 ;
      LAYER met4 ;
        RECT 74.260000 91.405000 74.580000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 91.815000 74.580000 92.135000 ;
      LAYER met4 ;
        RECT 74.260000 91.815000 74.580000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 92.225000 74.580000 92.545000 ;
      LAYER met4 ;
        RECT 74.260000 92.225000 74.580000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260000 92.635000 74.580000 92.955000 ;
      LAYER met4 ;
        RECT 74.260000 92.635000 74.580000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 17.800000 74.625000 18.120000 ;
      LAYER met4 ;
        RECT 74.305000 17.800000 74.625000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 18.230000 74.625000 18.550000 ;
      LAYER met4 ;
        RECT 74.305000 18.230000 74.625000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 18.660000 74.625000 18.980000 ;
      LAYER met4 ;
        RECT 74.305000 18.660000 74.625000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 19.090000 74.625000 19.410000 ;
      LAYER met4 ;
        RECT 74.305000 19.090000 74.625000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 19.520000 74.625000 19.840000 ;
      LAYER met4 ;
        RECT 74.305000 19.520000 74.625000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 19.950000 74.625000 20.270000 ;
      LAYER met4 ;
        RECT 74.305000 19.950000 74.625000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 20.380000 74.625000 20.700000 ;
      LAYER met4 ;
        RECT 74.305000 20.380000 74.625000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 20.810000 74.625000 21.130000 ;
      LAYER met4 ;
        RECT 74.305000 20.810000 74.625000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 21.240000 74.625000 21.560000 ;
      LAYER met4 ;
        RECT 74.305000 21.240000 74.625000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 21.670000 74.625000 21.990000 ;
      LAYER met4 ;
        RECT 74.305000 21.670000 74.625000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 22.100000 74.625000 22.420000 ;
      LAYER met4 ;
        RECT 74.305000 22.100000 74.625000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 82.795000 8.375000 83.115000 ;
      LAYER met4 ;
        RECT 8.055000 82.795000 8.375000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 83.205000 8.375000 83.525000 ;
      LAYER met4 ;
        RECT 8.055000 83.205000 8.375000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 83.615000 8.375000 83.935000 ;
      LAYER met4 ;
        RECT 8.055000 83.615000 8.375000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 84.025000 8.375000 84.345000 ;
      LAYER met4 ;
        RECT 8.055000 84.025000 8.375000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 84.435000 8.375000 84.755000 ;
      LAYER met4 ;
        RECT 8.055000 84.435000 8.375000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 84.845000 8.375000 85.165000 ;
      LAYER met4 ;
        RECT 8.055000 84.845000 8.375000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 85.255000 8.375000 85.575000 ;
      LAYER met4 ;
        RECT 8.055000 85.255000 8.375000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 85.665000 8.375000 85.985000 ;
      LAYER met4 ;
        RECT 8.055000 85.665000 8.375000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 86.075000 8.375000 86.395000 ;
      LAYER met4 ;
        RECT 8.055000 86.075000 8.375000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 86.485000 8.375000 86.805000 ;
      LAYER met4 ;
        RECT 8.055000 86.485000 8.375000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 86.895000 8.375000 87.215000 ;
      LAYER met4 ;
        RECT 8.055000 86.895000 8.375000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 87.305000 8.375000 87.625000 ;
      LAYER met4 ;
        RECT 8.055000 87.305000 8.375000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 87.715000 8.375000 88.035000 ;
      LAYER met4 ;
        RECT 8.055000 87.715000 8.375000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 88.125000 8.375000 88.445000 ;
      LAYER met4 ;
        RECT 8.055000 88.125000 8.375000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 88.535000 8.375000 88.855000 ;
      LAYER met4 ;
        RECT 8.055000 88.535000 8.375000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 88.945000 8.375000 89.265000 ;
      LAYER met4 ;
        RECT 8.055000 88.945000 8.375000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 89.355000 8.375000 89.675000 ;
      LAYER met4 ;
        RECT 8.055000 89.355000 8.375000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 89.765000 8.375000 90.085000 ;
      LAYER met4 ;
        RECT 8.055000 89.765000 8.375000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 90.175000 8.375000 90.495000 ;
      LAYER met4 ;
        RECT 8.055000 90.175000 8.375000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 90.585000 8.375000 90.905000 ;
      LAYER met4 ;
        RECT 8.055000 90.585000 8.375000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 90.995000 8.375000 91.315000 ;
      LAYER met4 ;
        RECT 8.055000 90.995000 8.375000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 91.405000 8.375000 91.725000 ;
      LAYER met4 ;
        RECT 8.055000 91.405000 8.375000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 91.815000 8.375000 92.135000 ;
      LAYER met4 ;
        RECT 8.055000 91.815000 8.375000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 92.225000 8.375000 92.545000 ;
      LAYER met4 ;
        RECT 8.055000 92.225000 8.375000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055000 92.635000 8.375000 92.955000 ;
      LAYER met4 ;
        RECT 8.055000 92.635000 8.375000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325000 17.800000 8.645000 18.120000 ;
      LAYER met4 ;
        RECT 8.325000 17.800000 8.645000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325000 18.230000 8.645000 18.550000 ;
      LAYER met4 ;
        RECT 8.325000 18.230000 8.645000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325000 18.660000 8.645000 18.980000 ;
      LAYER met4 ;
        RECT 8.325000 18.660000 8.645000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325000 19.090000 8.645000 19.410000 ;
      LAYER met4 ;
        RECT 8.325000 19.090000 8.645000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325000 19.520000 8.645000 19.840000 ;
      LAYER met4 ;
        RECT 8.325000 19.520000 8.645000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325000 19.950000 8.645000 20.270000 ;
      LAYER met4 ;
        RECT 8.325000 19.950000 8.645000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325000 20.380000 8.645000 20.700000 ;
      LAYER met4 ;
        RECT 8.325000 20.380000 8.645000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325000 20.810000 8.645000 21.130000 ;
      LAYER met4 ;
        RECT 8.325000 20.810000 8.645000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325000 21.240000 8.645000 21.560000 ;
      LAYER met4 ;
        RECT 8.325000 21.240000 8.645000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325000 21.670000 8.645000 21.990000 ;
      LAYER met4 ;
        RECT 8.325000 21.670000 8.645000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325000 22.100000 8.645000 22.420000 ;
      LAYER met4 ;
        RECT 8.325000 22.100000 8.645000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 68.065000 8.705000 68.385000 ;
      LAYER met4 ;
        RECT 8.385000 68.065000 8.705000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 68.475000 8.705000 68.795000 ;
      LAYER met4 ;
        RECT 8.385000 68.475000 8.705000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 68.885000 8.705000 69.205000 ;
      LAYER met4 ;
        RECT 8.385000 68.885000 8.705000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 69.295000 8.705000 69.615000 ;
      LAYER met4 ;
        RECT 8.385000 69.295000 8.705000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 69.705000 8.705000 70.025000 ;
      LAYER met4 ;
        RECT 8.385000 69.705000 8.705000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 70.115000 8.705000 70.435000 ;
      LAYER met4 ;
        RECT 8.385000 70.115000 8.705000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 70.525000 8.705000 70.845000 ;
      LAYER met4 ;
        RECT 8.385000 70.525000 8.705000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 70.935000 8.705000 71.255000 ;
      LAYER met4 ;
        RECT 8.385000 70.935000 8.705000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 71.345000 8.705000 71.665000 ;
      LAYER met4 ;
        RECT 8.385000 71.345000 8.705000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 71.755000 8.705000 72.075000 ;
      LAYER met4 ;
        RECT 8.385000 71.755000 8.705000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 72.165000 8.705000 72.485000 ;
      LAYER met4 ;
        RECT 8.385000 72.165000 8.705000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 72.575000 8.705000 72.895000 ;
      LAYER met4 ;
        RECT 8.385000 72.575000 8.705000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 72.985000 8.705000 73.305000 ;
      LAYER met4 ;
        RECT 8.385000 72.985000 8.705000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 73.390000 8.705000 73.710000 ;
      LAYER met4 ;
        RECT 8.385000 73.390000 8.705000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 73.795000 8.705000 74.115000 ;
      LAYER met4 ;
        RECT 8.385000 73.795000 8.705000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 74.200000 8.705000 74.520000 ;
      LAYER met4 ;
        RECT 8.385000 74.200000 8.705000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 74.605000 8.705000 74.925000 ;
      LAYER met4 ;
        RECT 8.385000 74.605000 8.705000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 75.010000 8.705000 75.330000 ;
      LAYER met4 ;
        RECT 8.385000 75.010000 8.705000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 75.415000 8.705000 75.735000 ;
      LAYER met4 ;
        RECT 8.385000 75.415000 8.705000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 75.820000 8.705000 76.140000 ;
      LAYER met4 ;
        RECT 8.385000 75.820000 8.705000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 76.225000 8.705000 76.545000 ;
      LAYER met4 ;
        RECT 8.385000 76.225000 8.705000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 76.630000 8.705000 76.950000 ;
      LAYER met4 ;
        RECT 8.385000 76.630000 8.705000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 77.035000 8.705000 77.355000 ;
      LAYER met4 ;
        RECT 8.385000 77.035000 8.705000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 77.440000 8.705000 77.760000 ;
      LAYER met4 ;
        RECT 8.385000 77.440000 8.705000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 77.845000 8.705000 78.165000 ;
      LAYER met4 ;
        RECT 8.385000 77.845000 8.705000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 78.250000 8.705000 78.570000 ;
      LAYER met4 ;
        RECT 8.385000 78.250000 8.705000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 78.655000 8.705000 78.975000 ;
      LAYER met4 ;
        RECT 8.385000 78.655000 8.705000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 79.060000 8.705000 79.380000 ;
      LAYER met4 ;
        RECT 8.385000 79.060000 8.705000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 79.465000 8.705000 79.785000 ;
      LAYER met4 ;
        RECT 8.385000 79.465000 8.705000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 79.870000 8.705000 80.190000 ;
      LAYER met4 ;
        RECT 8.385000 79.870000 8.705000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 80.275000 8.705000 80.595000 ;
      LAYER met4 ;
        RECT 8.385000 80.275000 8.705000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 80.680000 8.705000 81.000000 ;
      LAYER met4 ;
        RECT 8.385000 80.680000 8.705000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 81.085000 8.705000 81.405000 ;
      LAYER met4 ;
        RECT 8.385000 81.085000 8.705000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 81.490000 8.705000 81.810000 ;
      LAYER met4 ;
        RECT 8.385000 81.490000 8.705000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 81.895000 8.705000 82.215000 ;
      LAYER met4 ;
        RECT 8.385000 81.895000 8.705000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385000 82.300000 8.705000 82.620000 ;
      LAYER met4 ;
        RECT 8.385000 82.300000 8.705000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 82.795000 8.785000 83.115000 ;
      LAYER met4 ;
        RECT 8.465000 82.795000 8.785000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 83.205000 8.785000 83.525000 ;
      LAYER met4 ;
        RECT 8.465000 83.205000 8.785000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 83.615000 8.785000 83.935000 ;
      LAYER met4 ;
        RECT 8.465000 83.615000 8.785000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 84.025000 8.785000 84.345000 ;
      LAYER met4 ;
        RECT 8.465000 84.025000 8.785000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 84.435000 8.785000 84.755000 ;
      LAYER met4 ;
        RECT 8.465000 84.435000 8.785000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 84.845000 8.785000 85.165000 ;
      LAYER met4 ;
        RECT 8.465000 84.845000 8.785000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 85.255000 8.785000 85.575000 ;
      LAYER met4 ;
        RECT 8.465000 85.255000 8.785000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 85.665000 8.785000 85.985000 ;
      LAYER met4 ;
        RECT 8.465000 85.665000 8.785000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 86.075000 8.785000 86.395000 ;
      LAYER met4 ;
        RECT 8.465000 86.075000 8.785000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 86.485000 8.785000 86.805000 ;
      LAYER met4 ;
        RECT 8.465000 86.485000 8.785000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 86.895000 8.785000 87.215000 ;
      LAYER met4 ;
        RECT 8.465000 86.895000 8.785000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 87.305000 8.785000 87.625000 ;
      LAYER met4 ;
        RECT 8.465000 87.305000 8.785000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 87.715000 8.785000 88.035000 ;
      LAYER met4 ;
        RECT 8.465000 87.715000 8.785000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 88.125000 8.785000 88.445000 ;
      LAYER met4 ;
        RECT 8.465000 88.125000 8.785000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 88.535000 8.785000 88.855000 ;
      LAYER met4 ;
        RECT 8.465000 88.535000 8.785000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 88.945000 8.785000 89.265000 ;
      LAYER met4 ;
        RECT 8.465000 88.945000 8.785000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 89.355000 8.785000 89.675000 ;
      LAYER met4 ;
        RECT 8.465000 89.355000 8.785000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 89.765000 8.785000 90.085000 ;
      LAYER met4 ;
        RECT 8.465000 89.765000 8.785000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 90.175000 8.785000 90.495000 ;
      LAYER met4 ;
        RECT 8.465000 90.175000 8.785000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 90.585000 8.785000 90.905000 ;
      LAYER met4 ;
        RECT 8.465000 90.585000 8.785000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 90.995000 8.785000 91.315000 ;
      LAYER met4 ;
        RECT 8.465000 90.995000 8.785000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 91.405000 8.785000 91.725000 ;
      LAYER met4 ;
        RECT 8.465000 91.405000 8.785000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 91.815000 8.785000 92.135000 ;
      LAYER met4 ;
        RECT 8.465000 91.815000 8.785000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 92.225000 8.785000 92.545000 ;
      LAYER met4 ;
        RECT 8.465000 92.225000 8.785000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465000 92.635000 8.785000 92.955000 ;
      LAYER met4 ;
        RECT 8.465000 92.635000 8.785000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730000 17.800000 9.050000 18.120000 ;
      LAYER met4 ;
        RECT 8.730000 17.800000 9.050000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730000 18.230000 9.050000 18.550000 ;
      LAYER met4 ;
        RECT 8.730000 18.230000 9.050000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730000 18.660000 9.050000 18.980000 ;
      LAYER met4 ;
        RECT 8.730000 18.660000 9.050000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730000 19.090000 9.050000 19.410000 ;
      LAYER met4 ;
        RECT 8.730000 19.090000 9.050000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730000 19.520000 9.050000 19.840000 ;
      LAYER met4 ;
        RECT 8.730000 19.520000 9.050000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730000 19.950000 9.050000 20.270000 ;
      LAYER met4 ;
        RECT 8.730000 19.950000 9.050000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730000 20.380000 9.050000 20.700000 ;
      LAYER met4 ;
        RECT 8.730000 20.380000 9.050000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730000 20.810000 9.050000 21.130000 ;
      LAYER met4 ;
        RECT 8.730000 20.810000 9.050000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730000 21.240000 9.050000 21.560000 ;
      LAYER met4 ;
        RECT 8.730000 21.240000 9.050000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730000 21.670000 9.050000 21.990000 ;
      LAYER met4 ;
        RECT 8.730000 21.670000 9.050000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730000 22.100000 9.050000 22.420000 ;
      LAYER met4 ;
        RECT 8.730000 22.100000 9.050000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 68.065000 9.105000 68.385000 ;
      LAYER met4 ;
        RECT 8.785000 68.065000 9.105000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 68.475000 9.105000 68.795000 ;
      LAYER met4 ;
        RECT 8.785000 68.475000 9.105000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 68.885000 9.105000 69.205000 ;
      LAYER met4 ;
        RECT 8.785000 68.885000 9.105000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 69.295000 9.105000 69.615000 ;
      LAYER met4 ;
        RECT 8.785000 69.295000 9.105000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 69.705000 9.105000 70.025000 ;
      LAYER met4 ;
        RECT 8.785000 69.705000 9.105000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 70.115000 9.105000 70.435000 ;
      LAYER met4 ;
        RECT 8.785000 70.115000 9.105000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 70.525000 9.105000 70.845000 ;
      LAYER met4 ;
        RECT 8.785000 70.525000 9.105000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 70.935000 9.105000 71.255000 ;
      LAYER met4 ;
        RECT 8.785000 70.935000 9.105000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 71.345000 9.105000 71.665000 ;
      LAYER met4 ;
        RECT 8.785000 71.345000 9.105000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 71.755000 9.105000 72.075000 ;
      LAYER met4 ;
        RECT 8.785000 71.755000 9.105000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 72.165000 9.105000 72.485000 ;
      LAYER met4 ;
        RECT 8.785000 72.165000 9.105000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 72.575000 9.105000 72.895000 ;
      LAYER met4 ;
        RECT 8.785000 72.575000 9.105000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 72.985000 9.105000 73.305000 ;
      LAYER met4 ;
        RECT 8.785000 72.985000 9.105000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 73.390000 9.105000 73.710000 ;
      LAYER met4 ;
        RECT 8.785000 73.390000 9.105000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 73.795000 9.105000 74.115000 ;
      LAYER met4 ;
        RECT 8.785000 73.795000 9.105000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 74.200000 9.105000 74.520000 ;
      LAYER met4 ;
        RECT 8.785000 74.200000 9.105000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 74.605000 9.105000 74.925000 ;
      LAYER met4 ;
        RECT 8.785000 74.605000 9.105000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 75.010000 9.105000 75.330000 ;
      LAYER met4 ;
        RECT 8.785000 75.010000 9.105000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 75.415000 9.105000 75.735000 ;
      LAYER met4 ;
        RECT 8.785000 75.415000 9.105000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 75.820000 9.105000 76.140000 ;
      LAYER met4 ;
        RECT 8.785000 75.820000 9.105000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 76.225000 9.105000 76.545000 ;
      LAYER met4 ;
        RECT 8.785000 76.225000 9.105000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 76.630000 9.105000 76.950000 ;
      LAYER met4 ;
        RECT 8.785000 76.630000 9.105000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 77.035000 9.105000 77.355000 ;
      LAYER met4 ;
        RECT 8.785000 77.035000 9.105000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 77.440000 9.105000 77.760000 ;
      LAYER met4 ;
        RECT 8.785000 77.440000 9.105000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 77.845000 9.105000 78.165000 ;
      LAYER met4 ;
        RECT 8.785000 77.845000 9.105000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 78.250000 9.105000 78.570000 ;
      LAYER met4 ;
        RECT 8.785000 78.250000 9.105000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 78.655000 9.105000 78.975000 ;
      LAYER met4 ;
        RECT 8.785000 78.655000 9.105000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 79.060000 9.105000 79.380000 ;
      LAYER met4 ;
        RECT 8.785000 79.060000 9.105000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 79.465000 9.105000 79.785000 ;
      LAYER met4 ;
        RECT 8.785000 79.465000 9.105000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 79.870000 9.105000 80.190000 ;
      LAYER met4 ;
        RECT 8.785000 79.870000 9.105000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 80.275000 9.105000 80.595000 ;
      LAYER met4 ;
        RECT 8.785000 80.275000 9.105000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 80.680000 9.105000 81.000000 ;
      LAYER met4 ;
        RECT 8.785000 80.680000 9.105000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 81.085000 9.105000 81.405000 ;
      LAYER met4 ;
        RECT 8.785000 81.085000 9.105000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 81.490000 9.105000 81.810000 ;
      LAYER met4 ;
        RECT 8.785000 81.490000 9.105000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 81.895000 9.105000 82.215000 ;
      LAYER met4 ;
        RECT 8.785000 81.895000 9.105000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785000 82.300000 9.105000 82.620000 ;
      LAYER met4 ;
        RECT 8.785000 82.300000 9.105000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 82.795000 9.195000 83.115000 ;
      LAYER met4 ;
        RECT 8.875000 82.795000 9.195000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 83.205000 9.195000 83.525000 ;
      LAYER met4 ;
        RECT 8.875000 83.205000 9.195000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 83.615000 9.195000 83.935000 ;
      LAYER met4 ;
        RECT 8.875000 83.615000 9.195000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 84.025000 9.195000 84.345000 ;
      LAYER met4 ;
        RECT 8.875000 84.025000 9.195000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 84.435000 9.195000 84.755000 ;
      LAYER met4 ;
        RECT 8.875000 84.435000 9.195000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 84.845000 9.195000 85.165000 ;
      LAYER met4 ;
        RECT 8.875000 84.845000 9.195000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 85.255000 9.195000 85.575000 ;
      LAYER met4 ;
        RECT 8.875000 85.255000 9.195000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 85.665000 9.195000 85.985000 ;
      LAYER met4 ;
        RECT 8.875000 85.665000 9.195000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 86.075000 9.195000 86.395000 ;
      LAYER met4 ;
        RECT 8.875000 86.075000 9.195000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 86.485000 9.195000 86.805000 ;
      LAYER met4 ;
        RECT 8.875000 86.485000 9.195000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 86.895000 9.195000 87.215000 ;
      LAYER met4 ;
        RECT 8.875000 86.895000 9.195000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 87.305000 9.195000 87.625000 ;
      LAYER met4 ;
        RECT 8.875000 87.305000 9.195000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 87.715000 9.195000 88.035000 ;
      LAYER met4 ;
        RECT 8.875000 87.715000 9.195000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 88.125000 9.195000 88.445000 ;
      LAYER met4 ;
        RECT 8.875000 88.125000 9.195000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 88.535000 9.195000 88.855000 ;
      LAYER met4 ;
        RECT 8.875000 88.535000 9.195000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 88.945000 9.195000 89.265000 ;
      LAYER met4 ;
        RECT 8.875000 88.945000 9.195000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 89.355000 9.195000 89.675000 ;
      LAYER met4 ;
        RECT 8.875000 89.355000 9.195000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 89.765000 9.195000 90.085000 ;
      LAYER met4 ;
        RECT 8.875000 89.765000 9.195000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 90.175000 9.195000 90.495000 ;
      LAYER met4 ;
        RECT 8.875000 90.175000 9.195000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 90.585000 9.195000 90.905000 ;
      LAYER met4 ;
        RECT 8.875000 90.585000 9.195000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 90.995000 9.195000 91.315000 ;
      LAYER met4 ;
        RECT 8.875000 90.995000 9.195000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 91.405000 9.195000 91.725000 ;
      LAYER met4 ;
        RECT 8.875000 91.405000 9.195000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 91.815000 9.195000 92.135000 ;
      LAYER met4 ;
        RECT 8.875000 91.815000 9.195000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 92.225000 9.195000 92.545000 ;
      LAYER met4 ;
        RECT 8.875000 92.225000 9.195000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875000 92.635000 9.195000 92.955000 ;
      LAYER met4 ;
        RECT 8.875000 92.635000 9.195000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135000 17.800000 9.455000 18.120000 ;
      LAYER met4 ;
        RECT 9.135000 17.800000 9.455000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135000 18.230000 9.455000 18.550000 ;
      LAYER met4 ;
        RECT 9.135000 18.230000 9.455000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135000 18.660000 9.455000 18.980000 ;
      LAYER met4 ;
        RECT 9.135000 18.660000 9.455000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135000 19.090000 9.455000 19.410000 ;
      LAYER met4 ;
        RECT 9.135000 19.090000 9.455000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135000 19.520000 9.455000 19.840000 ;
      LAYER met4 ;
        RECT 9.135000 19.520000 9.455000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135000 19.950000 9.455000 20.270000 ;
      LAYER met4 ;
        RECT 9.135000 19.950000 9.455000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135000 20.380000 9.455000 20.700000 ;
      LAYER met4 ;
        RECT 9.135000 20.380000 9.455000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135000 20.810000 9.455000 21.130000 ;
      LAYER met4 ;
        RECT 9.135000 20.810000 9.455000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135000 21.240000 9.455000 21.560000 ;
      LAYER met4 ;
        RECT 9.135000 21.240000 9.455000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135000 21.670000 9.455000 21.990000 ;
      LAYER met4 ;
        RECT 9.135000 21.670000 9.455000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135000 22.100000 9.455000 22.420000 ;
      LAYER met4 ;
        RECT 9.135000 22.100000 9.455000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 68.065000 9.505000 68.385000 ;
      LAYER met4 ;
        RECT 9.185000 68.065000 9.505000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 68.475000 9.505000 68.795000 ;
      LAYER met4 ;
        RECT 9.185000 68.475000 9.505000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 68.885000 9.505000 69.205000 ;
      LAYER met4 ;
        RECT 9.185000 68.885000 9.505000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 69.295000 9.505000 69.615000 ;
      LAYER met4 ;
        RECT 9.185000 69.295000 9.505000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 69.705000 9.505000 70.025000 ;
      LAYER met4 ;
        RECT 9.185000 69.705000 9.505000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 70.115000 9.505000 70.435000 ;
      LAYER met4 ;
        RECT 9.185000 70.115000 9.505000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 70.525000 9.505000 70.845000 ;
      LAYER met4 ;
        RECT 9.185000 70.525000 9.505000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 70.935000 9.505000 71.255000 ;
      LAYER met4 ;
        RECT 9.185000 70.935000 9.505000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 71.345000 9.505000 71.665000 ;
      LAYER met4 ;
        RECT 9.185000 71.345000 9.505000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 71.755000 9.505000 72.075000 ;
      LAYER met4 ;
        RECT 9.185000 71.755000 9.505000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 72.165000 9.505000 72.485000 ;
      LAYER met4 ;
        RECT 9.185000 72.165000 9.505000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 72.575000 9.505000 72.895000 ;
      LAYER met4 ;
        RECT 9.185000 72.575000 9.505000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 72.985000 9.505000 73.305000 ;
      LAYER met4 ;
        RECT 9.185000 72.985000 9.505000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 73.390000 9.505000 73.710000 ;
      LAYER met4 ;
        RECT 9.185000 73.390000 9.505000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 73.795000 9.505000 74.115000 ;
      LAYER met4 ;
        RECT 9.185000 73.795000 9.505000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 74.200000 9.505000 74.520000 ;
      LAYER met4 ;
        RECT 9.185000 74.200000 9.505000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 74.605000 9.505000 74.925000 ;
      LAYER met4 ;
        RECT 9.185000 74.605000 9.505000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 75.010000 9.505000 75.330000 ;
      LAYER met4 ;
        RECT 9.185000 75.010000 9.505000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 75.415000 9.505000 75.735000 ;
      LAYER met4 ;
        RECT 9.185000 75.415000 9.505000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 75.820000 9.505000 76.140000 ;
      LAYER met4 ;
        RECT 9.185000 75.820000 9.505000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 76.225000 9.505000 76.545000 ;
      LAYER met4 ;
        RECT 9.185000 76.225000 9.505000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 76.630000 9.505000 76.950000 ;
      LAYER met4 ;
        RECT 9.185000 76.630000 9.505000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 77.035000 9.505000 77.355000 ;
      LAYER met4 ;
        RECT 9.185000 77.035000 9.505000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 77.440000 9.505000 77.760000 ;
      LAYER met4 ;
        RECT 9.185000 77.440000 9.505000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 77.845000 9.505000 78.165000 ;
      LAYER met4 ;
        RECT 9.185000 77.845000 9.505000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 78.250000 9.505000 78.570000 ;
      LAYER met4 ;
        RECT 9.185000 78.250000 9.505000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 78.655000 9.505000 78.975000 ;
      LAYER met4 ;
        RECT 9.185000 78.655000 9.505000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 79.060000 9.505000 79.380000 ;
      LAYER met4 ;
        RECT 9.185000 79.060000 9.505000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 79.465000 9.505000 79.785000 ;
      LAYER met4 ;
        RECT 9.185000 79.465000 9.505000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 79.870000 9.505000 80.190000 ;
      LAYER met4 ;
        RECT 9.185000 79.870000 9.505000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 80.275000 9.505000 80.595000 ;
      LAYER met4 ;
        RECT 9.185000 80.275000 9.505000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 80.680000 9.505000 81.000000 ;
      LAYER met4 ;
        RECT 9.185000 80.680000 9.505000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 81.085000 9.505000 81.405000 ;
      LAYER met4 ;
        RECT 9.185000 81.085000 9.505000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 81.490000 9.505000 81.810000 ;
      LAYER met4 ;
        RECT 9.185000 81.490000 9.505000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 81.895000 9.505000 82.215000 ;
      LAYER met4 ;
        RECT 9.185000 81.895000 9.505000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185000 82.300000 9.505000 82.620000 ;
      LAYER met4 ;
        RECT 9.185000 82.300000 9.505000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 82.795000 9.605000 83.115000 ;
      LAYER met4 ;
        RECT 9.285000 82.795000 9.605000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 83.205000 9.605000 83.525000 ;
      LAYER met4 ;
        RECT 9.285000 83.205000 9.605000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 83.615000 9.605000 83.935000 ;
      LAYER met4 ;
        RECT 9.285000 83.615000 9.605000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 84.025000 9.605000 84.345000 ;
      LAYER met4 ;
        RECT 9.285000 84.025000 9.605000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 84.435000 9.605000 84.755000 ;
      LAYER met4 ;
        RECT 9.285000 84.435000 9.605000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 84.845000 9.605000 85.165000 ;
      LAYER met4 ;
        RECT 9.285000 84.845000 9.605000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 85.255000 9.605000 85.575000 ;
      LAYER met4 ;
        RECT 9.285000 85.255000 9.605000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 85.665000 9.605000 85.985000 ;
      LAYER met4 ;
        RECT 9.285000 85.665000 9.605000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 86.075000 9.605000 86.395000 ;
      LAYER met4 ;
        RECT 9.285000 86.075000 9.605000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 86.485000 9.605000 86.805000 ;
      LAYER met4 ;
        RECT 9.285000 86.485000 9.605000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 86.895000 9.605000 87.215000 ;
      LAYER met4 ;
        RECT 9.285000 86.895000 9.605000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 87.305000 9.605000 87.625000 ;
      LAYER met4 ;
        RECT 9.285000 87.305000 9.605000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 87.715000 9.605000 88.035000 ;
      LAYER met4 ;
        RECT 9.285000 87.715000 9.605000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 88.125000 9.605000 88.445000 ;
      LAYER met4 ;
        RECT 9.285000 88.125000 9.605000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 88.535000 9.605000 88.855000 ;
      LAYER met4 ;
        RECT 9.285000 88.535000 9.605000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 88.945000 9.605000 89.265000 ;
      LAYER met4 ;
        RECT 9.285000 88.945000 9.605000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 89.355000 9.605000 89.675000 ;
      LAYER met4 ;
        RECT 9.285000 89.355000 9.605000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 89.765000 9.605000 90.085000 ;
      LAYER met4 ;
        RECT 9.285000 89.765000 9.605000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 90.175000 9.605000 90.495000 ;
      LAYER met4 ;
        RECT 9.285000 90.175000 9.605000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 90.585000 9.605000 90.905000 ;
      LAYER met4 ;
        RECT 9.285000 90.585000 9.605000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 90.995000 9.605000 91.315000 ;
      LAYER met4 ;
        RECT 9.285000 90.995000 9.605000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 91.405000 9.605000 91.725000 ;
      LAYER met4 ;
        RECT 9.285000 91.405000 9.605000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 91.815000 9.605000 92.135000 ;
      LAYER met4 ;
        RECT 9.285000 91.815000 9.605000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 92.225000 9.605000 92.545000 ;
      LAYER met4 ;
        RECT 9.285000 92.225000 9.605000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285000 92.635000 9.605000 92.955000 ;
      LAYER met4 ;
        RECT 9.285000 92.635000 9.605000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540000 17.800000 9.860000 18.120000 ;
      LAYER met4 ;
        RECT 9.540000 17.800000 9.860000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540000 18.230000 9.860000 18.550000 ;
      LAYER met4 ;
        RECT 9.540000 18.230000 9.860000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540000 18.660000 9.860000 18.980000 ;
      LAYER met4 ;
        RECT 9.540000 18.660000 9.860000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540000 19.090000 9.860000 19.410000 ;
      LAYER met4 ;
        RECT 9.540000 19.090000 9.860000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540000 19.520000 9.860000 19.840000 ;
      LAYER met4 ;
        RECT 9.540000 19.520000 9.860000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540000 19.950000 9.860000 20.270000 ;
      LAYER met4 ;
        RECT 9.540000 19.950000 9.860000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540000 20.380000 9.860000 20.700000 ;
      LAYER met4 ;
        RECT 9.540000 20.380000 9.860000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540000 20.810000 9.860000 21.130000 ;
      LAYER met4 ;
        RECT 9.540000 20.810000 9.860000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540000 21.240000 9.860000 21.560000 ;
      LAYER met4 ;
        RECT 9.540000 21.240000 9.860000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540000 21.670000 9.860000 21.990000 ;
      LAYER met4 ;
        RECT 9.540000 21.670000 9.860000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540000 22.100000 9.860000 22.420000 ;
      LAYER met4 ;
        RECT 9.540000 22.100000 9.860000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 68.065000 9.905000 68.385000 ;
      LAYER met4 ;
        RECT 9.585000 68.065000 9.905000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 68.475000 9.905000 68.795000 ;
      LAYER met4 ;
        RECT 9.585000 68.475000 9.905000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 68.885000 9.905000 69.205000 ;
      LAYER met4 ;
        RECT 9.585000 68.885000 9.905000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 69.295000 9.905000 69.615000 ;
      LAYER met4 ;
        RECT 9.585000 69.295000 9.905000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 69.705000 9.905000 70.025000 ;
      LAYER met4 ;
        RECT 9.585000 69.705000 9.905000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 70.115000 9.905000 70.435000 ;
      LAYER met4 ;
        RECT 9.585000 70.115000 9.905000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 70.525000 9.905000 70.845000 ;
      LAYER met4 ;
        RECT 9.585000 70.525000 9.905000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 70.935000 9.905000 71.255000 ;
      LAYER met4 ;
        RECT 9.585000 70.935000 9.905000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 71.345000 9.905000 71.665000 ;
      LAYER met4 ;
        RECT 9.585000 71.345000 9.905000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 71.755000 9.905000 72.075000 ;
      LAYER met4 ;
        RECT 9.585000 71.755000 9.905000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 72.165000 9.905000 72.485000 ;
      LAYER met4 ;
        RECT 9.585000 72.165000 9.905000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 72.575000 9.905000 72.895000 ;
      LAYER met4 ;
        RECT 9.585000 72.575000 9.905000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 72.985000 9.905000 73.305000 ;
      LAYER met4 ;
        RECT 9.585000 72.985000 9.905000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 73.390000 9.905000 73.710000 ;
      LAYER met4 ;
        RECT 9.585000 73.390000 9.905000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 73.795000 9.905000 74.115000 ;
      LAYER met4 ;
        RECT 9.585000 73.795000 9.905000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 74.200000 9.905000 74.520000 ;
      LAYER met4 ;
        RECT 9.585000 74.200000 9.905000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 74.605000 9.905000 74.925000 ;
      LAYER met4 ;
        RECT 9.585000 74.605000 9.905000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 75.010000 9.905000 75.330000 ;
      LAYER met4 ;
        RECT 9.585000 75.010000 9.905000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 75.415000 9.905000 75.735000 ;
      LAYER met4 ;
        RECT 9.585000 75.415000 9.905000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 75.820000 9.905000 76.140000 ;
      LAYER met4 ;
        RECT 9.585000 75.820000 9.905000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 76.225000 9.905000 76.545000 ;
      LAYER met4 ;
        RECT 9.585000 76.225000 9.905000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 76.630000 9.905000 76.950000 ;
      LAYER met4 ;
        RECT 9.585000 76.630000 9.905000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 77.035000 9.905000 77.355000 ;
      LAYER met4 ;
        RECT 9.585000 77.035000 9.905000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 77.440000 9.905000 77.760000 ;
      LAYER met4 ;
        RECT 9.585000 77.440000 9.905000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 77.845000 9.905000 78.165000 ;
      LAYER met4 ;
        RECT 9.585000 77.845000 9.905000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 78.250000 9.905000 78.570000 ;
      LAYER met4 ;
        RECT 9.585000 78.250000 9.905000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 78.655000 9.905000 78.975000 ;
      LAYER met4 ;
        RECT 9.585000 78.655000 9.905000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 79.060000 9.905000 79.380000 ;
      LAYER met4 ;
        RECT 9.585000 79.060000 9.905000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 79.465000 9.905000 79.785000 ;
      LAYER met4 ;
        RECT 9.585000 79.465000 9.905000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 79.870000 9.905000 80.190000 ;
      LAYER met4 ;
        RECT 9.585000 79.870000 9.905000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 80.275000 9.905000 80.595000 ;
      LAYER met4 ;
        RECT 9.585000 80.275000 9.905000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 80.680000 9.905000 81.000000 ;
      LAYER met4 ;
        RECT 9.585000 80.680000 9.905000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 81.085000 9.905000 81.405000 ;
      LAYER met4 ;
        RECT 9.585000 81.085000 9.905000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 81.490000 9.905000 81.810000 ;
      LAYER met4 ;
        RECT 9.585000 81.490000 9.905000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 81.895000 9.905000 82.215000 ;
      LAYER met4 ;
        RECT 9.585000 81.895000 9.905000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585000 82.300000 9.905000 82.620000 ;
      LAYER met4 ;
        RECT 9.585000 82.300000 9.905000 82.620000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 82.795000 10.015000 83.115000 ;
      LAYER met4 ;
        RECT 9.695000 82.795000 10.015000 83.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 83.205000 10.015000 83.525000 ;
      LAYER met4 ;
        RECT 9.695000 83.205000 10.015000 83.525000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 83.615000 10.015000 83.935000 ;
      LAYER met4 ;
        RECT 9.695000 83.615000 10.015000 83.935000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 84.025000 10.015000 84.345000 ;
      LAYER met4 ;
        RECT 9.695000 84.025000 10.015000 84.345000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 84.435000 10.015000 84.755000 ;
      LAYER met4 ;
        RECT 9.695000 84.435000 10.015000 84.755000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 84.845000 10.015000 85.165000 ;
      LAYER met4 ;
        RECT 9.695000 84.845000 10.015000 85.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 85.255000 10.015000 85.575000 ;
      LAYER met4 ;
        RECT 9.695000 85.255000 10.015000 85.575000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 85.665000 10.015000 85.985000 ;
      LAYER met4 ;
        RECT 9.695000 85.665000 10.015000 85.985000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 86.075000 10.015000 86.395000 ;
      LAYER met4 ;
        RECT 9.695000 86.075000 10.015000 86.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 86.485000 10.015000 86.805000 ;
      LAYER met4 ;
        RECT 9.695000 86.485000 10.015000 86.805000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 86.895000 10.015000 87.215000 ;
      LAYER met4 ;
        RECT 9.695000 86.895000 10.015000 87.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 87.305000 10.015000 87.625000 ;
      LAYER met4 ;
        RECT 9.695000 87.305000 10.015000 87.625000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 87.715000 10.015000 88.035000 ;
      LAYER met4 ;
        RECT 9.695000 87.715000 10.015000 88.035000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 88.125000 10.015000 88.445000 ;
      LAYER met4 ;
        RECT 9.695000 88.125000 10.015000 88.445000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 88.535000 10.015000 88.855000 ;
      LAYER met4 ;
        RECT 9.695000 88.535000 10.015000 88.855000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 88.945000 10.015000 89.265000 ;
      LAYER met4 ;
        RECT 9.695000 88.945000 10.015000 89.265000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 89.355000 10.015000 89.675000 ;
      LAYER met4 ;
        RECT 9.695000 89.355000 10.015000 89.675000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 89.765000 10.015000 90.085000 ;
      LAYER met4 ;
        RECT 9.695000 89.765000 10.015000 90.085000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 90.175000 10.015000 90.495000 ;
      LAYER met4 ;
        RECT 9.695000 90.175000 10.015000 90.495000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 90.585000 10.015000 90.905000 ;
      LAYER met4 ;
        RECT 9.695000 90.585000 10.015000 90.905000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 90.995000 10.015000 91.315000 ;
      LAYER met4 ;
        RECT 9.695000 90.995000 10.015000 91.315000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 91.405000 10.015000 91.725000 ;
      LAYER met4 ;
        RECT 9.695000 91.405000 10.015000 91.725000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 91.815000 10.015000 92.135000 ;
      LAYER met4 ;
        RECT 9.695000 91.815000 10.015000 92.135000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 92.225000 10.015000 92.545000 ;
      LAYER met4 ;
        RECT 9.695000 92.225000 10.015000 92.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695000 92.635000 10.015000 92.955000 ;
      LAYER met4 ;
        RECT 9.695000 92.635000 10.015000 92.955000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945000 17.800000 10.265000 18.120000 ;
      LAYER met4 ;
        RECT 9.945000 17.800000 10.265000 18.120000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945000 18.230000 10.265000 18.550000 ;
      LAYER met4 ;
        RECT 9.945000 18.230000 10.265000 18.550000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945000 18.660000 10.265000 18.980000 ;
      LAYER met4 ;
        RECT 9.945000 18.660000 10.265000 18.980000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945000 19.090000 10.265000 19.410000 ;
      LAYER met4 ;
        RECT 9.945000 19.090000 10.265000 19.410000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945000 19.520000 10.265000 19.840000 ;
      LAYER met4 ;
        RECT 9.945000 19.520000 10.265000 19.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945000 19.950000 10.265000 20.270000 ;
      LAYER met4 ;
        RECT 9.945000 19.950000 10.265000 20.270000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945000 20.380000 10.265000 20.700000 ;
      LAYER met4 ;
        RECT 9.945000 20.380000 10.265000 20.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945000 20.810000 10.265000 21.130000 ;
      LAYER met4 ;
        RECT 9.945000 20.810000 10.265000 21.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945000 21.240000 10.265000 21.560000 ;
      LAYER met4 ;
        RECT 9.945000 21.240000 10.265000 21.560000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945000 21.670000 10.265000 21.990000 ;
      LAYER met4 ;
        RECT 9.945000 21.670000 10.265000 21.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945000 22.100000 10.265000 22.420000 ;
      LAYER met4 ;
        RECT 9.945000 22.100000 10.265000 22.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 68.065000 10.305000 68.385000 ;
      LAYER met4 ;
        RECT 9.985000 68.065000 10.305000 68.385000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 68.475000 10.305000 68.795000 ;
      LAYER met4 ;
        RECT 9.985000 68.475000 10.305000 68.795000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 68.885000 10.305000 69.205000 ;
      LAYER met4 ;
        RECT 9.985000 68.885000 10.305000 69.205000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 69.295000 10.305000 69.615000 ;
      LAYER met4 ;
        RECT 9.985000 69.295000 10.305000 69.615000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 69.705000 10.305000 70.025000 ;
      LAYER met4 ;
        RECT 9.985000 69.705000 10.305000 70.025000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 70.115000 10.305000 70.435000 ;
      LAYER met4 ;
        RECT 9.985000 70.115000 10.305000 70.435000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 70.525000 10.305000 70.845000 ;
      LAYER met4 ;
        RECT 9.985000 70.525000 10.305000 70.845000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 70.935000 10.305000 71.255000 ;
      LAYER met4 ;
        RECT 9.985000 70.935000 10.305000 71.255000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 71.345000 10.305000 71.665000 ;
      LAYER met4 ;
        RECT 9.985000 71.345000 10.305000 71.665000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 71.755000 10.305000 72.075000 ;
      LAYER met4 ;
        RECT 9.985000 71.755000 10.305000 72.075000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 72.165000 10.305000 72.485000 ;
      LAYER met4 ;
        RECT 9.985000 72.165000 10.305000 72.485000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 72.575000 10.305000 72.895000 ;
      LAYER met4 ;
        RECT 9.985000 72.575000 10.305000 72.895000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 72.985000 10.305000 73.305000 ;
      LAYER met4 ;
        RECT 9.985000 72.985000 10.305000 73.305000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 73.390000 10.305000 73.710000 ;
      LAYER met4 ;
        RECT 9.985000 73.390000 10.305000 73.710000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 73.795000 10.305000 74.115000 ;
      LAYER met4 ;
        RECT 9.985000 73.795000 10.305000 74.115000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 74.200000 10.305000 74.520000 ;
      LAYER met4 ;
        RECT 9.985000 74.200000 10.305000 74.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 74.605000 10.305000 74.925000 ;
      LAYER met4 ;
        RECT 9.985000 74.605000 10.305000 74.925000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 75.010000 10.305000 75.330000 ;
      LAYER met4 ;
        RECT 9.985000 75.010000 10.305000 75.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 75.415000 10.305000 75.735000 ;
      LAYER met4 ;
        RECT 9.985000 75.415000 10.305000 75.735000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 75.820000 10.305000 76.140000 ;
      LAYER met4 ;
        RECT 9.985000 75.820000 10.305000 76.140000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 76.225000 10.305000 76.545000 ;
      LAYER met4 ;
        RECT 9.985000 76.225000 10.305000 76.545000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 76.630000 10.305000 76.950000 ;
      LAYER met4 ;
        RECT 9.985000 76.630000 10.305000 76.950000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 77.035000 10.305000 77.355000 ;
      LAYER met4 ;
        RECT 9.985000 77.035000 10.305000 77.355000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 77.440000 10.305000 77.760000 ;
      LAYER met4 ;
        RECT 9.985000 77.440000 10.305000 77.760000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 77.845000 10.305000 78.165000 ;
      LAYER met4 ;
        RECT 9.985000 77.845000 10.305000 78.165000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 78.250000 10.305000 78.570000 ;
      LAYER met4 ;
        RECT 9.985000 78.250000 10.305000 78.570000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 78.655000 10.305000 78.975000 ;
      LAYER met4 ;
        RECT 9.985000 78.655000 10.305000 78.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 79.060000 10.305000 79.380000 ;
      LAYER met4 ;
        RECT 9.985000 79.060000 10.305000 79.380000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 79.465000 10.305000 79.785000 ;
      LAYER met4 ;
        RECT 9.985000 79.465000 10.305000 79.785000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 79.870000 10.305000 80.190000 ;
      LAYER met4 ;
        RECT 9.985000 79.870000 10.305000 80.190000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 80.275000 10.305000 80.595000 ;
      LAYER met4 ;
        RECT 9.985000 80.275000 10.305000 80.595000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 80.680000 10.305000 81.000000 ;
      LAYER met4 ;
        RECT 9.985000 80.680000 10.305000 81.000000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 81.085000 10.305000 81.405000 ;
      LAYER met4 ;
        RECT 9.985000 81.085000 10.305000 81.405000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 81.490000 10.305000 81.810000 ;
      LAYER met4 ;
        RECT 9.985000 81.490000 10.305000 81.810000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 81.895000 10.305000 82.215000 ;
      LAYER met4 ;
        RECT 9.985000 81.895000 10.305000 82.215000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985000 82.300000 10.305000 82.620000 ;
      LAYER met4 ;
        RECT 9.985000 82.300000 10.305000 82.620000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.630000 62.100000 0.950000 62.420000 ;
      LAYER met4 ;
        RECT 0.630000 62.100000 0.950000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 62.510000 0.950000 62.830000 ;
      LAYER met4 ;
        RECT 0.630000 62.510000 0.950000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 62.920000 0.950000 63.240000 ;
      LAYER met4 ;
        RECT 0.630000 62.920000 0.950000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 63.330000 0.950000 63.650000 ;
      LAYER met4 ;
        RECT 0.630000 63.330000 0.950000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 63.740000 0.950000 64.060000 ;
      LAYER met4 ;
        RECT 0.630000 63.740000 0.950000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 64.150000 0.950000 64.470000 ;
      LAYER met4 ;
        RECT 0.630000 64.150000 0.950000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 64.560000 0.950000 64.880000 ;
      LAYER met4 ;
        RECT 0.630000 64.560000 0.950000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 64.970000 0.950000 65.290000 ;
      LAYER met4 ;
        RECT 0.630000 64.970000 0.950000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 65.380000 0.950000 65.700000 ;
      LAYER met4 ;
        RECT 0.630000 65.380000 0.950000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 65.790000 0.950000 66.110000 ;
      LAYER met4 ;
        RECT 0.630000 65.790000 0.950000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 66.200000 0.950000 66.520000 ;
      LAYER met4 ;
        RECT 0.630000 66.200000 0.950000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035000 62.100000 1.355000 62.420000 ;
      LAYER met4 ;
        RECT 1.035000 62.100000 1.355000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035000 62.510000 1.355000 62.830000 ;
      LAYER met4 ;
        RECT 1.035000 62.510000 1.355000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035000 62.920000 1.355000 63.240000 ;
      LAYER met4 ;
        RECT 1.035000 62.920000 1.355000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035000 63.330000 1.355000 63.650000 ;
      LAYER met4 ;
        RECT 1.035000 63.330000 1.355000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035000 63.740000 1.355000 64.060000 ;
      LAYER met4 ;
        RECT 1.035000 63.740000 1.355000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035000 64.150000 1.355000 64.470000 ;
      LAYER met4 ;
        RECT 1.035000 64.150000 1.355000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035000 64.560000 1.355000 64.880000 ;
      LAYER met4 ;
        RECT 1.035000 64.560000 1.355000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035000 64.970000 1.355000 65.290000 ;
      LAYER met4 ;
        RECT 1.035000 64.970000 1.355000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035000 65.380000 1.355000 65.700000 ;
      LAYER met4 ;
        RECT 1.035000 65.380000 1.355000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035000 65.790000 1.355000 66.110000 ;
      LAYER met4 ;
        RECT 1.035000 65.790000 1.355000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035000 66.200000 1.355000 66.520000 ;
      LAYER met4 ;
        RECT 1.035000 66.200000 1.355000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440000 62.100000 1.760000 62.420000 ;
      LAYER met4 ;
        RECT 1.440000 62.100000 1.760000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440000 62.510000 1.760000 62.830000 ;
      LAYER met4 ;
        RECT 1.440000 62.510000 1.760000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440000 62.920000 1.760000 63.240000 ;
      LAYER met4 ;
        RECT 1.440000 62.920000 1.760000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440000 63.330000 1.760000 63.650000 ;
      LAYER met4 ;
        RECT 1.440000 63.330000 1.760000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440000 63.740000 1.760000 64.060000 ;
      LAYER met4 ;
        RECT 1.440000 63.740000 1.760000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440000 64.150000 1.760000 64.470000 ;
      LAYER met4 ;
        RECT 1.440000 64.150000 1.760000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440000 64.560000 1.760000 64.880000 ;
      LAYER met4 ;
        RECT 1.440000 64.560000 1.760000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440000 64.970000 1.760000 65.290000 ;
      LAYER met4 ;
        RECT 1.440000 64.970000 1.760000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440000 65.380000 1.760000 65.700000 ;
      LAYER met4 ;
        RECT 1.440000 65.380000 1.760000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440000 65.790000 1.760000 66.110000 ;
      LAYER met4 ;
        RECT 1.440000 65.790000 1.760000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440000 66.200000 1.760000 66.520000 ;
      LAYER met4 ;
        RECT 1.440000 66.200000 1.760000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845000 62.100000 2.165000 62.420000 ;
      LAYER met4 ;
        RECT 1.845000 62.100000 2.165000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845000 62.510000 2.165000 62.830000 ;
      LAYER met4 ;
        RECT 1.845000 62.510000 2.165000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845000 62.920000 2.165000 63.240000 ;
      LAYER met4 ;
        RECT 1.845000 62.920000 2.165000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845000 63.330000 2.165000 63.650000 ;
      LAYER met4 ;
        RECT 1.845000 63.330000 2.165000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845000 63.740000 2.165000 64.060000 ;
      LAYER met4 ;
        RECT 1.845000 63.740000 2.165000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845000 64.150000 2.165000 64.470000 ;
      LAYER met4 ;
        RECT 1.845000 64.150000 2.165000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845000 64.560000 2.165000 64.880000 ;
      LAYER met4 ;
        RECT 1.845000 64.560000 2.165000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845000 64.970000 2.165000 65.290000 ;
      LAYER met4 ;
        RECT 1.845000 64.970000 2.165000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845000 65.380000 2.165000 65.700000 ;
      LAYER met4 ;
        RECT 1.845000 65.380000 2.165000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845000 65.790000 2.165000 66.110000 ;
      LAYER met4 ;
        RECT 1.845000 65.790000 2.165000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845000 66.200000 2.165000 66.520000 ;
      LAYER met4 ;
        RECT 1.845000 66.200000 2.165000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350000 62.100000 10.670000 62.420000 ;
      LAYER met4 ;
        RECT 10.350000 62.100000 10.670000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350000 62.510000 10.670000 62.830000 ;
      LAYER met4 ;
        RECT 10.350000 62.510000 10.670000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350000 62.920000 10.670000 63.240000 ;
      LAYER met4 ;
        RECT 10.350000 62.920000 10.670000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350000 63.330000 10.670000 63.650000 ;
      LAYER met4 ;
        RECT 10.350000 63.330000 10.670000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350000 63.740000 10.670000 64.060000 ;
      LAYER met4 ;
        RECT 10.350000 63.740000 10.670000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350000 64.150000 10.670000 64.470000 ;
      LAYER met4 ;
        RECT 10.350000 64.150000 10.670000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350000 64.560000 10.670000 64.880000 ;
      LAYER met4 ;
        RECT 10.350000 64.560000 10.670000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350000 64.970000 10.670000 65.290000 ;
      LAYER met4 ;
        RECT 10.350000 64.970000 10.670000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350000 65.380000 10.670000 65.700000 ;
      LAYER met4 ;
        RECT 10.350000 65.380000 10.670000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350000 65.790000 10.670000 66.110000 ;
      LAYER met4 ;
        RECT 10.350000 65.790000 10.670000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350000 66.200000 10.670000 66.520000 ;
      LAYER met4 ;
        RECT 10.350000 66.200000 10.670000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755000 62.100000 11.075000 62.420000 ;
      LAYER met4 ;
        RECT 10.755000 62.100000 11.075000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755000 62.510000 11.075000 62.830000 ;
      LAYER met4 ;
        RECT 10.755000 62.510000 11.075000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755000 62.920000 11.075000 63.240000 ;
      LAYER met4 ;
        RECT 10.755000 62.920000 11.075000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755000 63.330000 11.075000 63.650000 ;
      LAYER met4 ;
        RECT 10.755000 63.330000 11.075000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755000 63.740000 11.075000 64.060000 ;
      LAYER met4 ;
        RECT 10.755000 63.740000 11.075000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755000 64.150000 11.075000 64.470000 ;
      LAYER met4 ;
        RECT 10.755000 64.150000 11.075000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755000 64.560000 11.075000 64.880000 ;
      LAYER met4 ;
        RECT 10.755000 64.560000 11.075000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755000 64.970000 11.075000 65.290000 ;
      LAYER met4 ;
        RECT 10.755000 64.970000 11.075000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755000 65.380000 11.075000 65.700000 ;
      LAYER met4 ;
        RECT 10.755000 65.380000 11.075000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755000 65.790000 11.075000 66.110000 ;
      LAYER met4 ;
        RECT 10.755000 65.790000 11.075000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755000 66.200000 11.075000 66.520000 ;
      LAYER met4 ;
        RECT 10.755000 66.200000 11.075000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160000 62.100000 11.480000 62.420000 ;
      LAYER met4 ;
        RECT 11.160000 62.100000 11.480000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160000 62.510000 11.480000 62.830000 ;
      LAYER met4 ;
        RECT 11.160000 62.510000 11.480000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160000 62.920000 11.480000 63.240000 ;
      LAYER met4 ;
        RECT 11.160000 62.920000 11.480000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160000 63.330000 11.480000 63.650000 ;
      LAYER met4 ;
        RECT 11.160000 63.330000 11.480000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160000 63.740000 11.480000 64.060000 ;
      LAYER met4 ;
        RECT 11.160000 63.740000 11.480000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160000 64.150000 11.480000 64.470000 ;
      LAYER met4 ;
        RECT 11.160000 64.150000 11.480000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160000 64.560000 11.480000 64.880000 ;
      LAYER met4 ;
        RECT 11.160000 64.560000 11.480000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160000 64.970000 11.480000 65.290000 ;
      LAYER met4 ;
        RECT 11.160000 64.970000 11.480000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160000 65.380000 11.480000 65.700000 ;
      LAYER met4 ;
        RECT 11.160000 65.380000 11.480000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160000 65.790000 11.480000 66.110000 ;
      LAYER met4 ;
        RECT 11.160000 65.790000 11.480000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160000 66.200000 11.480000 66.520000 ;
      LAYER met4 ;
        RECT 11.160000 66.200000 11.480000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565000 62.100000 11.885000 62.420000 ;
      LAYER met4 ;
        RECT 11.565000 62.100000 11.885000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565000 62.510000 11.885000 62.830000 ;
      LAYER met4 ;
        RECT 11.565000 62.510000 11.885000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565000 62.920000 11.885000 63.240000 ;
      LAYER met4 ;
        RECT 11.565000 62.920000 11.885000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565000 63.330000 11.885000 63.650000 ;
      LAYER met4 ;
        RECT 11.565000 63.330000 11.885000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565000 63.740000 11.885000 64.060000 ;
      LAYER met4 ;
        RECT 11.565000 63.740000 11.885000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565000 64.150000 11.885000 64.470000 ;
      LAYER met4 ;
        RECT 11.565000 64.150000 11.885000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565000 64.560000 11.885000 64.880000 ;
      LAYER met4 ;
        RECT 11.565000 64.560000 11.885000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565000 64.970000 11.885000 65.290000 ;
      LAYER met4 ;
        RECT 11.565000 64.970000 11.885000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565000 65.380000 11.885000 65.700000 ;
      LAYER met4 ;
        RECT 11.565000 65.380000 11.885000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565000 65.790000 11.885000 66.110000 ;
      LAYER met4 ;
        RECT 11.565000 65.790000 11.885000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565000 66.200000 11.885000 66.520000 ;
      LAYER met4 ;
        RECT 11.565000 66.200000 11.885000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970000 62.100000 12.290000 62.420000 ;
      LAYER met4 ;
        RECT 11.970000 62.100000 12.290000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970000 62.510000 12.290000 62.830000 ;
      LAYER met4 ;
        RECT 11.970000 62.510000 12.290000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970000 62.920000 12.290000 63.240000 ;
      LAYER met4 ;
        RECT 11.970000 62.920000 12.290000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970000 63.330000 12.290000 63.650000 ;
      LAYER met4 ;
        RECT 11.970000 63.330000 12.290000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970000 63.740000 12.290000 64.060000 ;
      LAYER met4 ;
        RECT 11.970000 63.740000 12.290000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970000 64.150000 12.290000 64.470000 ;
      LAYER met4 ;
        RECT 11.970000 64.150000 12.290000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970000 64.560000 12.290000 64.880000 ;
      LAYER met4 ;
        RECT 11.970000 64.560000 12.290000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970000 64.970000 12.290000 65.290000 ;
      LAYER met4 ;
        RECT 11.970000 64.970000 12.290000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970000 65.380000 12.290000 65.700000 ;
      LAYER met4 ;
        RECT 11.970000 65.380000 12.290000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970000 65.790000 12.290000 66.110000 ;
      LAYER met4 ;
        RECT 11.970000 65.790000 12.290000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970000 66.200000 12.290000 66.520000 ;
      LAYER met4 ;
        RECT 11.970000 66.200000 12.290000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375000 62.100000 12.695000 62.420000 ;
      LAYER met4 ;
        RECT 12.375000 62.100000 12.695000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375000 62.510000 12.695000 62.830000 ;
      LAYER met4 ;
        RECT 12.375000 62.510000 12.695000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375000 62.920000 12.695000 63.240000 ;
      LAYER met4 ;
        RECT 12.375000 62.920000 12.695000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375000 63.330000 12.695000 63.650000 ;
      LAYER met4 ;
        RECT 12.375000 63.330000 12.695000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375000 63.740000 12.695000 64.060000 ;
      LAYER met4 ;
        RECT 12.375000 63.740000 12.695000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375000 64.150000 12.695000 64.470000 ;
      LAYER met4 ;
        RECT 12.375000 64.150000 12.695000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375000 64.560000 12.695000 64.880000 ;
      LAYER met4 ;
        RECT 12.375000 64.560000 12.695000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375000 64.970000 12.695000 65.290000 ;
      LAYER met4 ;
        RECT 12.375000 64.970000 12.695000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375000 65.380000 12.695000 65.700000 ;
      LAYER met4 ;
        RECT 12.375000 65.380000 12.695000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375000 65.790000 12.695000 66.110000 ;
      LAYER met4 ;
        RECT 12.375000 65.790000 12.695000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375000 66.200000 12.695000 66.520000 ;
      LAYER met4 ;
        RECT 12.375000 66.200000 12.695000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 62.100000 13.100000 62.420000 ;
      LAYER met4 ;
        RECT 12.780000 62.100000 13.100000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 62.510000 13.100000 62.830000 ;
      LAYER met4 ;
        RECT 12.780000 62.510000 13.100000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 62.920000 13.100000 63.240000 ;
      LAYER met4 ;
        RECT 12.780000 62.920000 13.100000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 63.330000 13.100000 63.650000 ;
      LAYER met4 ;
        RECT 12.780000 63.330000 13.100000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 63.740000 13.100000 64.060000 ;
      LAYER met4 ;
        RECT 12.780000 63.740000 13.100000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 64.150000 13.100000 64.470000 ;
      LAYER met4 ;
        RECT 12.780000 64.150000 13.100000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 64.560000 13.100000 64.880000 ;
      LAYER met4 ;
        RECT 12.780000 64.560000 13.100000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 64.970000 13.100000 65.290000 ;
      LAYER met4 ;
        RECT 12.780000 64.970000 13.100000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 65.380000 13.100000 65.700000 ;
      LAYER met4 ;
        RECT 12.780000 65.380000 13.100000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 65.790000 13.100000 66.110000 ;
      LAYER met4 ;
        RECT 12.780000 65.790000 13.100000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780000 66.200000 13.100000 66.520000 ;
      LAYER met4 ;
        RECT 12.780000 66.200000 13.100000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 62.100000 13.505000 62.420000 ;
      LAYER met4 ;
        RECT 13.185000 62.100000 13.505000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 62.510000 13.505000 62.830000 ;
      LAYER met4 ;
        RECT 13.185000 62.510000 13.505000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 62.920000 13.505000 63.240000 ;
      LAYER met4 ;
        RECT 13.185000 62.920000 13.505000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 63.330000 13.505000 63.650000 ;
      LAYER met4 ;
        RECT 13.185000 63.330000 13.505000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 63.740000 13.505000 64.060000 ;
      LAYER met4 ;
        RECT 13.185000 63.740000 13.505000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 64.150000 13.505000 64.470000 ;
      LAYER met4 ;
        RECT 13.185000 64.150000 13.505000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 64.560000 13.505000 64.880000 ;
      LAYER met4 ;
        RECT 13.185000 64.560000 13.505000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 64.970000 13.505000 65.290000 ;
      LAYER met4 ;
        RECT 13.185000 64.970000 13.505000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 65.380000 13.505000 65.700000 ;
      LAYER met4 ;
        RECT 13.185000 65.380000 13.505000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 65.790000 13.505000 66.110000 ;
      LAYER met4 ;
        RECT 13.185000 65.790000 13.505000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185000 66.200000 13.505000 66.520000 ;
      LAYER met4 ;
        RECT 13.185000 66.200000 13.505000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590000 62.100000 13.910000 62.420000 ;
      LAYER met4 ;
        RECT 13.590000 62.100000 13.910000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590000 62.510000 13.910000 62.830000 ;
      LAYER met4 ;
        RECT 13.590000 62.510000 13.910000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590000 62.920000 13.910000 63.240000 ;
      LAYER met4 ;
        RECT 13.590000 62.920000 13.910000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590000 63.330000 13.910000 63.650000 ;
      LAYER met4 ;
        RECT 13.590000 63.330000 13.910000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590000 63.740000 13.910000 64.060000 ;
      LAYER met4 ;
        RECT 13.590000 63.740000 13.910000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590000 64.150000 13.910000 64.470000 ;
      LAYER met4 ;
        RECT 13.590000 64.150000 13.910000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590000 64.560000 13.910000 64.880000 ;
      LAYER met4 ;
        RECT 13.590000 64.560000 13.910000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590000 64.970000 13.910000 65.290000 ;
      LAYER met4 ;
        RECT 13.590000 64.970000 13.910000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590000 65.380000 13.910000 65.700000 ;
      LAYER met4 ;
        RECT 13.590000 65.380000 13.910000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590000 65.790000 13.910000 66.110000 ;
      LAYER met4 ;
        RECT 13.590000 65.790000 13.910000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590000 66.200000 13.910000 66.520000 ;
      LAYER met4 ;
        RECT 13.590000 66.200000 13.910000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995000 62.100000 14.315000 62.420000 ;
      LAYER met4 ;
        RECT 13.995000 62.100000 14.315000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995000 62.510000 14.315000 62.830000 ;
      LAYER met4 ;
        RECT 13.995000 62.510000 14.315000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995000 62.920000 14.315000 63.240000 ;
      LAYER met4 ;
        RECT 13.995000 62.920000 14.315000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995000 63.330000 14.315000 63.650000 ;
      LAYER met4 ;
        RECT 13.995000 63.330000 14.315000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995000 63.740000 14.315000 64.060000 ;
      LAYER met4 ;
        RECT 13.995000 63.740000 14.315000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995000 64.150000 14.315000 64.470000 ;
      LAYER met4 ;
        RECT 13.995000 64.150000 14.315000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995000 64.560000 14.315000 64.880000 ;
      LAYER met4 ;
        RECT 13.995000 64.560000 14.315000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995000 64.970000 14.315000 65.290000 ;
      LAYER met4 ;
        RECT 13.995000 64.970000 14.315000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995000 65.380000 14.315000 65.700000 ;
      LAYER met4 ;
        RECT 13.995000 65.380000 14.315000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995000 65.790000 14.315000 66.110000 ;
      LAYER met4 ;
        RECT 13.995000 65.790000 14.315000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995000 66.200000 14.315000 66.520000 ;
      LAYER met4 ;
        RECT 13.995000 66.200000 14.315000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400000 62.100000 14.720000 62.420000 ;
      LAYER met4 ;
        RECT 14.400000 62.100000 14.720000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400000 62.510000 14.720000 62.830000 ;
      LAYER met4 ;
        RECT 14.400000 62.510000 14.720000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400000 62.920000 14.720000 63.240000 ;
      LAYER met4 ;
        RECT 14.400000 62.920000 14.720000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400000 63.330000 14.720000 63.650000 ;
      LAYER met4 ;
        RECT 14.400000 63.330000 14.720000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400000 63.740000 14.720000 64.060000 ;
      LAYER met4 ;
        RECT 14.400000 63.740000 14.720000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400000 64.150000 14.720000 64.470000 ;
      LAYER met4 ;
        RECT 14.400000 64.150000 14.720000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400000 64.560000 14.720000 64.880000 ;
      LAYER met4 ;
        RECT 14.400000 64.560000 14.720000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400000 64.970000 14.720000 65.290000 ;
      LAYER met4 ;
        RECT 14.400000 64.970000 14.720000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400000 65.380000 14.720000 65.700000 ;
      LAYER met4 ;
        RECT 14.400000 65.380000 14.720000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400000 65.790000 14.720000 66.110000 ;
      LAYER met4 ;
        RECT 14.400000 65.790000 14.720000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400000 66.200000 14.720000 66.520000 ;
      LAYER met4 ;
        RECT 14.400000 66.200000 14.720000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805000 62.100000 15.125000 62.420000 ;
      LAYER met4 ;
        RECT 14.805000 62.100000 15.125000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805000 62.510000 15.125000 62.830000 ;
      LAYER met4 ;
        RECT 14.805000 62.510000 15.125000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805000 62.920000 15.125000 63.240000 ;
      LAYER met4 ;
        RECT 14.805000 62.920000 15.125000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805000 63.330000 15.125000 63.650000 ;
      LAYER met4 ;
        RECT 14.805000 63.330000 15.125000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805000 63.740000 15.125000 64.060000 ;
      LAYER met4 ;
        RECT 14.805000 63.740000 15.125000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805000 64.150000 15.125000 64.470000 ;
      LAYER met4 ;
        RECT 14.805000 64.150000 15.125000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805000 64.560000 15.125000 64.880000 ;
      LAYER met4 ;
        RECT 14.805000 64.560000 15.125000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805000 64.970000 15.125000 65.290000 ;
      LAYER met4 ;
        RECT 14.805000 64.970000 15.125000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805000 65.380000 15.125000 65.700000 ;
      LAYER met4 ;
        RECT 14.805000 65.380000 15.125000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805000 65.790000 15.125000 66.110000 ;
      LAYER met4 ;
        RECT 14.805000 65.790000 15.125000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805000 66.200000 15.125000 66.520000 ;
      LAYER met4 ;
        RECT 14.805000 66.200000 15.125000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210000 62.100000 15.530000 62.420000 ;
      LAYER met4 ;
        RECT 15.210000 62.100000 15.530000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210000 62.510000 15.530000 62.830000 ;
      LAYER met4 ;
        RECT 15.210000 62.510000 15.530000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210000 62.920000 15.530000 63.240000 ;
      LAYER met4 ;
        RECT 15.210000 62.920000 15.530000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210000 63.330000 15.530000 63.650000 ;
      LAYER met4 ;
        RECT 15.210000 63.330000 15.530000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210000 63.740000 15.530000 64.060000 ;
      LAYER met4 ;
        RECT 15.210000 63.740000 15.530000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210000 64.150000 15.530000 64.470000 ;
      LAYER met4 ;
        RECT 15.210000 64.150000 15.530000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210000 64.560000 15.530000 64.880000 ;
      LAYER met4 ;
        RECT 15.210000 64.560000 15.530000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210000 64.970000 15.530000 65.290000 ;
      LAYER met4 ;
        RECT 15.210000 64.970000 15.530000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210000 65.380000 15.530000 65.700000 ;
      LAYER met4 ;
        RECT 15.210000 65.380000 15.530000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210000 65.790000 15.530000 66.110000 ;
      LAYER met4 ;
        RECT 15.210000 65.790000 15.530000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210000 66.200000 15.530000 66.520000 ;
      LAYER met4 ;
        RECT 15.210000 66.200000 15.530000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615000 62.100000 15.935000 62.420000 ;
      LAYER met4 ;
        RECT 15.615000 62.100000 15.935000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615000 62.510000 15.935000 62.830000 ;
      LAYER met4 ;
        RECT 15.615000 62.510000 15.935000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615000 62.920000 15.935000 63.240000 ;
      LAYER met4 ;
        RECT 15.615000 62.920000 15.935000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615000 63.330000 15.935000 63.650000 ;
      LAYER met4 ;
        RECT 15.615000 63.330000 15.935000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615000 63.740000 15.935000 64.060000 ;
      LAYER met4 ;
        RECT 15.615000 63.740000 15.935000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615000 64.150000 15.935000 64.470000 ;
      LAYER met4 ;
        RECT 15.615000 64.150000 15.935000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615000 64.560000 15.935000 64.880000 ;
      LAYER met4 ;
        RECT 15.615000 64.560000 15.935000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615000 64.970000 15.935000 65.290000 ;
      LAYER met4 ;
        RECT 15.615000 64.970000 15.935000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615000 65.380000 15.935000 65.700000 ;
      LAYER met4 ;
        RECT 15.615000 65.380000 15.935000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615000 65.790000 15.935000 66.110000 ;
      LAYER met4 ;
        RECT 15.615000 65.790000 15.935000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615000 66.200000 15.935000 66.520000 ;
      LAYER met4 ;
        RECT 15.615000 66.200000 15.935000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020000 62.100000 16.340000 62.420000 ;
      LAYER met4 ;
        RECT 16.020000 62.100000 16.340000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020000 62.510000 16.340000 62.830000 ;
      LAYER met4 ;
        RECT 16.020000 62.510000 16.340000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020000 62.920000 16.340000 63.240000 ;
      LAYER met4 ;
        RECT 16.020000 62.920000 16.340000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020000 63.330000 16.340000 63.650000 ;
      LAYER met4 ;
        RECT 16.020000 63.330000 16.340000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020000 63.740000 16.340000 64.060000 ;
      LAYER met4 ;
        RECT 16.020000 63.740000 16.340000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020000 64.150000 16.340000 64.470000 ;
      LAYER met4 ;
        RECT 16.020000 64.150000 16.340000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020000 64.560000 16.340000 64.880000 ;
      LAYER met4 ;
        RECT 16.020000 64.560000 16.340000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020000 64.970000 16.340000 65.290000 ;
      LAYER met4 ;
        RECT 16.020000 64.970000 16.340000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020000 65.380000 16.340000 65.700000 ;
      LAYER met4 ;
        RECT 16.020000 65.380000 16.340000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020000 65.790000 16.340000 66.110000 ;
      LAYER met4 ;
        RECT 16.020000 65.790000 16.340000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020000 66.200000 16.340000 66.520000 ;
      LAYER met4 ;
        RECT 16.020000 66.200000 16.340000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425000 62.100000 16.745000 62.420000 ;
      LAYER met4 ;
        RECT 16.425000 62.100000 16.745000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425000 62.510000 16.745000 62.830000 ;
      LAYER met4 ;
        RECT 16.425000 62.510000 16.745000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425000 62.920000 16.745000 63.240000 ;
      LAYER met4 ;
        RECT 16.425000 62.920000 16.745000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425000 63.330000 16.745000 63.650000 ;
      LAYER met4 ;
        RECT 16.425000 63.330000 16.745000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425000 63.740000 16.745000 64.060000 ;
      LAYER met4 ;
        RECT 16.425000 63.740000 16.745000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425000 64.150000 16.745000 64.470000 ;
      LAYER met4 ;
        RECT 16.425000 64.150000 16.745000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425000 64.560000 16.745000 64.880000 ;
      LAYER met4 ;
        RECT 16.425000 64.560000 16.745000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425000 64.970000 16.745000 65.290000 ;
      LAYER met4 ;
        RECT 16.425000 64.970000 16.745000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425000 65.380000 16.745000 65.700000 ;
      LAYER met4 ;
        RECT 16.425000 65.380000 16.745000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425000 65.790000 16.745000 66.110000 ;
      LAYER met4 ;
        RECT 16.425000 65.790000 16.745000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425000 66.200000 16.745000 66.520000 ;
      LAYER met4 ;
        RECT 16.425000 66.200000 16.745000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830000 62.100000 17.150000 62.420000 ;
      LAYER met4 ;
        RECT 16.830000 62.100000 17.150000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830000 62.510000 17.150000 62.830000 ;
      LAYER met4 ;
        RECT 16.830000 62.510000 17.150000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830000 62.920000 17.150000 63.240000 ;
      LAYER met4 ;
        RECT 16.830000 62.920000 17.150000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830000 63.330000 17.150000 63.650000 ;
      LAYER met4 ;
        RECT 16.830000 63.330000 17.150000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830000 63.740000 17.150000 64.060000 ;
      LAYER met4 ;
        RECT 16.830000 63.740000 17.150000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830000 64.150000 17.150000 64.470000 ;
      LAYER met4 ;
        RECT 16.830000 64.150000 17.150000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830000 64.560000 17.150000 64.880000 ;
      LAYER met4 ;
        RECT 16.830000 64.560000 17.150000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830000 64.970000 17.150000 65.290000 ;
      LAYER met4 ;
        RECT 16.830000 64.970000 17.150000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830000 65.380000 17.150000 65.700000 ;
      LAYER met4 ;
        RECT 16.830000 65.380000 17.150000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830000 65.790000 17.150000 66.110000 ;
      LAYER met4 ;
        RECT 16.830000 65.790000 17.150000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830000 66.200000 17.150000 66.520000 ;
      LAYER met4 ;
        RECT 16.830000 66.200000 17.150000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235000 62.100000 17.555000 62.420000 ;
      LAYER met4 ;
        RECT 17.235000 62.100000 17.555000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235000 62.510000 17.555000 62.830000 ;
      LAYER met4 ;
        RECT 17.235000 62.510000 17.555000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235000 62.920000 17.555000 63.240000 ;
      LAYER met4 ;
        RECT 17.235000 62.920000 17.555000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235000 63.330000 17.555000 63.650000 ;
      LAYER met4 ;
        RECT 17.235000 63.330000 17.555000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235000 63.740000 17.555000 64.060000 ;
      LAYER met4 ;
        RECT 17.235000 63.740000 17.555000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235000 64.150000 17.555000 64.470000 ;
      LAYER met4 ;
        RECT 17.235000 64.150000 17.555000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235000 64.560000 17.555000 64.880000 ;
      LAYER met4 ;
        RECT 17.235000 64.560000 17.555000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235000 64.970000 17.555000 65.290000 ;
      LAYER met4 ;
        RECT 17.235000 64.970000 17.555000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235000 65.380000 17.555000 65.700000 ;
      LAYER met4 ;
        RECT 17.235000 65.380000 17.555000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235000 65.790000 17.555000 66.110000 ;
      LAYER met4 ;
        RECT 17.235000 65.790000 17.555000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235000 66.200000 17.555000 66.520000 ;
      LAYER met4 ;
        RECT 17.235000 66.200000 17.555000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640000 62.100000 17.960000 62.420000 ;
      LAYER met4 ;
        RECT 17.640000 62.100000 17.960000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640000 62.510000 17.960000 62.830000 ;
      LAYER met4 ;
        RECT 17.640000 62.510000 17.960000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640000 62.920000 17.960000 63.240000 ;
      LAYER met4 ;
        RECT 17.640000 62.920000 17.960000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640000 63.330000 17.960000 63.650000 ;
      LAYER met4 ;
        RECT 17.640000 63.330000 17.960000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640000 63.740000 17.960000 64.060000 ;
      LAYER met4 ;
        RECT 17.640000 63.740000 17.960000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640000 64.150000 17.960000 64.470000 ;
      LAYER met4 ;
        RECT 17.640000 64.150000 17.960000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640000 64.560000 17.960000 64.880000 ;
      LAYER met4 ;
        RECT 17.640000 64.560000 17.960000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640000 64.970000 17.960000 65.290000 ;
      LAYER met4 ;
        RECT 17.640000 64.970000 17.960000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640000 65.380000 17.960000 65.700000 ;
      LAYER met4 ;
        RECT 17.640000 65.380000 17.960000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640000 65.790000 17.960000 66.110000 ;
      LAYER met4 ;
        RECT 17.640000 65.790000 17.960000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640000 66.200000 17.960000 66.520000 ;
      LAYER met4 ;
        RECT 17.640000 66.200000 17.960000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 62.100000 18.365000 62.420000 ;
      LAYER met4 ;
        RECT 18.045000 62.100000 18.365000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 62.510000 18.365000 62.830000 ;
      LAYER met4 ;
        RECT 18.045000 62.510000 18.365000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 62.920000 18.365000 63.240000 ;
      LAYER met4 ;
        RECT 18.045000 62.920000 18.365000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 63.330000 18.365000 63.650000 ;
      LAYER met4 ;
        RECT 18.045000 63.330000 18.365000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 63.740000 18.365000 64.060000 ;
      LAYER met4 ;
        RECT 18.045000 63.740000 18.365000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 64.150000 18.365000 64.470000 ;
      LAYER met4 ;
        RECT 18.045000 64.150000 18.365000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 64.560000 18.365000 64.880000 ;
      LAYER met4 ;
        RECT 18.045000 64.560000 18.365000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 64.970000 18.365000 65.290000 ;
      LAYER met4 ;
        RECT 18.045000 64.970000 18.365000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 65.380000 18.365000 65.700000 ;
      LAYER met4 ;
        RECT 18.045000 65.380000 18.365000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 65.790000 18.365000 66.110000 ;
      LAYER met4 ;
        RECT 18.045000 65.790000 18.365000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045000 66.200000 18.365000 66.520000 ;
      LAYER met4 ;
        RECT 18.045000 66.200000 18.365000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450000 62.100000 18.770000 62.420000 ;
      LAYER met4 ;
        RECT 18.450000 62.100000 18.770000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450000 62.510000 18.770000 62.830000 ;
      LAYER met4 ;
        RECT 18.450000 62.510000 18.770000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450000 62.920000 18.770000 63.240000 ;
      LAYER met4 ;
        RECT 18.450000 62.920000 18.770000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450000 63.330000 18.770000 63.650000 ;
      LAYER met4 ;
        RECT 18.450000 63.330000 18.770000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450000 63.740000 18.770000 64.060000 ;
      LAYER met4 ;
        RECT 18.450000 63.740000 18.770000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450000 64.150000 18.770000 64.470000 ;
      LAYER met4 ;
        RECT 18.450000 64.150000 18.770000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450000 64.560000 18.770000 64.880000 ;
      LAYER met4 ;
        RECT 18.450000 64.560000 18.770000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450000 64.970000 18.770000 65.290000 ;
      LAYER met4 ;
        RECT 18.450000 64.970000 18.770000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450000 65.380000 18.770000 65.700000 ;
      LAYER met4 ;
        RECT 18.450000 65.380000 18.770000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450000 65.790000 18.770000 66.110000 ;
      LAYER met4 ;
        RECT 18.450000 65.790000 18.770000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450000 66.200000 18.770000 66.520000 ;
      LAYER met4 ;
        RECT 18.450000 66.200000 18.770000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855000 62.100000 19.175000 62.420000 ;
      LAYER met4 ;
        RECT 18.855000 62.100000 19.175000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855000 62.510000 19.175000 62.830000 ;
      LAYER met4 ;
        RECT 18.855000 62.510000 19.175000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855000 62.920000 19.175000 63.240000 ;
      LAYER met4 ;
        RECT 18.855000 62.920000 19.175000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855000 63.330000 19.175000 63.650000 ;
      LAYER met4 ;
        RECT 18.855000 63.330000 19.175000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855000 63.740000 19.175000 64.060000 ;
      LAYER met4 ;
        RECT 18.855000 63.740000 19.175000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855000 64.150000 19.175000 64.470000 ;
      LAYER met4 ;
        RECT 18.855000 64.150000 19.175000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855000 64.560000 19.175000 64.880000 ;
      LAYER met4 ;
        RECT 18.855000 64.560000 19.175000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855000 64.970000 19.175000 65.290000 ;
      LAYER met4 ;
        RECT 18.855000 64.970000 19.175000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855000 65.380000 19.175000 65.700000 ;
      LAYER met4 ;
        RECT 18.855000 65.380000 19.175000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855000 65.790000 19.175000 66.110000 ;
      LAYER met4 ;
        RECT 18.855000 65.790000 19.175000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855000 66.200000 19.175000 66.520000 ;
      LAYER met4 ;
        RECT 18.855000 66.200000 19.175000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260000 62.100000 19.580000 62.420000 ;
      LAYER met4 ;
        RECT 19.260000 62.100000 19.580000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260000 62.510000 19.580000 62.830000 ;
      LAYER met4 ;
        RECT 19.260000 62.510000 19.580000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260000 62.920000 19.580000 63.240000 ;
      LAYER met4 ;
        RECT 19.260000 62.920000 19.580000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260000 63.330000 19.580000 63.650000 ;
      LAYER met4 ;
        RECT 19.260000 63.330000 19.580000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260000 63.740000 19.580000 64.060000 ;
      LAYER met4 ;
        RECT 19.260000 63.740000 19.580000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260000 64.150000 19.580000 64.470000 ;
      LAYER met4 ;
        RECT 19.260000 64.150000 19.580000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260000 64.560000 19.580000 64.880000 ;
      LAYER met4 ;
        RECT 19.260000 64.560000 19.580000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260000 64.970000 19.580000 65.290000 ;
      LAYER met4 ;
        RECT 19.260000 64.970000 19.580000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260000 65.380000 19.580000 65.700000 ;
      LAYER met4 ;
        RECT 19.260000 65.380000 19.580000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260000 65.790000 19.580000 66.110000 ;
      LAYER met4 ;
        RECT 19.260000 65.790000 19.580000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260000 66.200000 19.580000 66.520000 ;
      LAYER met4 ;
        RECT 19.260000 66.200000 19.580000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665000 62.100000 19.985000 62.420000 ;
      LAYER met4 ;
        RECT 19.665000 62.100000 19.985000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665000 62.510000 19.985000 62.830000 ;
      LAYER met4 ;
        RECT 19.665000 62.510000 19.985000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665000 62.920000 19.985000 63.240000 ;
      LAYER met4 ;
        RECT 19.665000 62.920000 19.985000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665000 63.330000 19.985000 63.650000 ;
      LAYER met4 ;
        RECT 19.665000 63.330000 19.985000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665000 63.740000 19.985000 64.060000 ;
      LAYER met4 ;
        RECT 19.665000 63.740000 19.985000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665000 64.150000 19.985000 64.470000 ;
      LAYER met4 ;
        RECT 19.665000 64.150000 19.985000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665000 64.560000 19.985000 64.880000 ;
      LAYER met4 ;
        RECT 19.665000 64.560000 19.985000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665000 64.970000 19.985000 65.290000 ;
      LAYER met4 ;
        RECT 19.665000 64.970000 19.985000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665000 65.380000 19.985000 65.700000 ;
      LAYER met4 ;
        RECT 19.665000 65.380000 19.985000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665000 65.790000 19.985000 66.110000 ;
      LAYER met4 ;
        RECT 19.665000 65.790000 19.985000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665000 66.200000 19.985000 66.520000 ;
      LAYER met4 ;
        RECT 19.665000 66.200000 19.985000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250000 62.100000 2.570000 62.420000 ;
      LAYER met4 ;
        RECT 2.250000 62.100000 2.570000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250000 62.510000 2.570000 62.830000 ;
      LAYER met4 ;
        RECT 2.250000 62.510000 2.570000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250000 62.920000 2.570000 63.240000 ;
      LAYER met4 ;
        RECT 2.250000 62.920000 2.570000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250000 63.330000 2.570000 63.650000 ;
      LAYER met4 ;
        RECT 2.250000 63.330000 2.570000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250000 63.740000 2.570000 64.060000 ;
      LAYER met4 ;
        RECT 2.250000 63.740000 2.570000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250000 64.150000 2.570000 64.470000 ;
      LAYER met4 ;
        RECT 2.250000 64.150000 2.570000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250000 64.560000 2.570000 64.880000 ;
      LAYER met4 ;
        RECT 2.250000 64.560000 2.570000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250000 64.970000 2.570000 65.290000 ;
      LAYER met4 ;
        RECT 2.250000 64.970000 2.570000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250000 65.380000 2.570000 65.700000 ;
      LAYER met4 ;
        RECT 2.250000 65.380000 2.570000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250000 65.790000 2.570000 66.110000 ;
      LAYER met4 ;
        RECT 2.250000 65.790000 2.570000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250000 66.200000 2.570000 66.520000 ;
      LAYER met4 ;
        RECT 2.250000 66.200000 2.570000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655000 62.100000 2.975000 62.420000 ;
      LAYER met4 ;
        RECT 2.655000 62.100000 2.975000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655000 62.510000 2.975000 62.830000 ;
      LAYER met4 ;
        RECT 2.655000 62.510000 2.975000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655000 62.920000 2.975000 63.240000 ;
      LAYER met4 ;
        RECT 2.655000 62.920000 2.975000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655000 63.330000 2.975000 63.650000 ;
      LAYER met4 ;
        RECT 2.655000 63.330000 2.975000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655000 63.740000 2.975000 64.060000 ;
      LAYER met4 ;
        RECT 2.655000 63.740000 2.975000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655000 64.150000 2.975000 64.470000 ;
      LAYER met4 ;
        RECT 2.655000 64.150000 2.975000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655000 64.560000 2.975000 64.880000 ;
      LAYER met4 ;
        RECT 2.655000 64.560000 2.975000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655000 64.970000 2.975000 65.290000 ;
      LAYER met4 ;
        RECT 2.655000 64.970000 2.975000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655000 65.380000 2.975000 65.700000 ;
      LAYER met4 ;
        RECT 2.655000 65.380000 2.975000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655000 65.790000 2.975000 66.110000 ;
      LAYER met4 ;
        RECT 2.655000 65.790000 2.975000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655000 66.200000 2.975000 66.520000 ;
      LAYER met4 ;
        RECT 2.655000 66.200000 2.975000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070000 62.100000 20.390000 62.420000 ;
      LAYER met4 ;
        RECT 20.070000 62.100000 20.390000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070000 62.510000 20.390000 62.830000 ;
      LAYER met4 ;
        RECT 20.070000 62.510000 20.390000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070000 62.920000 20.390000 63.240000 ;
      LAYER met4 ;
        RECT 20.070000 62.920000 20.390000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070000 63.330000 20.390000 63.650000 ;
      LAYER met4 ;
        RECT 20.070000 63.330000 20.390000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070000 63.740000 20.390000 64.060000 ;
      LAYER met4 ;
        RECT 20.070000 63.740000 20.390000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070000 64.150000 20.390000 64.470000 ;
      LAYER met4 ;
        RECT 20.070000 64.150000 20.390000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070000 64.560000 20.390000 64.880000 ;
      LAYER met4 ;
        RECT 20.070000 64.560000 20.390000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070000 64.970000 20.390000 65.290000 ;
      LAYER met4 ;
        RECT 20.070000 64.970000 20.390000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070000 65.380000 20.390000 65.700000 ;
      LAYER met4 ;
        RECT 20.070000 65.380000 20.390000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070000 65.790000 20.390000 66.110000 ;
      LAYER met4 ;
        RECT 20.070000 65.790000 20.390000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070000 66.200000 20.390000 66.520000 ;
      LAYER met4 ;
        RECT 20.070000 66.200000 20.390000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475000 62.100000 20.795000 62.420000 ;
      LAYER met4 ;
        RECT 20.475000 62.100000 20.795000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475000 62.510000 20.795000 62.830000 ;
      LAYER met4 ;
        RECT 20.475000 62.510000 20.795000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475000 62.920000 20.795000 63.240000 ;
      LAYER met4 ;
        RECT 20.475000 62.920000 20.795000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475000 63.330000 20.795000 63.650000 ;
      LAYER met4 ;
        RECT 20.475000 63.330000 20.795000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475000 63.740000 20.795000 64.060000 ;
      LAYER met4 ;
        RECT 20.475000 63.740000 20.795000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475000 64.150000 20.795000 64.470000 ;
      LAYER met4 ;
        RECT 20.475000 64.150000 20.795000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475000 64.560000 20.795000 64.880000 ;
      LAYER met4 ;
        RECT 20.475000 64.560000 20.795000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475000 64.970000 20.795000 65.290000 ;
      LAYER met4 ;
        RECT 20.475000 64.970000 20.795000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475000 65.380000 20.795000 65.700000 ;
      LAYER met4 ;
        RECT 20.475000 65.380000 20.795000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475000 65.790000 20.795000 66.110000 ;
      LAYER met4 ;
        RECT 20.475000 65.790000 20.795000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475000 66.200000 20.795000 66.520000 ;
      LAYER met4 ;
        RECT 20.475000 66.200000 20.795000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880000 62.100000 21.200000 62.420000 ;
      LAYER met4 ;
        RECT 20.880000 62.100000 21.200000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880000 62.510000 21.200000 62.830000 ;
      LAYER met4 ;
        RECT 20.880000 62.510000 21.200000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880000 62.920000 21.200000 63.240000 ;
      LAYER met4 ;
        RECT 20.880000 62.920000 21.200000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880000 63.330000 21.200000 63.650000 ;
      LAYER met4 ;
        RECT 20.880000 63.330000 21.200000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880000 63.740000 21.200000 64.060000 ;
      LAYER met4 ;
        RECT 20.880000 63.740000 21.200000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880000 64.150000 21.200000 64.470000 ;
      LAYER met4 ;
        RECT 20.880000 64.150000 21.200000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880000 64.560000 21.200000 64.880000 ;
      LAYER met4 ;
        RECT 20.880000 64.560000 21.200000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880000 64.970000 21.200000 65.290000 ;
      LAYER met4 ;
        RECT 20.880000 64.970000 21.200000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880000 65.380000 21.200000 65.700000 ;
      LAYER met4 ;
        RECT 20.880000 65.380000 21.200000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880000 65.790000 21.200000 66.110000 ;
      LAYER met4 ;
        RECT 20.880000 65.790000 21.200000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880000 66.200000 21.200000 66.520000 ;
      LAYER met4 ;
        RECT 20.880000 66.200000 21.200000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285000 62.100000 21.605000 62.420000 ;
      LAYER met4 ;
        RECT 21.285000 62.100000 21.605000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285000 62.510000 21.605000 62.830000 ;
      LAYER met4 ;
        RECT 21.285000 62.510000 21.605000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285000 62.920000 21.605000 63.240000 ;
      LAYER met4 ;
        RECT 21.285000 62.920000 21.605000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285000 63.330000 21.605000 63.650000 ;
      LAYER met4 ;
        RECT 21.285000 63.330000 21.605000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285000 63.740000 21.605000 64.060000 ;
      LAYER met4 ;
        RECT 21.285000 63.740000 21.605000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285000 64.150000 21.605000 64.470000 ;
      LAYER met4 ;
        RECT 21.285000 64.150000 21.605000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285000 64.560000 21.605000 64.880000 ;
      LAYER met4 ;
        RECT 21.285000 64.560000 21.605000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285000 64.970000 21.605000 65.290000 ;
      LAYER met4 ;
        RECT 21.285000 64.970000 21.605000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285000 65.380000 21.605000 65.700000 ;
      LAYER met4 ;
        RECT 21.285000 65.380000 21.605000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285000 65.790000 21.605000 66.110000 ;
      LAYER met4 ;
        RECT 21.285000 65.790000 21.605000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285000 66.200000 21.605000 66.520000 ;
      LAYER met4 ;
        RECT 21.285000 66.200000 21.605000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690000 62.100000 22.010000 62.420000 ;
      LAYER met4 ;
        RECT 21.690000 62.100000 22.010000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690000 62.510000 22.010000 62.830000 ;
      LAYER met4 ;
        RECT 21.690000 62.510000 22.010000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690000 62.920000 22.010000 63.240000 ;
      LAYER met4 ;
        RECT 21.690000 62.920000 22.010000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690000 63.330000 22.010000 63.650000 ;
      LAYER met4 ;
        RECT 21.690000 63.330000 22.010000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690000 63.740000 22.010000 64.060000 ;
      LAYER met4 ;
        RECT 21.690000 63.740000 22.010000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690000 64.150000 22.010000 64.470000 ;
      LAYER met4 ;
        RECT 21.690000 64.150000 22.010000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690000 64.560000 22.010000 64.880000 ;
      LAYER met4 ;
        RECT 21.690000 64.560000 22.010000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690000 64.970000 22.010000 65.290000 ;
      LAYER met4 ;
        RECT 21.690000 64.970000 22.010000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690000 65.380000 22.010000 65.700000 ;
      LAYER met4 ;
        RECT 21.690000 65.380000 22.010000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690000 65.790000 22.010000 66.110000 ;
      LAYER met4 ;
        RECT 21.690000 65.790000 22.010000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690000 66.200000 22.010000 66.520000 ;
      LAYER met4 ;
        RECT 21.690000 66.200000 22.010000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100000 62.100000 22.420000 62.420000 ;
      LAYER met4 ;
        RECT 22.100000 62.100000 22.420000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100000 62.510000 22.420000 62.830000 ;
      LAYER met4 ;
        RECT 22.100000 62.510000 22.420000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100000 62.920000 22.420000 63.240000 ;
      LAYER met4 ;
        RECT 22.100000 62.920000 22.420000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100000 63.330000 22.420000 63.650000 ;
      LAYER met4 ;
        RECT 22.100000 63.330000 22.420000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100000 63.740000 22.420000 64.060000 ;
      LAYER met4 ;
        RECT 22.100000 63.740000 22.420000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100000 64.150000 22.420000 64.470000 ;
      LAYER met4 ;
        RECT 22.100000 64.150000 22.420000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100000 64.560000 22.420000 64.880000 ;
      LAYER met4 ;
        RECT 22.100000 64.560000 22.420000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100000 64.970000 22.420000 65.290000 ;
      LAYER met4 ;
        RECT 22.100000 64.970000 22.420000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100000 65.380000 22.420000 65.700000 ;
      LAYER met4 ;
        RECT 22.100000 65.380000 22.420000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100000 65.790000 22.420000 66.110000 ;
      LAYER met4 ;
        RECT 22.100000 65.790000 22.420000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100000 66.200000 22.420000 66.520000 ;
      LAYER met4 ;
        RECT 22.100000 66.200000 22.420000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510000 62.100000 22.830000 62.420000 ;
      LAYER met4 ;
        RECT 22.510000 62.100000 22.830000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510000 62.510000 22.830000 62.830000 ;
      LAYER met4 ;
        RECT 22.510000 62.510000 22.830000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510000 62.920000 22.830000 63.240000 ;
      LAYER met4 ;
        RECT 22.510000 62.920000 22.830000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510000 63.330000 22.830000 63.650000 ;
      LAYER met4 ;
        RECT 22.510000 63.330000 22.830000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510000 63.740000 22.830000 64.060000 ;
      LAYER met4 ;
        RECT 22.510000 63.740000 22.830000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510000 64.150000 22.830000 64.470000 ;
      LAYER met4 ;
        RECT 22.510000 64.150000 22.830000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510000 64.560000 22.830000 64.880000 ;
      LAYER met4 ;
        RECT 22.510000 64.560000 22.830000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510000 64.970000 22.830000 65.290000 ;
      LAYER met4 ;
        RECT 22.510000 64.970000 22.830000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510000 65.380000 22.830000 65.700000 ;
      LAYER met4 ;
        RECT 22.510000 65.380000 22.830000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510000 65.790000 22.830000 66.110000 ;
      LAYER met4 ;
        RECT 22.510000 65.790000 22.830000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510000 66.200000 22.830000 66.520000 ;
      LAYER met4 ;
        RECT 22.510000 66.200000 22.830000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920000 62.100000 23.240000 62.420000 ;
      LAYER met4 ;
        RECT 22.920000 62.100000 23.240000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920000 62.510000 23.240000 62.830000 ;
      LAYER met4 ;
        RECT 22.920000 62.510000 23.240000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920000 62.920000 23.240000 63.240000 ;
      LAYER met4 ;
        RECT 22.920000 62.920000 23.240000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920000 63.330000 23.240000 63.650000 ;
      LAYER met4 ;
        RECT 22.920000 63.330000 23.240000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920000 63.740000 23.240000 64.060000 ;
      LAYER met4 ;
        RECT 22.920000 63.740000 23.240000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920000 64.150000 23.240000 64.470000 ;
      LAYER met4 ;
        RECT 22.920000 64.150000 23.240000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920000 64.560000 23.240000 64.880000 ;
      LAYER met4 ;
        RECT 22.920000 64.560000 23.240000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920000 64.970000 23.240000 65.290000 ;
      LAYER met4 ;
        RECT 22.920000 64.970000 23.240000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920000 65.380000 23.240000 65.700000 ;
      LAYER met4 ;
        RECT 22.920000 65.380000 23.240000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920000 65.790000 23.240000 66.110000 ;
      LAYER met4 ;
        RECT 22.920000 65.790000 23.240000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920000 66.200000 23.240000 66.520000 ;
      LAYER met4 ;
        RECT 22.920000 66.200000 23.240000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330000 62.100000 23.650000 62.420000 ;
      LAYER met4 ;
        RECT 23.330000 62.100000 23.650000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330000 62.510000 23.650000 62.830000 ;
      LAYER met4 ;
        RECT 23.330000 62.510000 23.650000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330000 62.920000 23.650000 63.240000 ;
      LAYER met4 ;
        RECT 23.330000 62.920000 23.650000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330000 63.330000 23.650000 63.650000 ;
      LAYER met4 ;
        RECT 23.330000 63.330000 23.650000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330000 63.740000 23.650000 64.060000 ;
      LAYER met4 ;
        RECT 23.330000 63.740000 23.650000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330000 64.150000 23.650000 64.470000 ;
      LAYER met4 ;
        RECT 23.330000 64.150000 23.650000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330000 64.560000 23.650000 64.880000 ;
      LAYER met4 ;
        RECT 23.330000 64.560000 23.650000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330000 64.970000 23.650000 65.290000 ;
      LAYER met4 ;
        RECT 23.330000 64.970000 23.650000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330000 65.380000 23.650000 65.700000 ;
      LAYER met4 ;
        RECT 23.330000 65.380000 23.650000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330000 65.790000 23.650000 66.110000 ;
      LAYER met4 ;
        RECT 23.330000 65.790000 23.650000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330000 66.200000 23.650000 66.520000 ;
      LAYER met4 ;
        RECT 23.330000 66.200000 23.650000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740000 62.100000 24.060000 62.420000 ;
      LAYER met4 ;
        RECT 23.740000 62.100000 24.060000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740000 62.510000 24.060000 62.830000 ;
      LAYER met4 ;
        RECT 23.740000 62.510000 24.060000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740000 62.920000 24.060000 63.240000 ;
      LAYER met4 ;
        RECT 23.740000 62.920000 24.060000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740000 63.330000 24.060000 63.650000 ;
      LAYER met4 ;
        RECT 23.740000 63.330000 24.060000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740000 63.740000 24.060000 64.060000 ;
      LAYER met4 ;
        RECT 23.740000 63.740000 24.060000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740000 64.150000 24.060000 64.470000 ;
      LAYER met4 ;
        RECT 23.740000 64.150000 24.060000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740000 64.560000 24.060000 64.880000 ;
      LAYER met4 ;
        RECT 23.740000 64.560000 24.060000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740000 64.970000 24.060000 65.290000 ;
      LAYER met4 ;
        RECT 23.740000 64.970000 24.060000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740000 65.380000 24.060000 65.700000 ;
      LAYER met4 ;
        RECT 23.740000 65.380000 24.060000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740000 65.790000 24.060000 66.110000 ;
      LAYER met4 ;
        RECT 23.740000 65.790000 24.060000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740000 66.200000 24.060000 66.520000 ;
      LAYER met4 ;
        RECT 23.740000 66.200000 24.060000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 62.100000 24.470000 62.420000 ;
      LAYER met4 ;
        RECT 24.150000 62.100000 24.470000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 62.510000 24.470000 62.830000 ;
      LAYER met4 ;
        RECT 24.150000 62.510000 24.470000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 62.920000 24.470000 63.240000 ;
      LAYER met4 ;
        RECT 24.150000 62.920000 24.470000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 63.330000 24.470000 63.650000 ;
      LAYER met4 ;
        RECT 24.150000 63.330000 24.470000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 63.740000 24.470000 64.060000 ;
      LAYER met4 ;
        RECT 24.150000 63.740000 24.470000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 64.150000 24.470000 64.470000 ;
      LAYER met4 ;
        RECT 24.150000 64.150000 24.470000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 64.560000 24.470000 64.880000 ;
      LAYER met4 ;
        RECT 24.150000 64.560000 24.470000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 64.970000 24.470000 65.290000 ;
      LAYER met4 ;
        RECT 24.150000 64.970000 24.470000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 65.380000 24.470000 65.700000 ;
      LAYER met4 ;
        RECT 24.150000 65.380000 24.470000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 65.790000 24.470000 66.110000 ;
      LAYER met4 ;
        RECT 24.150000 65.790000 24.470000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 66.200000 24.470000 66.520000 ;
      LAYER met4 ;
        RECT 24.150000 66.200000 24.470000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060000 62.100000 3.380000 62.420000 ;
      LAYER met4 ;
        RECT 3.060000 62.100000 3.380000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060000 62.510000 3.380000 62.830000 ;
      LAYER met4 ;
        RECT 3.060000 62.510000 3.380000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060000 62.920000 3.380000 63.240000 ;
      LAYER met4 ;
        RECT 3.060000 62.920000 3.380000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060000 63.330000 3.380000 63.650000 ;
      LAYER met4 ;
        RECT 3.060000 63.330000 3.380000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060000 63.740000 3.380000 64.060000 ;
      LAYER met4 ;
        RECT 3.060000 63.740000 3.380000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060000 64.150000 3.380000 64.470000 ;
      LAYER met4 ;
        RECT 3.060000 64.150000 3.380000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060000 64.560000 3.380000 64.880000 ;
      LAYER met4 ;
        RECT 3.060000 64.560000 3.380000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060000 64.970000 3.380000 65.290000 ;
      LAYER met4 ;
        RECT 3.060000 64.970000 3.380000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060000 65.380000 3.380000 65.700000 ;
      LAYER met4 ;
        RECT 3.060000 65.380000 3.380000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060000 65.790000 3.380000 66.110000 ;
      LAYER met4 ;
        RECT 3.060000 65.790000 3.380000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060000 66.200000 3.380000 66.520000 ;
      LAYER met4 ;
        RECT 3.060000 66.200000 3.380000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465000 62.100000 3.785000 62.420000 ;
      LAYER met4 ;
        RECT 3.465000 62.100000 3.785000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465000 62.510000 3.785000 62.830000 ;
      LAYER met4 ;
        RECT 3.465000 62.510000 3.785000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465000 62.920000 3.785000 63.240000 ;
      LAYER met4 ;
        RECT 3.465000 62.920000 3.785000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465000 63.330000 3.785000 63.650000 ;
      LAYER met4 ;
        RECT 3.465000 63.330000 3.785000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465000 63.740000 3.785000 64.060000 ;
      LAYER met4 ;
        RECT 3.465000 63.740000 3.785000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465000 64.150000 3.785000 64.470000 ;
      LAYER met4 ;
        RECT 3.465000 64.150000 3.785000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465000 64.560000 3.785000 64.880000 ;
      LAYER met4 ;
        RECT 3.465000 64.560000 3.785000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465000 64.970000 3.785000 65.290000 ;
      LAYER met4 ;
        RECT 3.465000 64.970000 3.785000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465000 65.380000 3.785000 65.700000 ;
      LAYER met4 ;
        RECT 3.465000 65.380000 3.785000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465000 65.790000 3.785000 66.110000 ;
      LAYER met4 ;
        RECT 3.465000 65.790000 3.785000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465000 66.200000 3.785000 66.520000 ;
      LAYER met4 ;
        RECT 3.465000 66.200000 3.785000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870000 62.100000 4.190000 62.420000 ;
      LAYER met4 ;
        RECT 3.870000 62.100000 4.190000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870000 62.510000 4.190000 62.830000 ;
      LAYER met4 ;
        RECT 3.870000 62.510000 4.190000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870000 62.920000 4.190000 63.240000 ;
      LAYER met4 ;
        RECT 3.870000 62.920000 4.190000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870000 63.330000 4.190000 63.650000 ;
      LAYER met4 ;
        RECT 3.870000 63.330000 4.190000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870000 63.740000 4.190000 64.060000 ;
      LAYER met4 ;
        RECT 3.870000 63.740000 4.190000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870000 64.150000 4.190000 64.470000 ;
      LAYER met4 ;
        RECT 3.870000 64.150000 4.190000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870000 64.560000 4.190000 64.880000 ;
      LAYER met4 ;
        RECT 3.870000 64.560000 4.190000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870000 64.970000 4.190000 65.290000 ;
      LAYER met4 ;
        RECT 3.870000 64.970000 4.190000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870000 65.380000 4.190000 65.700000 ;
      LAYER met4 ;
        RECT 3.870000 65.380000 4.190000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870000 65.790000 4.190000 66.110000 ;
      LAYER met4 ;
        RECT 3.870000 65.790000 4.190000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870000 66.200000 4.190000 66.520000 ;
      LAYER met4 ;
        RECT 3.870000 66.200000 4.190000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275000 62.100000 4.595000 62.420000 ;
      LAYER met4 ;
        RECT 4.275000 62.100000 4.595000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275000 62.510000 4.595000 62.830000 ;
      LAYER met4 ;
        RECT 4.275000 62.510000 4.595000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275000 62.920000 4.595000 63.240000 ;
      LAYER met4 ;
        RECT 4.275000 62.920000 4.595000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275000 63.330000 4.595000 63.650000 ;
      LAYER met4 ;
        RECT 4.275000 63.330000 4.595000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275000 63.740000 4.595000 64.060000 ;
      LAYER met4 ;
        RECT 4.275000 63.740000 4.595000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275000 64.150000 4.595000 64.470000 ;
      LAYER met4 ;
        RECT 4.275000 64.150000 4.595000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275000 64.560000 4.595000 64.880000 ;
      LAYER met4 ;
        RECT 4.275000 64.560000 4.595000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275000 64.970000 4.595000 65.290000 ;
      LAYER met4 ;
        RECT 4.275000 64.970000 4.595000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275000 65.380000 4.595000 65.700000 ;
      LAYER met4 ;
        RECT 4.275000 65.380000 4.595000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275000 65.790000 4.595000 66.110000 ;
      LAYER met4 ;
        RECT 4.275000 65.790000 4.595000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275000 66.200000 4.595000 66.520000 ;
      LAYER met4 ;
        RECT 4.275000 66.200000 4.595000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680000 62.100000 5.000000 62.420000 ;
      LAYER met4 ;
        RECT 4.680000 62.100000 5.000000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680000 62.510000 5.000000 62.830000 ;
      LAYER met4 ;
        RECT 4.680000 62.510000 5.000000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680000 62.920000 5.000000 63.240000 ;
      LAYER met4 ;
        RECT 4.680000 62.920000 5.000000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680000 63.330000 5.000000 63.650000 ;
      LAYER met4 ;
        RECT 4.680000 63.330000 5.000000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680000 63.740000 5.000000 64.060000 ;
      LAYER met4 ;
        RECT 4.680000 63.740000 5.000000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680000 64.150000 5.000000 64.470000 ;
      LAYER met4 ;
        RECT 4.680000 64.150000 5.000000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680000 64.560000 5.000000 64.880000 ;
      LAYER met4 ;
        RECT 4.680000 64.560000 5.000000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680000 64.970000 5.000000 65.290000 ;
      LAYER met4 ;
        RECT 4.680000 64.970000 5.000000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680000 65.380000 5.000000 65.700000 ;
      LAYER met4 ;
        RECT 4.680000 65.380000 5.000000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680000 65.790000 5.000000 66.110000 ;
      LAYER met4 ;
        RECT 4.680000 65.790000 5.000000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680000 66.200000 5.000000 66.520000 ;
      LAYER met4 ;
        RECT 4.680000 66.200000 5.000000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 62.100000 5.405000 62.420000 ;
      LAYER met4 ;
        RECT 5.085000 62.100000 5.405000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 62.510000 5.405000 62.830000 ;
      LAYER met4 ;
        RECT 5.085000 62.510000 5.405000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 62.920000 5.405000 63.240000 ;
      LAYER met4 ;
        RECT 5.085000 62.920000 5.405000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 63.330000 5.405000 63.650000 ;
      LAYER met4 ;
        RECT 5.085000 63.330000 5.405000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 63.740000 5.405000 64.060000 ;
      LAYER met4 ;
        RECT 5.085000 63.740000 5.405000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 64.150000 5.405000 64.470000 ;
      LAYER met4 ;
        RECT 5.085000 64.150000 5.405000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 64.560000 5.405000 64.880000 ;
      LAYER met4 ;
        RECT 5.085000 64.560000 5.405000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 64.970000 5.405000 65.290000 ;
      LAYER met4 ;
        RECT 5.085000 64.970000 5.405000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 65.380000 5.405000 65.700000 ;
      LAYER met4 ;
        RECT 5.085000 65.380000 5.405000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 65.790000 5.405000 66.110000 ;
      LAYER met4 ;
        RECT 5.085000 65.790000 5.405000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085000 66.200000 5.405000 66.520000 ;
      LAYER met4 ;
        RECT 5.085000 66.200000 5.405000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490000 62.100000 5.810000 62.420000 ;
      LAYER met4 ;
        RECT 5.490000 62.100000 5.810000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490000 62.510000 5.810000 62.830000 ;
      LAYER met4 ;
        RECT 5.490000 62.510000 5.810000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490000 62.920000 5.810000 63.240000 ;
      LAYER met4 ;
        RECT 5.490000 62.920000 5.810000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490000 63.330000 5.810000 63.650000 ;
      LAYER met4 ;
        RECT 5.490000 63.330000 5.810000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490000 63.740000 5.810000 64.060000 ;
      LAYER met4 ;
        RECT 5.490000 63.740000 5.810000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490000 64.150000 5.810000 64.470000 ;
      LAYER met4 ;
        RECT 5.490000 64.150000 5.810000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490000 64.560000 5.810000 64.880000 ;
      LAYER met4 ;
        RECT 5.490000 64.560000 5.810000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490000 64.970000 5.810000 65.290000 ;
      LAYER met4 ;
        RECT 5.490000 64.970000 5.810000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490000 65.380000 5.810000 65.700000 ;
      LAYER met4 ;
        RECT 5.490000 65.380000 5.810000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490000 65.790000 5.810000 66.110000 ;
      LAYER met4 ;
        RECT 5.490000 65.790000 5.810000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490000 66.200000 5.810000 66.520000 ;
      LAYER met4 ;
        RECT 5.490000 66.200000 5.810000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895000 62.100000 6.215000 62.420000 ;
      LAYER met4 ;
        RECT 5.895000 62.100000 6.215000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895000 62.510000 6.215000 62.830000 ;
      LAYER met4 ;
        RECT 5.895000 62.510000 6.215000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895000 62.920000 6.215000 63.240000 ;
      LAYER met4 ;
        RECT 5.895000 62.920000 6.215000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895000 63.330000 6.215000 63.650000 ;
      LAYER met4 ;
        RECT 5.895000 63.330000 6.215000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895000 63.740000 6.215000 64.060000 ;
      LAYER met4 ;
        RECT 5.895000 63.740000 6.215000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895000 64.150000 6.215000 64.470000 ;
      LAYER met4 ;
        RECT 5.895000 64.150000 6.215000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895000 64.560000 6.215000 64.880000 ;
      LAYER met4 ;
        RECT 5.895000 64.560000 6.215000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895000 64.970000 6.215000 65.290000 ;
      LAYER met4 ;
        RECT 5.895000 64.970000 6.215000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895000 65.380000 6.215000 65.700000 ;
      LAYER met4 ;
        RECT 5.895000 65.380000 6.215000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895000 65.790000 6.215000 66.110000 ;
      LAYER met4 ;
        RECT 5.895000 65.790000 6.215000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895000 66.200000 6.215000 66.520000 ;
      LAYER met4 ;
        RECT 5.895000 66.200000 6.215000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 62.100000 51.105000 62.420000 ;
      LAYER met4 ;
        RECT 50.785000 62.100000 51.105000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 62.510000 51.105000 62.830000 ;
      LAYER met4 ;
        RECT 50.785000 62.510000 51.105000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 62.920000 51.105000 63.240000 ;
      LAYER met4 ;
        RECT 50.785000 62.920000 51.105000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 63.330000 51.105000 63.650000 ;
      LAYER met4 ;
        RECT 50.785000 63.330000 51.105000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 63.740000 51.105000 64.060000 ;
      LAYER met4 ;
        RECT 50.785000 63.740000 51.105000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 64.150000 51.105000 64.470000 ;
      LAYER met4 ;
        RECT 50.785000 64.150000 51.105000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 64.560000 51.105000 64.880000 ;
      LAYER met4 ;
        RECT 50.785000 64.560000 51.105000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 64.970000 51.105000 65.290000 ;
      LAYER met4 ;
        RECT 50.785000 64.970000 51.105000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 65.380000 51.105000 65.700000 ;
      LAYER met4 ;
        RECT 50.785000 65.380000 51.105000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 65.790000 51.105000 66.110000 ;
      LAYER met4 ;
        RECT 50.785000 65.790000 51.105000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 66.200000 51.105000 66.520000 ;
      LAYER met4 ;
        RECT 50.785000 66.200000 51.105000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.190000 62.100000 51.510000 62.420000 ;
      LAYER met4 ;
        RECT 51.190000 62.100000 51.510000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.190000 62.510000 51.510000 62.830000 ;
      LAYER met4 ;
        RECT 51.190000 62.510000 51.510000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.190000 62.920000 51.510000 63.240000 ;
      LAYER met4 ;
        RECT 51.190000 62.920000 51.510000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.190000 63.330000 51.510000 63.650000 ;
      LAYER met4 ;
        RECT 51.190000 63.330000 51.510000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.190000 63.740000 51.510000 64.060000 ;
      LAYER met4 ;
        RECT 51.190000 63.740000 51.510000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.190000 64.150000 51.510000 64.470000 ;
      LAYER met4 ;
        RECT 51.190000 64.150000 51.510000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.190000 64.560000 51.510000 64.880000 ;
      LAYER met4 ;
        RECT 51.190000 64.560000 51.510000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.190000 64.970000 51.510000 65.290000 ;
      LAYER met4 ;
        RECT 51.190000 64.970000 51.510000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.190000 65.380000 51.510000 65.700000 ;
      LAYER met4 ;
        RECT 51.190000 65.380000 51.510000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.190000 65.790000 51.510000 66.110000 ;
      LAYER met4 ;
        RECT 51.190000 65.790000 51.510000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.190000 66.200000 51.510000 66.520000 ;
      LAYER met4 ;
        RECT 51.190000 66.200000 51.510000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.595000 62.100000 51.915000 62.420000 ;
      LAYER met4 ;
        RECT 51.595000 62.100000 51.915000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.595000 62.510000 51.915000 62.830000 ;
      LAYER met4 ;
        RECT 51.595000 62.510000 51.915000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.595000 62.920000 51.915000 63.240000 ;
      LAYER met4 ;
        RECT 51.595000 62.920000 51.915000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.595000 63.330000 51.915000 63.650000 ;
      LAYER met4 ;
        RECT 51.595000 63.330000 51.915000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.595000 63.740000 51.915000 64.060000 ;
      LAYER met4 ;
        RECT 51.595000 63.740000 51.915000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.595000 64.150000 51.915000 64.470000 ;
      LAYER met4 ;
        RECT 51.595000 64.150000 51.915000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.595000 64.560000 51.915000 64.880000 ;
      LAYER met4 ;
        RECT 51.595000 64.560000 51.915000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.595000 64.970000 51.915000 65.290000 ;
      LAYER met4 ;
        RECT 51.595000 64.970000 51.915000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.595000 65.380000 51.915000 65.700000 ;
      LAYER met4 ;
        RECT 51.595000 65.380000 51.915000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.595000 65.790000 51.915000 66.110000 ;
      LAYER met4 ;
        RECT 51.595000 65.790000 51.915000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.595000 66.200000 51.915000 66.520000 ;
      LAYER met4 ;
        RECT 51.595000 66.200000 51.915000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.000000 62.100000 52.320000 62.420000 ;
      LAYER met4 ;
        RECT 52.000000 62.100000 52.320000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.000000 62.510000 52.320000 62.830000 ;
      LAYER met4 ;
        RECT 52.000000 62.510000 52.320000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.000000 62.920000 52.320000 63.240000 ;
      LAYER met4 ;
        RECT 52.000000 62.920000 52.320000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.000000 63.330000 52.320000 63.650000 ;
      LAYER met4 ;
        RECT 52.000000 63.330000 52.320000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.000000 63.740000 52.320000 64.060000 ;
      LAYER met4 ;
        RECT 52.000000 63.740000 52.320000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.000000 64.150000 52.320000 64.470000 ;
      LAYER met4 ;
        RECT 52.000000 64.150000 52.320000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.000000 64.560000 52.320000 64.880000 ;
      LAYER met4 ;
        RECT 52.000000 64.560000 52.320000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.000000 64.970000 52.320000 65.290000 ;
      LAYER met4 ;
        RECT 52.000000 64.970000 52.320000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.000000 65.380000 52.320000 65.700000 ;
      LAYER met4 ;
        RECT 52.000000 65.380000 52.320000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.000000 65.790000 52.320000 66.110000 ;
      LAYER met4 ;
        RECT 52.000000 65.790000 52.320000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.000000 66.200000 52.320000 66.520000 ;
      LAYER met4 ;
        RECT 52.000000 66.200000 52.320000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 62.100000 52.725000 62.420000 ;
      LAYER met4 ;
        RECT 52.405000 62.100000 52.725000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 62.510000 52.725000 62.830000 ;
      LAYER met4 ;
        RECT 52.405000 62.510000 52.725000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 62.920000 52.725000 63.240000 ;
      LAYER met4 ;
        RECT 52.405000 62.920000 52.725000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 63.330000 52.725000 63.650000 ;
      LAYER met4 ;
        RECT 52.405000 63.330000 52.725000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 63.740000 52.725000 64.060000 ;
      LAYER met4 ;
        RECT 52.405000 63.740000 52.725000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 64.150000 52.725000 64.470000 ;
      LAYER met4 ;
        RECT 52.405000 64.150000 52.725000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 64.560000 52.725000 64.880000 ;
      LAYER met4 ;
        RECT 52.405000 64.560000 52.725000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 64.970000 52.725000 65.290000 ;
      LAYER met4 ;
        RECT 52.405000 64.970000 52.725000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 65.380000 52.725000 65.700000 ;
      LAYER met4 ;
        RECT 52.405000 65.380000 52.725000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 65.790000 52.725000 66.110000 ;
      LAYER met4 ;
        RECT 52.405000 65.790000 52.725000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405000 66.200000 52.725000 66.520000 ;
      LAYER met4 ;
        RECT 52.405000 66.200000 52.725000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.810000 62.100000 53.130000 62.420000 ;
      LAYER met4 ;
        RECT 52.810000 62.100000 53.130000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.810000 62.510000 53.130000 62.830000 ;
      LAYER met4 ;
        RECT 52.810000 62.510000 53.130000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.810000 62.920000 53.130000 63.240000 ;
      LAYER met4 ;
        RECT 52.810000 62.920000 53.130000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.810000 63.330000 53.130000 63.650000 ;
      LAYER met4 ;
        RECT 52.810000 63.330000 53.130000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.810000 63.740000 53.130000 64.060000 ;
      LAYER met4 ;
        RECT 52.810000 63.740000 53.130000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.810000 64.150000 53.130000 64.470000 ;
      LAYER met4 ;
        RECT 52.810000 64.150000 53.130000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.810000 64.560000 53.130000 64.880000 ;
      LAYER met4 ;
        RECT 52.810000 64.560000 53.130000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.810000 64.970000 53.130000 65.290000 ;
      LAYER met4 ;
        RECT 52.810000 64.970000 53.130000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.810000 65.380000 53.130000 65.700000 ;
      LAYER met4 ;
        RECT 52.810000 65.380000 53.130000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.810000 65.790000 53.130000 66.110000 ;
      LAYER met4 ;
        RECT 52.810000 65.790000 53.130000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.810000 66.200000 53.130000 66.520000 ;
      LAYER met4 ;
        RECT 52.810000 66.200000 53.130000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.215000 62.100000 53.535000 62.420000 ;
      LAYER met4 ;
        RECT 53.215000 62.100000 53.535000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.215000 62.510000 53.535000 62.830000 ;
      LAYER met4 ;
        RECT 53.215000 62.510000 53.535000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.215000 62.920000 53.535000 63.240000 ;
      LAYER met4 ;
        RECT 53.215000 62.920000 53.535000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.215000 63.330000 53.535000 63.650000 ;
      LAYER met4 ;
        RECT 53.215000 63.330000 53.535000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.215000 63.740000 53.535000 64.060000 ;
      LAYER met4 ;
        RECT 53.215000 63.740000 53.535000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.215000 64.150000 53.535000 64.470000 ;
      LAYER met4 ;
        RECT 53.215000 64.150000 53.535000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.215000 64.560000 53.535000 64.880000 ;
      LAYER met4 ;
        RECT 53.215000 64.560000 53.535000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.215000 64.970000 53.535000 65.290000 ;
      LAYER met4 ;
        RECT 53.215000 64.970000 53.535000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.215000 65.380000 53.535000 65.700000 ;
      LAYER met4 ;
        RECT 53.215000 65.380000 53.535000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.215000 65.790000 53.535000 66.110000 ;
      LAYER met4 ;
        RECT 53.215000 65.790000 53.535000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.215000 66.200000 53.535000 66.520000 ;
      LAYER met4 ;
        RECT 53.215000 66.200000 53.535000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.620000 62.100000 53.940000 62.420000 ;
      LAYER met4 ;
        RECT 53.620000 62.100000 53.940000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.620000 62.510000 53.940000 62.830000 ;
      LAYER met4 ;
        RECT 53.620000 62.510000 53.940000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.620000 62.920000 53.940000 63.240000 ;
      LAYER met4 ;
        RECT 53.620000 62.920000 53.940000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.620000 63.330000 53.940000 63.650000 ;
      LAYER met4 ;
        RECT 53.620000 63.330000 53.940000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.620000 63.740000 53.940000 64.060000 ;
      LAYER met4 ;
        RECT 53.620000 63.740000 53.940000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.620000 64.150000 53.940000 64.470000 ;
      LAYER met4 ;
        RECT 53.620000 64.150000 53.940000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.620000 64.560000 53.940000 64.880000 ;
      LAYER met4 ;
        RECT 53.620000 64.560000 53.940000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.620000 64.970000 53.940000 65.290000 ;
      LAYER met4 ;
        RECT 53.620000 64.970000 53.940000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.620000 65.380000 53.940000 65.700000 ;
      LAYER met4 ;
        RECT 53.620000 65.380000 53.940000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.620000 65.790000 53.940000 66.110000 ;
      LAYER met4 ;
        RECT 53.620000 65.790000 53.940000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.620000 66.200000 53.940000 66.520000 ;
      LAYER met4 ;
        RECT 53.620000 66.200000 53.940000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.025000 62.100000 54.345000 62.420000 ;
      LAYER met4 ;
        RECT 54.025000 62.100000 54.345000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.025000 62.510000 54.345000 62.830000 ;
      LAYER met4 ;
        RECT 54.025000 62.510000 54.345000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.025000 62.920000 54.345000 63.240000 ;
      LAYER met4 ;
        RECT 54.025000 62.920000 54.345000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.025000 63.330000 54.345000 63.650000 ;
      LAYER met4 ;
        RECT 54.025000 63.330000 54.345000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.025000 63.740000 54.345000 64.060000 ;
      LAYER met4 ;
        RECT 54.025000 63.740000 54.345000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.025000 64.150000 54.345000 64.470000 ;
      LAYER met4 ;
        RECT 54.025000 64.150000 54.345000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.025000 64.560000 54.345000 64.880000 ;
      LAYER met4 ;
        RECT 54.025000 64.560000 54.345000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.025000 64.970000 54.345000 65.290000 ;
      LAYER met4 ;
        RECT 54.025000 64.970000 54.345000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.025000 65.380000 54.345000 65.700000 ;
      LAYER met4 ;
        RECT 54.025000 65.380000 54.345000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.025000 65.790000 54.345000 66.110000 ;
      LAYER met4 ;
        RECT 54.025000 65.790000 54.345000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.025000 66.200000 54.345000 66.520000 ;
      LAYER met4 ;
        RECT 54.025000 66.200000 54.345000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.430000 62.100000 54.750000 62.420000 ;
      LAYER met4 ;
        RECT 54.430000 62.100000 54.750000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.430000 62.510000 54.750000 62.830000 ;
      LAYER met4 ;
        RECT 54.430000 62.510000 54.750000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.430000 62.920000 54.750000 63.240000 ;
      LAYER met4 ;
        RECT 54.430000 62.920000 54.750000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.430000 63.330000 54.750000 63.650000 ;
      LAYER met4 ;
        RECT 54.430000 63.330000 54.750000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.430000 63.740000 54.750000 64.060000 ;
      LAYER met4 ;
        RECT 54.430000 63.740000 54.750000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.430000 64.150000 54.750000 64.470000 ;
      LAYER met4 ;
        RECT 54.430000 64.150000 54.750000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.430000 64.560000 54.750000 64.880000 ;
      LAYER met4 ;
        RECT 54.430000 64.560000 54.750000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.430000 64.970000 54.750000 65.290000 ;
      LAYER met4 ;
        RECT 54.430000 64.970000 54.750000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.430000 65.380000 54.750000 65.700000 ;
      LAYER met4 ;
        RECT 54.430000 65.380000 54.750000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.430000 65.790000 54.750000 66.110000 ;
      LAYER met4 ;
        RECT 54.430000 65.790000 54.750000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.430000 66.200000 54.750000 66.520000 ;
      LAYER met4 ;
        RECT 54.430000 66.200000 54.750000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.835000 62.100000 55.155000 62.420000 ;
      LAYER met4 ;
        RECT 54.835000 62.100000 55.155000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.835000 62.510000 55.155000 62.830000 ;
      LAYER met4 ;
        RECT 54.835000 62.510000 55.155000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.835000 62.920000 55.155000 63.240000 ;
      LAYER met4 ;
        RECT 54.835000 62.920000 55.155000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.835000 63.330000 55.155000 63.650000 ;
      LAYER met4 ;
        RECT 54.835000 63.330000 55.155000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.835000 63.740000 55.155000 64.060000 ;
      LAYER met4 ;
        RECT 54.835000 63.740000 55.155000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.835000 64.150000 55.155000 64.470000 ;
      LAYER met4 ;
        RECT 54.835000 64.150000 55.155000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.835000 64.560000 55.155000 64.880000 ;
      LAYER met4 ;
        RECT 54.835000 64.560000 55.155000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.835000 64.970000 55.155000 65.290000 ;
      LAYER met4 ;
        RECT 54.835000 64.970000 55.155000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.835000 65.380000 55.155000 65.700000 ;
      LAYER met4 ;
        RECT 54.835000 65.380000 55.155000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.835000 65.790000 55.155000 66.110000 ;
      LAYER met4 ;
        RECT 54.835000 65.790000 55.155000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.835000 66.200000 55.155000 66.520000 ;
      LAYER met4 ;
        RECT 54.835000 66.200000 55.155000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.240000 62.100000 55.560000 62.420000 ;
      LAYER met4 ;
        RECT 55.240000 62.100000 55.560000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.240000 62.510000 55.560000 62.830000 ;
      LAYER met4 ;
        RECT 55.240000 62.510000 55.560000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.240000 62.920000 55.560000 63.240000 ;
      LAYER met4 ;
        RECT 55.240000 62.920000 55.560000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.240000 63.330000 55.560000 63.650000 ;
      LAYER met4 ;
        RECT 55.240000 63.330000 55.560000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.240000 63.740000 55.560000 64.060000 ;
      LAYER met4 ;
        RECT 55.240000 63.740000 55.560000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.240000 64.150000 55.560000 64.470000 ;
      LAYER met4 ;
        RECT 55.240000 64.150000 55.560000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.240000 64.560000 55.560000 64.880000 ;
      LAYER met4 ;
        RECT 55.240000 64.560000 55.560000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.240000 64.970000 55.560000 65.290000 ;
      LAYER met4 ;
        RECT 55.240000 64.970000 55.560000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.240000 65.380000 55.560000 65.700000 ;
      LAYER met4 ;
        RECT 55.240000 65.380000 55.560000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.240000 65.790000 55.560000 66.110000 ;
      LAYER met4 ;
        RECT 55.240000 65.790000 55.560000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.240000 66.200000 55.560000 66.520000 ;
      LAYER met4 ;
        RECT 55.240000 66.200000 55.560000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.645000 62.100000 55.965000 62.420000 ;
      LAYER met4 ;
        RECT 55.645000 62.100000 55.965000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.645000 62.510000 55.965000 62.830000 ;
      LAYER met4 ;
        RECT 55.645000 62.510000 55.965000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.645000 62.920000 55.965000 63.240000 ;
      LAYER met4 ;
        RECT 55.645000 62.920000 55.965000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.645000 63.330000 55.965000 63.650000 ;
      LAYER met4 ;
        RECT 55.645000 63.330000 55.965000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.645000 63.740000 55.965000 64.060000 ;
      LAYER met4 ;
        RECT 55.645000 63.740000 55.965000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.645000 64.150000 55.965000 64.470000 ;
      LAYER met4 ;
        RECT 55.645000 64.150000 55.965000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.645000 64.560000 55.965000 64.880000 ;
      LAYER met4 ;
        RECT 55.645000 64.560000 55.965000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.645000 64.970000 55.965000 65.290000 ;
      LAYER met4 ;
        RECT 55.645000 64.970000 55.965000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.645000 65.380000 55.965000 65.700000 ;
      LAYER met4 ;
        RECT 55.645000 65.380000 55.965000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.645000 65.790000 55.965000 66.110000 ;
      LAYER met4 ;
        RECT 55.645000 65.790000 55.965000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.645000 66.200000 55.965000 66.520000 ;
      LAYER met4 ;
        RECT 55.645000 66.200000 55.965000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.050000 62.100000 56.370000 62.420000 ;
      LAYER met4 ;
        RECT 56.050000 62.100000 56.370000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.050000 62.510000 56.370000 62.830000 ;
      LAYER met4 ;
        RECT 56.050000 62.510000 56.370000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.050000 62.920000 56.370000 63.240000 ;
      LAYER met4 ;
        RECT 56.050000 62.920000 56.370000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.050000 63.330000 56.370000 63.650000 ;
      LAYER met4 ;
        RECT 56.050000 63.330000 56.370000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.050000 63.740000 56.370000 64.060000 ;
      LAYER met4 ;
        RECT 56.050000 63.740000 56.370000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.050000 64.150000 56.370000 64.470000 ;
      LAYER met4 ;
        RECT 56.050000 64.150000 56.370000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.050000 64.560000 56.370000 64.880000 ;
      LAYER met4 ;
        RECT 56.050000 64.560000 56.370000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.050000 64.970000 56.370000 65.290000 ;
      LAYER met4 ;
        RECT 56.050000 64.970000 56.370000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.050000 65.380000 56.370000 65.700000 ;
      LAYER met4 ;
        RECT 56.050000 65.380000 56.370000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.050000 65.790000 56.370000 66.110000 ;
      LAYER met4 ;
        RECT 56.050000 65.790000 56.370000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.050000 66.200000 56.370000 66.520000 ;
      LAYER met4 ;
        RECT 56.050000 66.200000 56.370000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 62.100000 56.775000 62.420000 ;
      LAYER met4 ;
        RECT 56.455000 62.100000 56.775000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 62.510000 56.775000 62.830000 ;
      LAYER met4 ;
        RECT 56.455000 62.510000 56.775000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 62.920000 56.775000 63.240000 ;
      LAYER met4 ;
        RECT 56.455000 62.920000 56.775000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 63.330000 56.775000 63.650000 ;
      LAYER met4 ;
        RECT 56.455000 63.330000 56.775000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 63.740000 56.775000 64.060000 ;
      LAYER met4 ;
        RECT 56.455000 63.740000 56.775000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 64.150000 56.775000 64.470000 ;
      LAYER met4 ;
        RECT 56.455000 64.150000 56.775000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 64.560000 56.775000 64.880000 ;
      LAYER met4 ;
        RECT 56.455000 64.560000 56.775000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 64.970000 56.775000 65.290000 ;
      LAYER met4 ;
        RECT 56.455000 64.970000 56.775000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 65.380000 56.775000 65.700000 ;
      LAYER met4 ;
        RECT 56.455000 65.380000 56.775000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 65.790000 56.775000 66.110000 ;
      LAYER met4 ;
        RECT 56.455000 65.790000 56.775000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.455000 66.200000 56.775000 66.520000 ;
      LAYER met4 ;
        RECT 56.455000 66.200000 56.775000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.860000 62.100000 57.180000 62.420000 ;
      LAYER met4 ;
        RECT 56.860000 62.100000 57.180000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.860000 62.510000 57.180000 62.830000 ;
      LAYER met4 ;
        RECT 56.860000 62.510000 57.180000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.860000 62.920000 57.180000 63.240000 ;
      LAYER met4 ;
        RECT 56.860000 62.920000 57.180000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.860000 63.330000 57.180000 63.650000 ;
      LAYER met4 ;
        RECT 56.860000 63.330000 57.180000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.860000 63.740000 57.180000 64.060000 ;
      LAYER met4 ;
        RECT 56.860000 63.740000 57.180000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.860000 64.150000 57.180000 64.470000 ;
      LAYER met4 ;
        RECT 56.860000 64.150000 57.180000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.860000 64.560000 57.180000 64.880000 ;
      LAYER met4 ;
        RECT 56.860000 64.560000 57.180000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.860000 64.970000 57.180000 65.290000 ;
      LAYER met4 ;
        RECT 56.860000 64.970000 57.180000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.860000 65.380000 57.180000 65.700000 ;
      LAYER met4 ;
        RECT 56.860000 65.380000 57.180000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.860000 65.790000 57.180000 66.110000 ;
      LAYER met4 ;
        RECT 56.860000 65.790000 57.180000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.860000 66.200000 57.180000 66.520000 ;
      LAYER met4 ;
        RECT 56.860000 66.200000 57.180000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.265000 62.100000 57.585000 62.420000 ;
      LAYER met4 ;
        RECT 57.265000 62.100000 57.585000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.265000 62.510000 57.585000 62.830000 ;
      LAYER met4 ;
        RECT 57.265000 62.510000 57.585000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.265000 62.920000 57.585000 63.240000 ;
      LAYER met4 ;
        RECT 57.265000 62.920000 57.585000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.265000 63.330000 57.585000 63.650000 ;
      LAYER met4 ;
        RECT 57.265000 63.330000 57.585000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.265000 63.740000 57.585000 64.060000 ;
      LAYER met4 ;
        RECT 57.265000 63.740000 57.585000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.265000 64.150000 57.585000 64.470000 ;
      LAYER met4 ;
        RECT 57.265000 64.150000 57.585000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.265000 64.560000 57.585000 64.880000 ;
      LAYER met4 ;
        RECT 57.265000 64.560000 57.585000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.265000 64.970000 57.585000 65.290000 ;
      LAYER met4 ;
        RECT 57.265000 64.970000 57.585000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.265000 65.380000 57.585000 65.700000 ;
      LAYER met4 ;
        RECT 57.265000 65.380000 57.585000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.265000 65.790000 57.585000 66.110000 ;
      LAYER met4 ;
        RECT 57.265000 65.790000 57.585000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.265000 66.200000 57.585000 66.520000 ;
      LAYER met4 ;
        RECT 57.265000 66.200000 57.585000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.670000 62.100000 57.990000 62.420000 ;
      LAYER met4 ;
        RECT 57.670000 62.100000 57.990000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.670000 62.510000 57.990000 62.830000 ;
      LAYER met4 ;
        RECT 57.670000 62.510000 57.990000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.670000 62.920000 57.990000 63.240000 ;
      LAYER met4 ;
        RECT 57.670000 62.920000 57.990000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.670000 63.330000 57.990000 63.650000 ;
      LAYER met4 ;
        RECT 57.670000 63.330000 57.990000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.670000 63.740000 57.990000 64.060000 ;
      LAYER met4 ;
        RECT 57.670000 63.740000 57.990000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.670000 64.150000 57.990000 64.470000 ;
      LAYER met4 ;
        RECT 57.670000 64.150000 57.990000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.670000 64.560000 57.990000 64.880000 ;
      LAYER met4 ;
        RECT 57.670000 64.560000 57.990000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.670000 64.970000 57.990000 65.290000 ;
      LAYER met4 ;
        RECT 57.670000 64.970000 57.990000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.670000 65.380000 57.990000 65.700000 ;
      LAYER met4 ;
        RECT 57.670000 65.380000 57.990000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.670000 65.790000 57.990000 66.110000 ;
      LAYER met4 ;
        RECT 57.670000 65.790000 57.990000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.670000 66.200000 57.990000 66.520000 ;
      LAYER met4 ;
        RECT 57.670000 66.200000 57.990000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.075000 62.100000 58.395000 62.420000 ;
      LAYER met4 ;
        RECT 58.075000 62.100000 58.395000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.075000 62.510000 58.395000 62.830000 ;
      LAYER met4 ;
        RECT 58.075000 62.510000 58.395000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.075000 62.920000 58.395000 63.240000 ;
      LAYER met4 ;
        RECT 58.075000 62.920000 58.395000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.075000 63.330000 58.395000 63.650000 ;
      LAYER met4 ;
        RECT 58.075000 63.330000 58.395000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.075000 63.740000 58.395000 64.060000 ;
      LAYER met4 ;
        RECT 58.075000 63.740000 58.395000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.075000 64.150000 58.395000 64.470000 ;
      LAYER met4 ;
        RECT 58.075000 64.150000 58.395000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.075000 64.560000 58.395000 64.880000 ;
      LAYER met4 ;
        RECT 58.075000 64.560000 58.395000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.075000 64.970000 58.395000 65.290000 ;
      LAYER met4 ;
        RECT 58.075000 64.970000 58.395000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.075000 65.380000 58.395000 65.700000 ;
      LAYER met4 ;
        RECT 58.075000 65.380000 58.395000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.075000 65.790000 58.395000 66.110000 ;
      LAYER met4 ;
        RECT 58.075000 65.790000 58.395000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.075000 66.200000 58.395000 66.520000 ;
      LAYER met4 ;
        RECT 58.075000 66.200000 58.395000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 62.100000 58.800000 62.420000 ;
      LAYER met4 ;
        RECT 58.480000 62.100000 58.800000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 62.510000 58.800000 62.830000 ;
      LAYER met4 ;
        RECT 58.480000 62.510000 58.800000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 62.920000 58.800000 63.240000 ;
      LAYER met4 ;
        RECT 58.480000 62.920000 58.800000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 63.330000 58.800000 63.650000 ;
      LAYER met4 ;
        RECT 58.480000 63.330000 58.800000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 63.740000 58.800000 64.060000 ;
      LAYER met4 ;
        RECT 58.480000 63.740000 58.800000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 64.150000 58.800000 64.470000 ;
      LAYER met4 ;
        RECT 58.480000 64.150000 58.800000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 64.560000 58.800000 64.880000 ;
      LAYER met4 ;
        RECT 58.480000 64.560000 58.800000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 64.970000 58.800000 65.290000 ;
      LAYER met4 ;
        RECT 58.480000 64.970000 58.800000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 65.380000 58.800000 65.700000 ;
      LAYER met4 ;
        RECT 58.480000 65.380000 58.800000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 65.790000 58.800000 66.110000 ;
      LAYER met4 ;
        RECT 58.480000 65.790000 58.800000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480000 66.200000 58.800000 66.520000 ;
      LAYER met4 ;
        RECT 58.480000 66.200000 58.800000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.885000 62.100000 59.205000 62.420000 ;
      LAYER met4 ;
        RECT 58.885000 62.100000 59.205000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.885000 62.510000 59.205000 62.830000 ;
      LAYER met4 ;
        RECT 58.885000 62.510000 59.205000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.885000 62.920000 59.205000 63.240000 ;
      LAYER met4 ;
        RECT 58.885000 62.920000 59.205000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.885000 63.330000 59.205000 63.650000 ;
      LAYER met4 ;
        RECT 58.885000 63.330000 59.205000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.885000 63.740000 59.205000 64.060000 ;
      LAYER met4 ;
        RECT 58.885000 63.740000 59.205000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.885000 64.150000 59.205000 64.470000 ;
      LAYER met4 ;
        RECT 58.885000 64.150000 59.205000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.885000 64.560000 59.205000 64.880000 ;
      LAYER met4 ;
        RECT 58.885000 64.560000 59.205000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.885000 64.970000 59.205000 65.290000 ;
      LAYER met4 ;
        RECT 58.885000 64.970000 59.205000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.885000 65.380000 59.205000 65.700000 ;
      LAYER met4 ;
        RECT 58.885000 65.380000 59.205000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.885000 65.790000 59.205000 66.110000 ;
      LAYER met4 ;
        RECT 58.885000 65.790000 59.205000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.885000 66.200000 59.205000 66.520000 ;
      LAYER met4 ;
        RECT 58.885000 66.200000 59.205000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.290000 62.100000 59.610000 62.420000 ;
      LAYER met4 ;
        RECT 59.290000 62.100000 59.610000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.290000 62.510000 59.610000 62.830000 ;
      LAYER met4 ;
        RECT 59.290000 62.510000 59.610000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.290000 62.920000 59.610000 63.240000 ;
      LAYER met4 ;
        RECT 59.290000 62.920000 59.610000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.290000 63.330000 59.610000 63.650000 ;
      LAYER met4 ;
        RECT 59.290000 63.330000 59.610000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.290000 63.740000 59.610000 64.060000 ;
      LAYER met4 ;
        RECT 59.290000 63.740000 59.610000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.290000 64.150000 59.610000 64.470000 ;
      LAYER met4 ;
        RECT 59.290000 64.150000 59.610000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.290000 64.560000 59.610000 64.880000 ;
      LAYER met4 ;
        RECT 59.290000 64.560000 59.610000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.290000 64.970000 59.610000 65.290000 ;
      LAYER met4 ;
        RECT 59.290000 64.970000 59.610000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.290000 65.380000 59.610000 65.700000 ;
      LAYER met4 ;
        RECT 59.290000 65.380000 59.610000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.290000 65.790000 59.610000 66.110000 ;
      LAYER met4 ;
        RECT 59.290000 65.790000 59.610000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.290000 66.200000 59.610000 66.520000 ;
      LAYER met4 ;
        RECT 59.290000 66.200000 59.610000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.695000 62.100000 60.015000 62.420000 ;
      LAYER met4 ;
        RECT 59.695000 62.100000 60.015000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.695000 62.510000 60.015000 62.830000 ;
      LAYER met4 ;
        RECT 59.695000 62.510000 60.015000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.695000 62.920000 60.015000 63.240000 ;
      LAYER met4 ;
        RECT 59.695000 62.920000 60.015000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.695000 63.330000 60.015000 63.650000 ;
      LAYER met4 ;
        RECT 59.695000 63.330000 60.015000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.695000 63.740000 60.015000 64.060000 ;
      LAYER met4 ;
        RECT 59.695000 63.740000 60.015000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.695000 64.150000 60.015000 64.470000 ;
      LAYER met4 ;
        RECT 59.695000 64.150000 60.015000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.695000 64.560000 60.015000 64.880000 ;
      LAYER met4 ;
        RECT 59.695000 64.560000 60.015000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.695000 64.970000 60.015000 65.290000 ;
      LAYER met4 ;
        RECT 59.695000 64.970000 60.015000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.695000 65.380000 60.015000 65.700000 ;
      LAYER met4 ;
        RECT 59.695000 65.380000 60.015000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.695000 65.790000 60.015000 66.110000 ;
      LAYER met4 ;
        RECT 59.695000 65.790000 60.015000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.695000 66.200000 60.015000 66.520000 ;
      LAYER met4 ;
        RECT 59.695000 66.200000 60.015000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300000 62.100000 6.620000 62.420000 ;
      LAYER met4 ;
        RECT 6.300000 62.100000 6.620000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300000 62.510000 6.620000 62.830000 ;
      LAYER met4 ;
        RECT 6.300000 62.510000 6.620000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300000 62.920000 6.620000 63.240000 ;
      LAYER met4 ;
        RECT 6.300000 62.920000 6.620000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300000 63.330000 6.620000 63.650000 ;
      LAYER met4 ;
        RECT 6.300000 63.330000 6.620000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300000 63.740000 6.620000 64.060000 ;
      LAYER met4 ;
        RECT 6.300000 63.740000 6.620000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300000 64.150000 6.620000 64.470000 ;
      LAYER met4 ;
        RECT 6.300000 64.150000 6.620000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300000 64.560000 6.620000 64.880000 ;
      LAYER met4 ;
        RECT 6.300000 64.560000 6.620000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300000 64.970000 6.620000 65.290000 ;
      LAYER met4 ;
        RECT 6.300000 64.970000 6.620000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300000 65.380000 6.620000 65.700000 ;
      LAYER met4 ;
        RECT 6.300000 65.380000 6.620000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300000 65.790000 6.620000 66.110000 ;
      LAYER met4 ;
        RECT 6.300000 65.790000 6.620000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300000 66.200000 6.620000 66.520000 ;
      LAYER met4 ;
        RECT 6.300000 66.200000 6.620000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705000 62.100000 7.025000 62.420000 ;
      LAYER met4 ;
        RECT 6.705000 62.100000 7.025000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705000 62.510000 7.025000 62.830000 ;
      LAYER met4 ;
        RECT 6.705000 62.510000 7.025000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705000 62.920000 7.025000 63.240000 ;
      LAYER met4 ;
        RECT 6.705000 62.920000 7.025000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705000 63.330000 7.025000 63.650000 ;
      LAYER met4 ;
        RECT 6.705000 63.330000 7.025000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705000 63.740000 7.025000 64.060000 ;
      LAYER met4 ;
        RECT 6.705000 63.740000 7.025000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705000 64.150000 7.025000 64.470000 ;
      LAYER met4 ;
        RECT 6.705000 64.150000 7.025000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705000 64.560000 7.025000 64.880000 ;
      LAYER met4 ;
        RECT 6.705000 64.560000 7.025000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705000 64.970000 7.025000 65.290000 ;
      LAYER met4 ;
        RECT 6.705000 64.970000 7.025000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705000 65.380000 7.025000 65.700000 ;
      LAYER met4 ;
        RECT 6.705000 65.380000 7.025000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705000 65.790000 7.025000 66.110000 ;
      LAYER met4 ;
        RECT 6.705000 65.790000 7.025000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705000 66.200000 7.025000 66.520000 ;
      LAYER met4 ;
        RECT 6.705000 66.200000 7.025000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.100000 62.100000 60.420000 62.420000 ;
      LAYER met4 ;
        RECT 60.100000 62.100000 60.420000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.100000 62.510000 60.420000 62.830000 ;
      LAYER met4 ;
        RECT 60.100000 62.510000 60.420000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.100000 62.920000 60.420000 63.240000 ;
      LAYER met4 ;
        RECT 60.100000 62.920000 60.420000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.100000 63.330000 60.420000 63.650000 ;
      LAYER met4 ;
        RECT 60.100000 63.330000 60.420000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.100000 63.740000 60.420000 64.060000 ;
      LAYER met4 ;
        RECT 60.100000 63.740000 60.420000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.100000 64.150000 60.420000 64.470000 ;
      LAYER met4 ;
        RECT 60.100000 64.150000 60.420000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.100000 64.560000 60.420000 64.880000 ;
      LAYER met4 ;
        RECT 60.100000 64.560000 60.420000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.100000 64.970000 60.420000 65.290000 ;
      LAYER met4 ;
        RECT 60.100000 64.970000 60.420000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.100000 65.380000 60.420000 65.700000 ;
      LAYER met4 ;
        RECT 60.100000 65.380000 60.420000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.100000 65.790000 60.420000 66.110000 ;
      LAYER met4 ;
        RECT 60.100000 65.790000 60.420000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.100000 66.200000 60.420000 66.520000 ;
      LAYER met4 ;
        RECT 60.100000 66.200000 60.420000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 62.100000 60.825000 62.420000 ;
      LAYER met4 ;
        RECT 60.505000 62.100000 60.825000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 62.510000 60.825000 62.830000 ;
      LAYER met4 ;
        RECT 60.505000 62.510000 60.825000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 62.920000 60.825000 63.240000 ;
      LAYER met4 ;
        RECT 60.505000 62.920000 60.825000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 63.330000 60.825000 63.650000 ;
      LAYER met4 ;
        RECT 60.505000 63.330000 60.825000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 63.740000 60.825000 64.060000 ;
      LAYER met4 ;
        RECT 60.505000 63.740000 60.825000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 64.150000 60.825000 64.470000 ;
      LAYER met4 ;
        RECT 60.505000 64.150000 60.825000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 64.560000 60.825000 64.880000 ;
      LAYER met4 ;
        RECT 60.505000 64.560000 60.825000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 64.970000 60.825000 65.290000 ;
      LAYER met4 ;
        RECT 60.505000 64.970000 60.825000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 65.380000 60.825000 65.700000 ;
      LAYER met4 ;
        RECT 60.505000 65.380000 60.825000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 65.790000 60.825000 66.110000 ;
      LAYER met4 ;
        RECT 60.505000 65.790000 60.825000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.505000 66.200000 60.825000 66.520000 ;
      LAYER met4 ;
        RECT 60.505000 66.200000 60.825000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.910000 62.100000 61.230000 62.420000 ;
      LAYER met4 ;
        RECT 60.910000 62.100000 61.230000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.910000 62.510000 61.230000 62.830000 ;
      LAYER met4 ;
        RECT 60.910000 62.510000 61.230000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.910000 62.920000 61.230000 63.240000 ;
      LAYER met4 ;
        RECT 60.910000 62.920000 61.230000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.910000 63.330000 61.230000 63.650000 ;
      LAYER met4 ;
        RECT 60.910000 63.330000 61.230000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.910000 63.740000 61.230000 64.060000 ;
      LAYER met4 ;
        RECT 60.910000 63.740000 61.230000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.910000 64.150000 61.230000 64.470000 ;
      LAYER met4 ;
        RECT 60.910000 64.150000 61.230000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.910000 64.560000 61.230000 64.880000 ;
      LAYER met4 ;
        RECT 60.910000 64.560000 61.230000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.910000 64.970000 61.230000 65.290000 ;
      LAYER met4 ;
        RECT 60.910000 64.970000 61.230000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.910000 65.380000 61.230000 65.700000 ;
      LAYER met4 ;
        RECT 60.910000 65.380000 61.230000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.910000 65.790000 61.230000 66.110000 ;
      LAYER met4 ;
        RECT 60.910000 65.790000 61.230000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.910000 66.200000 61.230000 66.520000 ;
      LAYER met4 ;
        RECT 60.910000 66.200000 61.230000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.315000 62.100000 61.635000 62.420000 ;
      LAYER met4 ;
        RECT 61.315000 62.100000 61.635000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.315000 62.510000 61.635000 62.830000 ;
      LAYER met4 ;
        RECT 61.315000 62.510000 61.635000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.315000 62.920000 61.635000 63.240000 ;
      LAYER met4 ;
        RECT 61.315000 62.920000 61.635000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.315000 63.330000 61.635000 63.650000 ;
      LAYER met4 ;
        RECT 61.315000 63.330000 61.635000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.315000 63.740000 61.635000 64.060000 ;
      LAYER met4 ;
        RECT 61.315000 63.740000 61.635000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.315000 64.150000 61.635000 64.470000 ;
      LAYER met4 ;
        RECT 61.315000 64.150000 61.635000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.315000 64.560000 61.635000 64.880000 ;
      LAYER met4 ;
        RECT 61.315000 64.560000 61.635000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.315000 64.970000 61.635000 65.290000 ;
      LAYER met4 ;
        RECT 61.315000 64.970000 61.635000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.315000 65.380000 61.635000 65.700000 ;
      LAYER met4 ;
        RECT 61.315000 65.380000 61.635000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.315000 65.790000 61.635000 66.110000 ;
      LAYER met4 ;
        RECT 61.315000 65.790000 61.635000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.315000 66.200000 61.635000 66.520000 ;
      LAYER met4 ;
        RECT 61.315000 66.200000 61.635000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.720000 62.100000 62.040000 62.420000 ;
      LAYER met4 ;
        RECT 61.720000 62.100000 62.040000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.720000 62.510000 62.040000 62.830000 ;
      LAYER met4 ;
        RECT 61.720000 62.510000 62.040000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.720000 62.920000 62.040000 63.240000 ;
      LAYER met4 ;
        RECT 61.720000 62.920000 62.040000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.720000 63.330000 62.040000 63.650000 ;
      LAYER met4 ;
        RECT 61.720000 63.330000 62.040000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.720000 63.740000 62.040000 64.060000 ;
      LAYER met4 ;
        RECT 61.720000 63.740000 62.040000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.720000 64.150000 62.040000 64.470000 ;
      LAYER met4 ;
        RECT 61.720000 64.150000 62.040000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.720000 64.560000 62.040000 64.880000 ;
      LAYER met4 ;
        RECT 61.720000 64.560000 62.040000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.720000 64.970000 62.040000 65.290000 ;
      LAYER met4 ;
        RECT 61.720000 64.970000 62.040000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.720000 65.380000 62.040000 65.700000 ;
      LAYER met4 ;
        RECT 61.720000 65.380000 62.040000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.720000 65.790000 62.040000 66.110000 ;
      LAYER met4 ;
        RECT 61.720000 65.790000 62.040000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.720000 66.200000 62.040000 66.520000 ;
      LAYER met4 ;
        RECT 61.720000 66.200000 62.040000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.125000 62.100000 62.445000 62.420000 ;
      LAYER met4 ;
        RECT 62.125000 62.100000 62.445000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.125000 62.510000 62.445000 62.830000 ;
      LAYER met4 ;
        RECT 62.125000 62.510000 62.445000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.125000 62.920000 62.445000 63.240000 ;
      LAYER met4 ;
        RECT 62.125000 62.920000 62.445000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.125000 63.330000 62.445000 63.650000 ;
      LAYER met4 ;
        RECT 62.125000 63.330000 62.445000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.125000 63.740000 62.445000 64.060000 ;
      LAYER met4 ;
        RECT 62.125000 63.740000 62.445000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.125000 64.150000 62.445000 64.470000 ;
      LAYER met4 ;
        RECT 62.125000 64.150000 62.445000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.125000 64.560000 62.445000 64.880000 ;
      LAYER met4 ;
        RECT 62.125000 64.560000 62.445000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.125000 64.970000 62.445000 65.290000 ;
      LAYER met4 ;
        RECT 62.125000 64.970000 62.445000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.125000 65.380000 62.445000 65.700000 ;
      LAYER met4 ;
        RECT 62.125000 65.380000 62.445000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.125000 65.790000 62.445000 66.110000 ;
      LAYER met4 ;
        RECT 62.125000 65.790000 62.445000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.125000 66.200000 62.445000 66.520000 ;
      LAYER met4 ;
        RECT 62.125000 66.200000 62.445000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.530000 62.100000 62.850000 62.420000 ;
      LAYER met4 ;
        RECT 62.530000 62.100000 62.850000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.530000 62.510000 62.850000 62.830000 ;
      LAYER met4 ;
        RECT 62.530000 62.510000 62.850000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.530000 62.920000 62.850000 63.240000 ;
      LAYER met4 ;
        RECT 62.530000 62.920000 62.850000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.530000 63.330000 62.850000 63.650000 ;
      LAYER met4 ;
        RECT 62.530000 63.330000 62.850000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.530000 63.740000 62.850000 64.060000 ;
      LAYER met4 ;
        RECT 62.530000 63.740000 62.850000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.530000 64.150000 62.850000 64.470000 ;
      LAYER met4 ;
        RECT 62.530000 64.150000 62.850000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.530000 64.560000 62.850000 64.880000 ;
      LAYER met4 ;
        RECT 62.530000 64.560000 62.850000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.530000 64.970000 62.850000 65.290000 ;
      LAYER met4 ;
        RECT 62.530000 64.970000 62.850000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.530000 65.380000 62.850000 65.700000 ;
      LAYER met4 ;
        RECT 62.530000 65.380000 62.850000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.530000 65.790000 62.850000 66.110000 ;
      LAYER met4 ;
        RECT 62.530000 65.790000 62.850000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.530000 66.200000 62.850000 66.520000 ;
      LAYER met4 ;
        RECT 62.530000 66.200000 62.850000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.935000 62.100000 63.255000 62.420000 ;
      LAYER met4 ;
        RECT 62.935000 62.100000 63.255000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.935000 62.510000 63.255000 62.830000 ;
      LAYER met4 ;
        RECT 62.935000 62.510000 63.255000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.935000 62.920000 63.255000 63.240000 ;
      LAYER met4 ;
        RECT 62.935000 62.920000 63.255000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.935000 63.330000 63.255000 63.650000 ;
      LAYER met4 ;
        RECT 62.935000 63.330000 63.255000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.935000 63.740000 63.255000 64.060000 ;
      LAYER met4 ;
        RECT 62.935000 63.740000 63.255000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.935000 64.150000 63.255000 64.470000 ;
      LAYER met4 ;
        RECT 62.935000 64.150000 63.255000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.935000 64.560000 63.255000 64.880000 ;
      LAYER met4 ;
        RECT 62.935000 64.560000 63.255000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.935000 64.970000 63.255000 65.290000 ;
      LAYER met4 ;
        RECT 62.935000 64.970000 63.255000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.935000 65.380000 63.255000 65.700000 ;
      LAYER met4 ;
        RECT 62.935000 65.380000 63.255000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.935000 65.790000 63.255000 66.110000 ;
      LAYER met4 ;
        RECT 62.935000 65.790000 63.255000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.935000 66.200000 63.255000 66.520000 ;
      LAYER met4 ;
        RECT 62.935000 66.200000 63.255000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.340000 62.100000 63.660000 62.420000 ;
      LAYER met4 ;
        RECT 63.340000 62.100000 63.660000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.340000 62.510000 63.660000 62.830000 ;
      LAYER met4 ;
        RECT 63.340000 62.510000 63.660000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.340000 62.920000 63.660000 63.240000 ;
      LAYER met4 ;
        RECT 63.340000 62.920000 63.660000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.340000 63.330000 63.660000 63.650000 ;
      LAYER met4 ;
        RECT 63.340000 63.330000 63.660000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.340000 63.740000 63.660000 64.060000 ;
      LAYER met4 ;
        RECT 63.340000 63.740000 63.660000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.340000 64.150000 63.660000 64.470000 ;
      LAYER met4 ;
        RECT 63.340000 64.150000 63.660000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.340000 64.560000 63.660000 64.880000 ;
      LAYER met4 ;
        RECT 63.340000 64.560000 63.660000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.340000 64.970000 63.660000 65.290000 ;
      LAYER met4 ;
        RECT 63.340000 64.970000 63.660000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.340000 65.380000 63.660000 65.700000 ;
      LAYER met4 ;
        RECT 63.340000 65.380000 63.660000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.340000 65.790000 63.660000 66.110000 ;
      LAYER met4 ;
        RECT 63.340000 65.790000 63.660000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.340000 66.200000 63.660000 66.520000 ;
      LAYER met4 ;
        RECT 63.340000 66.200000 63.660000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.745000 62.100000 64.065000 62.420000 ;
      LAYER met4 ;
        RECT 63.745000 62.100000 64.065000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.745000 62.510000 64.065000 62.830000 ;
      LAYER met4 ;
        RECT 63.745000 62.510000 64.065000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.745000 62.920000 64.065000 63.240000 ;
      LAYER met4 ;
        RECT 63.745000 62.920000 64.065000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.745000 63.330000 64.065000 63.650000 ;
      LAYER met4 ;
        RECT 63.745000 63.330000 64.065000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.745000 63.740000 64.065000 64.060000 ;
      LAYER met4 ;
        RECT 63.745000 63.740000 64.065000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.745000 64.150000 64.065000 64.470000 ;
      LAYER met4 ;
        RECT 63.745000 64.150000 64.065000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.745000 64.560000 64.065000 64.880000 ;
      LAYER met4 ;
        RECT 63.745000 64.560000 64.065000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.745000 64.970000 64.065000 65.290000 ;
      LAYER met4 ;
        RECT 63.745000 64.970000 64.065000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.745000 65.380000 64.065000 65.700000 ;
      LAYER met4 ;
        RECT 63.745000 65.380000 64.065000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.745000 65.790000 64.065000 66.110000 ;
      LAYER met4 ;
        RECT 63.745000 65.790000 64.065000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.745000 66.200000 64.065000 66.520000 ;
      LAYER met4 ;
        RECT 63.745000 66.200000 64.065000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 62.100000 64.470000 62.420000 ;
      LAYER met4 ;
        RECT 64.150000 62.100000 64.470000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 62.510000 64.470000 62.830000 ;
      LAYER met4 ;
        RECT 64.150000 62.510000 64.470000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 62.920000 64.470000 63.240000 ;
      LAYER met4 ;
        RECT 64.150000 62.920000 64.470000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 63.330000 64.470000 63.650000 ;
      LAYER met4 ;
        RECT 64.150000 63.330000 64.470000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 63.740000 64.470000 64.060000 ;
      LAYER met4 ;
        RECT 64.150000 63.740000 64.470000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 64.150000 64.470000 64.470000 ;
      LAYER met4 ;
        RECT 64.150000 64.150000 64.470000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 64.560000 64.470000 64.880000 ;
      LAYER met4 ;
        RECT 64.150000 64.560000 64.470000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 64.970000 64.470000 65.290000 ;
      LAYER met4 ;
        RECT 64.150000 64.970000 64.470000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 65.380000 64.470000 65.700000 ;
      LAYER met4 ;
        RECT 64.150000 65.380000 64.470000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 65.790000 64.470000 66.110000 ;
      LAYER met4 ;
        RECT 64.150000 65.790000 64.470000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.150000 66.200000 64.470000 66.520000 ;
      LAYER met4 ;
        RECT 64.150000 66.200000 64.470000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.555000 62.100000 64.875000 62.420000 ;
      LAYER met4 ;
        RECT 64.555000 62.100000 64.875000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.555000 62.510000 64.875000 62.830000 ;
      LAYER met4 ;
        RECT 64.555000 62.510000 64.875000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.555000 62.920000 64.875000 63.240000 ;
      LAYER met4 ;
        RECT 64.555000 62.920000 64.875000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.555000 63.330000 64.875000 63.650000 ;
      LAYER met4 ;
        RECT 64.555000 63.330000 64.875000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.555000 63.740000 64.875000 64.060000 ;
      LAYER met4 ;
        RECT 64.555000 63.740000 64.875000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.555000 64.150000 64.875000 64.470000 ;
      LAYER met4 ;
        RECT 64.555000 64.150000 64.875000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.555000 64.560000 64.875000 64.880000 ;
      LAYER met4 ;
        RECT 64.555000 64.560000 64.875000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.555000 64.970000 64.875000 65.290000 ;
      LAYER met4 ;
        RECT 64.555000 64.970000 64.875000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.555000 65.380000 64.875000 65.700000 ;
      LAYER met4 ;
        RECT 64.555000 65.380000 64.875000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.555000 65.790000 64.875000 66.110000 ;
      LAYER met4 ;
        RECT 64.555000 65.790000 64.875000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.555000 66.200000 64.875000 66.520000 ;
      LAYER met4 ;
        RECT 64.555000 66.200000 64.875000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.960000 62.100000 65.280000 62.420000 ;
      LAYER met4 ;
        RECT 64.960000 62.100000 65.280000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.960000 62.510000 65.280000 62.830000 ;
      LAYER met4 ;
        RECT 64.960000 62.510000 65.280000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.960000 62.920000 65.280000 63.240000 ;
      LAYER met4 ;
        RECT 64.960000 62.920000 65.280000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.960000 63.330000 65.280000 63.650000 ;
      LAYER met4 ;
        RECT 64.960000 63.330000 65.280000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.960000 63.740000 65.280000 64.060000 ;
      LAYER met4 ;
        RECT 64.960000 63.740000 65.280000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.960000 64.150000 65.280000 64.470000 ;
      LAYER met4 ;
        RECT 64.960000 64.150000 65.280000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.960000 64.560000 65.280000 64.880000 ;
      LAYER met4 ;
        RECT 64.960000 64.560000 65.280000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.960000 64.970000 65.280000 65.290000 ;
      LAYER met4 ;
        RECT 64.960000 64.970000 65.280000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.960000 65.380000 65.280000 65.700000 ;
      LAYER met4 ;
        RECT 64.960000 65.380000 65.280000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.960000 65.790000 65.280000 66.110000 ;
      LAYER met4 ;
        RECT 64.960000 65.790000 65.280000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.960000 66.200000 65.280000 66.520000 ;
      LAYER met4 ;
        RECT 64.960000 66.200000 65.280000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.365000 62.100000 65.685000 62.420000 ;
      LAYER met4 ;
        RECT 65.365000 62.100000 65.685000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.365000 62.510000 65.685000 62.830000 ;
      LAYER met4 ;
        RECT 65.365000 62.510000 65.685000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.365000 62.920000 65.685000 63.240000 ;
      LAYER met4 ;
        RECT 65.365000 62.920000 65.685000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.365000 63.330000 65.685000 63.650000 ;
      LAYER met4 ;
        RECT 65.365000 63.330000 65.685000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.365000 63.740000 65.685000 64.060000 ;
      LAYER met4 ;
        RECT 65.365000 63.740000 65.685000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.365000 64.150000 65.685000 64.470000 ;
      LAYER met4 ;
        RECT 65.365000 64.150000 65.685000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.365000 64.560000 65.685000 64.880000 ;
      LAYER met4 ;
        RECT 65.365000 64.560000 65.685000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.365000 64.970000 65.685000 65.290000 ;
      LAYER met4 ;
        RECT 65.365000 64.970000 65.685000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.365000 65.380000 65.685000 65.700000 ;
      LAYER met4 ;
        RECT 65.365000 65.380000 65.685000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.365000 65.790000 65.685000 66.110000 ;
      LAYER met4 ;
        RECT 65.365000 65.790000 65.685000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.365000 66.200000 65.685000 66.520000 ;
      LAYER met4 ;
        RECT 65.365000 66.200000 65.685000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 62.100000 66.090000 62.420000 ;
      LAYER met4 ;
        RECT 65.770000 62.100000 66.090000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 62.510000 66.090000 62.830000 ;
      LAYER met4 ;
        RECT 65.770000 62.510000 66.090000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 62.920000 66.090000 63.240000 ;
      LAYER met4 ;
        RECT 65.770000 62.920000 66.090000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 63.330000 66.090000 63.650000 ;
      LAYER met4 ;
        RECT 65.770000 63.330000 66.090000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 63.740000 66.090000 64.060000 ;
      LAYER met4 ;
        RECT 65.770000 63.740000 66.090000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 64.150000 66.090000 64.470000 ;
      LAYER met4 ;
        RECT 65.770000 64.150000 66.090000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 64.560000 66.090000 64.880000 ;
      LAYER met4 ;
        RECT 65.770000 64.560000 66.090000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 64.970000 66.090000 65.290000 ;
      LAYER met4 ;
        RECT 65.770000 64.970000 66.090000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 65.380000 66.090000 65.700000 ;
      LAYER met4 ;
        RECT 65.770000 65.380000 66.090000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 65.790000 66.090000 66.110000 ;
      LAYER met4 ;
        RECT 65.770000 65.790000 66.090000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.770000 66.200000 66.090000 66.520000 ;
      LAYER met4 ;
        RECT 65.770000 66.200000 66.090000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.175000 62.100000 66.495000 62.420000 ;
      LAYER met4 ;
        RECT 66.175000 62.100000 66.495000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.175000 62.510000 66.495000 62.830000 ;
      LAYER met4 ;
        RECT 66.175000 62.510000 66.495000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.175000 62.920000 66.495000 63.240000 ;
      LAYER met4 ;
        RECT 66.175000 62.920000 66.495000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.175000 63.330000 66.495000 63.650000 ;
      LAYER met4 ;
        RECT 66.175000 63.330000 66.495000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.175000 63.740000 66.495000 64.060000 ;
      LAYER met4 ;
        RECT 66.175000 63.740000 66.495000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.175000 64.150000 66.495000 64.470000 ;
      LAYER met4 ;
        RECT 66.175000 64.150000 66.495000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.175000 64.560000 66.495000 64.880000 ;
      LAYER met4 ;
        RECT 66.175000 64.560000 66.495000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.175000 64.970000 66.495000 65.290000 ;
      LAYER met4 ;
        RECT 66.175000 64.970000 66.495000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.175000 65.380000 66.495000 65.700000 ;
      LAYER met4 ;
        RECT 66.175000 65.380000 66.495000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.175000 65.790000 66.495000 66.110000 ;
      LAYER met4 ;
        RECT 66.175000 65.790000 66.495000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.175000 66.200000 66.495000 66.520000 ;
      LAYER met4 ;
        RECT 66.175000 66.200000 66.495000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.580000 62.100000 66.900000 62.420000 ;
      LAYER met4 ;
        RECT 66.580000 62.100000 66.900000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.580000 62.510000 66.900000 62.830000 ;
      LAYER met4 ;
        RECT 66.580000 62.510000 66.900000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.580000 62.920000 66.900000 63.240000 ;
      LAYER met4 ;
        RECT 66.580000 62.920000 66.900000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.580000 63.330000 66.900000 63.650000 ;
      LAYER met4 ;
        RECT 66.580000 63.330000 66.900000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.580000 63.740000 66.900000 64.060000 ;
      LAYER met4 ;
        RECT 66.580000 63.740000 66.900000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.580000 64.150000 66.900000 64.470000 ;
      LAYER met4 ;
        RECT 66.580000 64.150000 66.900000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.580000 64.560000 66.900000 64.880000 ;
      LAYER met4 ;
        RECT 66.580000 64.560000 66.900000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.580000 64.970000 66.900000 65.290000 ;
      LAYER met4 ;
        RECT 66.580000 64.970000 66.900000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.580000 65.380000 66.900000 65.700000 ;
      LAYER met4 ;
        RECT 66.580000 65.380000 66.900000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.580000 65.790000 66.900000 66.110000 ;
      LAYER met4 ;
        RECT 66.580000 65.790000 66.900000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.580000 66.200000 66.900000 66.520000 ;
      LAYER met4 ;
        RECT 66.580000 66.200000 66.900000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.985000 62.100000 67.305000 62.420000 ;
      LAYER met4 ;
        RECT 66.985000 62.100000 67.305000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.985000 62.510000 67.305000 62.830000 ;
      LAYER met4 ;
        RECT 66.985000 62.510000 67.305000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.985000 62.920000 67.305000 63.240000 ;
      LAYER met4 ;
        RECT 66.985000 62.920000 67.305000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.985000 63.330000 67.305000 63.650000 ;
      LAYER met4 ;
        RECT 66.985000 63.330000 67.305000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.985000 63.740000 67.305000 64.060000 ;
      LAYER met4 ;
        RECT 66.985000 63.740000 67.305000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.985000 64.150000 67.305000 64.470000 ;
      LAYER met4 ;
        RECT 66.985000 64.150000 67.305000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.985000 64.560000 67.305000 64.880000 ;
      LAYER met4 ;
        RECT 66.985000 64.560000 67.305000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.985000 64.970000 67.305000 65.290000 ;
      LAYER met4 ;
        RECT 66.985000 64.970000 67.305000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.985000 65.380000 67.305000 65.700000 ;
      LAYER met4 ;
        RECT 66.985000 65.380000 67.305000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.985000 65.790000 67.305000 66.110000 ;
      LAYER met4 ;
        RECT 66.985000 65.790000 67.305000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.985000 66.200000 67.305000 66.520000 ;
      LAYER met4 ;
        RECT 66.985000 66.200000 67.305000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 62.100000 67.710000 62.420000 ;
      LAYER met4 ;
        RECT 67.390000 62.100000 67.710000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 62.510000 67.710000 62.830000 ;
      LAYER met4 ;
        RECT 67.390000 62.510000 67.710000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 62.920000 67.710000 63.240000 ;
      LAYER met4 ;
        RECT 67.390000 62.920000 67.710000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 63.330000 67.710000 63.650000 ;
      LAYER met4 ;
        RECT 67.390000 63.330000 67.710000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 63.740000 67.710000 64.060000 ;
      LAYER met4 ;
        RECT 67.390000 63.740000 67.710000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 64.150000 67.710000 64.470000 ;
      LAYER met4 ;
        RECT 67.390000 64.150000 67.710000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 64.560000 67.710000 64.880000 ;
      LAYER met4 ;
        RECT 67.390000 64.560000 67.710000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 64.970000 67.710000 65.290000 ;
      LAYER met4 ;
        RECT 67.390000 64.970000 67.710000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 65.380000 67.710000 65.700000 ;
      LAYER met4 ;
        RECT 67.390000 65.380000 67.710000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 65.790000 67.710000 66.110000 ;
      LAYER met4 ;
        RECT 67.390000 65.790000 67.710000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390000 66.200000 67.710000 66.520000 ;
      LAYER met4 ;
        RECT 67.390000 66.200000 67.710000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.795000 62.100000 68.115000 62.420000 ;
      LAYER met4 ;
        RECT 67.795000 62.100000 68.115000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.795000 62.510000 68.115000 62.830000 ;
      LAYER met4 ;
        RECT 67.795000 62.510000 68.115000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.795000 62.920000 68.115000 63.240000 ;
      LAYER met4 ;
        RECT 67.795000 62.920000 68.115000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.795000 63.330000 68.115000 63.650000 ;
      LAYER met4 ;
        RECT 67.795000 63.330000 68.115000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.795000 63.740000 68.115000 64.060000 ;
      LAYER met4 ;
        RECT 67.795000 63.740000 68.115000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.795000 64.150000 68.115000 64.470000 ;
      LAYER met4 ;
        RECT 67.795000 64.150000 68.115000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.795000 64.560000 68.115000 64.880000 ;
      LAYER met4 ;
        RECT 67.795000 64.560000 68.115000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.795000 64.970000 68.115000 65.290000 ;
      LAYER met4 ;
        RECT 67.795000 64.970000 68.115000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.795000 65.380000 68.115000 65.700000 ;
      LAYER met4 ;
        RECT 67.795000 65.380000 68.115000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.795000 65.790000 68.115000 66.110000 ;
      LAYER met4 ;
        RECT 67.795000 65.790000 68.115000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.795000 66.200000 68.115000 66.520000 ;
      LAYER met4 ;
        RECT 67.795000 66.200000 68.115000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.200000 62.100000 68.520000 62.420000 ;
      LAYER met4 ;
        RECT 68.200000 62.100000 68.520000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.200000 62.510000 68.520000 62.830000 ;
      LAYER met4 ;
        RECT 68.200000 62.510000 68.520000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.200000 62.920000 68.520000 63.240000 ;
      LAYER met4 ;
        RECT 68.200000 62.920000 68.520000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.200000 63.330000 68.520000 63.650000 ;
      LAYER met4 ;
        RECT 68.200000 63.330000 68.520000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.200000 63.740000 68.520000 64.060000 ;
      LAYER met4 ;
        RECT 68.200000 63.740000 68.520000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.200000 64.150000 68.520000 64.470000 ;
      LAYER met4 ;
        RECT 68.200000 64.150000 68.520000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.200000 64.560000 68.520000 64.880000 ;
      LAYER met4 ;
        RECT 68.200000 64.560000 68.520000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.200000 64.970000 68.520000 65.290000 ;
      LAYER met4 ;
        RECT 68.200000 64.970000 68.520000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.200000 65.380000 68.520000 65.700000 ;
      LAYER met4 ;
        RECT 68.200000 65.380000 68.520000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.200000 65.790000 68.520000 66.110000 ;
      LAYER met4 ;
        RECT 68.200000 65.790000 68.520000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.200000 66.200000 68.520000 66.520000 ;
      LAYER met4 ;
        RECT 68.200000 66.200000 68.520000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.605000 62.100000 68.925000 62.420000 ;
      LAYER met4 ;
        RECT 68.605000 62.100000 68.925000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.605000 62.510000 68.925000 62.830000 ;
      LAYER met4 ;
        RECT 68.605000 62.510000 68.925000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.605000 62.920000 68.925000 63.240000 ;
      LAYER met4 ;
        RECT 68.605000 62.920000 68.925000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.605000 63.330000 68.925000 63.650000 ;
      LAYER met4 ;
        RECT 68.605000 63.330000 68.925000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.605000 63.740000 68.925000 64.060000 ;
      LAYER met4 ;
        RECT 68.605000 63.740000 68.925000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.605000 64.150000 68.925000 64.470000 ;
      LAYER met4 ;
        RECT 68.605000 64.150000 68.925000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.605000 64.560000 68.925000 64.880000 ;
      LAYER met4 ;
        RECT 68.605000 64.560000 68.925000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.605000 64.970000 68.925000 65.290000 ;
      LAYER met4 ;
        RECT 68.605000 64.970000 68.925000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.605000 65.380000 68.925000 65.700000 ;
      LAYER met4 ;
        RECT 68.605000 65.380000 68.925000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.605000 65.790000 68.925000 66.110000 ;
      LAYER met4 ;
        RECT 68.605000 65.790000 68.925000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.605000 66.200000 68.925000 66.520000 ;
      LAYER met4 ;
        RECT 68.605000 66.200000 68.925000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010000 62.100000 69.330000 62.420000 ;
      LAYER met4 ;
        RECT 69.010000 62.100000 69.330000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010000 62.510000 69.330000 62.830000 ;
      LAYER met4 ;
        RECT 69.010000 62.510000 69.330000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010000 62.920000 69.330000 63.240000 ;
      LAYER met4 ;
        RECT 69.010000 62.920000 69.330000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010000 63.330000 69.330000 63.650000 ;
      LAYER met4 ;
        RECT 69.010000 63.330000 69.330000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010000 63.740000 69.330000 64.060000 ;
      LAYER met4 ;
        RECT 69.010000 63.740000 69.330000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010000 64.150000 69.330000 64.470000 ;
      LAYER met4 ;
        RECT 69.010000 64.150000 69.330000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010000 64.560000 69.330000 64.880000 ;
      LAYER met4 ;
        RECT 69.010000 64.560000 69.330000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010000 64.970000 69.330000 65.290000 ;
      LAYER met4 ;
        RECT 69.010000 64.970000 69.330000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010000 65.380000 69.330000 65.700000 ;
      LAYER met4 ;
        RECT 69.010000 65.380000 69.330000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010000 65.790000 69.330000 66.110000 ;
      LAYER met4 ;
        RECT 69.010000 65.790000 69.330000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010000 66.200000 69.330000 66.520000 ;
      LAYER met4 ;
        RECT 69.010000 66.200000 69.330000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.415000 62.100000 69.735000 62.420000 ;
      LAYER met4 ;
        RECT 69.415000 62.100000 69.735000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.415000 62.510000 69.735000 62.830000 ;
      LAYER met4 ;
        RECT 69.415000 62.510000 69.735000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.415000 62.920000 69.735000 63.240000 ;
      LAYER met4 ;
        RECT 69.415000 62.920000 69.735000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.415000 63.330000 69.735000 63.650000 ;
      LAYER met4 ;
        RECT 69.415000 63.330000 69.735000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.415000 63.740000 69.735000 64.060000 ;
      LAYER met4 ;
        RECT 69.415000 63.740000 69.735000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.415000 64.150000 69.735000 64.470000 ;
      LAYER met4 ;
        RECT 69.415000 64.150000 69.735000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.415000 64.560000 69.735000 64.880000 ;
      LAYER met4 ;
        RECT 69.415000 64.560000 69.735000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.415000 64.970000 69.735000 65.290000 ;
      LAYER met4 ;
        RECT 69.415000 64.970000 69.735000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.415000 65.380000 69.735000 65.700000 ;
      LAYER met4 ;
        RECT 69.415000 65.380000 69.735000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.415000 65.790000 69.735000 66.110000 ;
      LAYER met4 ;
        RECT 69.415000 65.790000 69.735000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.415000 66.200000 69.735000 66.520000 ;
      LAYER met4 ;
        RECT 69.415000 66.200000 69.735000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.820000 62.100000 70.140000 62.420000 ;
      LAYER met4 ;
        RECT 69.820000 62.100000 70.140000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.820000 62.510000 70.140000 62.830000 ;
      LAYER met4 ;
        RECT 69.820000 62.510000 70.140000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.820000 62.920000 70.140000 63.240000 ;
      LAYER met4 ;
        RECT 69.820000 62.920000 70.140000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.820000 63.330000 70.140000 63.650000 ;
      LAYER met4 ;
        RECT 69.820000 63.330000 70.140000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.820000 63.740000 70.140000 64.060000 ;
      LAYER met4 ;
        RECT 69.820000 63.740000 70.140000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.820000 64.150000 70.140000 64.470000 ;
      LAYER met4 ;
        RECT 69.820000 64.150000 70.140000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.820000 64.560000 70.140000 64.880000 ;
      LAYER met4 ;
        RECT 69.820000 64.560000 70.140000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.820000 64.970000 70.140000 65.290000 ;
      LAYER met4 ;
        RECT 69.820000 64.970000 70.140000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.820000 65.380000 70.140000 65.700000 ;
      LAYER met4 ;
        RECT 69.820000 65.380000 70.140000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.820000 65.790000 70.140000 66.110000 ;
      LAYER met4 ;
        RECT 69.820000 65.790000 70.140000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.820000 66.200000 70.140000 66.520000 ;
      LAYER met4 ;
        RECT 69.820000 66.200000 70.140000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110000 62.100000 7.430000 62.420000 ;
      LAYER met4 ;
        RECT 7.110000 62.100000 7.430000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110000 62.510000 7.430000 62.830000 ;
      LAYER met4 ;
        RECT 7.110000 62.510000 7.430000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110000 62.920000 7.430000 63.240000 ;
      LAYER met4 ;
        RECT 7.110000 62.920000 7.430000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110000 63.330000 7.430000 63.650000 ;
      LAYER met4 ;
        RECT 7.110000 63.330000 7.430000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110000 63.740000 7.430000 64.060000 ;
      LAYER met4 ;
        RECT 7.110000 63.740000 7.430000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110000 64.150000 7.430000 64.470000 ;
      LAYER met4 ;
        RECT 7.110000 64.150000 7.430000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110000 64.560000 7.430000 64.880000 ;
      LAYER met4 ;
        RECT 7.110000 64.560000 7.430000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110000 64.970000 7.430000 65.290000 ;
      LAYER met4 ;
        RECT 7.110000 64.970000 7.430000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110000 65.380000 7.430000 65.700000 ;
      LAYER met4 ;
        RECT 7.110000 65.380000 7.430000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110000 65.790000 7.430000 66.110000 ;
      LAYER met4 ;
        RECT 7.110000 65.790000 7.430000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110000 66.200000 7.430000 66.520000 ;
      LAYER met4 ;
        RECT 7.110000 66.200000 7.430000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515000 62.100000 7.835000 62.420000 ;
      LAYER met4 ;
        RECT 7.515000 62.100000 7.835000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515000 62.510000 7.835000 62.830000 ;
      LAYER met4 ;
        RECT 7.515000 62.510000 7.835000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515000 62.920000 7.835000 63.240000 ;
      LAYER met4 ;
        RECT 7.515000 62.920000 7.835000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515000 63.330000 7.835000 63.650000 ;
      LAYER met4 ;
        RECT 7.515000 63.330000 7.835000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515000 63.740000 7.835000 64.060000 ;
      LAYER met4 ;
        RECT 7.515000 63.740000 7.835000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515000 64.150000 7.835000 64.470000 ;
      LAYER met4 ;
        RECT 7.515000 64.150000 7.835000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515000 64.560000 7.835000 64.880000 ;
      LAYER met4 ;
        RECT 7.515000 64.560000 7.835000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515000 64.970000 7.835000 65.290000 ;
      LAYER met4 ;
        RECT 7.515000 64.970000 7.835000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515000 65.380000 7.835000 65.700000 ;
      LAYER met4 ;
        RECT 7.515000 65.380000 7.835000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515000 65.790000 7.835000 66.110000 ;
      LAYER met4 ;
        RECT 7.515000 65.790000 7.835000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515000 66.200000 7.835000 66.520000 ;
      LAYER met4 ;
        RECT 7.515000 66.200000 7.835000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920000 62.100000 8.240000 62.420000 ;
      LAYER met4 ;
        RECT 7.920000 62.100000 8.240000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920000 62.510000 8.240000 62.830000 ;
      LAYER met4 ;
        RECT 7.920000 62.510000 8.240000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920000 62.920000 8.240000 63.240000 ;
      LAYER met4 ;
        RECT 7.920000 62.920000 8.240000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920000 63.330000 8.240000 63.650000 ;
      LAYER met4 ;
        RECT 7.920000 63.330000 8.240000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920000 63.740000 8.240000 64.060000 ;
      LAYER met4 ;
        RECT 7.920000 63.740000 8.240000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920000 64.150000 8.240000 64.470000 ;
      LAYER met4 ;
        RECT 7.920000 64.150000 8.240000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920000 64.560000 8.240000 64.880000 ;
      LAYER met4 ;
        RECT 7.920000 64.560000 8.240000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920000 64.970000 8.240000 65.290000 ;
      LAYER met4 ;
        RECT 7.920000 64.970000 8.240000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920000 65.380000 8.240000 65.700000 ;
      LAYER met4 ;
        RECT 7.920000 65.380000 8.240000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920000 65.790000 8.240000 66.110000 ;
      LAYER met4 ;
        RECT 7.920000 65.790000 8.240000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920000 66.200000 8.240000 66.520000 ;
      LAYER met4 ;
        RECT 7.920000 66.200000 8.240000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.225000 62.100000 70.545000 62.420000 ;
      LAYER met4 ;
        RECT 70.225000 62.100000 70.545000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.225000 62.510000 70.545000 62.830000 ;
      LAYER met4 ;
        RECT 70.225000 62.510000 70.545000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.225000 62.920000 70.545000 63.240000 ;
      LAYER met4 ;
        RECT 70.225000 62.920000 70.545000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.225000 63.330000 70.545000 63.650000 ;
      LAYER met4 ;
        RECT 70.225000 63.330000 70.545000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.225000 63.740000 70.545000 64.060000 ;
      LAYER met4 ;
        RECT 70.225000 63.740000 70.545000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.225000 64.150000 70.545000 64.470000 ;
      LAYER met4 ;
        RECT 70.225000 64.150000 70.545000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.225000 64.560000 70.545000 64.880000 ;
      LAYER met4 ;
        RECT 70.225000 64.560000 70.545000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.225000 64.970000 70.545000 65.290000 ;
      LAYER met4 ;
        RECT 70.225000 64.970000 70.545000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.225000 65.380000 70.545000 65.700000 ;
      LAYER met4 ;
        RECT 70.225000 65.380000 70.545000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.225000 65.790000 70.545000 66.110000 ;
      LAYER met4 ;
        RECT 70.225000 65.790000 70.545000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.225000 66.200000 70.545000 66.520000 ;
      LAYER met4 ;
        RECT 70.225000 66.200000 70.545000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630000 62.100000 70.950000 62.420000 ;
      LAYER met4 ;
        RECT 70.630000 62.100000 70.950000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630000 62.510000 70.950000 62.830000 ;
      LAYER met4 ;
        RECT 70.630000 62.510000 70.950000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630000 62.920000 70.950000 63.240000 ;
      LAYER met4 ;
        RECT 70.630000 62.920000 70.950000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630000 63.330000 70.950000 63.650000 ;
      LAYER met4 ;
        RECT 70.630000 63.330000 70.950000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630000 63.740000 70.950000 64.060000 ;
      LAYER met4 ;
        RECT 70.630000 63.740000 70.950000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630000 64.150000 70.950000 64.470000 ;
      LAYER met4 ;
        RECT 70.630000 64.150000 70.950000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630000 64.560000 70.950000 64.880000 ;
      LAYER met4 ;
        RECT 70.630000 64.560000 70.950000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630000 64.970000 70.950000 65.290000 ;
      LAYER met4 ;
        RECT 70.630000 64.970000 70.950000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630000 65.380000 70.950000 65.700000 ;
      LAYER met4 ;
        RECT 70.630000 65.380000 70.950000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630000 65.790000 70.950000 66.110000 ;
      LAYER met4 ;
        RECT 70.630000 65.790000 70.950000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630000 66.200000 70.950000 66.520000 ;
      LAYER met4 ;
        RECT 70.630000 66.200000 70.950000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.035000 62.100000 71.355000 62.420000 ;
      LAYER met4 ;
        RECT 71.035000 62.100000 71.355000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.035000 62.510000 71.355000 62.830000 ;
      LAYER met4 ;
        RECT 71.035000 62.510000 71.355000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.035000 62.920000 71.355000 63.240000 ;
      LAYER met4 ;
        RECT 71.035000 62.920000 71.355000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.035000 63.330000 71.355000 63.650000 ;
      LAYER met4 ;
        RECT 71.035000 63.330000 71.355000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.035000 63.740000 71.355000 64.060000 ;
      LAYER met4 ;
        RECT 71.035000 63.740000 71.355000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.035000 64.150000 71.355000 64.470000 ;
      LAYER met4 ;
        RECT 71.035000 64.150000 71.355000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.035000 64.560000 71.355000 64.880000 ;
      LAYER met4 ;
        RECT 71.035000 64.560000 71.355000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.035000 64.970000 71.355000 65.290000 ;
      LAYER met4 ;
        RECT 71.035000 64.970000 71.355000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.035000 65.380000 71.355000 65.700000 ;
      LAYER met4 ;
        RECT 71.035000 65.380000 71.355000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.035000 65.790000 71.355000 66.110000 ;
      LAYER met4 ;
        RECT 71.035000 65.790000 71.355000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.035000 66.200000 71.355000 66.520000 ;
      LAYER met4 ;
        RECT 71.035000 66.200000 71.355000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 62.100000 71.760000 62.420000 ;
      LAYER met4 ;
        RECT 71.440000 62.100000 71.760000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 62.510000 71.760000 62.830000 ;
      LAYER met4 ;
        RECT 71.440000 62.510000 71.760000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 62.920000 71.760000 63.240000 ;
      LAYER met4 ;
        RECT 71.440000 62.920000 71.760000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 63.330000 71.760000 63.650000 ;
      LAYER met4 ;
        RECT 71.440000 63.330000 71.760000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 63.740000 71.760000 64.060000 ;
      LAYER met4 ;
        RECT 71.440000 63.740000 71.760000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 64.150000 71.760000 64.470000 ;
      LAYER met4 ;
        RECT 71.440000 64.150000 71.760000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 64.560000 71.760000 64.880000 ;
      LAYER met4 ;
        RECT 71.440000 64.560000 71.760000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 64.970000 71.760000 65.290000 ;
      LAYER met4 ;
        RECT 71.440000 64.970000 71.760000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 65.380000 71.760000 65.700000 ;
      LAYER met4 ;
        RECT 71.440000 65.380000 71.760000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 65.790000 71.760000 66.110000 ;
      LAYER met4 ;
        RECT 71.440000 65.790000 71.760000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440000 66.200000 71.760000 66.520000 ;
      LAYER met4 ;
        RECT 71.440000 66.200000 71.760000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.845000 62.100000 72.165000 62.420000 ;
      LAYER met4 ;
        RECT 71.845000 62.100000 72.165000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.845000 62.510000 72.165000 62.830000 ;
      LAYER met4 ;
        RECT 71.845000 62.510000 72.165000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.845000 62.920000 72.165000 63.240000 ;
      LAYER met4 ;
        RECT 71.845000 62.920000 72.165000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.845000 63.330000 72.165000 63.650000 ;
      LAYER met4 ;
        RECT 71.845000 63.330000 72.165000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.845000 63.740000 72.165000 64.060000 ;
      LAYER met4 ;
        RECT 71.845000 63.740000 72.165000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.845000 64.150000 72.165000 64.470000 ;
      LAYER met4 ;
        RECT 71.845000 64.150000 72.165000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.845000 64.560000 72.165000 64.880000 ;
      LAYER met4 ;
        RECT 71.845000 64.560000 72.165000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.845000 64.970000 72.165000 65.290000 ;
      LAYER met4 ;
        RECT 71.845000 64.970000 72.165000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.845000 65.380000 72.165000 65.700000 ;
      LAYER met4 ;
        RECT 71.845000 65.380000 72.165000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.845000 65.790000 72.165000 66.110000 ;
      LAYER met4 ;
        RECT 71.845000 65.790000 72.165000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.845000 66.200000 72.165000 66.520000 ;
      LAYER met4 ;
        RECT 71.845000 66.200000 72.165000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.255000 62.100000 72.575000 62.420000 ;
      LAYER met4 ;
        RECT 72.255000 62.100000 72.575000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.255000 62.510000 72.575000 62.830000 ;
      LAYER met4 ;
        RECT 72.255000 62.510000 72.575000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.255000 62.920000 72.575000 63.240000 ;
      LAYER met4 ;
        RECT 72.255000 62.920000 72.575000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.255000 63.330000 72.575000 63.650000 ;
      LAYER met4 ;
        RECT 72.255000 63.330000 72.575000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.255000 63.740000 72.575000 64.060000 ;
      LAYER met4 ;
        RECT 72.255000 63.740000 72.575000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.255000 64.150000 72.575000 64.470000 ;
      LAYER met4 ;
        RECT 72.255000 64.150000 72.575000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.255000 64.560000 72.575000 64.880000 ;
      LAYER met4 ;
        RECT 72.255000 64.560000 72.575000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.255000 64.970000 72.575000 65.290000 ;
      LAYER met4 ;
        RECT 72.255000 64.970000 72.575000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.255000 65.380000 72.575000 65.700000 ;
      LAYER met4 ;
        RECT 72.255000 65.380000 72.575000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.255000 65.790000 72.575000 66.110000 ;
      LAYER met4 ;
        RECT 72.255000 65.790000 72.575000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.255000 66.200000 72.575000 66.520000 ;
      LAYER met4 ;
        RECT 72.255000 66.200000 72.575000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.665000 62.100000 72.985000 62.420000 ;
      LAYER met4 ;
        RECT 72.665000 62.100000 72.985000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.665000 62.510000 72.985000 62.830000 ;
      LAYER met4 ;
        RECT 72.665000 62.510000 72.985000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.665000 62.920000 72.985000 63.240000 ;
      LAYER met4 ;
        RECT 72.665000 62.920000 72.985000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.665000 63.330000 72.985000 63.650000 ;
      LAYER met4 ;
        RECT 72.665000 63.330000 72.985000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.665000 63.740000 72.985000 64.060000 ;
      LAYER met4 ;
        RECT 72.665000 63.740000 72.985000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.665000 64.150000 72.985000 64.470000 ;
      LAYER met4 ;
        RECT 72.665000 64.150000 72.985000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.665000 64.560000 72.985000 64.880000 ;
      LAYER met4 ;
        RECT 72.665000 64.560000 72.985000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.665000 64.970000 72.985000 65.290000 ;
      LAYER met4 ;
        RECT 72.665000 64.970000 72.985000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.665000 65.380000 72.985000 65.700000 ;
      LAYER met4 ;
        RECT 72.665000 65.380000 72.985000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.665000 65.790000 72.985000 66.110000 ;
      LAYER met4 ;
        RECT 72.665000 65.790000 72.985000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.665000 66.200000 72.985000 66.520000 ;
      LAYER met4 ;
        RECT 72.665000 66.200000 72.985000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.075000 62.100000 73.395000 62.420000 ;
      LAYER met4 ;
        RECT 73.075000 62.100000 73.395000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.075000 62.510000 73.395000 62.830000 ;
      LAYER met4 ;
        RECT 73.075000 62.510000 73.395000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.075000 62.920000 73.395000 63.240000 ;
      LAYER met4 ;
        RECT 73.075000 62.920000 73.395000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.075000 63.330000 73.395000 63.650000 ;
      LAYER met4 ;
        RECT 73.075000 63.330000 73.395000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.075000 63.740000 73.395000 64.060000 ;
      LAYER met4 ;
        RECT 73.075000 63.740000 73.395000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.075000 64.150000 73.395000 64.470000 ;
      LAYER met4 ;
        RECT 73.075000 64.150000 73.395000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.075000 64.560000 73.395000 64.880000 ;
      LAYER met4 ;
        RECT 73.075000 64.560000 73.395000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.075000 64.970000 73.395000 65.290000 ;
      LAYER met4 ;
        RECT 73.075000 64.970000 73.395000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.075000 65.380000 73.395000 65.700000 ;
      LAYER met4 ;
        RECT 73.075000 65.380000 73.395000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.075000 65.790000 73.395000 66.110000 ;
      LAYER met4 ;
        RECT 73.075000 65.790000 73.395000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.075000 66.200000 73.395000 66.520000 ;
      LAYER met4 ;
        RECT 73.075000 66.200000 73.395000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.485000 62.100000 73.805000 62.420000 ;
      LAYER met4 ;
        RECT 73.485000 62.100000 73.805000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.485000 62.510000 73.805000 62.830000 ;
      LAYER met4 ;
        RECT 73.485000 62.510000 73.805000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.485000 62.920000 73.805000 63.240000 ;
      LAYER met4 ;
        RECT 73.485000 62.920000 73.805000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.485000 63.330000 73.805000 63.650000 ;
      LAYER met4 ;
        RECT 73.485000 63.330000 73.805000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.485000 63.740000 73.805000 64.060000 ;
      LAYER met4 ;
        RECT 73.485000 63.740000 73.805000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.485000 64.150000 73.805000 64.470000 ;
      LAYER met4 ;
        RECT 73.485000 64.150000 73.805000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.485000 64.560000 73.805000 64.880000 ;
      LAYER met4 ;
        RECT 73.485000 64.560000 73.805000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.485000 64.970000 73.805000 65.290000 ;
      LAYER met4 ;
        RECT 73.485000 64.970000 73.805000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.485000 65.380000 73.805000 65.700000 ;
      LAYER met4 ;
        RECT 73.485000 65.380000 73.805000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.485000 65.790000 73.805000 66.110000 ;
      LAYER met4 ;
        RECT 73.485000 65.790000 73.805000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.485000 66.200000 73.805000 66.520000 ;
      LAYER met4 ;
        RECT 73.485000 66.200000 73.805000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.895000 62.100000 74.215000 62.420000 ;
      LAYER met4 ;
        RECT 73.895000 62.100000 74.215000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.895000 62.510000 74.215000 62.830000 ;
      LAYER met4 ;
        RECT 73.895000 62.510000 74.215000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.895000 62.920000 74.215000 63.240000 ;
      LAYER met4 ;
        RECT 73.895000 62.920000 74.215000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.895000 63.330000 74.215000 63.650000 ;
      LAYER met4 ;
        RECT 73.895000 63.330000 74.215000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.895000 63.740000 74.215000 64.060000 ;
      LAYER met4 ;
        RECT 73.895000 63.740000 74.215000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.895000 64.150000 74.215000 64.470000 ;
      LAYER met4 ;
        RECT 73.895000 64.150000 74.215000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.895000 64.560000 74.215000 64.880000 ;
      LAYER met4 ;
        RECT 73.895000 64.560000 74.215000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.895000 64.970000 74.215000 65.290000 ;
      LAYER met4 ;
        RECT 73.895000 64.970000 74.215000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.895000 65.380000 74.215000 65.700000 ;
      LAYER met4 ;
        RECT 73.895000 65.380000 74.215000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.895000 65.790000 74.215000 66.110000 ;
      LAYER met4 ;
        RECT 73.895000 65.790000 74.215000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.895000 66.200000 74.215000 66.520000 ;
      LAYER met4 ;
        RECT 73.895000 66.200000 74.215000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 62.100000 74.625000 62.420000 ;
      LAYER met4 ;
        RECT 74.305000 62.100000 74.625000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 62.510000 74.625000 62.830000 ;
      LAYER met4 ;
        RECT 74.305000 62.510000 74.625000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 62.920000 74.625000 63.240000 ;
      LAYER met4 ;
        RECT 74.305000 62.920000 74.625000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 63.330000 74.625000 63.650000 ;
      LAYER met4 ;
        RECT 74.305000 63.330000 74.625000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 63.740000 74.625000 64.060000 ;
      LAYER met4 ;
        RECT 74.305000 63.740000 74.625000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 64.150000 74.625000 64.470000 ;
      LAYER met4 ;
        RECT 74.305000 64.150000 74.625000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 64.560000 74.625000 64.880000 ;
      LAYER met4 ;
        RECT 74.305000 64.560000 74.625000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 64.970000 74.625000 65.290000 ;
      LAYER met4 ;
        RECT 74.305000 64.970000 74.625000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 65.380000 74.625000 65.700000 ;
      LAYER met4 ;
        RECT 74.305000 65.380000 74.625000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 65.790000 74.625000 66.110000 ;
      LAYER met4 ;
        RECT 74.305000 65.790000 74.625000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 66.200000 74.625000 66.520000 ;
      LAYER met4 ;
        RECT 74.305000 66.200000 74.625000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325000 62.100000 8.645000 62.420000 ;
      LAYER met4 ;
        RECT 8.325000 62.100000 8.645000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325000 62.510000 8.645000 62.830000 ;
      LAYER met4 ;
        RECT 8.325000 62.510000 8.645000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325000 62.920000 8.645000 63.240000 ;
      LAYER met4 ;
        RECT 8.325000 62.920000 8.645000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325000 63.330000 8.645000 63.650000 ;
      LAYER met4 ;
        RECT 8.325000 63.330000 8.645000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325000 63.740000 8.645000 64.060000 ;
      LAYER met4 ;
        RECT 8.325000 63.740000 8.645000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325000 64.150000 8.645000 64.470000 ;
      LAYER met4 ;
        RECT 8.325000 64.150000 8.645000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325000 64.560000 8.645000 64.880000 ;
      LAYER met4 ;
        RECT 8.325000 64.560000 8.645000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325000 64.970000 8.645000 65.290000 ;
      LAYER met4 ;
        RECT 8.325000 64.970000 8.645000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325000 65.380000 8.645000 65.700000 ;
      LAYER met4 ;
        RECT 8.325000 65.380000 8.645000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325000 65.790000 8.645000 66.110000 ;
      LAYER met4 ;
        RECT 8.325000 65.790000 8.645000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325000 66.200000 8.645000 66.520000 ;
      LAYER met4 ;
        RECT 8.325000 66.200000 8.645000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730000 62.100000 9.050000 62.420000 ;
      LAYER met4 ;
        RECT 8.730000 62.100000 9.050000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730000 62.510000 9.050000 62.830000 ;
      LAYER met4 ;
        RECT 8.730000 62.510000 9.050000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730000 62.920000 9.050000 63.240000 ;
      LAYER met4 ;
        RECT 8.730000 62.920000 9.050000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730000 63.330000 9.050000 63.650000 ;
      LAYER met4 ;
        RECT 8.730000 63.330000 9.050000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730000 63.740000 9.050000 64.060000 ;
      LAYER met4 ;
        RECT 8.730000 63.740000 9.050000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730000 64.150000 9.050000 64.470000 ;
      LAYER met4 ;
        RECT 8.730000 64.150000 9.050000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730000 64.560000 9.050000 64.880000 ;
      LAYER met4 ;
        RECT 8.730000 64.560000 9.050000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730000 64.970000 9.050000 65.290000 ;
      LAYER met4 ;
        RECT 8.730000 64.970000 9.050000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730000 65.380000 9.050000 65.700000 ;
      LAYER met4 ;
        RECT 8.730000 65.380000 9.050000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730000 65.790000 9.050000 66.110000 ;
      LAYER met4 ;
        RECT 8.730000 65.790000 9.050000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730000 66.200000 9.050000 66.520000 ;
      LAYER met4 ;
        RECT 8.730000 66.200000 9.050000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135000 62.100000 9.455000 62.420000 ;
      LAYER met4 ;
        RECT 9.135000 62.100000 9.455000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135000 62.510000 9.455000 62.830000 ;
      LAYER met4 ;
        RECT 9.135000 62.510000 9.455000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135000 62.920000 9.455000 63.240000 ;
      LAYER met4 ;
        RECT 9.135000 62.920000 9.455000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135000 63.330000 9.455000 63.650000 ;
      LAYER met4 ;
        RECT 9.135000 63.330000 9.455000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135000 63.740000 9.455000 64.060000 ;
      LAYER met4 ;
        RECT 9.135000 63.740000 9.455000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135000 64.150000 9.455000 64.470000 ;
      LAYER met4 ;
        RECT 9.135000 64.150000 9.455000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135000 64.560000 9.455000 64.880000 ;
      LAYER met4 ;
        RECT 9.135000 64.560000 9.455000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135000 64.970000 9.455000 65.290000 ;
      LAYER met4 ;
        RECT 9.135000 64.970000 9.455000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135000 65.380000 9.455000 65.700000 ;
      LAYER met4 ;
        RECT 9.135000 65.380000 9.455000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135000 65.790000 9.455000 66.110000 ;
      LAYER met4 ;
        RECT 9.135000 65.790000 9.455000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135000 66.200000 9.455000 66.520000 ;
      LAYER met4 ;
        RECT 9.135000 66.200000 9.455000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540000 62.100000 9.860000 62.420000 ;
      LAYER met4 ;
        RECT 9.540000 62.100000 9.860000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540000 62.510000 9.860000 62.830000 ;
      LAYER met4 ;
        RECT 9.540000 62.510000 9.860000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540000 62.920000 9.860000 63.240000 ;
      LAYER met4 ;
        RECT 9.540000 62.920000 9.860000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540000 63.330000 9.860000 63.650000 ;
      LAYER met4 ;
        RECT 9.540000 63.330000 9.860000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540000 63.740000 9.860000 64.060000 ;
      LAYER met4 ;
        RECT 9.540000 63.740000 9.860000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540000 64.150000 9.860000 64.470000 ;
      LAYER met4 ;
        RECT 9.540000 64.150000 9.860000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540000 64.560000 9.860000 64.880000 ;
      LAYER met4 ;
        RECT 9.540000 64.560000 9.860000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540000 64.970000 9.860000 65.290000 ;
      LAYER met4 ;
        RECT 9.540000 64.970000 9.860000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540000 65.380000 9.860000 65.700000 ;
      LAYER met4 ;
        RECT 9.540000 65.380000 9.860000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540000 65.790000 9.860000 66.110000 ;
      LAYER met4 ;
        RECT 9.540000 65.790000 9.860000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540000 66.200000 9.860000 66.520000 ;
      LAYER met4 ;
        RECT 9.540000 66.200000 9.860000 66.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945000 62.100000 10.265000 62.420000 ;
      LAYER met4 ;
        RECT 9.945000 62.100000 10.265000 62.420000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945000 62.510000 10.265000 62.830000 ;
      LAYER met4 ;
        RECT 9.945000 62.510000 10.265000 62.830000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945000 62.920000 10.265000 63.240000 ;
      LAYER met4 ;
        RECT 9.945000 62.920000 10.265000 63.240000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945000 63.330000 10.265000 63.650000 ;
      LAYER met4 ;
        RECT 9.945000 63.330000 10.265000 63.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945000 63.740000 10.265000 64.060000 ;
      LAYER met4 ;
        RECT 9.945000 63.740000 10.265000 64.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945000 64.150000 10.265000 64.470000 ;
      LAYER met4 ;
        RECT 9.945000 64.150000 10.265000 64.470000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945000 64.560000 10.265000 64.880000 ;
      LAYER met4 ;
        RECT 9.945000 64.560000 10.265000 64.880000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945000 64.970000 10.265000 65.290000 ;
      LAYER met4 ;
        RECT 9.945000 64.970000 10.265000 65.290000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945000 65.380000 10.265000 65.700000 ;
      LAYER met4 ;
        RECT 9.945000 65.380000 10.265000 65.700000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945000 65.790000 10.265000 66.110000 ;
      LAYER met4 ;
        RECT 9.945000 65.790000 10.265000 66.110000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945000 66.200000 10.265000 66.520000 ;
      LAYER met4 ;
        RECT 9.945000 66.200000 10.265000 66.520000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met3 ;
      RECT 0.595000 17.790000 74.660000 92.960000 ;
    LAYER met4 ;
      RECT 0.000000  0.035000 75.000000  45.965000 ;
      RECT 0.000000 49.745000 75.000000  50.725000 ;
      RECT 0.000000 54.505000 75.000000 198.000000 ;
    LAYER met5 ;
      RECT 0.000000  0.135000 72.130000  13.035000 ;
      RECT 0.000000 13.035000 72.435000  17.885000 ;
      RECT 0.000000 17.885000 75.000000  22.335000 ;
      RECT 0.000000 22.335000 72.130000  34.835000 ;
      RECT 0.000000 34.835000 75.000000  38.085000 ;
      RECT 0.000000 38.085000 72.130000  62.185000 ;
      RECT 0.000000 62.185000 75.000000 198.000000 ;
  END
END sky130_fd_io__overlay_vddio_lvc
END LIBRARY
