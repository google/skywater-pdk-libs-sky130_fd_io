# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sky130_fd_io__top_vrefcapv2
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 17.28 BY 200 ;
  SYMMETRY X Y R90 ;

  PIN cneg
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 3.475 0 6.475 0.83 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.475 0 13.475 0.83 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.475 196.705 13.475 198.91 ;
        RECT 10.475 195.825 13.475 195.895 ;
        RECT 10.405 195.895 13.475 195.965 ;
        RECT 10.335 195.965 13.475 196.035 ;
        RECT 10.265 196.035 13.475 196.105 ;
        RECT 10.195 196.105 13.475 196.175 ;
        RECT 10.125 196.175 13.475 196.245 ;
        RECT 10.055 196.245 13.475 196.315 ;
        RECT 9.985 196.315 13.475 196.385 ;
        RECT 9.915 196.385 13.475 196.455 ;
        RECT 9.845 196.455 13.475 196.525 ;
        RECT 9.775 196.525 13.475 196.595 ;
        RECT 9.705 196.595 13.475 196.665 ;
        RECT 9.635 196.665 13.475 196.705 ;
        RECT 3.475 195.825 6.475 195.895 ;
        RECT 3.475 195.895 6.545 195.965 ;
        RECT 3.475 195.965 6.615 196.035 ;
        RECT 3.475 196.035 6.685 196.105 ;
        RECT 3.475 196.105 6.755 196.175 ;
        RECT 3.475 196.175 6.825 196.245 ;
        RECT 3.475 196.245 6.895 196.315 ;
        RECT 3.475 196.315 6.965 196.385 ;
        RECT 3.475 196.385 7.035 196.455 ;
        RECT 3.475 196.455 7.105 196.525 ;
        RECT 3.475 196.525 7.175 196.595 ;
        RECT 3.475 196.595 7.245 196.665 ;
        RECT 3.475 196.665 7.315 196.705 ;
        RECT 10.475 0 13.475 195.825 ;
        RECT 3.475 0 6.475 195.825 ;
    END
  END cneg

  PIN cpos
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 7.475 0 9.475 0.83 ;
    END
    PORT
      LAYER met2 ;
        RECT 7.475 0 9.475 195.315 ;
    END
  END cpos

  PIN amuxbus_a
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0 53.125 17.28 56.105 ;
    END
    ANTENNAPARTIALMETALSIDEAREA 18.816 LAYER met4 ;
  END amuxbus_a

  PIN amuxbus_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0 48.365 17.28 51.345 ;
    END
    ANTENNAPARTIALMETALSIDEAREA 18.816 LAYER met4 ;
  END amuxbus_b

  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 41.685 17.28 46.135 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 41.585 17.28 46.235 ;
    END
  END vssd

  PIN vdda
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 15.035 17.28 18.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 14.935 17.28 18.385 ;
    END
  END vdda

  PIN vswitch
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 31.985 17.28 35.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 31.885 17.28 35.335 ;
    END
  END vswitch

  PIN vcchib
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 2.135 17.28 7.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 2.035 17.28 7.485 ;
    END
  END vcchib

  PIN vssa
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 36.835 17.28 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0 47.735 17.28 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 36.735 17.28 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 47.735 17.28 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 51.645 17.28 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 56.405 17.28 56.735 ;
    END
  END vssa

  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 8.985 17.28 13.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 8.885 17.28 13.535 ;
    END
  END vccd

  PIN vssio_q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 58.335 17.28 62.585 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 58.235 17.28 62.685 ;
    END
  END vssio_q

  PIN vddio
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 19.885 17.28 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 0 70.035 17.28 94.985 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 19.785 17.28 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 70.035 17.28 95 ;
    END
  END vddio

  PIN vddio_q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 64.185 17.28 68.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 64.085 17.28 68.535 ;
    END
  END vddio_q

  PIN vssio
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 25.935 17.28 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0 175.785 17.28 200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 25.835 17.28 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0 175.785 17.28 200 ;
    END
  END vssio
  OBS
    LAYER li1 ;
      RECT 13.275 174.38 13.445 184.11 ;
      RECT 14.455 163.73 14.625 173.46 ;
      RECT 14.455 153.01 14.625 162.74 ;
      RECT 14.455 142.43 14.625 152.16 ;
      RECT 14.455 131.71 14.625 141.44 ;
      RECT 14.455 185.09 14.625 194.82 ;
      RECT 14.455 174.38 14.625 184.11 ;
      RECT 5.015 57.23 5.185 66.96 ;
      RECT 3.835 57.23 4.005 66.96 ;
      RECT 5.015 67.81 5.185 77.54 ;
      RECT 3.835 67.81 4.005 77.54 ;
      RECT 6.195 110.41 6.365 120.14 ;
      RECT 7.375 110.41 7.545 120.14 ;
      RECT 6.195 99.83 6.365 109.56 ;
      RECT 7.375 99.83 7.545 109.56 ;
      RECT 6.195 89.11 6.365 98.84 ;
      RECT 7.375 89.11 7.545 98.84 ;
      RECT 7.375 46.51 7.545 56.24 ;
      RECT 6.195 46.51 6.365 56.24 ;
      RECT 6.195 121.13 6.365 130.86 ;
      RECT 7.375 121.13 7.545 130.86 ;
      RECT 7.375 78.53 7.545 88.26 ;
      RECT 6.195 78.53 6.365 88.26 ;
      RECT 7.375 57.23 7.545 66.96 ;
      RECT 6.195 57.23 6.365 66.96 ;
      RECT 7.375 67.81 7.545 77.54 ;
      RECT 6.195 67.81 6.365 77.54 ;
      RECT 8.555 110.41 8.725 120.14 ;
      RECT 9.735 110.41 9.905 120.14 ;
      RECT 10.915 110.41 11.085 120.14 ;
      RECT 8.555 99.83 8.725 109.56 ;
      RECT 9.735 99.83 9.905 109.56 ;
      RECT 10.915 99.83 11.085 109.56 ;
      RECT 8.555 89.11 8.725 98.84 ;
      RECT 9.735 89.11 9.905 98.84 ;
      RECT 10.915 89.11 11.085 98.84 ;
      RECT 10.915 46.51 11.085 56.24 ;
      RECT 9.735 46.51 9.905 56.24 ;
      RECT 8.555 46.51 8.725 56.24 ;
      RECT 8.555 121.13 8.725 130.86 ;
      RECT 9.735 121.13 9.905 130.86 ;
      RECT 10.915 121.13 11.085 130.86 ;
      RECT 10.915 78.53 11.085 88.26 ;
      RECT 9.735 78.53 9.905 88.26 ;
      RECT 8.555 78.53 8.725 88.26 ;
      RECT 10.915 57.23 11.085 66.96 ;
      RECT 9.735 57.23 9.905 66.96 ;
      RECT 8.555 57.23 8.725 66.96 ;
      RECT 10.915 67.81 11.085 77.54 ;
      RECT 9.735 67.81 9.905 77.54 ;
      RECT 8.555 67.81 8.725 77.54 ;
      RECT 12.095 110.41 12.265 120.14 ;
      RECT 13.275 110.41 13.445 120.14 ;
      RECT 12.095 99.83 12.265 109.56 ;
      RECT 13.275 99.83 13.445 109.56 ;
      RECT 12.095 89.11 12.265 98.84 ;
      RECT 13.275 89.11 13.445 98.84 ;
      RECT 13.275 46.51 13.445 56.24 ;
      RECT 12.095 46.51 12.265 56.24 ;
      RECT 12.095 121.13 12.265 130.86 ;
      RECT 13.275 121.13 13.445 130.86 ;
      RECT 13.275 78.53 13.445 88.26 ;
      RECT 12.095 78.53 12.265 88.26 ;
      RECT 13.275 57.23 13.445 66.96 ;
      RECT 12.095 57.23 12.265 66.96 ;
      RECT 13.275 67.81 13.445 77.54 ;
      RECT 12.095 67.81 12.265 77.54 ;
      RECT 14.455 121.13 14.625 130.86 ;
      RECT 14.455 110.41 14.625 120.14 ;
      RECT 14.455 99.83 14.625 109.56 ;
      RECT 14.455 89.11 14.625 98.84 ;
      RECT 14.455 46.51 14.625 56.24 ;
      RECT 14.455 78.53 14.625 88.26 ;
      RECT 14.455 57.23 14.625 66.96 ;
      RECT 14.455 67.81 14.625 77.54 ;
      RECT 2.655 153.01 2.825 162.74 ;
      RECT 2.655 142.43 2.825 152.16 ;
      RECT 2.655 131.71 2.825 141.44 ;
      RECT 2.655 185.09 2.825 194.82 ;
      RECT 2.655 174.38 2.825 184.11 ;
      RECT 2.655 163.73 2.825 173.46 ;
      RECT 3.835 153.01 4.005 162.74 ;
      RECT 5.015 153.01 5.185 162.74 ;
      RECT 3.835 142.43 4.005 152.16 ;
      RECT 5.015 142.43 5.185 152.16 ;
      RECT 3.835 131.71 4.005 141.44 ;
      RECT 5.015 131.71 5.185 141.44 ;
      RECT 3.835 185.09 4.005 194.82 ;
      RECT 5.015 185.09 5.185 194.82 ;
      RECT 3.835 174.38 4.005 184.11 ;
      RECT 5.015 174.38 5.185 184.11 ;
      RECT 3.835 163.73 4.005 173.46 ;
      RECT 5.015 163.73 5.185 173.46 ;
      RECT 7.375 163.73 7.545 173.46 ;
      RECT 6.195 153.01 6.365 162.74 ;
      RECT 7.375 153.01 7.545 162.74 ;
      RECT 6.195 142.43 6.365 152.16 ;
      RECT 7.375 142.43 7.545 152.16 ;
      RECT 6.195 131.71 6.365 141.44 ;
      RECT 7.375 131.71 7.545 141.44 ;
      RECT 6.195 185.09 6.365 194.82 ;
      RECT 7.375 185.09 7.545 194.82 ;
      RECT 6.195 174.38 6.365 184.11 ;
      RECT 7.375 174.38 7.545 184.11 ;
      RECT 6.195 163.73 6.365 173.46 ;
      RECT 8.555 163.73 8.725 173.46 ;
      RECT 9.735 163.73 9.905 173.46 ;
      RECT 10.915 163.73 11.085 173.46 ;
      RECT 8.555 153.01 8.725 162.74 ;
      RECT 9.735 153.01 9.905 162.74 ;
      RECT 10.915 153.01 11.085 162.74 ;
      RECT 8.555 142.43 8.725 152.16 ;
      RECT 9.735 142.43 9.905 152.16 ;
      RECT 10.915 142.43 11.085 152.16 ;
      RECT 8.555 131.71 8.725 141.44 ;
      RECT 9.735 131.71 9.905 141.44 ;
      RECT 10.915 131.71 11.085 141.44 ;
      RECT 8.555 185.09 8.725 194.82 ;
      RECT 8.555 174.38 8.725 184.11 ;
      RECT 9.735 185.09 9.905 194.82 ;
      RECT 10.915 185.09 11.085 194.82 ;
      RECT 9.735 174.38 9.905 184.11 ;
      RECT 10.915 174.38 11.085 184.11 ;
      RECT 12.095 163.73 12.265 173.46 ;
      RECT 13.275 163.73 13.445 173.46 ;
      RECT 12.095 153.01 12.265 162.74 ;
      RECT 13.275 153.01 13.445 162.74 ;
      RECT 12.095 142.43 12.265 152.16 ;
      RECT 13.275 142.43 13.445 152.16 ;
      RECT 12.095 131.71 12.265 141.44 ;
      RECT 13.275 131.71 13.445 141.44 ;
      RECT 12.095 185.09 12.265 194.82 ;
      RECT 13.275 185.09 13.445 194.82 ;
      RECT 12.095 174.38 12.265 184.11 ;
      RECT 2.88 88.6 14.4 88.77 ;
      RECT 2.88 14.05 14.4 14.22 ;
      RECT 2.88 24.7 14.4 24.87 ;
      RECT 2.88 35.35 14.4 35.52 ;
      RECT 2.88 46 14.4 46.17 ;
      RECT 2.88 56.65 14.4 56.82 ;
      RECT 2.88 67.3 14.4 67.47 ;
      RECT 2.88 77.95 14.4 78.12 ;
      RECT 1.865 195.655 15.415 195.955 ;
      RECT 15.115 2.9 15.415 195.655 ;
      RECT 1.865 2.6 15.415 2.9 ;
      RECT 1.865 2.9 2.165 195.655 ;
      RECT 2.88 195.1 14.4 195.27 ;
      RECT 2.88 3.4 14.4 3.57 ;
      RECT 2.88 184.45 14.4 184.62 ;
      RECT 2.88 141.85 14.4 142.02 ;
      RECT 2.88 152.5 14.4 152.67 ;
      RECT 2.88 163.15 14.4 163.32 ;
      RECT 2.88 173.8 14.4 173.97 ;
      RECT 2.88 131.2 14.4 131.37 ;
      RECT 2.88 120.55 14.4 120.72 ;
      RECT 2.88 109.9 14.4 110.07 ;
      RECT 2.88 99.25 14.4 99.42 ;
      RECT 0.6 199.17 16.68 199.4 ;
      RECT 0.6 0.83 0.83 199.17 ;
      RECT 16.45 0.83 16.68 199.17 ;
      RECT 0.6 0.6 16.68 0.83 ;
      RECT 2.655 35.93 2.825 45.66 ;
      RECT 2.655 14.63 2.825 24.36 ;
      RECT 2.655 25.21 2.825 34.94 ;
      RECT 2.655 3.87 2.825 13.6 ;
      RECT 5.015 35.93 5.185 45.66 ;
      RECT 3.835 35.93 4.005 45.66 ;
      RECT 5.015 14.63 5.185 24.36 ;
      RECT 3.835 14.63 4.005 24.36 ;
      RECT 5.015 25.21 5.185 34.94 ;
      RECT 3.835 25.21 4.005 34.94 ;
      RECT 5.015 3.87 5.185 13.6 ;
      RECT 3.835 3.87 4.005 13.6 ;
      RECT 7.375 35.93 7.545 45.66 ;
      RECT 6.195 35.93 6.365 45.66 ;
      RECT 7.375 14.63 7.545 24.36 ;
      RECT 6.195 14.63 6.365 24.36 ;
      RECT 7.375 25.21 7.545 34.94 ;
      RECT 6.195 25.21 6.365 34.94 ;
      RECT 7.375 3.87 7.545 13.6 ;
      RECT 6.195 3.87 6.365 13.6 ;
      RECT 10.915 35.93 11.085 45.66 ;
      RECT 9.735 35.93 9.905 45.66 ;
      RECT 8.555 35.93 8.725 45.66 ;
      RECT 10.915 14.63 11.085 24.36 ;
      RECT 9.735 14.63 9.905 24.36 ;
      RECT 8.555 14.63 8.725 24.36 ;
      RECT 10.915 25.21 11.085 34.94 ;
      RECT 9.735 25.21 9.905 34.94 ;
      RECT 8.555 25.21 8.725 34.94 ;
      RECT 10.915 3.87 11.085 13.6 ;
      RECT 9.735 3.87 9.905 13.6 ;
      RECT 8.555 3.87 8.725 13.6 ;
      RECT 13.275 35.93 13.445 45.66 ;
      RECT 12.095 35.93 12.265 45.66 ;
      RECT 13.275 14.63 13.445 24.36 ;
      RECT 12.095 14.63 12.265 24.36 ;
      RECT 13.275 25.21 13.445 34.94 ;
      RECT 12.095 25.21 12.265 34.94 ;
      RECT 13.275 3.87 13.445 13.6 ;
      RECT 12.095 3.87 12.265 13.6 ;
      RECT 14.455 35.93 14.625 45.66 ;
      RECT 14.455 25.21 14.625 34.94 ;
      RECT 14.455 3.83 14.625 13.56 ;
      RECT 14.455 14.63 14.625 24.36 ;
      RECT 2.655 110.41 2.825 120.14 ;
      RECT 2.655 99.83 2.825 109.56 ;
      RECT 2.655 89.11 2.825 98.84 ;
      RECT 2.655 46.51 2.825 56.24 ;
      RECT 2.655 121.13 2.825 130.86 ;
      RECT 2.655 78.53 2.825 88.26 ;
      RECT 2.655 57.23 2.825 66.96 ;
      RECT 2.655 67.81 2.825 77.54 ;
      RECT 3.835 110.41 4.005 120.14 ;
      RECT 5.015 110.41 5.185 120.14 ;
      RECT 3.835 99.83 4.005 109.56 ;
      RECT 5.015 99.83 5.185 109.56 ;
      RECT 3.835 89.11 4.005 98.84 ;
      RECT 5.015 89.11 5.185 98.84 ;
      RECT 5.015 46.51 5.185 56.24 ;
      RECT 3.835 46.51 4.005 56.24 ;
      RECT 3.835 121.13 4.005 130.86 ;
      RECT 5.015 121.13 5.185 130.86 ;
      RECT 5.015 78.53 5.185 88.26 ;
      RECT 3.835 78.53 4.005 88.26 ;
    LAYER met4 ;
      RECT 0 46.635 17.28 47.435 ;
      RECT 0 57.035 17.28 57.835 ;
      RECT 0 24.835 17.28 25.435 ;
      RECT 0 18.785 17.28 19.385 ;
      RECT 0 46.635 17.28 47.335 ;
      RECT 0 57.135 17.28 57.835 ;
      RECT 0 13.935 17.28 14.535 ;
      RECT 0 30.885 17.28 31.485 ;
      RECT 0 35.735 17.28 36.335 ;
      RECT 0 40.585 17.28 41.185 ;
      RECT 0 68.935 17.28 69.635 ;
      RECT 0 63.085 17.28 63.685 ;
      RECT 0 0 17.28 1.635 ;
      RECT 0 7.885 17.28 8.485 ;
      RECT 0 95.4 17.28 175.385 ;
    LAYER met3 ;
      RECT 0 0 3.175 1.13 ;
      RECT 0 1.13 17.28 200 ;
      RECT 6.775 0 7.175 1.13 ;
      RECT 9.775 0 10.175 1.13 ;
      RECT 13.775 0 17.28 1.13 ;
      RECT 13.875 0 17.28 4.235 ;
      RECT 0 1.23 17.28 200 ;
      RECT 0 0 3.075 4.235 ;
    LAYER met2 ;
      RECT 0 199.19 17.28 200 ;
      RECT 0 0 3.335 191.755 ;
      RECT 3.195 191.755 3.335 191.895 ;
      RECT 6.615 0 7.335 195.175 ;
      RECT 6.615 195.175 7.335 195.315 ;
      RECT 6.755 195.315 7.335 195.455 ;
      RECT 6.755 195.455 10.195 195.71 ;
      RECT 6.755 195.71 9.48 196.425 ;
      RECT 7.865 196.425 8.945 196.565 ;
      RECT 9.615 195.315 10.195 195.455 ;
      RECT 9.615 195.175 10.195 195.315 ;
      RECT 9.615 0 10.335 195.175 ;
      RECT 13.615 0 17.28 191.755 ;
      RECT 3.195 199.19 13.755 200 ;
      RECT 0 0 3.195 200 ;
      RECT 13.755 0 17.28 200 ;
      RECT 6.755 195.595 10.195 195.71 ;
      RECT 6.755 0 7.195 195.595 ;
      RECT 9.755 0 10.195 195.595 ;
      RECT 6.825 195.71 10.125 195.78 ;
      RECT 6.895 195.78 10.055 195.85 ;
      RECT 6.965 195.85 9.985 195.92 ;
      RECT 7.035 195.92 9.915 195.99 ;
      RECT 7.105 195.99 9.845 196.06 ;
      RECT 7.175 196.06 9.775 196.13 ;
      RECT 7.245 196.13 9.705 196.2 ;
      RECT 7.315 196.2 9.635 196.27 ;
      RECT 7.385 196.27 9.565 196.34 ;
      RECT 7.455 196.34 9.495 196.41 ;
      RECT 7.47 196.41 9.48 196.425 ;
    LAYER met5 ;
      RECT 0 0 17.28 1.335 ;
      RECT 0 95.785 17.28 174.985 ;
    LAYER met1 ;
      RECT 0 0 17.28 200 ;
  END
END sky130_fd_io__top_vrefcapv2
  
END LIBRARY
