# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__top_gpio_ovtv2
  CLASS BLOCK ;
  FOREIGN sky130_fd_io__top_gpio_ovtv2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  140.0000 BY  200.0000 ;
  SYMMETRY R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.930000 53.125000 140.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.710000 48.365000 140.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN ANALOG_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.115000 0.000000 8.445000 14.070000 ;
    END
  END ANALOG_EN
  PIN ANALOG_POL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 65.235000 0.000000 65.565000 1.165000 ;
    END
  END ANALOG_POL
  PIN ANALOG_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 51.655000 0.000000 51.985000 8.060000 ;
    END
  END ANALOG_SEL
  PIN DM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.125000 0.000000 129.455000 20.955000 ;
    END
  END DM[0]
  PIN DM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 128.275000 0.000000 128.605000 20.180000 ;
    END
  END DM[1]
  PIN DM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.395000 0.000000 108.725000 20.640000 ;
    END
  END DM[2]
  PIN ENABLE_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.135000 0.000000 22.465000 30.150000 ;
    END
  END ENABLE_H
  PIN ENABLE_INP_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 7.110000 0.000000 7.440000 0.670000 ;
    END
  END ENABLE_INP_H
  PIN ENABLE_VDDA_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.770000 0.000000 9.100000 7.915000 ;
    END
  END ENABLE_VDDA_H
  PIN ENABLE_VDDIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 95.845000 0.000000 96.215000 20.755000 ;
    END
  END ENABLE_VDDIO
  PIN ENABLE_VSWITCH_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 5.765000 0.000000 6.365000 12.470000 ;
    END
  END ENABLE_VSWITCH_H
  PIN HLD_H_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 19.635000 0.000000 19.965000 17.985000 ;
    END
  END HLD_H_N
  PIN HLD_OVR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 27.355000 0.000000 27.685000 14.055000 ;
    END
  END HLD_OVR
  PIN HYS_TRIM
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 45.355000 0.000000 45.685000 8.060000 ;
    END
  END HYS_TRIM
  PIN IB_MODE_SEL[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 86.815000 0.000000 87.145000 20.980000 ;
    END
  END IB_MODE_SEL[0]
  PIN IB_MODE_SEL[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 66.935000 0.000000 67.265000 20.980000 ;
    END
  END IB_MODE_SEL[1]
  PIN IN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 20.380000 0.000000 20.710000 11.310000 ;
    END
  END IN
  PIN INP_DIS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 107.545000 0.000000 107.875000 8.060000 ;
    END
  END INP_DIS
  PIN IN_H
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 24.380000 0.000000 24.710000 0.940000 ;
    END
  END IN_H
  PIN OE_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 124.445000 0.000000 124.775000 8.060000 ;
    END
  END OE_N
  PIN OUT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.125000 0.000000 74.455000 14.865000 ;
    END
  END OUT
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 17.930000 117.530000 86.325000 162.905000 ;
    END
  END PAD
  PIN PAD_A_ESD_0_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.600000 0.000000 2.200000 5.470000 ;
    END
  END PAD_A_ESD_0_H
  PIN PAD_A_ESD_1_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.330000 0.000000 0.930000 71.380000 ;
    END
  END PAD_A_ESD_1_H
  PIN PAD_A_NOESD_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2.885000 0.000000 3.485000 5.900000 ;
    END
  END PAD_A_NOESD_H
  PIN SLEW_CTL[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 66.085000 0.000000 66.415000 20.980000 ;
    END
  END SLEW_CTL[0]
  PIN SLEW_CTL[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.205000 0.000000 46.535000 20.980000 ;
    END
  END SLEW_CTL[1]
  PIN SLOW
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 125.140000 0.000000 125.470000 11.965000 ;
    END
  END SLOW
  PIN TIE_HI_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.975000 0.000000 130.305000 61.655000 ;
    END
  END TIE_HI_ESD
  PIN TIE_LO_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.290000 0.000000 115.890000 39.035000 ;
    END
  END TIE_LO_ESD
  PIN VINREF
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 44.035000 0.000000 44.365000 4.885000 ;
    END
  END VINREF
  PIN VTRIP_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 87.665000 0.000000 87.995000 20.980000 ;
    END
  END VTRIP_SEL
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 138.730000 8.985000 140.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 138.730000 2.135000 140.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 139.035000 15.035000 140.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 138.730000 70.035000 140.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 138.730000 64.185000 140.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 138.730000 47.735000 140.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 138.730000 41.685000 140.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 138.730000 25.935000 140.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 138.730000 58.335000 140.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 138.730000 31.985000 140.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT 0.230000 0.200000 140.000000 199.780000 ;
    LAYER met1 ;
      RECT 0.080000 0.000000 140.000000 199.810000 ;
    LAYER met2 ;
      RECT 0.080000 0.000000 140.000000 199.955000 ;
    LAYER met3 ;
      RECT   0.330000 71.780000 140.000000 199.715000 ;
      RECT   1.330000  5.870000   2.485000   6.300000 ;
      RECT   1.330000  6.300000   5.365000  12.870000 ;
      RECT   1.330000 12.870000   7.715000  14.470000 ;
      RECT   1.330000 14.470000  19.235000  18.385000 ;
      RECT   1.330000 18.385000  21.735000  30.550000 ;
      RECT   1.330000 30.550000 114.890000  39.435000 ;
      RECT   1.330000 39.435000 129.575000  62.055000 ;
      RECT   1.330000 62.055000 140.000000  71.780000 ;
      RECT   3.885000  0.000000   5.365000   6.300000 ;
      RECT   6.765000  1.070000   7.715000  12.870000 ;
      RECT   8.845000  8.315000  19.235000  14.470000 ;
      RECT   9.500000  0.000000  19.235000   8.315000 ;
      RECT  20.365000 11.710000  21.735000  18.385000 ;
      RECT  21.110000  0.000000  21.735000  11.710000 ;
      RECT  22.865000  0.000000  23.980000   1.340000 ;
      RECT  22.865000  1.340000  26.955000  14.455000 ;
      RECT  22.865000 14.455000  45.805000  21.380000 ;
      RECT  22.865000 21.380000 114.890000  30.550000 ;
      RECT  25.110000  0.000000  26.955000   1.340000 ;
      RECT  28.085000  0.000000  43.635000   5.285000 ;
      RECT  28.085000  5.285000  44.955000   8.460000 ;
      RECT  28.085000  8.460000  45.805000  14.455000 ;
      RECT  44.765000  0.000000  44.955000   5.285000 ;
      RECT  46.935000  0.000000  51.255000   8.460000 ;
      RECT  46.935000  8.460000  65.685000  21.380000 ;
      RECT  52.385000  0.000000  64.835000   1.565000 ;
      RECT  52.385000  1.565000  65.685000   8.460000 ;
      RECT  67.665000  0.000000  73.725000  15.265000 ;
      RECT  67.665000 15.265000  86.415000  21.380000 ;
      RECT  74.855000  0.000000  86.415000  15.265000 ;
      RECT  88.395000  0.000000  95.445000  21.155000 ;
      RECT  88.395000 21.155000 114.890000  21.380000 ;
      RECT  96.615000  0.000000 107.145000   8.460000 ;
      RECT  96.615000  8.460000 107.995000  21.040000 ;
      RECT  96.615000 21.040000 114.890000  21.155000 ;
      RECT 109.125000  0.000000 114.890000  21.040000 ;
      RECT 116.290000  0.000000 124.045000   8.460000 ;
      RECT 116.290000  8.460000 124.740000  12.365000 ;
      RECT 116.290000 12.365000 127.875000  20.580000 ;
      RECT 116.290000 20.580000 128.725000  21.355000 ;
      RECT 116.290000 21.355000 129.575000  39.435000 ;
      RECT 125.870000  0.000000 127.875000  12.365000 ;
      RECT 130.705000  0.000000 140.000000  62.055000 ;
    LAYER met4 ;
      RECT 0.000000  1.160000 140.000000  47.965000 ;
      RECT 0.000000 47.965000  99.310000  51.745000 ;
      RECT 0.000000 51.745000 140.000000  52.725000 ;
      RECT 0.000000 52.725000  48.530000  56.505000 ;
      RECT 0.000000 56.505000 140.000000 200.000000 ;
    LAYER met5 ;
      RECT  0.000000   2.135000 137.130000  15.035000 ;
      RECT  0.000000  15.035000 137.435000  19.885000 ;
      RECT  0.000000  19.885000 140.000000  24.335000 ;
      RECT  0.000000  24.335000 137.130000  36.835000 ;
      RECT  0.000000  36.835000 140.000000  40.085000 ;
      RECT  0.000000  40.085000 137.130000  96.585000 ;
      RECT  0.000000  96.585000 140.000000 115.930000 ;
      RECT  0.000000 115.930000  16.330000 164.505000 ;
      RECT  0.000000 164.505000 140.000000 200.000000 ;
      RECT 87.925000 115.930000 140.000000 164.505000 ;
  END
END sky130_fd_io__top_gpio_ovtv2
END LIBRARY
