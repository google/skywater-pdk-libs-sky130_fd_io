/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_IO__TOP_SIO_MACRO_PP_SYMBOL_V
`define SKY130_FD_IO__TOP_SIO_MACRO_PP_SYMBOL_V

/**
 * top_sio_macro: sky130_fd_io__sio_macro consists of two SIO cells
 *                and a reference generator cell.
 *
 * Verilog stub (with power pins) for graphical symbol definition
 * generation.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_io__top_sio_macro (
           //# {{data|Data Signals}}
           input        DFT_REFGEN      ,
           input  [1:0] SLOW            ,
           output [1:0] IN              ,
           input  [1:0] INP_DIS         ,
           output [1:0] IN_H            ,
           input  [1:0] OUT             ,
           inout  [1:0] PAD             ,
           inout  [1:0] PAD_A_ESD_0_H   ,
           inout  [1:0] PAD_A_ESD_1_H   ,
           inout  [1:0] PAD_A_NOESD_H   ,

           //# {{control|Control Signals}}
           inout        AMUXBUS_A       ,
           inout        AMUXBUS_B       ,
           input  [2:0] DM0             ,
           input  [2:0] DM1             ,
           input        ENABLE_H        ,
           input        ENABLE_VDDA_H   ,
           input  [1:0] HLD_H_N         ,
           input        HLD_H_N_REFGEN  ,
           input  [1:0] HLD_OVR         ,
           input  [1:0] IBUF_SEL        ,
           input        IBUF_SEL_REFGEN ,
           input  [1:0] OE_N            ,

           //# {{power|Power}}
           input  [2:0] VOH_SEL         ,
           input  [1:0] VREF_SEL        ,
           input  [1:0] VREG_EN         ,
           input        VREG_EN_REFGEN  ,
           input  [1:0] VTRIP_SEL       ,
           input        VTRIP_SEL_REFGEN,
           inout        VSWITCH         ,
           inout        VCCD            ,
           inout        VCCHIB          ,
           inout        VDDA            ,
           inout        VDDIO           ,
           inout        VDDIO_Q         ,
           inout        VINREF_DFT      ,
           input        VOHREF          ,
           inout        VOUTREF_DFT     ,
           inout        VSSA            ,
           inout        VSSD            ,
           inout        VSSIO           ,
           inout        VSSIO_Q         ,
           output [1:0] TIE_LO_ESD
       );
endmodule

`default_nettype wire
`endif  // SKY130_FD_IO__TOP_SIO_MACRO_PP_SYMBOL_V
