# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_io__overlay_vssa_lvc
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 198 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 1.270000 54.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 1.270000 49.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 6.885000 1.270000 11.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 6.885000 75.000000 11.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 6.985000 1.270000 11.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 0.035000 1.270000 5.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 0.035000 75.000000 5.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 0.135000 1.270000 5.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 12.935000 0.965000 16.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 12.935000 75.000000 16.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 13.035000 0.965000 16.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 13.035000 75.000000 16.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 17.785000 1.270000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 68.035000 1.270000 93.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 17.785000 75.000000 22.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 68.035000 75.000000 93.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 17.885000 1.270000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 68.035000 1.270000 92.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 17.885000 75.000000 22.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 62.085000 1.270000 66.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 62.085000 75.000000 66.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 62.185000 1.270000 66.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.500000 34.740000 24.400000 38.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500000 49.650000 24.400000 50.820000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000 34.740000 74.655000 38.180000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755000 49.650000 74.655000 50.820000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 34.735000 24.375000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 45.735000 1.270000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 49.645000 24.375000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 54.405000 1.270000 54.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.780000 34.735000 75.000000 38.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.780000 49.645000 75.000000 50.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 45.735000 75.000000 46.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 54.405000 75.000000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 34.840000 1.270000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 45.735000 1.270000 54.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 34.840000 75.000000 38.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.590000 34.820000  0.790000 35.020000 ;
        RECT  0.590000 35.260000  0.790000 35.460000 ;
        RECT  0.590000 35.700000  0.790000 35.900000 ;
        RECT  0.590000 36.140000  0.790000 36.340000 ;
        RECT  0.590000 36.580000  0.790000 36.780000 ;
        RECT  0.590000 37.020000  0.790000 37.220000 ;
        RECT  0.590000 37.460000  0.790000 37.660000 ;
        RECT  0.590000 37.900000  0.790000 38.100000 ;
        RECT  0.590000 49.715000  0.790000 49.915000 ;
        RECT  0.590000 50.135000  0.790000 50.335000 ;
        RECT  0.590000 50.555000  0.790000 50.755000 ;
        RECT  1.000000 34.820000  1.200000 35.020000 ;
        RECT  1.000000 35.260000  1.200000 35.460000 ;
        RECT  1.000000 35.700000  1.200000 35.900000 ;
        RECT  1.000000 36.140000  1.200000 36.340000 ;
        RECT  1.000000 36.580000  1.200000 36.780000 ;
        RECT  1.000000 37.020000  1.200000 37.220000 ;
        RECT  1.000000 37.460000  1.200000 37.660000 ;
        RECT  1.000000 37.900000  1.200000 38.100000 ;
        RECT  1.000000 49.715000  1.200000 49.915000 ;
        RECT  1.000000 50.135000  1.200000 50.335000 ;
        RECT  1.000000 50.555000  1.200000 50.755000 ;
        RECT  1.410000 34.820000  1.610000 35.020000 ;
        RECT  1.410000 35.260000  1.610000 35.460000 ;
        RECT  1.410000 35.700000  1.610000 35.900000 ;
        RECT  1.410000 36.140000  1.610000 36.340000 ;
        RECT  1.410000 36.580000  1.610000 36.780000 ;
        RECT  1.410000 37.020000  1.610000 37.220000 ;
        RECT  1.410000 37.460000  1.610000 37.660000 ;
        RECT  1.410000 37.900000  1.610000 38.100000 ;
        RECT  1.410000 49.715000  1.610000 49.915000 ;
        RECT  1.410000 50.135000  1.610000 50.335000 ;
        RECT  1.410000 50.555000  1.610000 50.755000 ;
        RECT  1.820000 34.820000  2.020000 35.020000 ;
        RECT  1.820000 35.260000  2.020000 35.460000 ;
        RECT  1.820000 35.700000  2.020000 35.900000 ;
        RECT  1.820000 36.140000  2.020000 36.340000 ;
        RECT  1.820000 36.580000  2.020000 36.780000 ;
        RECT  1.820000 37.020000  2.020000 37.220000 ;
        RECT  1.820000 37.460000  2.020000 37.660000 ;
        RECT  1.820000 37.900000  2.020000 38.100000 ;
        RECT  1.820000 49.715000  2.020000 49.915000 ;
        RECT  1.820000 50.135000  2.020000 50.335000 ;
        RECT  1.820000 50.555000  2.020000 50.755000 ;
        RECT  2.230000 34.820000  2.430000 35.020000 ;
        RECT  2.230000 35.260000  2.430000 35.460000 ;
        RECT  2.230000 35.700000  2.430000 35.900000 ;
        RECT  2.230000 36.140000  2.430000 36.340000 ;
        RECT  2.230000 36.580000  2.430000 36.780000 ;
        RECT  2.230000 37.020000  2.430000 37.220000 ;
        RECT  2.230000 37.460000  2.430000 37.660000 ;
        RECT  2.230000 37.900000  2.430000 38.100000 ;
        RECT  2.230000 49.715000  2.430000 49.915000 ;
        RECT  2.230000 50.135000  2.430000 50.335000 ;
        RECT  2.230000 50.555000  2.430000 50.755000 ;
        RECT  2.640000 34.820000  2.840000 35.020000 ;
        RECT  2.640000 35.260000  2.840000 35.460000 ;
        RECT  2.640000 35.700000  2.840000 35.900000 ;
        RECT  2.640000 36.140000  2.840000 36.340000 ;
        RECT  2.640000 36.580000  2.840000 36.780000 ;
        RECT  2.640000 37.020000  2.840000 37.220000 ;
        RECT  2.640000 37.460000  2.840000 37.660000 ;
        RECT  2.640000 37.900000  2.840000 38.100000 ;
        RECT  2.640000 49.715000  2.840000 49.915000 ;
        RECT  2.640000 50.135000  2.840000 50.335000 ;
        RECT  2.640000 50.555000  2.840000 50.755000 ;
        RECT  3.050000 34.820000  3.250000 35.020000 ;
        RECT  3.050000 35.260000  3.250000 35.460000 ;
        RECT  3.050000 35.700000  3.250000 35.900000 ;
        RECT  3.050000 36.140000  3.250000 36.340000 ;
        RECT  3.050000 36.580000  3.250000 36.780000 ;
        RECT  3.050000 37.020000  3.250000 37.220000 ;
        RECT  3.050000 37.460000  3.250000 37.660000 ;
        RECT  3.050000 37.900000  3.250000 38.100000 ;
        RECT  3.050000 49.715000  3.250000 49.915000 ;
        RECT  3.050000 50.135000  3.250000 50.335000 ;
        RECT  3.050000 50.555000  3.250000 50.755000 ;
        RECT  3.455000 34.820000  3.655000 35.020000 ;
        RECT  3.455000 35.260000  3.655000 35.460000 ;
        RECT  3.455000 35.700000  3.655000 35.900000 ;
        RECT  3.455000 36.140000  3.655000 36.340000 ;
        RECT  3.455000 36.580000  3.655000 36.780000 ;
        RECT  3.455000 37.020000  3.655000 37.220000 ;
        RECT  3.455000 37.460000  3.655000 37.660000 ;
        RECT  3.455000 37.900000  3.655000 38.100000 ;
        RECT  3.455000 49.715000  3.655000 49.915000 ;
        RECT  3.455000 50.135000  3.655000 50.335000 ;
        RECT  3.455000 50.555000  3.655000 50.755000 ;
        RECT  3.860000 34.820000  4.060000 35.020000 ;
        RECT  3.860000 35.260000  4.060000 35.460000 ;
        RECT  3.860000 35.700000  4.060000 35.900000 ;
        RECT  3.860000 36.140000  4.060000 36.340000 ;
        RECT  3.860000 36.580000  4.060000 36.780000 ;
        RECT  3.860000 37.020000  4.060000 37.220000 ;
        RECT  3.860000 37.460000  4.060000 37.660000 ;
        RECT  3.860000 37.900000  4.060000 38.100000 ;
        RECT  3.860000 49.715000  4.060000 49.915000 ;
        RECT  3.860000 50.135000  4.060000 50.335000 ;
        RECT  3.860000 50.555000  4.060000 50.755000 ;
        RECT  4.265000 34.820000  4.465000 35.020000 ;
        RECT  4.265000 35.260000  4.465000 35.460000 ;
        RECT  4.265000 35.700000  4.465000 35.900000 ;
        RECT  4.265000 36.140000  4.465000 36.340000 ;
        RECT  4.265000 36.580000  4.465000 36.780000 ;
        RECT  4.265000 37.020000  4.465000 37.220000 ;
        RECT  4.265000 37.460000  4.465000 37.660000 ;
        RECT  4.265000 37.900000  4.465000 38.100000 ;
        RECT  4.265000 49.715000  4.465000 49.915000 ;
        RECT  4.265000 50.135000  4.465000 50.335000 ;
        RECT  4.265000 50.555000  4.465000 50.755000 ;
        RECT  4.670000 34.820000  4.870000 35.020000 ;
        RECT  4.670000 35.260000  4.870000 35.460000 ;
        RECT  4.670000 35.700000  4.870000 35.900000 ;
        RECT  4.670000 36.140000  4.870000 36.340000 ;
        RECT  4.670000 36.580000  4.870000 36.780000 ;
        RECT  4.670000 37.020000  4.870000 37.220000 ;
        RECT  4.670000 37.460000  4.870000 37.660000 ;
        RECT  4.670000 37.900000  4.870000 38.100000 ;
        RECT  4.670000 49.715000  4.870000 49.915000 ;
        RECT  4.670000 50.135000  4.870000 50.335000 ;
        RECT  4.670000 50.555000  4.870000 50.755000 ;
        RECT  5.075000 34.820000  5.275000 35.020000 ;
        RECT  5.075000 35.260000  5.275000 35.460000 ;
        RECT  5.075000 35.700000  5.275000 35.900000 ;
        RECT  5.075000 36.140000  5.275000 36.340000 ;
        RECT  5.075000 36.580000  5.275000 36.780000 ;
        RECT  5.075000 37.020000  5.275000 37.220000 ;
        RECT  5.075000 37.460000  5.275000 37.660000 ;
        RECT  5.075000 37.900000  5.275000 38.100000 ;
        RECT  5.075000 49.715000  5.275000 49.915000 ;
        RECT  5.075000 50.135000  5.275000 50.335000 ;
        RECT  5.075000 50.555000  5.275000 50.755000 ;
        RECT  5.480000 34.820000  5.680000 35.020000 ;
        RECT  5.480000 35.260000  5.680000 35.460000 ;
        RECT  5.480000 35.700000  5.680000 35.900000 ;
        RECT  5.480000 36.140000  5.680000 36.340000 ;
        RECT  5.480000 36.580000  5.680000 36.780000 ;
        RECT  5.480000 37.020000  5.680000 37.220000 ;
        RECT  5.480000 37.460000  5.680000 37.660000 ;
        RECT  5.480000 37.900000  5.680000 38.100000 ;
        RECT  5.480000 49.715000  5.680000 49.915000 ;
        RECT  5.480000 50.135000  5.680000 50.335000 ;
        RECT  5.480000 50.555000  5.680000 50.755000 ;
        RECT  5.885000 34.820000  6.085000 35.020000 ;
        RECT  5.885000 35.260000  6.085000 35.460000 ;
        RECT  5.885000 35.700000  6.085000 35.900000 ;
        RECT  5.885000 36.140000  6.085000 36.340000 ;
        RECT  5.885000 36.580000  6.085000 36.780000 ;
        RECT  5.885000 37.020000  6.085000 37.220000 ;
        RECT  5.885000 37.460000  6.085000 37.660000 ;
        RECT  5.885000 37.900000  6.085000 38.100000 ;
        RECT  5.885000 49.715000  6.085000 49.915000 ;
        RECT  5.885000 50.135000  6.085000 50.335000 ;
        RECT  5.885000 50.555000  6.085000 50.755000 ;
        RECT  6.290000 34.820000  6.490000 35.020000 ;
        RECT  6.290000 35.260000  6.490000 35.460000 ;
        RECT  6.290000 35.700000  6.490000 35.900000 ;
        RECT  6.290000 36.140000  6.490000 36.340000 ;
        RECT  6.290000 36.580000  6.490000 36.780000 ;
        RECT  6.290000 37.020000  6.490000 37.220000 ;
        RECT  6.290000 37.460000  6.490000 37.660000 ;
        RECT  6.290000 37.900000  6.490000 38.100000 ;
        RECT  6.290000 49.715000  6.490000 49.915000 ;
        RECT  6.290000 50.135000  6.490000 50.335000 ;
        RECT  6.290000 50.555000  6.490000 50.755000 ;
        RECT  6.695000 34.820000  6.895000 35.020000 ;
        RECT  6.695000 35.260000  6.895000 35.460000 ;
        RECT  6.695000 35.700000  6.895000 35.900000 ;
        RECT  6.695000 36.140000  6.895000 36.340000 ;
        RECT  6.695000 36.580000  6.895000 36.780000 ;
        RECT  6.695000 37.020000  6.895000 37.220000 ;
        RECT  6.695000 37.460000  6.895000 37.660000 ;
        RECT  6.695000 37.900000  6.895000 38.100000 ;
        RECT  6.695000 49.715000  6.895000 49.915000 ;
        RECT  6.695000 50.135000  6.895000 50.335000 ;
        RECT  6.695000 50.555000  6.895000 50.755000 ;
        RECT  7.100000 34.820000  7.300000 35.020000 ;
        RECT  7.100000 35.260000  7.300000 35.460000 ;
        RECT  7.100000 35.700000  7.300000 35.900000 ;
        RECT  7.100000 36.140000  7.300000 36.340000 ;
        RECT  7.100000 36.580000  7.300000 36.780000 ;
        RECT  7.100000 37.020000  7.300000 37.220000 ;
        RECT  7.100000 37.460000  7.300000 37.660000 ;
        RECT  7.100000 37.900000  7.300000 38.100000 ;
        RECT  7.100000 49.715000  7.300000 49.915000 ;
        RECT  7.100000 50.135000  7.300000 50.335000 ;
        RECT  7.100000 50.555000  7.300000 50.755000 ;
        RECT  7.505000 34.820000  7.705000 35.020000 ;
        RECT  7.505000 35.260000  7.705000 35.460000 ;
        RECT  7.505000 35.700000  7.705000 35.900000 ;
        RECT  7.505000 36.140000  7.705000 36.340000 ;
        RECT  7.505000 36.580000  7.705000 36.780000 ;
        RECT  7.505000 37.020000  7.705000 37.220000 ;
        RECT  7.505000 37.460000  7.705000 37.660000 ;
        RECT  7.505000 37.900000  7.705000 38.100000 ;
        RECT  7.505000 49.715000  7.705000 49.915000 ;
        RECT  7.505000 50.135000  7.705000 50.335000 ;
        RECT  7.505000 50.555000  7.705000 50.755000 ;
        RECT  7.910000 34.820000  8.110000 35.020000 ;
        RECT  7.910000 35.260000  8.110000 35.460000 ;
        RECT  7.910000 35.700000  8.110000 35.900000 ;
        RECT  7.910000 36.140000  8.110000 36.340000 ;
        RECT  7.910000 36.580000  8.110000 36.780000 ;
        RECT  7.910000 37.020000  8.110000 37.220000 ;
        RECT  7.910000 37.460000  8.110000 37.660000 ;
        RECT  7.910000 37.900000  8.110000 38.100000 ;
        RECT  7.910000 49.715000  8.110000 49.915000 ;
        RECT  7.910000 50.135000  8.110000 50.335000 ;
        RECT  7.910000 50.555000  8.110000 50.755000 ;
        RECT  8.315000 34.820000  8.515000 35.020000 ;
        RECT  8.315000 35.260000  8.515000 35.460000 ;
        RECT  8.315000 35.700000  8.515000 35.900000 ;
        RECT  8.315000 36.140000  8.515000 36.340000 ;
        RECT  8.315000 36.580000  8.515000 36.780000 ;
        RECT  8.315000 37.020000  8.515000 37.220000 ;
        RECT  8.315000 37.460000  8.515000 37.660000 ;
        RECT  8.315000 37.900000  8.515000 38.100000 ;
        RECT  8.315000 49.715000  8.515000 49.915000 ;
        RECT  8.315000 50.135000  8.515000 50.335000 ;
        RECT  8.315000 50.555000  8.515000 50.755000 ;
        RECT  8.720000 34.820000  8.920000 35.020000 ;
        RECT  8.720000 35.260000  8.920000 35.460000 ;
        RECT  8.720000 35.700000  8.920000 35.900000 ;
        RECT  8.720000 36.140000  8.920000 36.340000 ;
        RECT  8.720000 36.580000  8.920000 36.780000 ;
        RECT  8.720000 37.020000  8.920000 37.220000 ;
        RECT  8.720000 37.460000  8.920000 37.660000 ;
        RECT  8.720000 37.900000  8.920000 38.100000 ;
        RECT  8.720000 49.715000  8.920000 49.915000 ;
        RECT  8.720000 50.135000  8.920000 50.335000 ;
        RECT  8.720000 50.555000  8.920000 50.755000 ;
        RECT  9.125000 34.820000  9.325000 35.020000 ;
        RECT  9.125000 35.260000  9.325000 35.460000 ;
        RECT  9.125000 35.700000  9.325000 35.900000 ;
        RECT  9.125000 36.140000  9.325000 36.340000 ;
        RECT  9.125000 36.580000  9.325000 36.780000 ;
        RECT  9.125000 37.020000  9.325000 37.220000 ;
        RECT  9.125000 37.460000  9.325000 37.660000 ;
        RECT  9.125000 37.900000  9.325000 38.100000 ;
        RECT  9.125000 49.715000  9.325000 49.915000 ;
        RECT  9.125000 50.135000  9.325000 50.335000 ;
        RECT  9.125000 50.555000  9.325000 50.755000 ;
        RECT  9.530000 34.820000  9.730000 35.020000 ;
        RECT  9.530000 35.260000  9.730000 35.460000 ;
        RECT  9.530000 35.700000  9.730000 35.900000 ;
        RECT  9.530000 36.140000  9.730000 36.340000 ;
        RECT  9.530000 36.580000  9.730000 36.780000 ;
        RECT  9.530000 37.020000  9.730000 37.220000 ;
        RECT  9.530000 37.460000  9.730000 37.660000 ;
        RECT  9.530000 37.900000  9.730000 38.100000 ;
        RECT  9.530000 49.715000  9.730000 49.915000 ;
        RECT  9.530000 50.135000  9.730000 50.335000 ;
        RECT  9.530000 50.555000  9.730000 50.755000 ;
        RECT  9.935000 34.820000 10.135000 35.020000 ;
        RECT  9.935000 35.260000 10.135000 35.460000 ;
        RECT  9.935000 35.700000 10.135000 35.900000 ;
        RECT  9.935000 36.140000 10.135000 36.340000 ;
        RECT  9.935000 36.580000 10.135000 36.780000 ;
        RECT  9.935000 37.020000 10.135000 37.220000 ;
        RECT  9.935000 37.460000 10.135000 37.660000 ;
        RECT  9.935000 37.900000 10.135000 38.100000 ;
        RECT  9.935000 49.715000 10.135000 49.915000 ;
        RECT  9.935000 50.135000 10.135000 50.335000 ;
        RECT  9.935000 50.555000 10.135000 50.755000 ;
        RECT 10.340000 34.820000 10.540000 35.020000 ;
        RECT 10.340000 35.260000 10.540000 35.460000 ;
        RECT 10.340000 35.700000 10.540000 35.900000 ;
        RECT 10.340000 36.140000 10.540000 36.340000 ;
        RECT 10.340000 36.580000 10.540000 36.780000 ;
        RECT 10.340000 37.020000 10.540000 37.220000 ;
        RECT 10.340000 37.460000 10.540000 37.660000 ;
        RECT 10.340000 37.900000 10.540000 38.100000 ;
        RECT 10.340000 49.715000 10.540000 49.915000 ;
        RECT 10.340000 50.135000 10.540000 50.335000 ;
        RECT 10.340000 50.555000 10.540000 50.755000 ;
        RECT 10.745000 34.820000 10.945000 35.020000 ;
        RECT 10.745000 35.260000 10.945000 35.460000 ;
        RECT 10.745000 35.700000 10.945000 35.900000 ;
        RECT 10.745000 36.140000 10.945000 36.340000 ;
        RECT 10.745000 36.580000 10.945000 36.780000 ;
        RECT 10.745000 37.020000 10.945000 37.220000 ;
        RECT 10.745000 37.460000 10.945000 37.660000 ;
        RECT 10.745000 37.900000 10.945000 38.100000 ;
        RECT 10.745000 49.715000 10.945000 49.915000 ;
        RECT 10.745000 50.135000 10.945000 50.335000 ;
        RECT 10.745000 50.555000 10.945000 50.755000 ;
        RECT 11.150000 34.820000 11.350000 35.020000 ;
        RECT 11.150000 35.260000 11.350000 35.460000 ;
        RECT 11.150000 35.700000 11.350000 35.900000 ;
        RECT 11.150000 36.140000 11.350000 36.340000 ;
        RECT 11.150000 36.580000 11.350000 36.780000 ;
        RECT 11.150000 37.020000 11.350000 37.220000 ;
        RECT 11.150000 37.460000 11.350000 37.660000 ;
        RECT 11.150000 37.900000 11.350000 38.100000 ;
        RECT 11.150000 49.715000 11.350000 49.915000 ;
        RECT 11.150000 50.135000 11.350000 50.335000 ;
        RECT 11.150000 50.555000 11.350000 50.755000 ;
        RECT 11.555000 34.820000 11.755000 35.020000 ;
        RECT 11.555000 35.260000 11.755000 35.460000 ;
        RECT 11.555000 35.700000 11.755000 35.900000 ;
        RECT 11.555000 36.140000 11.755000 36.340000 ;
        RECT 11.555000 36.580000 11.755000 36.780000 ;
        RECT 11.555000 37.020000 11.755000 37.220000 ;
        RECT 11.555000 37.460000 11.755000 37.660000 ;
        RECT 11.555000 37.900000 11.755000 38.100000 ;
        RECT 11.555000 49.715000 11.755000 49.915000 ;
        RECT 11.555000 50.135000 11.755000 50.335000 ;
        RECT 11.555000 50.555000 11.755000 50.755000 ;
        RECT 11.960000 34.820000 12.160000 35.020000 ;
        RECT 11.960000 35.260000 12.160000 35.460000 ;
        RECT 11.960000 35.700000 12.160000 35.900000 ;
        RECT 11.960000 36.140000 12.160000 36.340000 ;
        RECT 11.960000 36.580000 12.160000 36.780000 ;
        RECT 11.960000 37.020000 12.160000 37.220000 ;
        RECT 11.960000 37.460000 12.160000 37.660000 ;
        RECT 11.960000 37.900000 12.160000 38.100000 ;
        RECT 11.960000 49.715000 12.160000 49.915000 ;
        RECT 11.960000 50.135000 12.160000 50.335000 ;
        RECT 11.960000 50.555000 12.160000 50.755000 ;
        RECT 12.365000 34.820000 12.565000 35.020000 ;
        RECT 12.365000 35.260000 12.565000 35.460000 ;
        RECT 12.365000 35.700000 12.565000 35.900000 ;
        RECT 12.365000 36.140000 12.565000 36.340000 ;
        RECT 12.365000 36.580000 12.565000 36.780000 ;
        RECT 12.365000 37.020000 12.565000 37.220000 ;
        RECT 12.365000 37.460000 12.565000 37.660000 ;
        RECT 12.365000 37.900000 12.565000 38.100000 ;
        RECT 12.365000 49.715000 12.565000 49.915000 ;
        RECT 12.365000 50.135000 12.565000 50.335000 ;
        RECT 12.365000 50.555000 12.565000 50.755000 ;
        RECT 12.770000 34.820000 12.970000 35.020000 ;
        RECT 12.770000 35.260000 12.970000 35.460000 ;
        RECT 12.770000 35.700000 12.970000 35.900000 ;
        RECT 12.770000 36.140000 12.970000 36.340000 ;
        RECT 12.770000 36.580000 12.970000 36.780000 ;
        RECT 12.770000 37.020000 12.970000 37.220000 ;
        RECT 12.770000 37.460000 12.970000 37.660000 ;
        RECT 12.770000 37.900000 12.970000 38.100000 ;
        RECT 12.770000 49.715000 12.970000 49.915000 ;
        RECT 12.770000 50.135000 12.970000 50.335000 ;
        RECT 12.770000 50.555000 12.970000 50.755000 ;
        RECT 13.175000 34.820000 13.375000 35.020000 ;
        RECT 13.175000 35.260000 13.375000 35.460000 ;
        RECT 13.175000 35.700000 13.375000 35.900000 ;
        RECT 13.175000 36.140000 13.375000 36.340000 ;
        RECT 13.175000 36.580000 13.375000 36.780000 ;
        RECT 13.175000 37.020000 13.375000 37.220000 ;
        RECT 13.175000 37.460000 13.375000 37.660000 ;
        RECT 13.175000 37.900000 13.375000 38.100000 ;
        RECT 13.175000 49.715000 13.375000 49.915000 ;
        RECT 13.175000 50.135000 13.375000 50.335000 ;
        RECT 13.175000 50.555000 13.375000 50.755000 ;
        RECT 13.580000 34.820000 13.780000 35.020000 ;
        RECT 13.580000 35.260000 13.780000 35.460000 ;
        RECT 13.580000 35.700000 13.780000 35.900000 ;
        RECT 13.580000 36.140000 13.780000 36.340000 ;
        RECT 13.580000 36.580000 13.780000 36.780000 ;
        RECT 13.580000 37.020000 13.780000 37.220000 ;
        RECT 13.580000 37.460000 13.780000 37.660000 ;
        RECT 13.580000 37.900000 13.780000 38.100000 ;
        RECT 13.580000 49.715000 13.780000 49.915000 ;
        RECT 13.580000 50.135000 13.780000 50.335000 ;
        RECT 13.580000 50.555000 13.780000 50.755000 ;
        RECT 13.985000 34.820000 14.185000 35.020000 ;
        RECT 13.985000 35.260000 14.185000 35.460000 ;
        RECT 13.985000 35.700000 14.185000 35.900000 ;
        RECT 13.985000 36.140000 14.185000 36.340000 ;
        RECT 13.985000 36.580000 14.185000 36.780000 ;
        RECT 13.985000 37.020000 14.185000 37.220000 ;
        RECT 13.985000 37.460000 14.185000 37.660000 ;
        RECT 13.985000 37.900000 14.185000 38.100000 ;
        RECT 13.985000 49.715000 14.185000 49.915000 ;
        RECT 13.985000 50.135000 14.185000 50.335000 ;
        RECT 13.985000 50.555000 14.185000 50.755000 ;
        RECT 14.390000 34.820000 14.590000 35.020000 ;
        RECT 14.390000 35.260000 14.590000 35.460000 ;
        RECT 14.390000 35.700000 14.590000 35.900000 ;
        RECT 14.390000 36.140000 14.590000 36.340000 ;
        RECT 14.390000 36.580000 14.590000 36.780000 ;
        RECT 14.390000 37.020000 14.590000 37.220000 ;
        RECT 14.390000 37.460000 14.590000 37.660000 ;
        RECT 14.390000 37.900000 14.590000 38.100000 ;
        RECT 14.390000 49.715000 14.590000 49.915000 ;
        RECT 14.390000 50.135000 14.590000 50.335000 ;
        RECT 14.390000 50.555000 14.590000 50.755000 ;
        RECT 14.795000 34.820000 14.995000 35.020000 ;
        RECT 14.795000 35.260000 14.995000 35.460000 ;
        RECT 14.795000 35.700000 14.995000 35.900000 ;
        RECT 14.795000 36.140000 14.995000 36.340000 ;
        RECT 14.795000 36.580000 14.995000 36.780000 ;
        RECT 14.795000 37.020000 14.995000 37.220000 ;
        RECT 14.795000 37.460000 14.995000 37.660000 ;
        RECT 14.795000 37.900000 14.995000 38.100000 ;
        RECT 14.795000 49.715000 14.995000 49.915000 ;
        RECT 14.795000 50.135000 14.995000 50.335000 ;
        RECT 14.795000 50.555000 14.995000 50.755000 ;
        RECT 15.200000 34.820000 15.400000 35.020000 ;
        RECT 15.200000 35.260000 15.400000 35.460000 ;
        RECT 15.200000 35.700000 15.400000 35.900000 ;
        RECT 15.200000 36.140000 15.400000 36.340000 ;
        RECT 15.200000 36.580000 15.400000 36.780000 ;
        RECT 15.200000 37.020000 15.400000 37.220000 ;
        RECT 15.200000 37.460000 15.400000 37.660000 ;
        RECT 15.200000 37.900000 15.400000 38.100000 ;
        RECT 15.200000 49.715000 15.400000 49.915000 ;
        RECT 15.200000 50.135000 15.400000 50.335000 ;
        RECT 15.200000 50.555000 15.400000 50.755000 ;
        RECT 15.605000 34.820000 15.805000 35.020000 ;
        RECT 15.605000 35.260000 15.805000 35.460000 ;
        RECT 15.605000 35.700000 15.805000 35.900000 ;
        RECT 15.605000 36.140000 15.805000 36.340000 ;
        RECT 15.605000 36.580000 15.805000 36.780000 ;
        RECT 15.605000 37.020000 15.805000 37.220000 ;
        RECT 15.605000 37.460000 15.805000 37.660000 ;
        RECT 15.605000 37.900000 15.805000 38.100000 ;
        RECT 15.605000 49.715000 15.805000 49.915000 ;
        RECT 15.605000 50.135000 15.805000 50.335000 ;
        RECT 15.605000 50.555000 15.805000 50.755000 ;
        RECT 16.010000 34.820000 16.210000 35.020000 ;
        RECT 16.010000 35.260000 16.210000 35.460000 ;
        RECT 16.010000 35.700000 16.210000 35.900000 ;
        RECT 16.010000 36.140000 16.210000 36.340000 ;
        RECT 16.010000 36.580000 16.210000 36.780000 ;
        RECT 16.010000 37.020000 16.210000 37.220000 ;
        RECT 16.010000 37.460000 16.210000 37.660000 ;
        RECT 16.010000 37.900000 16.210000 38.100000 ;
        RECT 16.010000 49.715000 16.210000 49.915000 ;
        RECT 16.010000 50.135000 16.210000 50.335000 ;
        RECT 16.010000 50.555000 16.210000 50.755000 ;
        RECT 16.415000 34.820000 16.615000 35.020000 ;
        RECT 16.415000 35.260000 16.615000 35.460000 ;
        RECT 16.415000 35.700000 16.615000 35.900000 ;
        RECT 16.415000 36.140000 16.615000 36.340000 ;
        RECT 16.415000 36.580000 16.615000 36.780000 ;
        RECT 16.415000 37.020000 16.615000 37.220000 ;
        RECT 16.415000 37.460000 16.615000 37.660000 ;
        RECT 16.415000 37.900000 16.615000 38.100000 ;
        RECT 16.415000 49.715000 16.615000 49.915000 ;
        RECT 16.415000 50.135000 16.615000 50.335000 ;
        RECT 16.415000 50.555000 16.615000 50.755000 ;
        RECT 16.820000 34.820000 17.020000 35.020000 ;
        RECT 16.820000 35.260000 17.020000 35.460000 ;
        RECT 16.820000 35.700000 17.020000 35.900000 ;
        RECT 16.820000 36.140000 17.020000 36.340000 ;
        RECT 16.820000 36.580000 17.020000 36.780000 ;
        RECT 16.820000 37.020000 17.020000 37.220000 ;
        RECT 16.820000 37.460000 17.020000 37.660000 ;
        RECT 16.820000 37.900000 17.020000 38.100000 ;
        RECT 16.820000 49.715000 17.020000 49.915000 ;
        RECT 16.820000 50.135000 17.020000 50.335000 ;
        RECT 16.820000 50.555000 17.020000 50.755000 ;
        RECT 17.225000 34.820000 17.425000 35.020000 ;
        RECT 17.225000 35.260000 17.425000 35.460000 ;
        RECT 17.225000 35.700000 17.425000 35.900000 ;
        RECT 17.225000 36.140000 17.425000 36.340000 ;
        RECT 17.225000 36.580000 17.425000 36.780000 ;
        RECT 17.225000 37.020000 17.425000 37.220000 ;
        RECT 17.225000 37.460000 17.425000 37.660000 ;
        RECT 17.225000 37.900000 17.425000 38.100000 ;
        RECT 17.225000 49.715000 17.425000 49.915000 ;
        RECT 17.225000 50.135000 17.425000 50.335000 ;
        RECT 17.225000 50.555000 17.425000 50.755000 ;
        RECT 17.630000 34.820000 17.830000 35.020000 ;
        RECT 17.630000 35.260000 17.830000 35.460000 ;
        RECT 17.630000 35.700000 17.830000 35.900000 ;
        RECT 17.630000 36.140000 17.830000 36.340000 ;
        RECT 17.630000 36.580000 17.830000 36.780000 ;
        RECT 17.630000 37.020000 17.830000 37.220000 ;
        RECT 17.630000 37.460000 17.830000 37.660000 ;
        RECT 17.630000 37.900000 17.830000 38.100000 ;
        RECT 17.630000 49.715000 17.830000 49.915000 ;
        RECT 17.630000 50.135000 17.830000 50.335000 ;
        RECT 17.630000 50.555000 17.830000 50.755000 ;
        RECT 18.035000 34.820000 18.235000 35.020000 ;
        RECT 18.035000 35.260000 18.235000 35.460000 ;
        RECT 18.035000 35.700000 18.235000 35.900000 ;
        RECT 18.035000 36.140000 18.235000 36.340000 ;
        RECT 18.035000 36.580000 18.235000 36.780000 ;
        RECT 18.035000 37.020000 18.235000 37.220000 ;
        RECT 18.035000 37.460000 18.235000 37.660000 ;
        RECT 18.035000 37.900000 18.235000 38.100000 ;
        RECT 18.035000 49.715000 18.235000 49.915000 ;
        RECT 18.035000 50.135000 18.235000 50.335000 ;
        RECT 18.035000 50.555000 18.235000 50.755000 ;
        RECT 18.440000 34.820000 18.640000 35.020000 ;
        RECT 18.440000 35.260000 18.640000 35.460000 ;
        RECT 18.440000 35.700000 18.640000 35.900000 ;
        RECT 18.440000 36.140000 18.640000 36.340000 ;
        RECT 18.440000 36.580000 18.640000 36.780000 ;
        RECT 18.440000 37.020000 18.640000 37.220000 ;
        RECT 18.440000 37.460000 18.640000 37.660000 ;
        RECT 18.440000 37.900000 18.640000 38.100000 ;
        RECT 18.440000 49.715000 18.640000 49.915000 ;
        RECT 18.440000 50.135000 18.640000 50.335000 ;
        RECT 18.440000 50.555000 18.640000 50.755000 ;
        RECT 18.845000 34.820000 19.045000 35.020000 ;
        RECT 18.845000 35.260000 19.045000 35.460000 ;
        RECT 18.845000 35.700000 19.045000 35.900000 ;
        RECT 18.845000 36.140000 19.045000 36.340000 ;
        RECT 18.845000 36.580000 19.045000 36.780000 ;
        RECT 18.845000 37.020000 19.045000 37.220000 ;
        RECT 18.845000 37.460000 19.045000 37.660000 ;
        RECT 18.845000 37.900000 19.045000 38.100000 ;
        RECT 18.845000 49.715000 19.045000 49.915000 ;
        RECT 18.845000 50.135000 19.045000 50.335000 ;
        RECT 18.845000 50.555000 19.045000 50.755000 ;
        RECT 19.250000 34.820000 19.450000 35.020000 ;
        RECT 19.250000 35.260000 19.450000 35.460000 ;
        RECT 19.250000 35.700000 19.450000 35.900000 ;
        RECT 19.250000 36.140000 19.450000 36.340000 ;
        RECT 19.250000 36.580000 19.450000 36.780000 ;
        RECT 19.250000 37.020000 19.450000 37.220000 ;
        RECT 19.250000 37.460000 19.450000 37.660000 ;
        RECT 19.250000 37.900000 19.450000 38.100000 ;
        RECT 19.250000 49.715000 19.450000 49.915000 ;
        RECT 19.250000 50.135000 19.450000 50.335000 ;
        RECT 19.250000 50.555000 19.450000 50.755000 ;
        RECT 19.655000 34.820000 19.855000 35.020000 ;
        RECT 19.655000 35.260000 19.855000 35.460000 ;
        RECT 19.655000 35.700000 19.855000 35.900000 ;
        RECT 19.655000 36.140000 19.855000 36.340000 ;
        RECT 19.655000 36.580000 19.855000 36.780000 ;
        RECT 19.655000 37.020000 19.855000 37.220000 ;
        RECT 19.655000 37.460000 19.855000 37.660000 ;
        RECT 19.655000 37.900000 19.855000 38.100000 ;
        RECT 19.655000 49.715000 19.855000 49.915000 ;
        RECT 19.655000 50.135000 19.855000 50.335000 ;
        RECT 19.655000 50.555000 19.855000 50.755000 ;
        RECT 20.060000 34.820000 20.260000 35.020000 ;
        RECT 20.060000 35.260000 20.260000 35.460000 ;
        RECT 20.060000 35.700000 20.260000 35.900000 ;
        RECT 20.060000 36.140000 20.260000 36.340000 ;
        RECT 20.060000 36.580000 20.260000 36.780000 ;
        RECT 20.060000 37.020000 20.260000 37.220000 ;
        RECT 20.060000 37.460000 20.260000 37.660000 ;
        RECT 20.060000 37.900000 20.260000 38.100000 ;
        RECT 20.060000 49.715000 20.260000 49.915000 ;
        RECT 20.060000 50.135000 20.260000 50.335000 ;
        RECT 20.060000 50.555000 20.260000 50.755000 ;
        RECT 20.465000 34.820000 20.665000 35.020000 ;
        RECT 20.465000 35.260000 20.665000 35.460000 ;
        RECT 20.465000 35.700000 20.665000 35.900000 ;
        RECT 20.465000 36.140000 20.665000 36.340000 ;
        RECT 20.465000 36.580000 20.665000 36.780000 ;
        RECT 20.465000 37.020000 20.665000 37.220000 ;
        RECT 20.465000 37.460000 20.665000 37.660000 ;
        RECT 20.465000 37.900000 20.665000 38.100000 ;
        RECT 20.465000 49.715000 20.665000 49.915000 ;
        RECT 20.465000 50.135000 20.665000 50.335000 ;
        RECT 20.465000 50.555000 20.665000 50.755000 ;
        RECT 20.870000 34.820000 21.070000 35.020000 ;
        RECT 20.870000 35.260000 21.070000 35.460000 ;
        RECT 20.870000 35.700000 21.070000 35.900000 ;
        RECT 20.870000 36.140000 21.070000 36.340000 ;
        RECT 20.870000 36.580000 21.070000 36.780000 ;
        RECT 20.870000 37.020000 21.070000 37.220000 ;
        RECT 20.870000 37.460000 21.070000 37.660000 ;
        RECT 20.870000 37.900000 21.070000 38.100000 ;
        RECT 20.870000 49.715000 21.070000 49.915000 ;
        RECT 20.870000 50.135000 21.070000 50.335000 ;
        RECT 20.870000 50.555000 21.070000 50.755000 ;
        RECT 21.275000 34.820000 21.475000 35.020000 ;
        RECT 21.275000 35.260000 21.475000 35.460000 ;
        RECT 21.275000 35.700000 21.475000 35.900000 ;
        RECT 21.275000 36.140000 21.475000 36.340000 ;
        RECT 21.275000 36.580000 21.475000 36.780000 ;
        RECT 21.275000 37.020000 21.475000 37.220000 ;
        RECT 21.275000 37.460000 21.475000 37.660000 ;
        RECT 21.275000 37.900000 21.475000 38.100000 ;
        RECT 21.275000 49.715000 21.475000 49.915000 ;
        RECT 21.275000 50.135000 21.475000 50.335000 ;
        RECT 21.275000 50.555000 21.475000 50.755000 ;
        RECT 21.680000 34.820000 21.880000 35.020000 ;
        RECT 21.680000 35.260000 21.880000 35.460000 ;
        RECT 21.680000 35.700000 21.880000 35.900000 ;
        RECT 21.680000 36.140000 21.880000 36.340000 ;
        RECT 21.680000 36.580000 21.880000 36.780000 ;
        RECT 21.680000 37.020000 21.880000 37.220000 ;
        RECT 21.680000 37.460000 21.880000 37.660000 ;
        RECT 21.680000 37.900000 21.880000 38.100000 ;
        RECT 21.680000 49.715000 21.880000 49.915000 ;
        RECT 21.680000 50.135000 21.880000 50.335000 ;
        RECT 21.680000 50.555000 21.880000 50.755000 ;
        RECT 22.085000 34.820000 22.285000 35.020000 ;
        RECT 22.085000 35.260000 22.285000 35.460000 ;
        RECT 22.085000 35.700000 22.285000 35.900000 ;
        RECT 22.085000 36.140000 22.285000 36.340000 ;
        RECT 22.085000 36.580000 22.285000 36.780000 ;
        RECT 22.085000 37.020000 22.285000 37.220000 ;
        RECT 22.085000 37.460000 22.285000 37.660000 ;
        RECT 22.085000 37.900000 22.285000 38.100000 ;
        RECT 22.085000 49.715000 22.285000 49.915000 ;
        RECT 22.085000 50.135000 22.285000 50.335000 ;
        RECT 22.085000 50.555000 22.285000 50.755000 ;
        RECT 22.490000 34.820000 22.690000 35.020000 ;
        RECT 22.490000 35.260000 22.690000 35.460000 ;
        RECT 22.490000 35.700000 22.690000 35.900000 ;
        RECT 22.490000 36.140000 22.690000 36.340000 ;
        RECT 22.490000 36.580000 22.690000 36.780000 ;
        RECT 22.490000 37.020000 22.690000 37.220000 ;
        RECT 22.490000 37.460000 22.690000 37.660000 ;
        RECT 22.490000 37.900000 22.690000 38.100000 ;
        RECT 22.490000 49.715000 22.690000 49.915000 ;
        RECT 22.490000 50.135000 22.690000 50.335000 ;
        RECT 22.490000 50.555000 22.690000 50.755000 ;
        RECT 22.895000 34.820000 23.095000 35.020000 ;
        RECT 22.895000 35.260000 23.095000 35.460000 ;
        RECT 22.895000 35.700000 23.095000 35.900000 ;
        RECT 22.895000 36.140000 23.095000 36.340000 ;
        RECT 22.895000 36.580000 23.095000 36.780000 ;
        RECT 22.895000 37.020000 23.095000 37.220000 ;
        RECT 22.895000 37.460000 23.095000 37.660000 ;
        RECT 22.895000 37.900000 23.095000 38.100000 ;
        RECT 22.895000 49.715000 23.095000 49.915000 ;
        RECT 22.895000 50.135000 23.095000 50.335000 ;
        RECT 22.895000 50.555000 23.095000 50.755000 ;
        RECT 23.300000 34.820000 23.500000 35.020000 ;
        RECT 23.300000 35.260000 23.500000 35.460000 ;
        RECT 23.300000 35.700000 23.500000 35.900000 ;
        RECT 23.300000 36.140000 23.500000 36.340000 ;
        RECT 23.300000 36.580000 23.500000 36.780000 ;
        RECT 23.300000 37.020000 23.500000 37.220000 ;
        RECT 23.300000 37.460000 23.500000 37.660000 ;
        RECT 23.300000 37.900000 23.500000 38.100000 ;
        RECT 23.300000 49.715000 23.500000 49.915000 ;
        RECT 23.300000 50.135000 23.500000 50.335000 ;
        RECT 23.300000 50.555000 23.500000 50.755000 ;
        RECT 23.705000 34.820000 23.905000 35.020000 ;
        RECT 23.705000 35.260000 23.905000 35.460000 ;
        RECT 23.705000 35.700000 23.905000 35.900000 ;
        RECT 23.705000 36.140000 23.905000 36.340000 ;
        RECT 23.705000 36.580000 23.905000 36.780000 ;
        RECT 23.705000 37.020000 23.905000 37.220000 ;
        RECT 23.705000 37.460000 23.905000 37.660000 ;
        RECT 23.705000 37.900000 23.905000 38.100000 ;
        RECT 23.705000 49.715000 23.905000 49.915000 ;
        RECT 23.705000 50.135000 23.905000 50.335000 ;
        RECT 23.705000 50.555000 23.905000 50.755000 ;
        RECT 24.110000 34.820000 24.310000 35.020000 ;
        RECT 24.110000 35.260000 24.310000 35.460000 ;
        RECT 24.110000 35.700000 24.310000 35.900000 ;
        RECT 24.110000 36.140000 24.310000 36.340000 ;
        RECT 24.110000 36.580000 24.310000 36.780000 ;
        RECT 24.110000 37.020000 24.310000 37.220000 ;
        RECT 24.110000 37.460000 24.310000 37.660000 ;
        RECT 24.110000 37.900000 24.310000 38.100000 ;
        RECT 24.110000 49.715000 24.310000 49.915000 ;
        RECT 24.110000 50.135000 24.310000 50.335000 ;
        RECT 24.110000 50.555000 24.310000 50.755000 ;
        RECT 50.845000 34.820000 51.045000 35.020000 ;
        RECT 50.845000 35.260000 51.045000 35.460000 ;
        RECT 50.845000 35.700000 51.045000 35.900000 ;
        RECT 50.845000 36.140000 51.045000 36.340000 ;
        RECT 50.845000 36.580000 51.045000 36.780000 ;
        RECT 50.845000 37.020000 51.045000 37.220000 ;
        RECT 50.845000 37.460000 51.045000 37.660000 ;
        RECT 50.845000 37.900000 51.045000 38.100000 ;
        RECT 50.845000 49.715000 51.045000 49.915000 ;
        RECT 50.845000 50.135000 51.045000 50.335000 ;
        RECT 50.845000 50.555000 51.045000 50.755000 ;
        RECT 51.255000 34.820000 51.455000 35.020000 ;
        RECT 51.255000 35.260000 51.455000 35.460000 ;
        RECT 51.255000 35.700000 51.455000 35.900000 ;
        RECT 51.255000 36.140000 51.455000 36.340000 ;
        RECT 51.255000 36.580000 51.455000 36.780000 ;
        RECT 51.255000 37.020000 51.455000 37.220000 ;
        RECT 51.255000 37.460000 51.455000 37.660000 ;
        RECT 51.255000 37.900000 51.455000 38.100000 ;
        RECT 51.255000 49.715000 51.455000 49.915000 ;
        RECT 51.255000 50.135000 51.455000 50.335000 ;
        RECT 51.255000 50.555000 51.455000 50.755000 ;
        RECT 51.665000 34.820000 51.865000 35.020000 ;
        RECT 51.665000 35.260000 51.865000 35.460000 ;
        RECT 51.665000 35.700000 51.865000 35.900000 ;
        RECT 51.665000 36.140000 51.865000 36.340000 ;
        RECT 51.665000 36.580000 51.865000 36.780000 ;
        RECT 51.665000 37.020000 51.865000 37.220000 ;
        RECT 51.665000 37.460000 51.865000 37.660000 ;
        RECT 51.665000 37.900000 51.865000 38.100000 ;
        RECT 51.665000 49.715000 51.865000 49.915000 ;
        RECT 51.665000 50.135000 51.865000 50.335000 ;
        RECT 51.665000 50.555000 51.865000 50.755000 ;
        RECT 52.075000 34.820000 52.275000 35.020000 ;
        RECT 52.075000 35.260000 52.275000 35.460000 ;
        RECT 52.075000 35.700000 52.275000 35.900000 ;
        RECT 52.075000 36.140000 52.275000 36.340000 ;
        RECT 52.075000 36.580000 52.275000 36.780000 ;
        RECT 52.075000 37.020000 52.275000 37.220000 ;
        RECT 52.075000 37.460000 52.275000 37.660000 ;
        RECT 52.075000 37.900000 52.275000 38.100000 ;
        RECT 52.075000 49.715000 52.275000 49.915000 ;
        RECT 52.075000 50.135000 52.275000 50.335000 ;
        RECT 52.075000 50.555000 52.275000 50.755000 ;
        RECT 52.485000 34.820000 52.685000 35.020000 ;
        RECT 52.485000 35.260000 52.685000 35.460000 ;
        RECT 52.485000 35.700000 52.685000 35.900000 ;
        RECT 52.485000 36.140000 52.685000 36.340000 ;
        RECT 52.485000 36.580000 52.685000 36.780000 ;
        RECT 52.485000 37.020000 52.685000 37.220000 ;
        RECT 52.485000 37.460000 52.685000 37.660000 ;
        RECT 52.485000 37.900000 52.685000 38.100000 ;
        RECT 52.485000 49.715000 52.685000 49.915000 ;
        RECT 52.485000 50.135000 52.685000 50.335000 ;
        RECT 52.485000 50.555000 52.685000 50.755000 ;
        RECT 52.895000 34.820000 53.095000 35.020000 ;
        RECT 52.895000 35.260000 53.095000 35.460000 ;
        RECT 52.895000 35.700000 53.095000 35.900000 ;
        RECT 52.895000 36.140000 53.095000 36.340000 ;
        RECT 52.895000 36.580000 53.095000 36.780000 ;
        RECT 52.895000 37.020000 53.095000 37.220000 ;
        RECT 52.895000 37.460000 53.095000 37.660000 ;
        RECT 52.895000 37.900000 53.095000 38.100000 ;
        RECT 52.895000 49.715000 53.095000 49.915000 ;
        RECT 52.895000 50.135000 53.095000 50.335000 ;
        RECT 52.895000 50.555000 53.095000 50.755000 ;
        RECT 53.305000 34.820000 53.505000 35.020000 ;
        RECT 53.305000 35.260000 53.505000 35.460000 ;
        RECT 53.305000 35.700000 53.505000 35.900000 ;
        RECT 53.305000 36.140000 53.505000 36.340000 ;
        RECT 53.305000 36.580000 53.505000 36.780000 ;
        RECT 53.305000 37.020000 53.505000 37.220000 ;
        RECT 53.305000 37.460000 53.505000 37.660000 ;
        RECT 53.305000 37.900000 53.505000 38.100000 ;
        RECT 53.305000 49.715000 53.505000 49.915000 ;
        RECT 53.305000 50.135000 53.505000 50.335000 ;
        RECT 53.305000 50.555000 53.505000 50.755000 ;
        RECT 53.710000 34.820000 53.910000 35.020000 ;
        RECT 53.710000 35.260000 53.910000 35.460000 ;
        RECT 53.710000 35.700000 53.910000 35.900000 ;
        RECT 53.710000 36.140000 53.910000 36.340000 ;
        RECT 53.710000 36.580000 53.910000 36.780000 ;
        RECT 53.710000 37.020000 53.910000 37.220000 ;
        RECT 53.710000 37.460000 53.910000 37.660000 ;
        RECT 53.710000 37.900000 53.910000 38.100000 ;
        RECT 53.710000 49.715000 53.910000 49.915000 ;
        RECT 53.710000 50.135000 53.910000 50.335000 ;
        RECT 53.710000 50.555000 53.910000 50.755000 ;
        RECT 54.115000 34.820000 54.315000 35.020000 ;
        RECT 54.115000 35.260000 54.315000 35.460000 ;
        RECT 54.115000 35.700000 54.315000 35.900000 ;
        RECT 54.115000 36.140000 54.315000 36.340000 ;
        RECT 54.115000 36.580000 54.315000 36.780000 ;
        RECT 54.115000 37.020000 54.315000 37.220000 ;
        RECT 54.115000 37.460000 54.315000 37.660000 ;
        RECT 54.115000 37.900000 54.315000 38.100000 ;
        RECT 54.115000 49.715000 54.315000 49.915000 ;
        RECT 54.115000 50.135000 54.315000 50.335000 ;
        RECT 54.115000 50.555000 54.315000 50.755000 ;
        RECT 54.520000 34.820000 54.720000 35.020000 ;
        RECT 54.520000 35.260000 54.720000 35.460000 ;
        RECT 54.520000 35.700000 54.720000 35.900000 ;
        RECT 54.520000 36.140000 54.720000 36.340000 ;
        RECT 54.520000 36.580000 54.720000 36.780000 ;
        RECT 54.520000 37.020000 54.720000 37.220000 ;
        RECT 54.520000 37.460000 54.720000 37.660000 ;
        RECT 54.520000 37.900000 54.720000 38.100000 ;
        RECT 54.520000 49.715000 54.720000 49.915000 ;
        RECT 54.520000 50.135000 54.720000 50.335000 ;
        RECT 54.520000 50.555000 54.720000 50.755000 ;
        RECT 54.925000 34.820000 55.125000 35.020000 ;
        RECT 54.925000 35.260000 55.125000 35.460000 ;
        RECT 54.925000 35.700000 55.125000 35.900000 ;
        RECT 54.925000 36.140000 55.125000 36.340000 ;
        RECT 54.925000 36.580000 55.125000 36.780000 ;
        RECT 54.925000 37.020000 55.125000 37.220000 ;
        RECT 54.925000 37.460000 55.125000 37.660000 ;
        RECT 54.925000 37.900000 55.125000 38.100000 ;
        RECT 54.925000 49.715000 55.125000 49.915000 ;
        RECT 54.925000 50.135000 55.125000 50.335000 ;
        RECT 54.925000 50.555000 55.125000 50.755000 ;
        RECT 55.330000 34.820000 55.530000 35.020000 ;
        RECT 55.330000 35.260000 55.530000 35.460000 ;
        RECT 55.330000 35.700000 55.530000 35.900000 ;
        RECT 55.330000 36.140000 55.530000 36.340000 ;
        RECT 55.330000 36.580000 55.530000 36.780000 ;
        RECT 55.330000 37.020000 55.530000 37.220000 ;
        RECT 55.330000 37.460000 55.530000 37.660000 ;
        RECT 55.330000 37.900000 55.530000 38.100000 ;
        RECT 55.330000 49.715000 55.530000 49.915000 ;
        RECT 55.330000 50.135000 55.530000 50.335000 ;
        RECT 55.330000 50.555000 55.530000 50.755000 ;
        RECT 55.735000 34.820000 55.935000 35.020000 ;
        RECT 55.735000 35.260000 55.935000 35.460000 ;
        RECT 55.735000 35.700000 55.935000 35.900000 ;
        RECT 55.735000 36.140000 55.935000 36.340000 ;
        RECT 55.735000 36.580000 55.935000 36.780000 ;
        RECT 55.735000 37.020000 55.935000 37.220000 ;
        RECT 55.735000 37.460000 55.935000 37.660000 ;
        RECT 55.735000 37.900000 55.935000 38.100000 ;
        RECT 55.735000 49.715000 55.935000 49.915000 ;
        RECT 55.735000 50.135000 55.935000 50.335000 ;
        RECT 55.735000 50.555000 55.935000 50.755000 ;
        RECT 56.140000 34.820000 56.340000 35.020000 ;
        RECT 56.140000 35.260000 56.340000 35.460000 ;
        RECT 56.140000 35.700000 56.340000 35.900000 ;
        RECT 56.140000 36.140000 56.340000 36.340000 ;
        RECT 56.140000 36.580000 56.340000 36.780000 ;
        RECT 56.140000 37.020000 56.340000 37.220000 ;
        RECT 56.140000 37.460000 56.340000 37.660000 ;
        RECT 56.140000 37.900000 56.340000 38.100000 ;
        RECT 56.140000 49.715000 56.340000 49.915000 ;
        RECT 56.140000 50.135000 56.340000 50.335000 ;
        RECT 56.140000 50.555000 56.340000 50.755000 ;
        RECT 56.545000 34.820000 56.745000 35.020000 ;
        RECT 56.545000 35.260000 56.745000 35.460000 ;
        RECT 56.545000 35.700000 56.745000 35.900000 ;
        RECT 56.545000 36.140000 56.745000 36.340000 ;
        RECT 56.545000 36.580000 56.745000 36.780000 ;
        RECT 56.545000 37.020000 56.745000 37.220000 ;
        RECT 56.545000 37.460000 56.745000 37.660000 ;
        RECT 56.545000 37.900000 56.745000 38.100000 ;
        RECT 56.545000 49.715000 56.745000 49.915000 ;
        RECT 56.545000 50.135000 56.745000 50.335000 ;
        RECT 56.545000 50.555000 56.745000 50.755000 ;
        RECT 56.950000 34.820000 57.150000 35.020000 ;
        RECT 56.950000 35.260000 57.150000 35.460000 ;
        RECT 56.950000 35.700000 57.150000 35.900000 ;
        RECT 56.950000 36.140000 57.150000 36.340000 ;
        RECT 56.950000 36.580000 57.150000 36.780000 ;
        RECT 56.950000 37.020000 57.150000 37.220000 ;
        RECT 56.950000 37.460000 57.150000 37.660000 ;
        RECT 56.950000 37.900000 57.150000 38.100000 ;
        RECT 56.950000 49.715000 57.150000 49.915000 ;
        RECT 56.950000 50.135000 57.150000 50.335000 ;
        RECT 56.950000 50.555000 57.150000 50.755000 ;
        RECT 57.355000 34.820000 57.555000 35.020000 ;
        RECT 57.355000 35.260000 57.555000 35.460000 ;
        RECT 57.355000 35.700000 57.555000 35.900000 ;
        RECT 57.355000 36.140000 57.555000 36.340000 ;
        RECT 57.355000 36.580000 57.555000 36.780000 ;
        RECT 57.355000 37.020000 57.555000 37.220000 ;
        RECT 57.355000 37.460000 57.555000 37.660000 ;
        RECT 57.355000 37.900000 57.555000 38.100000 ;
        RECT 57.355000 49.715000 57.555000 49.915000 ;
        RECT 57.355000 50.135000 57.555000 50.335000 ;
        RECT 57.355000 50.555000 57.555000 50.755000 ;
        RECT 57.760000 34.820000 57.960000 35.020000 ;
        RECT 57.760000 35.260000 57.960000 35.460000 ;
        RECT 57.760000 35.700000 57.960000 35.900000 ;
        RECT 57.760000 36.140000 57.960000 36.340000 ;
        RECT 57.760000 36.580000 57.960000 36.780000 ;
        RECT 57.760000 37.020000 57.960000 37.220000 ;
        RECT 57.760000 37.460000 57.960000 37.660000 ;
        RECT 57.760000 37.900000 57.960000 38.100000 ;
        RECT 57.760000 49.715000 57.960000 49.915000 ;
        RECT 57.760000 50.135000 57.960000 50.335000 ;
        RECT 57.760000 50.555000 57.960000 50.755000 ;
        RECT 58.165000 34.820000 58.365000 35.020000 ;
        RECT 58.165000 35.260000 58.365000 35.460000 ;
        RECT 58.165000 35.700000 58.365000 35.900000 ;
        RECT 58.165000 36.140000 58.365000 36.340000 ;
        RECT 58.165000 36.580000 58.365000 36.780000 ;
        RECT 58.165000 37.020000 58.365000 37.220000 ;
        RECT 58.165000 37.460000 58.365000 37.660000 ;
        RECT 58.165000 37.900000 58.365000 38.100000 ;
        RECT 58.165000 49.715000 58.365000 49.915000 ;
        RECT 58.165000 50.135000 58.365000 50.335000 ;
        RECT 58.165000 50.555000 58.365000 50.755000 ;
        RECT 58.570000 34.820000 58.770000 35.020000 ;
        RECT 58.570000 35.260000 58.770000 35.460000 ;
        RECT 58.570000 35.700000 58.770000 35.900000 ;
        RECT 58.570000 36.140000 58.770000 36.340000 ;
        RECT 58.570000 36.580000 58.770000 36.780000 ;
        RECT 58.570000 37.020000 58.770000 37.220000 ;
        RECT 58.570000 37.460000 58.770000 37.660000 ;
        RECT 58.570000 37.900000 58.770000 38.100000 ;
        RECT 58.570000 49.715000 58.770000 49.915000 ;
        RECT 58.570000 50.135000 58.770000 50.335000 ;
        RECT 58.570000 50.555000 58.770000 50.755000 ;
        RECT 58.975000 34.820000 59.175000 35.020000 ;
        RECT 58.975000 35.260000 59.175000 35.460000 ;
        RECT 58.975000 35.700000 59.175000 35.900000 ;
        RECT 58.975000 36.140000 59.175000 36.340000 ;
        RECT 58.975000 36.580000 59.175000 36.780000 ;
        RECT 58.975000 37.020000 59.175000 37.220000 ;
        RECT 58.975000 37.460000 59.175000 37.660000 ;
        RECT 58.975000 37.900000 59.175000 38.100000 ;
        RECT 58.975000 49.715000 59.175000 49.915000 ;
        RECT 58.975000 50.135000 59.175000 50.335000 ;
        RECT 58.975000 50.555000 59.175000 50.755000 ;
        RECT 59.380000 34.820000 59.580000 35.020000 ;
        RECT 59.380000 35.260000 59.580000 35.460000 ;
        RECT 59.380000 35.700000 59.580000 35.900000 ;
        RECT 59.380000 36.140000 59.580000 36.340000 ;
        RECT 59.380000 36.580000 59.580000 36.780000 ;
        RECT 59.380000 37.020000 59.580000 37.220000 ;
        RECT 59.380000 37.460000 59.580000 37.660000 ;
        RECT 59.380000 37.900000 59.580000 38.100000 ;
        RECT 59.380000 49.715000 59.580000 49.915000 ;
        RECT 59.380000 50.135000 59.580000 50.335000 ;
        RECT 59.380000 50.555000 59.580000 50.755000 ;
        RECT 59.785000 34.820000 59.985000 35.020000 ;
        RECT 59.785000 35.260000 59.985000 35.460000 ;
        RECT 59.785000 35.700000 59.985000 35.900000 ;
        RECT 59.785000 36.140000 59.985000 36.340000 ;
        RECT 59.785000 36.580000 59.985000 36.780000 ;
        RECT 59.785000 37.020000 59.985000 37.220000 ;
        RECT 59.785000 37.460000 59.985000 37.660000 ;
        RECT 59.785000 37.900000 59.985000 38.100000 ;
        RECT 59.785000 49.715000 59.985000 49.915000 ;
        RECT 59.785000 50.135000 59.985000 50.335000 ;
        RECT 59.785000 50.555000 59.985000 50.755000 ;
        RECT 60.190000 34.820000 60.390000 35.020000 ;
        RECT 60.190000 35.260000 60.390000 35.460000 ;
        RECT 60.190000 35.700000 60.390000 35.900000 ;
        RECT 60.190000 36.140000 60.390000 36.340000 ;
        RECT 60.190000 36.580000 60.390000 36.780000 ;
        RECT 60.190000 37.020000 60.390000 37.220000 ;
        RECT 60.190000 37.460000 60.390000 37.660000 ;
        RECT 60.190000 37.900000 60.390000 38.100000 ;
        RECT 60.190000 49.715000 60.390000 49.915000 ;
        RECT 60.190000 50.135000 60.390000 50.335000 ;
        RECT 60.190000 50.555000 60.390000 50.755000 ;
        RECT 60.595000 34.820000 60.795000 35.020000 ;
        RECT 60.595000 35.260000 60.795000 35.460000 ;
        RECT 60.595000 35.700000 60.795000 35.900000 ;
        RECT 60.595000 36.140000 60.795000 36.340000 ;
        RECT 60.595000 36.580000 60.795000 36.780000 ;
        RECT 60.595000 37.020000 60.795000 37.220000 ;
        RECT 60.595000 37.460000 60.795000 37.660000 ;
        RECT 60.595000 37.900000 60.795000 38.100000 ;
        RECT 60.595000 49.715000 60.795000 49.915000 ;
        RECT 60.595000 50.135000 60.795000 50.335000 ;
        RECT 60.595000 50.555000 60.795000 50.755000 ;
        RECT 61.000000 34.820000 61.200000 35.020000 ;
        RECT 61.000000 35.260000 61.200000 35.460000 ;
        RECT 61.000000 35.700000 61.200000 35.900000 ;
        RECT 61.000000 36.140000 61.200000 36.340000 ;
        RECT 61.000000 36.580000 61.200000 36.780000 ;
        RECT 61.000000 37.020000 61.200000 37.220000 ;
        RECT 61.000000 37.460000 61.200000 37.660000 ;
        RECT 61.000000 37.900000 61.200000 38.100000 ;
        RECT 61.000000 49.715000 61.200000 49.915000 ;
        RECT 61.000000 50.135000 61.200000 50.335000 ;
        RECT 61.000000 50.555000 61.200000 50.755000 ;
        RECT 61.405000 34.820000 61.605000 35.020000 ;
        RECT 61.405000 35.260000 61.605000 35.460000 ;
        RECT 61.405000 35.700000 61.605000 35.900000 ;
        RECT 61.405000 36.140000 61.605000 36.340000 ;
        RECT 61.405000 36.580000 61.605000 36.780000 ;
        RECT 61.405000 37.020000 61.605000 37.220000 ;
        RECT 61.405000 37.460000 61.605000 37.660000 ;
        RECT 61.405000 37.900000 61.605000 38.100000 ;
        RECT 61.405000 49.715000 61.605000 49.915000 ;
        RECT 61.405000 50.135000 61.605000 50.335000 ;
        RECT 61.405000 50.555000 61.605000 50.755000 ;
        RECT 61.810000 34.820000 62.010000 35.020000 ;
        RECT 61.810000 35.260000 62.010000 35.460000 ;
        RECT 61.810000 35.700000 62.010000 35.900000 ;
        RECT 61.810000 36.140000 62.010000 36.340000 ;
        RECT 61.810000 36.580000 62.010000 36.780000 ;
        RECT 61.810000 37.020000 62.010000 37.220000 ;
        RECT 61.810000 37.460000 62.010000 37.660000 ;
        RECT 61.810000 37.900000 62.010000 38.100000 ;
        RECT 61.810000 49.715000 62.010000 49.915000 ;
        RECT 61.810000 50.135000 62.010000 50.335000 ;
        RECT 61.810000 50.555000 62.010000 50.755000 ;
        RECT 62.215000 34.820000 62.415000 35.020000 ;
        RECT 62.215000 35.260000 62.415000 35.460000 ;
        RECT 62.215000 35.700000 62.415000 35.900000 ;
        RECT 62.215000 36.140000 62.415000 36.340000 ;
        RECT 62.215000 36.580000 62.415000 36.780000 ;
        RECT 62.215000 37.020000 62.415000 37.220000 ;
        RECT 62.215000 37.460000 62.415000 37.660000 ;
        RECT 62.215000 37.900000 62.415000 38.100000 ;
        RECT 62.215000 49.715000 62.415000 49.915000 ;
        RECT 62.215000 50.135000 62.415000 50.335000 ;
        RECT 62.215000 50.555000 62.415000 50.755000 ;
        RECT 62.620000 34.820000 62.820000 35.020000 ;
        RECT 62.620000 35.260000 62.820000 35.460000 ;
        RECT 62.620000 35.700000 62.820000 35.900000 ;
        RECT 62.620000 36.140000 62.820000 36.340000 ;
        RECT 62.620000 36.580000 62.820000 36.780000 ;
        RECT 62.620000 37.020000 62.820000 37.220000 ;
        RECT 62.620000 37.460000 62.820000 37.660000 ;
        RECT 62.620000 37.900000 62.820000 38.100000 ;
        RECT 62.620000 49.715000 62.820000 49.915000 ;
        RECT 62.620000 50.135000 62.820000 50.335000 ;
        RECT 62.620000 50.555000 62.820000 50.755000 ;
        RECT 63.025000 34.820000 63.225000 35.020000 ;
        RECT 63.025000 35.260000 63.225000 35.460000 ;
        RECT 63.025000 35.700000 63.225000 35.900000 ;
        RECT 63.025000 36.140000 63.225000 36.340000 ;
        RECT 63.025000 36.580000 63.225000 36.780000 ;
        RECT 63.025000 37.020000 63.225000 37.220000 ;
        RECT 63.025000 37.460000 63.225000 37.660000 ;
        RECT 63.025000 37.900000 63.225000 38.100000 ;
        RECT 63.025000 49.715000 63.225000 49.915000 ;
        RECT 63.025000 50.135000 63.225000 50.335000 ;
        RECT 63.025000 50.555000 63.225000 50.755000 ;
        RECT 63.430000 34.820000 63.630000 35.020000 ;
        RECT 63.430000 35.260000 63.630000 35.460000 ;
        RECT 63.430000 35.700000 63.630000 35.900000 ;
        RECT 63.430000 36.140000 63.630000 36.340000 ;
        RECT 63.430000 36.580000 63.630000 36.780000 ;
        RECT 63.430000 37.020000 63.630000 37.220000 ;
        RECT 63.430000 37.460000 63.630000 37.660000 ;
        RECT 63.430000 37.900000 63.630000 38.100000 ;
        RECT 63.430000 49.715000 63.630000 49.915000 ;
        RECT 63.430000 50.135000 63.630000 50.335000 ;
        RECT 63.430000 50.555000 63.630000 50.755000 ;
        RECT 63.835000 34.820000 64.035000 35.020000 ;
        RECT 63.835000 35.260000 64.035000 35.460000 ;
        RECT 63.835000 35.700000 64.035000 35.900000 ;
        RECT 63.835000 36.140000 64.035000 36.340000 ;
        RECT 63.835000 36.580000 64.035000 36.780000 ;
        RECT 63.835000 37.020000 64.035000 37.220000 ;
        RECT 63.835000 37.460000 64.035000 37.660000 ;
        RECT 63.835000 37.900000 64.035000 38.100000 ;
        RECT 63.835000 49.715000 64.035000 49.915000 ;
        RECT 63.835000 50.135000 64.035000 50.335000 ;
        RECT 63.835000 50.555000 64.035000 50.755000 ;
        RECT 64.240000 34.820000 64.440000 35.020000 ;
        RECT 64.240000 35.260000 64.440000 35.460000 ;
        RECT 64.240000 35.700000 64.440000 35.900000 ;
        RECT 64.240000 36.140000 64.440000 36.340000 ;
        RECT 64.240000 36.580000 64.440000 36.780000 ;
        RECT 64.240000 37.020000 64.440000 37.220000 ;
        RECT 64.240000 37.460000 64.440000 37.660000 ;
        RECT 64.240000 37.900000 64.440000 38.100000 ;
        RECT 64.240000 49.715000 64.440000 49.915000 ;
        RECT 64.240000 50.135000 64.440000 50.335000 ;
        RECT 64.240000 50.555000 64.440000 50.755000 ;
        RECT 64.645000 34.820000 64.845000 35.020000 ;
        RECT 64.645000 35.260000 64.845000 35.460000 ;
        RECT 64.645000 35.700000 64.845000 35.900000 ;
        RECT 64.645000 36.140000 64.845000 36.340000 ;
        RECT 64.645000 36.580000 64.845000 36.780000 ;
        RECT 64.645000 37.020000 64.845000 37.220000 ;
        RECT 64.645000 37.460000 64.845000 37.660000 ;
        RECT 64.645000 37.900000 64.845000 38.100000 ;
        RECT 64.645000 49.715000 64.845000 49.915000 ;
        RECT 64.645000 50.135000 64.845000 50.335000 ;
        RECT 64.645000 50.555000 64.845000 50.755000 ;
        RECT 65.050000 34.820000 65.250000 35.020000 ;
        RECT 65.050000 35.260000 65.250000 35.460000 ;
        RECT 65.050000 35.700000 65.250000 35.900000 ;
        RECT 65.050000 36.140000 65.250000 36.340000 ;
        RECT 65.050000 36.580000 65.250000 36.780000 ;
        RECT 65.050000 37.020000 65.250000 37.220000 ;
        RECT 65.050000 37.460000 65.250000 37.660000 ;
        RECT 65.050000 37.900000 65.250000 38.100000 ;
        RECT 65.050000 49.715000 65.250000 49.915000 ;
        RECT 65.050000 50.135000 65.250000 50.335000 ;
        RECT 65.050000 50.555000 65.250000 50.755000 ;
        RECT 65.455000 34.820000 65.655000 35.020000 ;
        RECT 65.455000 35.260000 65.655000 35.460000 ;
        RECT 65.455000 35.700000 65.655000 35.900000 ;
        RECT 65.455000 36.140000 65.655000 36.340000 ;
        RECT 65.455000 36.580000 65.655000 36.780000 ;
        RECT 65.455000 37.020000 65.655000 37.220000 ;
        RECT 65.455000 37.460000 65.655000 37.660000 ;
        RECT 65.455000 37.900000 65.655000 38.100000 ;
        RECT 65.455000 49.715000 65.655000 49.915000 ;
        RECT 65.455000 50.135000 65.655000 50.335000 ;
        RECT 65.455000 50.555000 65.655000 50.755000 ;
        RECT 65.860000 34.820000 66.060000 35.020000 ;
        RECT 65.860000 35.260000 66.060000 35.460000 ;
        RECT 65.860000 35.700000 66.060000 35.900000 ;
        RECT 65.860000 36.140000 66.060000 36.340000 ;
        RECT 65.860000 36.580000 66.060000 36.780000 ;
        RECT 65.860000 37.020000 66.060000 37.220000 ;
        RECT 65.860000 37.460000 66.060000 37.660000 ;
        RECT 65.860000 37.900000 66.060000 38.100000 ;
        RECT 65.860000 49.715000 66.060000 49.915000 ;
        RECT 65.860000 50.135000 66.060000 50.335000 ;
        RECT 65.860000 50.555000 66.060000 50.755000 ;
        RECT 66.265000 34.820000 66.465000 35.020000 ;
        RECT 66.265000 35.260000 66.465000 35.460000 ;
        RECT 66.265000 35.700000 66.465000 35.900000 ;
        RECT 66.265000 36.140000 66.465000 36.340000 ;
        RECT 66.265000 36.580000 66.465000 36.780000 ;
        RECT 66.265000 37.020000 66.465000 37.220000 ;
        RECT 66.265000 37.460000 66.465000 37.660000 ;
        RECT 66.265000 37.900000 66.465000 38.100000 ;
        RECT 66.265000 49.715000 66.465000 49.915000 ;
        RECT 66.265000 50.135000 66.465000 50.335000 ;
        RECT 66.265000 50.555000 66.465000 50.755000 ;
        RECT 66.670000 34.820000 66.870000 35.020000 ;
        RECT 66.670000 35.260000 66.870000 35.460000 ;
        RECT 66.670000 35.700000 66.870000 35.900000 ;
        RECT 66.670000 36.140000 66.870000 36.340000 ;
        RECT 66.670000 36.580000 66.870000 36.780000 ;
        RECT 66.670000 37.020000 66.870000 37.220000 ;
        RECT 66.670000 37.460000 66.870000 37.660000 ;
        RECT 66.670000 37.900000 66.870000 38.100000 ;
        RECT 66.670000 49.715000 66.870000 49.915000 ;
        RECT 66.670000 50.135000 66.870000 50.335000 ;
        RECT 66.670000 50.555000 66.870000 50.755000 ;
        RECT 67.075000 34.820000 67.275000 35.020000 ;
        RECT 67.075000 35.260000 67.275000 35.460000 ;
        RECT 67.075000 35.700000 67.275000 35.900000 ;
        RECT 67.075000 36.140000 67.275000 36.340000 ;
        RECT 67.075000 36.580000 67.275000 36.780000 ;
        RECT 67.075000 37.020000 67.275000 37.220000 ;
        RECT 67.075000 37.460000 67.275000 37.660000 ;
        RECT 67.075000 37.900000 67.275000 38.100000 ;
        RECT 67.075000 49.715000 67.275000 49.915000 ;
        RECT 67.075000 50.135000 67.275000 50.335000 ;
        RECT 67.075000 50.555000 67.275000 50.755000 ;
        RECT 67.480000 34.820000 67.680000 35.020000 ;
        RECT 67.480000 35.260000 67.680000 35.460000 ;
        RECT 67.480000 35.700000 67.680000 35.900000 ;
        RECT 67.480000 36.140000 67.680000 36.340000 ;
        RECT 67.480000 36.580000 67.680000 36.780000 ;
        RECT 67.480000 37.020000 67.680000 37.220000 ;
        RECT 67.480000 37.460000 67.680000 37.660000 ;
        RECT 67.480000 37.900000 67.680000 38.100000 ;
        RECT 67.480000 49.715000 67.680000 49.915000 ;
        RECT 67.480000 50.135000 67.680000 50.335000 ;
        RECT 67.480000 50.555000 67.680000 50.755000 ;
        RECT 67.885000 34.820000 68.085000 35.020000 ;
        RECT 67.885000 35.260000 68.085000 35.460000 ;
        RECT 67.885000 35.700000 68.085000 35.900000 ;
        RECT 67.885000 36.140000 68.085000 36.340000 ;
        RECT 67.885000 36.580000 68.085000 36.780000 ;
        RECT 67.885000 37.020000 68.085000 37.220000 ;
        RECT 67.885000 37.460000 68.085000 37.660000 ;
        RECT 67.885000 37.900000 68.085000 38.100000 ;
        RECT 67.885000 49.715000 68.085000 49.915000 ;
        RECT 67.885000 50.135000 68.085000 50.335000 ;
        RECT 67.885000 50.555000 68.085000 50.755000 ;
        RECT 68.290000 34.820000 68.490000 35.020000 ;
        RECT 68.290000 35.260000 68.490000 35.460000 ;
        RECT 68.290000 35.700000 68.490000 35.900000 ;
        RECT 68.290000 36.140000 68.490000 36.340000 ;
        RECT 68.290000 36.580000 68.490000 36.780000 ;
        RECT 68.290000 37.020000 68.490000 37.220000 ;
        RECT 68.290000 37.460000 68.490000 37.660000 ;
        RECT 68.290000 37.900000 68.490000 38.100000 ;
        RECT 68.290000 49.715000 68.490000 49.915000 ;
        RECT 68.290000 50.135000 68.490000 50.335000 ;
        RECT 68.290000 50.555000 68.490000 50.755000 ;
        RECT 68.695000 34.820000 68.895000 35.020000 ;
        RECT 68.695000 35.260000 68.895000 35.460000 ;
        RECT 68.695000 35.700000 68.895000 35.900000 ;
        RECT 68.695000 36.140000 68.895000 36.340000 ;
        RECT 68.695000 36.580000 68.895000 36.780000 ;
        RECT 68.695000 37.020000 68.895000 37.220000 ;
        RECT 68.695000 37.460000 68.895000 37.660000 ;
        RECT 68.695000 37.900000 68.895000 38.100000 ;
        RECT 68.695000 49.715000 68.895000 49.915000 ;
        RECT 68.695000 50.135000 68.895000 50.335000 ;
        RECT 68.695000 50.555000 68.895000 50.755000 ;
        RECT 69.100000 34.820000 69.300000 35.020000 ;
        RECT 69.100000 35.260000 69.300000 35.460000 ;
        RECT 69.100000 35.700000 69.300000 35.900000 ;
        RECT 69.100000 36.140000 69.300000 36.340000 ;
        RECT 69.100000 36.580000 69.300000 36.780000 ;
        RECT 69.100000 37.020000 69.300000 37.220000 ;
        RECT 69.100000 37.460000 69.300000 37.660000 ;
        RECT 69.100000 37.900000 69.300000 38.100000 ;
        RECT 69.100000 49.715000 69.300000 49.915000 ;
        RECT 69.100000 50.135000 69.300000 50.335000 ;
        RECT 69.100000 50.555000 69.300000 50.755000 ;
        RECT 69.505000 34.820000 69.705000 35.020000 ;
        RECT 69.505000 35.260000 69.705000 35.460000 ;
        RECT 69.505000 35.700000 69.705000 35.900000 ;
        RECT 69.505000 36.140000 69.705000 36.340000 ;
        RECT 69.505000 36.580000 69.705000 36.780000 ;
        RECT 69.505000 37.020000 69.705000 37.220000 ;
        RECT 69.505000 37.460000 69.705000 37.660000 ;
        RECT 69.505000 37.900000 69.705000 38.100000 ;
        RECT 69.505000 49.715000 69.705000 49.915000 ;
        RECT 69.505000 50.135000 69.705000 50.335000 ;
        RECT 69.505000 50.555000 69.705000 50.755000 ;
        RECT 69.910000 34.820000 70.110000 35.020000 ;
        RECT 69.910000 35.260000 70.110000 35.460000 ;
        RECT 69.910000 35.700000 70.110000 35.900000 ;
        RECT 69.910000 36.140000 70.110000 36.340000 ;
        RECT 69.910000 36.580000 70.110000 36.780000 ;
        RECT 69.910000 37.020000 70.110000 37.220000 ;
        RECT 69.910000 37.460000 70.110000 37.660000 ;
        RECT 69.910000 37.900000 70.110000 38.100000 ;
        RECT 69.910000 49.715000 70.110000 49.915000 ;
        RECT 69.910000 50.135000 70.110000 50.335000 ;
        RECT 69.910000 50.555000 70.110000 50.755000 ;
        RECT 70.315000 34.820000 70.515000 35.020000 ;
        RECT 70.315000 35.260000 70.515000 35.460000 ;
        RECT 70.315000 35.700000 70.515000 35.900000 ;
        RECT 70.315000 36.140000 70.515000 36.340000 ;
        RECT 70.315000 36.580000 70.515000 36.780000 ;
        RECT 70.315000 37.020000 70.515000 37.220000 ;
        RECT 70.315000 37.460000 70.515000 37.660000 ;
        RECT 70.315000 37.900000 70.515000 38.100000 ;
        RECT 70.315000 49.715000 70.515000 49.915000 ;
        RECT 70.315000 50.135000 70.515000 50.335000 ;
        RECT 70.315000 50.555000 70.515000 50.755000 ;
        RECT 70.720000 34.820000 70.920000 35.020000 ;
        RECT 70.720000 35.260000 70.920000 35.460000 ;
        RECT 70.720000 35.700000 70.920000 35.900000 ;
        RECT 70.720000 36.140000 70.920000 36.340000 ;
        RECT 70.720000 36.580000 70.920000 36.780000 ;
        RECT 70.720000 37.020000 70.920000 37.220000 ;
        RECT 70.720000 37.460000 70.920000 37.660000 ;
        RECT 70.720000 37.900000 70.920000 38.100000 ;
        RECT 70.720000 49.715000 70.920000 49.915000 ;
        RECT 70.720000 50.135000 70.920000 50.335000 ;
        RECT 70.720000 50.555000 70.920000 50.755000 ;
        RECT 71.125000 34.820000 71.325000 35.020000 ;
        RECT 71.125000 35.260000 71.325000 35.460000 ;
        RECT 71.125000 35.700000 71.325000 35.900000 ;
        RECT 71.125000 36.140000 71.325000 36.340000 ;
        RECT 71.125000 36.580000 71.325000 36.780000 ;
        RECT 71.125000 37.020000 71.325000 37.220000 ;
        RECT 71.125000 37.460000 71.325000 37.660000 ;
        RECT 71.125000 37.900000 71.325000 38.100000 ;
        RECT 71.125000 49.715000 71.325000 49.915000 ;
        RECT 71.125000 50.135000 71.325000 50.335000 ;
        RECT 71.125000 50.555000 71.325000 50.755000 ;
        RECT 71.530000 34.820000 71.730000 35.020000 ;
        RECT 71.530000 35.260000 71.730000 35.460000 ;
        RECT 71.530000 35.700000 71.730000 35.900000 ;
        RECT 71.530000 36.140000 71.730000 36.340000 ;
        RECT 71.530000 36.580000 71.730000 36.780000 ;
        RECT 71.530000 37.020000 71.730000 37.220000 ;
        RECT 71.530000 37.460000 71.730000 37.660000 ;
        RECT 71.530000 37.900000 71.730000 38.100000 ;
        RECT 71.530000 49.715000 71.730000 49.915000 ;
        RECT 71.530000 50.135000 71.730000 50.335000 ;
        RECT 71.530000 50.555000 71.730000 50.755000 ;
        RECT 71.935000 34.820000 72.135000 35.020000 ;
        RECT 71.935000 35.260000 72.135000 35.460000 ;
        RECT 71.935000 35.700000 72.135000 35.900000 ;
        RECT 71.935000 36.140000 72.135000 36.340000 ;
        RECT 71.935000 36.580000 72.135000 36.780000 ;
        RECT 71.935000 37.020000 72.135000 37.220000 ;
        RECT 71.935000 37.460000 72.135000 37.660000 ;
        RECT 71.935000 37.900000 72.135000 38.100000 ;
        RECT 71.935000 49.715000 72.135000 49.915000 ;
        RECT 71.935000 50.135000 72.135000 50.335000 ;
        RECT 71.935000 50.555000 72.135000 50.755000 ;
        RECT 72.340000 34.820000 72.540000 35.020000 ;
        RECT 72.340000 35.260000 72.540000 35.460000 ;
        RECT 72.340000 35.700000 72.540000 35.900000 ;
        RECT 72.340000 36.140000 72.540000 36.340000 ;
        RECT 72.340000 36.580000 72.540000 36.780000 ;
        RECT 72.340000 37.020000 72.540000 37.220000 ;
        RECT 72.340000 37.460000 72.540000 37.660000 ;
        RECT 72.340000 37.900000 72.540000 38.100000 ;
        RECT 72.340000 49.715000 72.540000 49.915000 ;
        RECT 72.340000 50.135000 72.540000 50.335000 ;
        RECT 72.340000 50.555000 72.540000 50.755000 ;
        RECT 72.745000 34.820000 72.945000 35.020000 ;
        RECT 72.745000 35.260000 72.945000 35.460000 ;
        RECT 72.745000 35.700000 72.945000 35.900000 ;
        RECT 72.745000 36.140000 72.945000 36.340000 ;
        RECT 72.745000 36.580000 72.945000 36.780000 ;
        RECT 72.745000 37.020000 72.945000 37.220000 ;
        RECT 72.745000 37.460000 72.945000 37.660000 ;
        RECT 72.745000 37.900000 72.945000 38.100000 ;
        RECT 72.745000 49.715000 72.945000 49.915000 ;
        RECT 72.745000 50.135000 72.945000 50.335000 ;
        RECT 72.745000 50.555000 72.945000 50.755000 ;
        RECT 73.150000 34.820000 73.350000 35.020000 ;
        RECT 73.150000 35.260000 73.350000 35.460000 ;
        RECT 73.150000 35.700000 73.350000 35.900000 ;
        RECT 73.150000 36.140000 73.350000 36.340000 ;
        RECT 73.150000 36.580000 73.350000 36.780000 ;
        RECT 73.150000 37.020000 73.350000 37.220000 ;
        RECT 73.150000 37.460000 73.350000 37.660000 ;
        RECT 73.150000 37.900000 73.350000 38.100000 ;
        RECT 73.150000 49.715000 73.350000 49.915000 ;
        RECT 73.150000 50.135000 73.350000 50.335000 ;
        RECT 73.150000 50.555000 73.350000 50.755000 ;
        RECT 73.555000 34.820000 73.755000 35.020000 ;
        RECT 73.555000 35.260000 73.755000 35.460000 ;
        RECT 73.555000 35.700000 73.755000 35.900000 ;
        RECT 73.555000 36.140000 73.755000 36.340000 ;
        RECT 73.555000 36.580000 73.755000 36.780000 ;
        RECT 73.555000 37.020000 73.755000 37.220000 ;
        RECT 73.555000 37.460000 73.755000 37.660000 ;
        RECT 73.555000 37.900000 73.755000 38.100000 ;
        RECT 73.555000 49.715000 73.755000 49.915000 ;
        RECT 73.555000 50.135000 73.755000 50.335000 ;
        RECT 73.555000 50.555000 73.755000 50.755000 ;
        RECT 73.960000 34.820000 74.160000 35.020000 ;
        RECT 73.960000 35.260000 74.160000 35.460000 ;
        RECT 73.960000 35.700000 74.160000 35.900000 ;
        RECT 73.960000 36.140000 74.160000 36.340000 ;
        RECT 73.960000 36.580000 74.160000 36.780000 ;
        RECT 73.960000 37.020000 74.160000 37.220000 ;
        RECT 73.960000 37.460000 74.160000 37.660000 ;
        RECT 73.960000 37.900000 74.160000 38.100000 ;
        RECT 73.960000 49.715000 74.160000 49.915000 ;
        RECT 73.960000 50.135000 74.160000 50.335000 ;
        RECT 73.960000 50.555000 74.160000 50.755000 ;
        RECT 74.365000 34.820000 74.565000 35.020000 ;
        RECT 74.365000 35.260000 74.565000 35.460000 ;
        RECT 74.365000 35.700000 74.565000 35.900000 ;
        RECT 74.365000 36.140000 74.565000 36.340000 ;
        RECT 74.365000 36.580000 74.565000 36.780000 ;
        RECT 74.365000 37.020000 74.565000 37.220000 ;
        RECT 74.365000 37.460000 74.565000 37.660000 ;
        RECT 74.365000 37.900000 74.565000 38.100000 ;
        RECT 74.365000 49.715000 74.565000 49.915000 ;
        RECT 74.365000 50.135000 74.565000 50.335000 ;
        RECT 74.365000 50.555000 74.565000 50.755000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 39.585000 1.270000 44.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 39.585000 75.000000 44.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 39.685000 1.270000 44.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 23.835000 1.270000 28.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 23.835000 75.000000 28.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 173.785000 1.270000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 23.935000 1.270000 28.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 173.785000 75.000000 198.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 56.235000 1.270000 60.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.235000 75.000000 60.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 56.335000 1.270000 60.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 29.885000 1.270000 33.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 29.885000 75.000000 33.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 29.985000 1.270000 33.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 198.000000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 75.000000 198.000000 ;
    LAYER met3 ;
      RECT  0.000000  0.000000 75.000000  34.340000 ;
      RECT  0.000000 38.580000 75.000000  49.250000 ;
      RECT  0.000000 51.220000 75.000000 198.000000 ;
      RECT 24.800000  0.000000 50.355000 198.000000 ;
      RECT 24.800000  0.000000 50.355000 198.000000 ;
      RECT 24.800000 34.340000 50.355000  38.580000 ;
      RECT 24.800000 49.250000 50.355000  51.220000 ;
    LAYER met4 ;
      RECT  0.000000   5.885000  1.670000   6.485000 ;
      RECT  0.000000  11.935000  1.365000  12.535000 ;
      RECT  0.000000  16.785000  1.365000  17.385000 ;
      RECT  0.000000  22.835000  1.670000  23.435000 ;
      RECT  0.000000  28.885000  1.670000  29.485000 ;
      RECT  0.000000  33.735000  1.670000  34.335000 ;
      RECT  0.000000  38.585000  1.670000  39.185000 ;
      RECT  0.000000  44.635000  1.670000  45.335000 ;
      RECT  0.000000  55.135000  1.670000  55.835000 ;
      RECT  0.000000  61.085000  1.670000  61.685000 ;
      RECT  0.000000  66.935000  1.670000  67.635000 ;
      RECT  0.000000  93.400000 75.000000 173.385000 ;
      RECT  1.365000  11.935000 73.635000  17.385000 ;
      RECT  1.365000  11.935000 73.635000  17.385000 ;
      RECT  1.670000   0.000000 73.330000  11.935000 ;
      RECT  1.670000   0.000000 73.330000  34.335000 ;
      RECT  1.670000   0.000000 73.330000  34.335000 ;
      RECT  1.670000   0.000000 73.330000  34.335000 ;
      RECT  1.670000   0.000000 73.330000  34.335000 ;
      RECT  1.670000   0.000000 73.330000  34.335000 ;
      RECT  1.670000  17.385000 73.330000  34.335000 ;
      RECT  1.670000  38.585000 73.330000  49.245000 ;
      RECT  1.670000  38.585000 73.330000  49.245000 ;
      RECT  1.670000  38.585000 73.330000  49.245000 ;
      RECT  1.670000  51.225000 73.330000  93.400000 ;
      RECT  1.670000  51.225000 73.330000 198.000000 ;
      RECT  1.670000  51.225000 73.330000 198.000000 ;
      RECT  1.670000  51.225000 73.330000 198.000000 ;
      RECT  1.670000  51.225000 73.330000 198.000000 ;
      RECT  1.670000  51.225000 73.330000 198.000000 ;
      RECT  1.670000 173.385000 73.330000 198.000000 ;
      RECT 24.775000   0.000000 50.380000  51.225000 ;
      RECT 24.775000   0.000000 50.380000 198.000000 ;
      RECT 24.775000  34.335000 50.380000  38.585000 ;
      RECT 24.775000  49.245000 50.380000  51.225000 ;
      RECT 73.330000   5.885000 75.000000   6.485000 ;
      RECT 73.330000  22.835000 75.000000  23.435000 ;
      RECT 73.330000  28.885000 75.000000  29.485000 ;
      RECT 73.330000  33.735000 75.000000  34.335000 ;
      RECT 73.330000  38.585000 75.000000  39.185000 ;
      RECT 73.330000  44.635000 75.000000  45.335000 ;
      RECT 73.330000  55.135000 75.000000  55.835000 ;
      RECT 73.330000  61.085000 75.000000  61.685000 ;
      RECT 73.330000  66.935000 75.000000  67.635000 ;
      RECT 73.635000  11.935000 75.000000  12.535000 ;
      RECT 73.635000  16.785000 75.000000  17.385000 ;
    LAYER met5 ;
      RECT 0.000000  93.785000 75.000000 172.985000 ;
      RECT 1.765000  12.235000 73.235000  17.085000 ;
      RECT 2.070000   0.000000 72.930000  12.235000 ;
      RECT 2.070000  17.085000 72.930000  93.785000 ;
      RECT 2.070000 172.985000 72.930000 198.000000 ;
  END
END sky130_fd_io__overlay_vssa_lvc
END LIBRARY
