# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_io__overlay_vssio_hvc
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 75 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 1.270000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 8.885000 75.000000 13.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.985000 1.270000 13.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 2.035000 75.000000 7.485000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2.135000 1.270000 7.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035000 14.935000 75.000000 18.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 15.035000 0.965000 18.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 1.270000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 19.785000 75.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 70.035000 75.000000 95.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 19.885000 1.270000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 70.035000 1.270000 94.985000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 19.885000 75.000000 24.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 1.270000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 64.085000 75.000000 68.535000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 64.185000 1.270000 68.435000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 1.270000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 1.270000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 36.735000 75.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 47.735000 75.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 51.645000 75.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 56.405000 75.000000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 36.840000 1.270000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 47.735000 1.270000 56.735000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 36.840000 75.000000 40.085000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 1.270000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 41.585000 75.000000 46.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 41.685000 1.270000 46.135000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT  0.495000 173.155000 13.500000 195.340000 ;
        RECT  0.495000 195.340000 13.500000 195.490000 ;
        RECT  0.495000 195.490000 13.650000 195.640000 ;
        RECT  0.495000 195.640000 13.800000 195.790000 ;
        RECT  0.495000 195.790000 13.950000 195.940000 ;
        RECT  0.495000 195.940000 14.100000 196.090000 ;
        RECT  0.495000 196.090000 14.250000 196.240000 ;
        RECT  0.495000 196.240000 14.400000 196.390000 ;
        RECT  0.495000 196.390000 14.550000 196.540000 ;
        RECT  0.495000 196.540000 14.700000 196.690000 ;
        RECT  0.495000 196.690000 14.850000 196.840000 ;
        RECT  0.495000 196.840000 15.000000 196.990000 ;
        RECT  0.495000 196.990000 15.150000 197.140000 ;
        RECT  0.495000 197.140000 15.300000 197.175000 ;
        RECT  0.495000 197.175000 74.290000 200.000000 ;
        RECT 59.700000 197.110000 74.290000 197.175000 ;
        RECT 59.850000 196.960000 74.290000 197.110000 ;
        RECT 60.000000 196.810000 74.290000 196.960000 ;
        RECT 60.150000 196.660000 74.290000 196.810000 ;
        RECT 60.300000 196.510000 74.290000 196.660000 ;
        RECT 60.450000 196.360000 74.290000 196.510000 ;
        RECT 60.600000 196.210000 74.290000 196.360000 ;
        RECT 60.750000 196.060000 74.290000 196.210000 ;
        RECT 60.900000 195.910000 74.290000 196.060000 ;
        RECT 61.050000 195.760000 74.290000 195.910000 ;
        RECT 61.200000 195.610000 74.290000 195.760000 ;
        RECT 61.350000 195.460000 74.290000 195.610000 ;
        RECT 61.500000 173.320000 74.290000 195.310000 ;
        RECT 61.500000 195.310000 74.290000 195.460000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.495000 25.840000 24.395000 30.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000 25.840000 74.290000 30.480000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000  1.270000 175.930000 ;
        RECT 0.000000 175.930000 13.475000 199.920000 ;
        RECT 0.000000 199.920000  1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 24.370000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 13.595000 196.230000 14.255000 196.970000 ;
    END
    PORT
      LAYER met4 ;
        RECT 13.630000 197.170000 61.325000 199.930000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.415000 25.835000 75.000000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.680000 196.230000 61.340000 196.970000 ;
    END
    PORT
      LAYER met4 ;
        RECT 61.505000 175.930000 75.000000 199.920000 ;
        RECT 73.730000 175.785000 75.000000 175.930000 ;
        RECT 73.730000 199.920000 75.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 25.935000 1.270000 30.385000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 175.785000 75.000000 200.000000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.585000  25.910000  0.785000  26.110000 ;
        RECT  0.585000  26.340000  0.785000  26.540000 ;
        RECT  0.585000  26.770000  0.785000  26.970000 ;
        RECT  0.585000  27.200000  0.785000  27.400000 ;
        RECT  0.585000  27.630000  0.785000  27.830000 ;
        RECT  0.585000  28.060000  0.785000  28.260000 ;
        RECT  0.585000  28.490000  0.785000  28.690000 ;
        RECT  0.585000  28.920000  0.785000  29.120000 ;
        RECT  0.585000  29.350000  0.785000  29.550000 ;
        RECT  0.585000  29.780000  0.785000  29.980000 ;
        RECT  0.585000  30.210000  0.785000  30.410000 ;
        RECT  0.685000 175.995000  0.885000 176.195000 ;
        RECT  0.685000 176.395000  0.885000 176.595000 ;
        RECT  0.685000 176.795000  0.885000 176.995000 ;
        RECT  0.685000 177.195000  0.885000 177.395000 ;
        RECT  0.685000 177.595000  0.885000 177.795000 ;
        RECT  0.685000 177.995000  0.885000 178.195000 ;
        RECT  0.685000 178.395000  0.885000 178.595000 ;
        RECT  0.685000 178.795000  0.885000 178.995000 ;
        RECT  0.685000 179.195000  0.885000 179.395000 ;
        RECT  0.685000 179.595000  0.885000 179.795000 ;
        RECT  0.685000 179.995000  0.885000 180.195000 ;
        RECT  0.685000 180.395000  0.885000 180.595000 ;
        RECT  0.685000 180.795000  0.885000 180.995000 ;
        RECT  0.685000 181.195000  0.885000 181.395000 ;
        RECT  0.685000 181.595000  0.885000 181.795000 ;
        RECT  0.685000 181.995000  0.885000 182.195000 ;
        RECT  0.685000 182.395000  0.885000 182.595000 ;
        RECT  0.685000 182.795000  0.885000 182.995000 ;
        RECT  0.685000 183.195000  0.885000 183.395000 ;
        RECT  0.685000 183.595000  0.885000 183.795000 ;
        RECT  0.685000 183.995000  0.885000 184.195000 ;
        RECT  0.685000 184.395000  0.885000 184.595000 ;
        RECT  0.685000 184.795000  0.885000 184.995000 ;
        RECT  0.685000 185.195000  0.885000 185.395000 ;
        RECT  0.685000 185.595000  0.885000 185.795000 ;
        RECT  0.685000 185.995000  0.885000 186.195000 ;
        RECT  0.685000 186.395000  0.885000 186.595000 ;
        RECT  0.685000 186.795000  0.885000 186.995000 ;
        RECT  0.685000 187.195000  0.885000 187.395000 ;
        RECT  0.685000 187.595000  0.885000 187.795000 ;
        RECT  0.685000 187.995000  0.885000 188.195000 ;
        RECT  0.685000 188.395000  0.885000 188.595000 ;
        RECT  0.685000 188.795000  0.885000 188.995000 ;
        RECT  0.685000 189.195000  0.885000 189.395000 ;
        RECT  0.685000 189.595000  0.885000 189.795000 ;
        RECT  0.685000 189.995000  0.885000 190.195000 ;
        RECT  0.685000 190.395000  0.885000 190.595000 ;
        RECT  0.685000 190.795000  0.885000 190.995000 ;
        RECT  0.685000 191.195000  0.885000 191.395000 ;
        RECT  0.685000 191.595000  0.885000 191.795000 ;
        RECT  0.685000 191.995000  0.885000 192.195000 ;
        RECT  0.685000 192.395000  0.885000 192.595000 ;
        RECT  0.685000 192.795000  0.885000 192.995000 ;
        RECT  0.685000 193.195000  0.885000 193.395000 ;
        RECT  0.685000 193.595000  0.885000 193.795000 ;
        RECT  0.685000 193.995000  0.885000 194.195000 ;
        RECT  0.685000 194.395000  0.885000 194.595000 ;
        RECT  0.685000 194.795000  0.885000 194.995000 ;
        RECT  0.685000 195.200000  0.885000 195.400000 ;
        RECT  0.685000 195.605000  0.885000 195.805000 ;
        RECT  0.685000 196.010000  0.885000 196.210000 ;
        RECT  0.685000 196.415000  0.885000 196.615000 ;
        RECT  0.685000 196.820000  0.885000 197.020000 ;
        RECT  0.685000 197.225000  0.885000 197.425000 ;
        RECT  0.685000 197.630000  0.885000 197.830000 ;
        RECT  0.685000 198.035000  0.885000 198.235000 ;
        RECT  0.685000 198.440000  0.885000 198.640000 ;
        RECT  0.685000 198.845000  0.885000 199.045000 ;
        RECT  0.685000 199.250000  0.885000 199.450000 ;
        RECT  0.685000 199.655000  0.885000 199.855000 ;
        RECT  0.995000  25.910000  1.195000  26.110000 ;
        RECT  0.995000  26.340000  1.195000  26.540000 ;
        RECT  0.995000  26.770000  1.195000  26.970000 ;
        RECT  0.995000  27.200000  1.195000  27.400000 ;
        RECT  0.995000  27.630000  1.195000  27.830000 ;
        RECT  0.995000  28.060000  1.195000  28.260000 ;
        RECT  0.995000  28.490000  1.195000  28.690000 ;
        RECT  0.995000  28.920000  1.195000  29.120000 ;
        RECT  0.995000  29.350000  1.195000  29.550000 ;
        RECT  0.995000  29.780000  1.195000  29.980000 ;
        RECT  0.995000  30.210000  1.195000  30.410000 ;
        RECT  1.085000 175.995000  1.285000 176.195000 ;
        RECT  1.085000 176.395000  1.285000 176.595000 ;
        RECT  1.085000 176.795000  1.285000 176.995000 ;
        RECT  1.085000 177.195000  1.285000 177.395000 ;
        RECT  1.085000 177.595000  1.285000 177.795000 ;
        RECT  1.085000 177.995000  1.285000 178.195000 ;
        RECT  1.085000 178.395000  1.285000 178.595000 ;
        RECT  1.085000 178.795000  1.285000 178.995000 ;
        RECT  1.085000 179.195000  1.285000 179.395000 ;
        RECT  1.085000 179.595000  1.285000 179.795000 ;
        RECT  1.085000 179.995000  1.285000 180.195000 ;
        RECT  1.085000 180.395000  1.285000 180.595000 ;
        RECT  1.085000 180.795000  1.285000 180.995000 ;
        RECT  1.085000 181.195000  1.285000 181.395000 ;
        RECT  1.085000 181.595000  1.285000 181.795000 ;
        RECT  1.085000 181.995000  1.285000 182.195000 ;
        RECT  1.085000 182.395000  1.285000 182.595000 ;
        RECT  1.085000 182.795000  1.285000 182.995000 ;
        RECT  1.085000 183.195000  1.285000 183.395000 ;
        RECT  1.085000 183.595000  1.285000 183.795000 ;
        RECT  1.085000 183.995000  1.285000 184.195000 ;
        RECT  1.085000 184.395000  1.285000 184.595000 ;
        RECT  1.085000 184.795000  1.285000 184.995000 ;
        RECT  1.085000 185.195000  1.285000 185.395000 ;
        RECT  1.085000 185.595000  1.285000 185.795000 ;
        RECT  1.085000 185.995000  1.285000 186.195000 ;
        RECT  1.085000 186.395000  1.285000 186.595000 ;
        RECT  1.085000 186.795000  1.285000 186.995000 ;
        RECT  1.085000 187.195000  1.285000 187.395000 ;
        RECT  1.085000 187.595000  1.285000 187.795000 ;
        RECT  1.085000 187.995000  1.285000 188.195000 ;
        RECT  1.085000 188.395000  1.285000 188.595000 ;
        RECT  1.085000 188.795000  1.285000 188.995000 ;
        RECT  1.085000 189.195000  1.285000 189.395000 ;
        RECT  1.085000 189.595000  1.285000 189.795000 ;
        RECT  1.085000 189.995000  1.285000 190.195000 ;
        RECT  1.085000 190.395000  1.285000 190.595000 ;
        RECT  1.085000 190.795000  1.285000 190.995000 ;
        RECT  1.085000 191.195000  1.285000 191.395000 ;
        RECT  1.085000 191.595000  1.285000 191.795000 ;
        RECT  1.085000 191.995000  1.285000 192.195000 ;
        RECT  1.085000 192.395000  1.285000 192.595000 ;
        RECT  1.085000 192.795000  1.285000 192.995000 ;
        RECT  1.085000 193.195000  1.285000 193.395000 ;
        RECT  1.085000 193.595000  1.285000 193.795000 ;
        RECT  1.085000 193.995000  1.285000 194.195000 ;
        RECT  1.085000 194.395000  1.285000 194.595000 ;
        RECT  1.085000 194.795000  1.285000 194.995000 ;
        RECT  1.085000 195.200000  1.285000 195.400000 ;
        RECT  1.085000 195.605000  1.285000 195.805000 ;
        RECT  1.085000 196.010000  1.285000 196.210000 ;
        RECT  1.085000 196.415000  1.285000 196.615000 ;
        RECT  1.085000 196.820000  1.285000 197.020000 ;
        RECT  1.085000 197.225000  1.285000 197.425000 ;
        RECT  1.085000 197.630000  1.285000 197.830000 ;
        RECT  1.085000 198.035000  1.285000 198.235000 ;
        RECT  1.085000 198.440000  1.285000 198.640000 ;
        RECT  1.085000 198.845000  1.285000 199.045000 ;
        RECT  1.085000 199.250000  1.285000 199.450000 ;
        RECT  1.085000 199.655000  1.285000 199.855000 ;
        RECT  1.405000  25.910000  1.605000  26.110000 ;
        RECT  1.405000  26.340000  1.605000  26.540000 ;
        RECT  1.405000  26.770000  1.605000  26.970000 ;
        RECT  1.405000  27.200000  1.605000  27.400000 ;
        RECT  1.405000  27.630000  1.605000  27.830000 ;
        RECT  1.405000  28.060000  1.605000  28.260000 ;
        RECT  1.405000  28.490000  1.605000  28.690000 ;
        RECT  1.405000  28.920000  1.605000  29.120000 ;
        RECT  1.405000  29.350000  1.605000  29.550000 ;
        RECT  1.405000  29.780000  1.605000  29.980000 ;
        RECT  1.405000  30.210000  1.605000  30.410000 ;
        RECT  1.485000 175.995000  1.685000 176.195000 ;
        RECT  1.485000 176.395000  1.685000 176.595000 ;
        RECT  1.485000 176.795000  1.685000 176.995000 ;
        RECT  1.485000 177.195000  1.685000 177.395000 ;
        RECT  1.485000 177.595000  1.685000 177.795000 ;
        RECT  1.485000 177.995000  1.685000 178.195000 ;
        RECT  1.485000 178.395000  1.685000 178.595000 ;
        RECT  1.485000 178.795000  1.685000 178.995000 ;
        RECT  1.485000 179.195000  1.685000 179.395000 ;
        RECT  1.485000 179.595000  1.685000 179.795000 ;
        RECT  1.485000 179.995000  1.685000 180.195000 ;
        RECT  1.485000 180.395000  1.685000 180.595000 ;
        RECT  1.485000 180.795000  1.685000 180.995000 ;
        RECT  1.485000 181.195000  1.685000 181.395000 ;
        RECT  1.485000 181.595000  1.685000 181.795000 ;
        RECT  1.485000 181.995000  1.685000 182.195000 ;
        RECT  1.485000 182.395000  1.685000 182.595000 ;
        RECT  1.485000 182.795000  1.685000 182.995000 ;
        RECT  1.485000 183.195000  1.685000 183.395000 ;
        RECT  1.485000 183.595000  1.685000 183.795000 ;
        RECT  1.485000 183.995000  1.685000 184.195000 ;
        RECT  1.485000 184.395000  1.685000 184.595000 ;
        RECT  1.485000 184.795000  1.685000 184.995000 ;
        RECT  1.485000 185.195000  1.685000 185.395000 ;
        RECT  1.485000 185.595000  1.685000 185.795000 ;
        RECT  1.485000 185.995000  1.685000 186.195000 ;
        RECT  1.485000 186.395000  1.685000 186.595000 ;
        RECT  1.485000 186.795000  1.685000 186.995000 ;
        RECT  1.485000 187.195000  1.685000 187.395000 ;
        RECT  1.485000 187.595000  1.685000 187.795000 ;
        RECT  1.485000 187.995000  1.685000 188.195000 ;
        RECT  1.485000 188.395000  1.685000 188.595000 ;
        RECT  1.485000 188.795000  1.685000 188.995000 ;
        RECT  1.485000 189.195000  1.685000 189.395000 ;
        RECT  1.485000 189.595000  1.685000 189.795000 ;
        RECT  1.485000 189.995000  1.685000 190.195000 ;
        RECT  1.485000 190.395000  1.685000 190.595000 ;
        RECT  1.485000 190.795000  1.685000 190.995000 ;
        RECT  1.485000 191.195000  1.685000 191.395000 ;
        RECT  1.485000 191.595000  1.685000 191.795000 ;
        RECT  1.485000 191.995000  1.685000 192.195000 ;
        RECT  1.485000 192.395000  1.685000 192.595000 ;
        RECT  1.485000 192.795000  1.685000 192.995000 ;
        RECT  1.485000 193.195000  1.685000 193.395000 ;
        RECT  1.485000 193.595000  1.685000 193.795000 ;
        RECT  1.485000 193.995000  1.685000 194.195000 ;
        RECT  1.485000 194.395000  1.685000 194.595000 ;
        RECT  1.485000 194.795000  1.685000 194.995000 ;
        RECT  1.485000 195.200000  1.685000 195.400000 ;
        RECT  1.485000 195.605000  1.685000 195.805000 ;
        RECT  1.485000 196.010000  1.685000 196.210000 ;
        RECT  1.485000 196.415000  1.685000 196.615000 ;
        RECT  1.485000 196.820000  1.685000 197.020000 ;
        RECT  1.485000 197.225000  1.685000 197.425000 ;
        RECT  1.485000 197.630000  1.685000 197.830000 ;
        RECT  1.485000 198.035000  1.685000 198.235000 ;
        RECT  1.485000 198.440000  1.685000 198.640000 ;
        RECT  1.485000 198.845000  1.685000 199.045000 ;
        RECT  1.485000 199.250000  1.685000 199.450000 ;
        RECT  1.485000 199.655000  1.685000 199.855000 ;
        RECT  1.815000  25.910000  2.015000  26.110000 ;
        RECT  1.815000  26.340000  2.015000  26.540000 ;
        RECT  1.815000  26.770000  2.015000  26.970000 ;
        RECT  1.815000  27.200000  2.015000  27.400000 ;
        RECT  1.815000  27.630000  2.015000  27.830000 ;
        RECT  1.815000  28.060000  2.015000  28.260000 ;
        RECT  1.815000  28.490000  2.015000  28.690000 ;
        RECT  1.815000  28.920000  2.015000  29.120000 ;
        RECT  1.815000  29.350000  2.015000  29.550000 ;
        RECT  1.815000  29.780000  2.015000  29.980000 ;
        RECT  1.815000  30.210000  2.015000  30.410000 ;
        RECT  1.885000 175.995000  2.085000 176.195000 ;
        RECT  1.885000 176.395000  2.085000 176.595000 ;
        RECT  1.885000 176.795000  2.085000 176.995000 ;
        RECT  1.885000 177.195000  2.085000 177.395000 ;
        RECT  1.885000 177.595000  2.085000 177.795000 ;
        RECT  1.885000 177.995000  2.085000 178.195000 ;
        RECT  1.885000 178.395000  2.085000 178.595000 ;
        RECT  1.885000 178.795000  2.085000 178.995000 ;
        RECT  1.885000 179.195000  2.085000 179.395000 ;
        RECT  1.885000 179.595000  2.085000 179.795000 ;
        RECT  1.885000 179.995000  2.085000 180.195000 ;
        RECT  1.885000 180.395000  2.085000 180.595000 ;
        RECT  1.885000 180.795000  2.085000 180.995000 ;
        RECT  1.885000 181.195000  2.085000 181.395000 ;
        RECT  1.885000 181.595000  2.085000 181.795000 ;
        RECT  1.885000 181.995000  2.085000 182.195000 ;
        RECT  1.885000 182.395000  2.085000 182.595000 ;
        RECT  1.885000 182.795000  2.085000 182.995000 ;
        RECT  1.885000 183.195000  2.085000 183.395000 ;
        RECT  1.885000 183.595000  2.085000 183.795000 ;
        RECT  1.885000 183.995000  2.085000 184.195000 ;
        RECT  1.885000 184.395000  2.085000 184.595000 ;
        RECT  1.885000 184.795000  2.085000 184.995000 ;
        RECT  1.885000 185.195000  2.085000 185.395000 ;
        RECT  1.885000 185.595000  2.085000 185.795000 ;
        RECT  1.885000 185.995000  2.085000 186.195000 ;
        RECT  1.885000 186.395000  2.085000 186.595000 ;
        RECT  1.885000 186.795000  2.085000 186.995000 ;
        RECT  1.885000 187.195000  2.085000 187.395000 ;
        RECT  1.885000 187.595000  2.085000 187.795000 ;
        RECT  1.885000 187.995000  2.085000 188.195000 ;
        RECT  1.885000 188.395000  2.085000 188.595000 ;
        RECT  1.885000 188.795000  2.085000 188.995000 ;
        RECT  1.885000 189.195000  2.085000 189.395000 ;
        RECT  1.885000 189.595000  2.085000 189.795000 ;
        RECT  1.885000 189.995000  2.085000 190.195000 ;
        RECT  1.885000 190.395000  2.085000 190.595000 ;
        RECT  1.885000 190.795000  2.085000 190.995000 ;
        RECT  1.885000 191.195000  2.085000 191.395000 ;
        RECT  1.885000 191.595000  2.085000 191.795000 ;
        RECT  1.885000 191.995000  2.085000 192.195000 ;
        RECT  1.885000 192.395000  2.085000 192.595000 ;
        RECT  1.885000 192.795000  2.085000 192.995000 ;
        RECT  1.885000 193.195000  2.085000 193.395000 ;
        RECT  1.885000 193.595000  2.085000 193.795000 ;
        RECT  1.885000 193.995000  2.085000 194.195000 ;
        RECT  1.885000 194.395000  2.085000 194.595000 ;
        RECT  1.885000 194.795000  2.085000 194.995000 ;
        RECT  1.885000 195.200000  2.085000 195.400000 ;
        RECT  1.885000 195.605000  2.085000 195.805000 ;
        RECT  1.885000 196.010000  2.085000 196.210000 ;
        RECT  1.885000 196.415000  2.085000 196.615000 ;
        RECT  1.885000 196.820000  2.085000 197.020000 ;
        RECT  1.885000 197.225000  2.085000 197.425000 ;
        RECT  1.885000 197.630000  2.085000 197.830000 ;
        RECT  1.885000 198.035000  2.085000 198.235000 ;
        RECT  1.885000 198.440000  2.085000 198.640000 ;
        RECT  1.885000 198.845000  2.085000 199.045000 ;
        RECT  1.885000 199.250000  2.085000 199.450000 ;
        RECT  1.885000 199.655000  2.085000 199.855000 ;
        RECT  2.225000  25.910000  2.425000  26.110000 ;
        RECT  2.225000  26.340000  2.425000  26.540000 ;
        RECT  2.225000  26.770000  2.425000  26.970000 ;
        RECT  2.225000  27.200000  2.425000  27.400000 ;
        RECT  2.225000  27.630000  2.425000  27.830000 ;
        RECT  2.225000  28.060000  2.425000  28.260000 ;
        RECT  2.225000  28.490000  2.425000  28.690000 ;
        RECT  2.225000  28.920000  2.425000  29.120000 ;
        RECT  2.225000  29.350000  2.425000  29.550000 ;
        RECT  2.225000  29.780000  2.425000  29.980000 ;
        RECT  2.225000  30.210000  2.425000  30.410000 ;
        RECT  2.285000 175.995000  2.485000 176.195000 ;
        RECT  2.285000 176.395000  2.485000 176.595000 ;
        RECT  2.285000 176.795000  2.485000 176.995000 ;
        RECT  2.285000 177.195000  2.485000 177.395000 ;
        RECT  2.285000 177.595000  2.485000 177.795000 ;
        RECT  2.285000 177.995000  2.485000 178.195000 ;
        RECT  2.285000 178.395000  2.485000 178.595000 ;
        RECT  2.285000 178.795000  2.485000 178.995000 ;
        RECT  2.285000 179.195000  2.485000 179.395000 ;
        RECT  2.285000 179.595000  2.485000 179.795000 ;
        RECT  2.285000 179.995000  2.485000 180.195000 ;
        RECT  2.285000 180.395000  2.485000 180.595000 ;
        RECT  2.285000 180.795000  2.485000 180.995000 ;
        RECT  2.285000 181.195000  2.485000 181.395000 ;
        RECT  2.285000 181.595000  2.485000 181.795000 ;
        RECT  2.285000 181.995000  2.485000 182.195000 ;
        RECT  2.285000 182.395000  2.485000 182.595000 ;
        RECT  2.285000 182.795000  2.485000 182.995000 ;
        RECT  2.285000 183.195000  2.485000 183.395000 ;
        RECT  2.285000 183.595000  2.485000 183.795000 ;
        RECT  2.285000 183.995000  2.485000 184.195000 ;
        RECT  2.285000 184.395000  2.485000 184.595000 ;
        RECT  2.285000 184.795000  2.485000 184.995000 ;
        RECT  2.285000 185.195000  2.485000 185.395000 ;
        RECT  2.285000 185.595000  2.485000 185.795000 ;
        RECT  2.285000 185.995000  2.485000 186.195000 ;
        RECT  2.285000 186.395000  2.485000 186.595000 ;
        RECT  2.285000 186.795000  2.485000 186.995000 ;
        RECT  2.285000 187.195000  2.485000 187.395000 ;
        RECT  2.285000 187.595000  2.485000 187.795000 ;
        RECT  2.285000 187.995000  2.485000 188.195000 ;
        RECT  2.285000 188.395000  2.485000 188.595000 ;
        RECT  2.285000 188.795000  2.485000 188.995000 ;
        RECT  2.285000 189.195000  2.485000 189.395000 ;
        RECT  2.285000 189.595000  2.485000 189.795000 ;
        RECT  2.285000 189.995000  2.485000 190.195000 ;
        RECT  2.285000 190.395000  2.485000 190.595000 ;
        RECT  2.285000 190.795000  2.485000 190.995000 ;
        RECT  2.285000 191.195000  2.485000 191.395000 ;
        RECT  2.285000 191.595000  2.485000 191.795000 ;
        RECT  2.285000 191.995000  2.485000 192.195000 ;
        RECT  2.285000 192.395000  2.485000 192.595000 ;
        RECT  2.285000 192.795000  2.485000 192.995000 ;
        RECT  2.285000 193.195000  2.485000 193.395000 ;
        RECT  2.285000 193.595000  2.485000 193.795000 ;
        RECT  2.285000 193.995000  2.485000 194.195000 ;
        RECT  2.285000 194.395000  2.485000 194.595000 ;
        RECT  2.285000 194.795000  2.485000 194.995000 ;
        RECT  2.285000 195.200000  2.485000 195.400000 ;
        RECT  2.285000 195.605000  2.485000 195.805000 ;
        RECT  2.285000 196.010000  2.485000 196.210000 ;
        RECT  2.285000 196.415000  2.485000 196.615000 ;
        RECT  2.285000 196.820000  2.485000 197.020000 ;
        RECT  2.285000 197.225000  2.485000 197.425000 ;
        RECT  2.285000 197.630000  2.485000 197.830000 ;
        RECT  2.285000 198.035000  2.485000 198.235000 ;
        RECT  2.285000 198.440000  2.485000 198.640000 ;
        RECT  2.285000 198.845000  2.485000 199.045000 ;
        RECT  2.285000 199.250000  2.485000 199.450000 ;
        RECT  2.285000 199.655000  2.485000 199.855000 ;
        RECT  2.635000  25.910000  2.835000  26.110000 ;
        RECT  2.635000  26.340000  2.835000  26.540000 ;
        RECT  2.635000  26.770000  2.835000  26.970000 ;
        RECT  2.635000  27.200000  2.835000  27.400000 ;
        RECT  2.635000  27.630000  2.835000  27.830000 ;
        RECT  2.635000  28.060000  2.835000  28.260000 ;
        RECT  2.635000  28.490000  2.835000  28.690000 ;
        RECT  2.635000  28.920000  2.835000  29.120000 ;
        RECT  2.635000  29.350000  2.835000  29.550000 ;
        RECT  2.635000  29.780000  2.835000  29.980000 ;
        RECT  2.635000  30.210000  2.835000  30.410000 ;
        RECT  2.685000 175.995000  2.885000 176.195000 ;
        RECT  2.685000 176.395000  2.885000 176.595000 ;
        RECT  2.685000 176.795000  2.885000 176.995000 ;
        RECT  2.685000 177.195000  2.885000 177.395000 ;
        RECT  2.685000 177.595000  2.885000 177.795000 ;
        RECT  2.685000 177.995000  2.885000 178.195000 ;
        RECT  2.685000 178.395000  2.885000 178.595000 ;
        RECT  2.685000 178.795000  2.885000 178.995000 ;
        RECT  2.685000 179.195000  2.885000 179.395000 ;
        RECT  2.685000 179.595000  2.885000 179.795000 ;
        RECT  2.685000 179.995000  2.885000 180.195000 ;
        RECT  2.685000 180.395000  2.885000 180.595000 ;
        RECT  2.685000 180.795000  2.885000 180.995000 ;
        RECT  2.685000 181.195000  2.885000 181.395000 ;
        RECT  2.685000 181.595000  2.885000 181.795000 ;
        RECT  2.685000 181.995000  2.885000 182.195000 ;
        RECT  2.685000 182.395000  2.885000 182.595000 ;
        RECT  2.685000 182.795000  2.885000 182.995000 ;
        RECT  2.685000 183.195000  2.885000 183.395000 ;
        RECT  2.685000 183.595000  2.885000 183.795000 ;
        RECT  2.685000 183.995000  2.885000 184.195000 ;
        RECT  2.685000 184.395000  2.885000 184.595000 ;
        RECT  2.685000 184.795000  2.885000 184.995000 ;
        RECT  2.685000 185.195000  2.885000 185.395000 ;
        RECT  2.685000 185.595000  2.885000 185.795000 ;
        RECT  2.685000 185.995000  2.885000 186.195000 ;
        RECT  2.685000 186.395000  2.885000 186.595000 ;
        RECT  2.685000 186.795000  2.885000 186.995000 ;
        RECT  2.685000 187.195000  2.885000 187.395000 ;
        RECT  2.685000 187.595000  2.885000 187.795000 ;
        RECT  2.685000 187.995000  2.885000 188.195000 ;
        RECT  2.685000 188.395000  2.885000 188.595000 ;
        RECT  2.685000 188.795000  2.885000 188.995000 ;
        RECT  2.685000 189.195000  2.885000 189.395000 ;
        RECT  2.685000 189.595000  2.885000 189.795000 ;
        RECT  2.685000 189.995000  2.885000 190.195000 ;
        RECT  2.685000 190.395000  2.885000 190.595000 ;
        RECT  2.685000 190.795000  2.885000 190.995000 ;
        RECT  2.685000 191.195000  2.885000 191.395000 ;
        RECT  2.685000 191.595000  2.885000 191.795000 ;
        RECT  2.685000 191.995000  2.885000 192.195000 ;
        RECT  2.685000 192.395000  2.885000 192.595000 ;
        RECT  2.685000 192.795000  2.885000 192.995000 ;
        RECT  2.685000 193.195000  2.885000 193.395000 ;
        RECT  2.685000 193.595000  2.885000 193.795000 ;
        RECT  2.685000 193.995000  2.885000 194.195000 ;
        RECT  2.685000 194.395000  2.885000 194.595000 ;
        RECT  2.685000 194.795000  2.885000 194.995000 ;
        RECT  2.685000 195.200000  2.885000 195.400000 ;
        RECT  2.685000 195.605000  2.885000 195.805000 ;
        RECT  2.685000 196.010000  2.885000 196.210000 ;
        RECT  2.685000 196.415000  2.885000 196.615000 ;
        RECT  2.685000 196.820000  2.885000 197.020000 ;
        RECT  2.685000 197.225000  2.885000 197.425000 ;
        RECT  2.685000 197.630000  2.885000 197.830000 ;
        RECT  2.685000 198.035000  2.885000 198.235000 ;
        RECT  2.685000 198.440000  2.885000 198.640000 ;
        RECT  2.685000 198.845000  2.885000 199.045000 ;
        RECT  2.685000 199.250000  2.885000 199.450000 ;
        RECT  2.685000 199.655000  2.885000 199.855000 ;
        RECT  3.045000  25.910000  3.245000  26.110000 ;
        RECT  3.045000  26.340000  3.245000  26.540000 ;
        RECT  3.045000  26.770000  3.245000  26.970000 ;
        RECT  3.045000  27.200000  3.245000  27.400000 ;
        RECT  3.045000  27.630000  3.245000  27.830000 ;
        RECT  3.045000  28.060000  3.245000  28.260000 ;
        RECT  3.045000  28.490000  3.245000  28.690000 ;
        RECT  3.045000  28.920000  3.245000  29.120000 ;
        RECT  3.045000  29.350000  3.245000  29.550000 ;
        RECT  3.045000  29.780000  3.245000  29.980000 ;
        RECT  3.045000  30.210000  3.245000  30.410000 ;
        RECT  3.085000 175.995000  3.285000 176.195000 ;
        RECT  3.085000 176.395000  3.285000 176.595000 ;
        RECT  3.085000 176.795000  3.285000 176.995000 ;
        RECT  3.085000 177.195000  3.285000 177.395000 ;
        RECT  3.085000 177.595000  3.285000 177.795000 ;
        RECT  3.085000 177.995000  3.285000 178.195000 ;
        RECT  3.085000 178.395000  3.285000 178.595000 ;
        RECT  3.085000 178.795000  3.285000 178.995000 ;
        RECT  3.085000 179.195000  3.285000 179.395000 ;
        RECT  3.085000 179.595000  3.285000 179.795000 ;
        RECT  3.085000 179.995000  3.285000 180.195000 ;
        RECT  3.085000 180.395000  3.285000 180.595000 ;
        RECT  3.085000 180.795000  3.285000 180.995000 ;
        RECT  3.085000 181.195000  3.285000 181.395000 ;
        RECT  3.085000 181.595000  3.285000 181.795000 ;
        RECT  3.085000 181.995000  3.285000 182.195000 ;
        RECT  3.085000 182.395000  3.285000 182.595000 ;
        RECT  3.085000 182.795000  3.285000 182.995000 ;
        RECT  3.085000 183.195000  3.285000 183.395000 ;
        RECT  3.085000 183.595000  3.285000 183.795000 ;
        RECT  3.085000 183.995000  3.285000 184.195000 ;
        RECT  3.085000 184.395000  3.285000 184.595000 ;
        RECT  3.085000 184.795000  3.285000 184.995000 ;
        RECT  3.085000 185.195000  3.285000 185.395000 ;
        RECT  3.085000 185.595000  3.285000 185.795000 ;
        RECT  3.085000 185.995000  3.285000 186.195000 ;
        RECT  3.085000 186.395000  3.285000 186.595000 ;
        RECT  3.085000 186.795000  3.285000 186.995000 ;
        RECT  3.085000 187.195000  3.285000 187.395000 ;
        RECT  3.085000 187.595000  3.285000 187.795000 ;
        RECT  3.085000 187.995000  3.285000 188.195000 ;
        RECT  3.085000 188.395000  3.285000 188.595000 ;
        RECT  3.085000 188.795000  3.285000 188.995000 ;
        RECT  3.085000 189.195000  3.285000 189.395000 ;
        RECT  3.085000 189.595000  3.285000 189.795000 ;
        RECT  3.085000 189.995000  3.285000 190.195000 ;
        RECT  3.085000 190.395000  3.285000 190.595000 ;
        RECT  3.085000 190.795000  3.285000 190.995000 ;
        RECT  3.085000 191.195000  3.285000 191.395000 ;
        RECT  3.085000 191.595000  3.285000 191.795000 ;
        RECT  3.085000 191.995000  3.285000 192.195000 ;
        RECT  3.085000 192.395000  3.285000 192.595000 ;
        RECT  3.085000 192.795000  3.285000 192.995000 ;
        RECT  3.085000 193.195000  3.285000 193.395000 ;
        RECT  3.085000 193.595000  3.285000 193.795000 ;
        RECT  3.085000 193.995000  3.285000 194.195000 ;
        RECT  3.085000 194.395000  3.285000 194.595000 ;
        RECT  3.085000 194.795000  3.285000 194.995000 ;
        RECT  3.085000 195.200000  3.285000 195.400000 ;
        RECT  3.085000 195.605000  3.285000 195.805000 ;
        RECT  3.085000 196.010000  3.285000 196.210000 ;
        RECT  3.085000 196.415000  3.285000 196.615000 ;
        RECT  3.085000 196.820000  3.285000 197.020000 ;
        RECT  3.085000 197.225000  3.285000 197.425000 ;
        RECT  3.085000 197.630000  3.285000 197.830000 ;
        RECT  3.085000 198.035000  3.285000 198.235000 ;
        RECT  3.085000 198.440000  3.285000 198.640000 ;
        RECT  3.085000 198.845000  3.285000 199.045000 ;
        RECT  3.085000 199.250000  3.285000 199.450000 ;
        RECT  3.085000 199.655000  3.285000 199.855000 ;
        RECT  3.450000  25.910000  3.650000  26.110000 ;
        RECT  3.450000  26.340000  3.650000  26.540000 ;
        RECT  3.450000  26.770000  3.650000  26.970000 ;
        RECT  3.450000  27.200000  3.650000  27.400000 ;
        RECT  3.450000  27.630000  3.650000  27.830000 ;
        RECT  3.450000  28.060000  3.650000  28.260000 ;
        RECT  3.450000  28.490000  3.650000  28.690000 ;
        RECT  3.450000  28.920000  3.650000  29.120000 ;
        RECT  3.450000  29.350000  3.650000  29.550000 ;
        RECT  3.450000  29.780000  3.650000  29.980000 ;
        RECT  3.450000  30.210000  3.650000  30.410000 ;
        RECT  3.485000 175.995000  3.685000 176.195000 ;
        RECT  3.485000 176.395000  3.685000 176.595000 ;
        RECT  3.485000 176.795000  3.685000 176.995000 ;
        RECT  3.485000 177.195000  3.685000 177.395000 ;
        RECT  3.485000 177.595000  3.685000 177.795000 ;
        RECT  3.485000 177.995000  3.685000 178.195000 ;
        RECT  3.485000 178.395000  3.685000 178.595000 ;
        RECT  3.485000 178.795000  3.685000 178.995000 ;
        RECT  3.485000 179.195000  3.685000 179.395000 ;
        RECT  3.485000 179.595000  3.685000 179.795000 ;
        RECT  3.485000 179.995000  3.685000 180.195000 ;
        RECT  3.485000 180.395000  3.685000 180.595000 ;
        RECT  3.485000 180.795000  3.685000 180.995000 ;
        RECT  3.485000 181.195000  3.685000 181.395000 ;
        RECT  3.485000 181.595000  3.685000 181.795000 ;
        RECT  3.485000 181.995000  3.685000 182.195000 ;
        RECT  3.485000 182.395000  3.685000 182.595000 ;
        RECT  3.485000 182.795000  3.685000 182.995000 ;
        RECT  3.485000 183.195000  3.685000 183.395000 ;
        RECT  3.485000 183.595000  3.685000 183.795000 ;
        RECT  3.485000 183.995000  3.685000 184.195000 ;
        RECT  3.485000 184.395000  3.685000 184.595000 ;
        RECT  3.485000 184.795000  3.685000 184.995000 ;
        RECT  3.485000 185.195000  3.685000 185.395000 ;
        RECT  3.485000 185.595000  3.685000 185.795000 ;
        RECT  3.485000 185.995000  3.685000 186.195000 ;
        RECT  3.485000 186.395000  3.685000 186.595000 ;
        RECT  3.485000 186.795000  3.685000 186.995000 ;
        RECT  3.485000 187.195000  3.685000 187.395000 ;
        RECT  3.485000 187.595000  3.685000 187.795000 ;
        RECT  3.485000 187.995000  3.685000 188.195000 ;
        RECT  3.485000 188.395000  3.685000 188.595000 ;
        RECT  3.485000 188.795000  3.685000 188.995000 ;
        RECT  3.485000 189.195000  3.685000 189.395000 ;
        RECT  3.485000 189.595000  3.685000 189.795000 ;
        RECT  3.485000 189.995000  3.685000 190.195000 ;
        RECT  3.485000 190.395000  3.685000 190.595000 ;
        RECT  3.485000 190.795000  3.685000 190.995000 ;
        RECT  3.485000 191.195000  3.685000 191.395000 ;
        RECT  3.485000 191.595000  3.685000 191.795000 ;
        RECT  3.485000 191.995000  3.685000 192.195000 ;
        RECT  3.485000 192.395000  3.685000 192.595000 ;
        RECT  3.485000 192.795000  3.685000 192.995000 ;
        RECT  3.485000 193.195000  3.685000 193.395000 ;
        RECT  3.485000 193.595000  3.685000 193.795000 ;
        RECT  3.485000 193.995000  3.685000 194.195000 ;
        RECT  3.485000 194.395000  3.685000 194.595000 ;
        RECT  3.485000 194.795000  3.685000 194.995000 ;
        RECT  3.485000 195.200000  3.685000 195.400000 ;
        RECT  3.485000 195.605000  3.685000 195.805000 ;
        RECT  3.485000 196.010000  3.685000 196.210000 ;
        RECT  3.485000 196.415000  3.685000 196.615000 ;
        RECT  3.485000 196.820000  3.685000 197.020000 ;
        RECT  3.485000 197.225000  3.685000 197.425000 ;
        RECT  3.485000 197.630000  3.685000 197.830000 ;
        RECT  3.485000 198.035000  3.685000 198.235000 ;
        RECT  3.485000 198.440000  3.685000 198.640000 ;
        RECT  3.485000 198.845000  3.685000 199.045000 ;
        RECT  3.485000 199.250000  3.685000 199.450000 ;
        RECT  3.485000 199.655000  3.685000 199.855000 ;
        RECT  3.855000  25.910000  4.055000  26.110000 ;
        RECT  3.855000  26.340000  4.055000  26.540000 ;
        RECT  3.855000  26.770000  4.055000  26.970000 ;
        RECT  3.855000  27.200000  4.055000  27.400000 ;
        RECT  3.855000  27.630000  4.055000  27.830000 ;
        RECT  3.855000  28.060000  4.055000  28.260000 ;
        RECT  3.855000  28.490000  4.055000  28.690000 ;
        RECT  3.855000  28.920000  4.055000  29.120000 ;
        RECT  3.855000  29.350000  4.055000  29.550000 ;
        RECT  3.855000  29.780000  4.055000  29.980000 ;
        RECT  3.855000  30.210000  4.055000  30.410000 ;
        RECT  3.885000 175.995000  4.085000 176.195000 ;
        RECT  3.885000 176.395000  4.085000 176.595000 ;
        RECT  3.885000 176.795000  4.085000 176.995000 ;
        RECT  3.885000 177.195000  4.085000 177.395000 ;
        RECT  3.885000 177.595000  4.085000 177.795000 ;
        RECT  3.885000 177.995000  4.085000 178.195000 ;
        RECT  3.885000 178.395000  4.085000 178.595000 ;
        RECT  3.885000 178.795000  4.085000 178.995000 ;
        RECT  3.885000 179.195000  4.085000 179.395000 ;
        RECT  3.885000 179.595000  4.085000 179.795000 ;
        RECT  3.885000 179.995000  4.085000 180.195000 ;
        RECT  3.885000 180.395000  4.085000 180.595000 ;
        RECT  3.885000 180.795000  4.085000 180.995000 ;
        RECT  3.885000 181.195000  4.085000 181.395000 ;
        RECT  3.885000 181.595000  4.085000 181.795000 ;
        RECT  3.885000 181.995000  4.085000 182.195000 ;
        RECT  3.885000 182.395000  4.085000 182.595000 ;
        RECT  3.885000 182.795000  4.085000 182.995000 ;
        RECT  3.885000 183.195000  4.085000 183.395000 ;
        RECT  3.885000 183.595000  4.085000 183.795000 ;
        RECT  3.885000 183.995000  4.085000 184.195000 ;
        RECT  3.885000 184.395000  4.085000 184.595000 ;
        RECT  3.885000 184.795000  4.085000 184.995000 ;
        RECT  3.885000 185.195000  4.085000 185.395000 ;
        RECT  3.885000 185.595000  4.085000 185.795000 ;
        RECT  3.885000 185.995000  4.085000 186.195000 ;
        RECT  3.885000 186.395000  4.085000 186.595000 ;
        RECT  3.885000 186.795000  4.085000 186.995000 ;
        RECT  3.885000 187.195000  4.085000 187.395000 ;
        RECT  3.885000 187.595000  4.085000 187.795000 ;
        RECT  3.885000 187.995000  4.085000 188.195000 ;
        RECT  3.885000 188.395000  4.085000 188.595000 ;
        RECT  3.885000 188.795000  4.085000 188.995000 ;
        RECT  3.885000 189.195000  4.085000 189.395000 ;
        RECT  3.885000 189.595000  4.085000 189.795000 ;
        RECT  3.885000 189.995000  4.085000 190.195000 ;
        RECT  3.885000 190.395000  4.085000 190.595000 ;
        RECT  3.885000 190.795000  4.085000 190.995000 ;
        RECT  3.885000 191.195000  4.085000 191.395000 ;
        RECT  3.885000 191.595000  4.085000 191.795000 ;
        RECT  3.885000 191.995000  4.085000 192.195000 ;
        RECT  3.885000 192.395000  4.085000 192.595000 ;
        RECT  3.885000 192.795000  4.085000 192.995000 ;
        RECT  3.885000 193.195000  4.085000 193.395000 ;
        RECT  3.885000 193.595000  4.085000 193.795000 ;
        RECT  3.885000 193.995000  4.085000 194.195000 ;
        RECT  3.885000 194.395000  4.085000 194.595000 ;
        RECT  3.885000 194.795000  4.085000 194.995000 ;
        RECT  3.885000 195.200000  4.085000 195.400000 ;
        RECT  3.885000 195.605000  4.085000 195.805000 ;
        RECT  3.885000 196.010000  4.085000 196.210000 ;
        RECT  3.885000 196.415000  4.085000 196.615000 ;
        RECT  3.885000 196.820000  4.085000 197.020000 ;
        RECT  3.885000 197.225000  4.085000 197.425000 ;
        RECT  3.885000 197.630000  4.085000 197.830000 ;
        RECT  3.885000 198.035000  4.085000 198.235000 ;
        RECT  3.885000 198.440000  4.085000 198.640000 ;
        RECT  3.885000 198.845000  4.085000 199.045000 ;
        RECT  3.885000 199.250000  4.085000 199.450000 ;
        RECT  3.885000 199.655000  4.085000 199.855000 ;
        RECT  4.260000  25.910000  4.460000  26.110000 ;
        RECT  4.260000  26.340000  4.460000  26.540000 ;
        RECT  4.260000  26.770000  4.460000  26.970000 ;
        RECT  4.260000  27.200000  4.460000  27.400000 ;
        RECT  4.260000  27.630000  4.460000  27.830000 ;
        RECT  4.260000  28.060000  4.460000  28.260000 ;
        RECT  4.260000  28.490000  4.460000  28.690000 ;
        RECT  4.260000  28.920000  4.460000  29.120000 ;
        RECT  4.260000  29.350000  4.460000  29.550000 ;
        RECT  4.260000  29.780000  4.460000  29.980000 ;
        RECT  4.260000  30.210000  4.460000  30.410000 ;
        RECT  4.285000 175.995000  4.485000 176.195000 ;
        RECT  4.285000 176.395000  4.485000 176.595000 ;
        RECT  4.285000 176.795000  4.485000 176.995000 ;
        RECT  4.285000 177.195000  4.485000 177.395000 ;
        RECT  4.285000 177.595000  4.485000 177.795000 ;
        RECT  4.285000 177.995000  4.485000 178.195000 ;
        RECT  4.285000 178.395000  4.485000 178.595000 ;
        RECT  4.285000 178.795000  4.485000 178.995000 ;
        RECT  4.285000 179.195000  4.485000 179.395000 ;
        RECT  4.285000 179.595000  4.485000 179.795000 ;
        RECT  4.285000 179.995000  4.485000 180.195000 ;
        RECT  4.285000 180.395000  4.485000 180.595000 ;
        RECT  4.285000 180.795000  4.485000 180.995000 ;
        RECT  4.285000 181.195000  4.485000 181.395000 ;
        RECT  4.285000 181.595000  4.485000 181.795000 ;
        RECT  4.285000 181.995000  4.485000 182.195000 ;
        RECT  4.285000 182.395000  4.485000 182.595000 ;
        RECT  4.285000 182.795000  4.485000 182.995000 ;
        RECT  4.285000 183.195000  4.485000 183.395000 ;
        RECT  4.285000 183.595000  4.485000 183.795000 ;
        RECT  4.285000 183.995000  4.485000 184.195000 ;
        RECT  4.285000 184.395000  4.485000 184.595000 ;
        RECT  4.285000 184.795000  4.485000 184.995000 ;
        RECT  4.285000 185.195000  4.485000 185.395000 ;
        RECT  4.285000 185.595000  4.485000 185.795000 ;
        RECT  4.285000 185.995000  4.485000 186.195000 ;
        RECT  4.285000 186.395000  4.485000 186.595000 ;
        RECT  4.285000 186.795000  4.485000 186.995000 ;
        RECT  4.285000 187.195000  4.485000 187.395000 ;
        RECT  4.285000 187.595000  4.485000 187.795000 ;
        RECT  4.285000 187.995000  4.485000 188.195000 ;
        RECT  4.285000 188.395000  4.485000 188.595000 ;
        RECT  4.285000 188.795000  4.485000 188.995000 ;
        RECT  4.285000 189.195000  4.485000 189.395000 ;
        RECT  4.285000 189.595000  4.485000 189.795000 ;
        RECT  4.285000 189.995000  4.485000 190.195000 ;
        RECT  4.285000 190.395000  4.485000 190.595000 ;
        RECT  4.285000 190.795000  4.485000 190.995000 ;
        RECT  4.285000 191.195000  4.485000 191.395000 ;
        RECT  4.285000 191.595000  4.485000 191.795000 ;
        RECT  4.285000 191.995000  4.485000 192.195000 ;
        RECT  4.285000 192.395000  4.485000 192.595000 ;
        RECT  4.285000 192.795000  4.485000 192.995000 ;
        RECT  4.285000 193.195000  4.485000 193.395000 ;
        RECT  4.285000 193.595000  4.485000 193.795000 ;
        RECT  4.285000 193.995000  4.485000 194.195000 ;
        RECT  4.285000 194.395000  4.485000 194.595000 ;
        RECT  4.285000 194.795000  4.485000 194.995000 ;
        RECT  4.285000 195.200000  4.485000 195.400000 ;
        RECT  4.285000 195.605000  4.485000 195.805000 ;
        RECT  4.285000 196.010000  4.485000 196.210000 ;
        RECT  4.285000 196.415000  4.485000 196.615000 ;
        RECT  4.285000 196.820000  4.485000 197.020000 ;
        RECT  4.285000 197.225000  4.485000 197.425000 ;
        RECT  4.285000 197.630000  4.485000 197.830000 ;
        RECT  4.285000 198.035000  4.485000 198.235000 ;
        RECT  4.285000 198.440000  4.485000 198.640000 ;
        RECT  4.285000 198.845000  4.485000 199.045000 ;
        RECT  4.285000 199.250000  4.485000 199.450000 ;
        RECT  4.285000 199.655000  4.485000 199.855000 ;
        RECT  4.665000  25.910000  4.865000  26.110000 ;
        RECT  4.665000  26.340000  4.865000  26.540000 ;
        RECT  4.665000  26.770000  4.865000  26.970000 ;
        RECT  4.665000  27.200000  4.865000  27.400000 ;
        RECT  4.665000  27.630000  4.865000  27.830000 ;
        RECT  4.665000  28.060000  4.865000  28.260000 ;
        RECT  4.665000  28.490000  4.865000  28.690000 ;
        RECT  4.665000  28.920000  4.865000  29.120000 ;
        RECT  4.665000  29.350000  4.865000  29.550000 ;
        RECT  4.665000  29.780000  4.865000  29.980000 ;
        RECT  4.665000  30.210000  4.865000  30.410000 ;
        RECT  4.685000 175.995000  4.885000 176.195000 ;
        RECT  4.685000 176.395000  4.885000 176.595000 ;
        RECT  4.685000 176.795000  4.885000 176.995000 ;
        RECT  4.685000 177.195000  4.885000 177.395000 ;
        RECT  4.685000 177.595000  4.885000 177.795000 ;
        RECT  4.685000 177.995000  4.885000 178.195000 ;
        RECT  4.685000 178.395000  4.885000 178.595000 ;
        RECT  4.685000 178.795000  4.885000 178.995000 ;
        RECT  4.685000 179.195000  4.885000 179.395000 ;
        RECT  4.685000 179.595000  4.885000 179.795000 ;
        RECT  4.685000 179.995000  4.885000 180.195000 ;
        RECT  4.685000 180.395000  4.885000 180.595000 ;
        RECT  4.685000 180.795000  4.885000 180.995000 ;
        RECT  4.685000 181.195000  4.885000 181.395000 ;
        RECT  4.685000 181.595000  4.885000 181.795000 ;
        RECT  4.685000 181.995000  4.885000 182.195000 ;
        RECT  4.685000 182.395000  4.885000 182.595000 ;
        RECT  4.685000 182.795000  4.885000 182.995000 ;
        RECT  4.685000 183.195000  4.885000 183.395000 ;
        RECT  4.685000 183.595000  4.885000 183.795000 ;
        RECT  4.685000 183.995000  4.885000 184.195000 ;
        RECT  4.685000 184.395000  4.885000 184.595000 ;
        RECT  4.685000 184.795000  4.885000 184.995000 ;
        RECT  4.685000 185.195000  4.885000 185.395000 ;
        RECT  4.685000 185.595000  4.885000 185.795000 ;
        RECT  4.685000 185.995000  4.885000 186.195000 ;
        RECT  4.685000 186.395000  4.885000 186.595000 ;
        RECT  4.685000 186.795000  4.885000 186.995000 ;
        RECT  4.685000 187.195000  4.885000 187.395000 ;
        RECT  4.685000 187.595000  4.885000 187.795000 ;
        RECT  4.685000 187.995000  4.885000 188.195000 ;
        RECT  4.685000 188.395000  4.885000 188.595000 ;
        RECT  4.685000 188.795000  4.885000 188.995000 ;
        RECT  4.685000 189.195000  4.885000 189.395000 ;
        RECT  4.685000 189.595000  4.885000 189.795000 ;
        RECT  4.685000 189.995000  4.885000 190.195000 ;
        RECT  4.685000 190.395000  4.885000 190.595000 ;
        RECT  4.685000 190.795000  4.885000 190.995000 ;
        RECT  4.685000 191.195000  4.885000 191.395000 ;
        RECT  4.685000 191.595000  4.885000 191.795000 ;
        RECT  4.685000 191.995000  4.885000 192.195000 ;
        RECT  4.685000 192.395000  4.885000 192.595000 ;
        RECT  4.685000 192.795000  4.885000 192.995000 ;
        RECT  4.685000 193.195000  4.885000 193.395000 ;
        RECT  4.685000 193.595000  4.885000 193.795000 ;
        RECT  4.685000 193.995000  4.885000 194.195000 ;
        RECT  4.685000 194.395000  4.885000 194.595000 ;
        RECT  4.685000 194.795000  4.885000 194.995000 ;
        RECT  4.685000 195.200000  4.885000 195.400000 ;
        RECT  4.685000 195.605000  4.885000 195.805000 ;
        RECT  4.685000 196.010000  4.885000 196.210000 ;
        RECT  4.685000 196.415000  4.885000 196.615000 ;
        RECT  4.685000 196.820000  4.885000 197.020000 ;
        RECT  4.685000 197.225000  4.885000 197.425000 ;
        RECT  4.685000 197.630000  4.885000 197.830000 ;
        RECT  4.685000 198.035000  4.885000 198.235000 ;
        RECT  4.685000 198.440000  4.885000 198.640000 ;
        RECT  4.685000 198.845000  4.885000 199.045000 ;
        RECT  4.685000 199.250000  4.885000 199.450000 ;
        RECT  4.685000 199.655000  4.885000 199.855000 ;
        RECT  5.070000  25.910000  5.270000  26.110000 ;
        RECT  5.070000  26.340000  5.270000  26.540000 ;
        RECT  5.070000  26.770000  5.270000  26.970000 ;
        RECT  5.070000  27.200000  5.270000  27.400000 ;
        RECT  5.070000  27.630000  5.270000  27.830000 ;
        RECT  5.070000  28.060000  5.270000  28.260000 ;
        RECT  5.070000  28.490000  5.270000  28.690000 ;
        RECT  5.070000  28.920000  5.270000  29.120000 ;
        RECT  5.070000  29.350000  5.270000  29.550000 ;
        RECT  5.070000  29.780000  5.270000  29.980000 ;
        RECT  5.070000  30.210000  5.270000  30.410000 ;
        RECT  5.085000 175.995000  5.285000 176.195000 ;
        RECT  5.085000 176.395000  5.285000 176.595000 ;
        RECT  5.085000 176.795000  5.285000 176.995000 ;
        RECT  5.085000 177.195000  5.285000 177.395000 ;
        RECT  5.085000 177.595000  5.285000 177.795000 ;
        RECT  5.085000 177.995000  5.285000 178.195000 ;
        RECT  5.085000 178.395000  5.285000 178.595000 ;
        RECT  5.085000 178.795000  5.285000 178.995000 ;
        RECT  5.085000 179.195000  5.285000 179.395000 ;
        RECT  5.085000 179.595000  5.285000 179.795000 ;
        RECT  5.085000 179.995000  5.285000 180.195000 ;
        RECT  5.085000 180.395000  5.285000 180.595000 ;
        RECT  5.085000 180.795000  5.285000 180.995000 ;
        RECT  5.085000 181.195000  5.285000 181.395000 ;
        RECT  5.085000 181.595000  5.285000 181.795000 ;
        RECT  5.085000 181.995000  5.285000 182.195000 ;
        RECT  5.085000 182.395000  5.285000 182.595000 ;
        RECT  5.085000 182.795000  5.285000 182.995000 ;
        RECT  5.085000 183.195000  5.285000 183.395000 ;
        RECT  5.085000 183.595000  5.285000 183.795000 ;
        RECT  5.085000 183.995000  5.285000 184.195000 ;
        RECT  5.085000 184.395000  5.285000 184.595000 ;
        RECT  5.085000 184.795000  5.285000 184.995000 ;
        RECT  5.085000 185.195000  5.285000 185.395000 ;
        RECT  5.085000 185.595000  5.285000 185.795000 ;
        RECT  5.085000 185.995000  5.285000 186.195000 ;
        RECT  5.085000 186.395000  5.285000 186.595000 ;
        RECT  5.085000 186.795000  5.285000 186.995000 ;
        RECT  5.085000 187.195000  5.285000 187.395000 ;
        RECT  5.085000 187.595000  5.285000 187.795000 ;
        RECT  5.085000 187.995000  5.285000 188.195000 ;
        RECT  5.085000 188.395000  5.285000 188.595000 ;
        RECT  5.085000 188.795000  5.285000 188.995000 ;
        RECT  5.085000 189.195000  5.285000 189.395000 ;
        RECT  5.085000 189.595000  5.285000 189.795000 ;
        RECT  5.085000 189.995000  5.285000 190.195000 ;
        RECT  5.085000 190.395000  5.285000 190.595000 ;
        RECT  5.085000 190.795000  5.285000 190.995000 ;
        RECT  5.085000 191.195000  5.285000 191.395000 ;
        RECT  5.085000 191.595000  5.285000 191.795000 ;
        RECT  5.085000 191.995000  5.285000 192.195000 ;
        RECT  5.085000 192.395000  5.285000 192.595000 ;
        RECT  5.085000 192.795000  5.285000 192.995000 ;
        RECT  5.085000 193.195000  5.285000 193.395000 ;
        RECT  5.085000 193.595000  5.285000 193.795000 ;
        RECT  5.085000 193.995000  5.285000 194.195000 ;
        RECT  5.085000 194.395000  5.285000 194.595000 ;
        RECT  5.085000 194.795000  5.285000 194.995000 ;
        RECT  5.085000 195.200000  5.285000 195.400000 ;
        RECT  5.085000 195.605000  5.285000 195.805000 ;
        RECT  5.085000 196.010000  5.285000 196.210000 ;
        RECT  5.085000 196.415000  5.285000 196.615000 ;
        RECT  5.085000 196.820000  5.285000 197.020000 ;
        RECT  5.085000 197.225000  5.285000 197.425000 ;
        RECT  5.085000 197.630000  5.285000 197.830000 ;
        RECT  5.085000 198.035000  5.285000 198.235000 ;
        RECT  5.085000 198.440000  5.285000 198.640000 ;
        RECT  5.085000 198.845000  5.285000 199.045000 ;
        RECT  5.085000 199.250000  5.285000 199.450000 ;
        RECT  5.085000 199.655000  5.285000 199.855000 ;
        RECT  5.475000  25.910000  5.675000  26.110000 ;
        RECT  5.475000  26.340000  5.675000  26.540000 ;
        RECT  5.475000  26.770000  5.675000  26.970000 ;
        RECT  5.475000  27.200000  5.675000  27.400000 ;
        RECT  5.475000  27.630000  5.675000  27.830000 ;
        RECT  5.475000  28.060000  5.675000  28.260000 ;
        RECT  5.475000  28.490000  5.675000  28.690000 ;
        RECT  5.475000  28.920000  5.675000  29.120000 ;
        RECT  5.475000  29.350000  5.675000  29.550000 ;
        RECT  5.475000  29.780000  5.675000  29.980000 ;
        RECT  5.475000  30.210000  5.675000  30.410000 ;
        RECT  5.485000 175.995000  5.685000 176.195000 ;
        RECT  5.485000 176.395000  5.685000 176.595000 ;
        RECT  5.485000 176.795000  5.685000 176.995000 ;
        RECT  5.485000 177.195000  5.685000 177.395000 ;
        RECT  5.485000 177.595000  5.685000 177.795000 ;
        RECT  5.485000 177.995000  5.685000 178.195000 ;
        RECT  5.485000 178.395000  5.685000 178.595000 ;
        RECT  5.485000 178.795000  5.685000 178.995000 ;
        RECT  5.485000 179.195000  5.685000 179.395000 ;
        RECT  5.485000 179.595000  5.685000 179.795000 ;
        RECT  5.485000 179.995000  5.685000 180.195000 ;
        RECT  5.485000 180.395000  5.685000 180.595000 ;
        RECT  5.485000 180.795000  5.685000 180.995000 ;
        RECT  5.485000 181.195000  5.685000 181.395000 ;
        RECT  5.485000 181.595000  5.685000 181.795000 ;
        RECT  5.485000 181.995000  5.685000 182.195000 ;
        RECT  5.485000 182.395000  5.685000 182.595000 ;
        RECT  5.485000 182.795000  5.685000 182.995000 ;
        RECT  5.485000 183.195000  5.685000 183.395000 ;
        RECT  5.485000 183.595000  5.685000 183.795000 ;
        RECT  5.485000 183.995000  5.685000 184.195000 ;
        RECT  5.485000 184.395000  5.685000 184.595000 ;
        RECT  5.485000 184.795000  5.685000 184.995000 ;
        RECT  5.485000 185.195000  5.685000 185.395000 ;
        RECT  5.485000 185.595000  5.685000 185.795000 ;
        RECT  5.485000 185.995000  5.685000 186.195000 ;
        RECT  5.485000 186.395000  5.685000 186.595000 ;
        RECT  5.485000 186.795000  5.685000 186.995000 ;
        RECT  5.485000 187.195000  5.685000 187.395000 ;
        RECT  5.485000 187.595000  5.685000 187.795000 ;
        RECT  5.485000 187.995000  5.685000 188.195000 ;
        RECT  5.485000 188.395000  5.685000 188.595000 ;
        RECT  5.485000 188.795000  5.685000 188.995000 ;
        RECT  5.485000 189.195000  5.685000 189.395000 ;
        RECT  5.485000 189.595000  5.685000 189.795000 ;
        RECT  5.485000 189.995000  5.685000 190.195000 ;
        RECT  5.485000 190.395000  5.685000 190.595000 ;
        RECT  5.485000 190.795000  5.685000 190.995000 ;
        RECT  5.485000 191.195000  5.685000 191.395000 ;
        RECT  5.485000 191.595000  5.685000 191.795000 ;
        RECT  5.485000 191.995000  5.685000 192.195000 ;
        RECT  5.485000 192.395000  5.685000 192.595000 ;
        RECT  5.485000 192.795000  5.685000 192.995000 ;
        RECT  5.485000 193.195000  5.685000 193.395000 ;
        RECT  5.485000 193.595000  5.685000 193.795000 ;
        RECT  5.485000 193.995000  5.685000 194.195000 ;
        RECT  5.485000 194.395000  5.685000 194.595000 ;
        RECT  5.485000 194.795000  5.685000 194.995000 ;
        RECT  5.485000 195.200000  5.685000 195.400000 ;
        RECT  5.485000 195.605000  5.685000 195.805000 ;
        RECT  5.485000 196.010000  5.685000 196.210000 ;
        RECT  5.485000 196.415000  5.685000 196.615000 ;
        RECT  5.485000 196.820000  5.685000 197.020000 ;
        RECT  5.485000 197.225000  5.685000 197.425000 ;
        RECT  5.485000 197.630000  5.685000 197.830000 ;
        RECT  5.485000 198.035000  5.685000 198.235000 ;
        RECT  5.485000 198.440000  5.685000 198.640000 ;
        RECT  5.485000 198.845000  5.685000 199.045000 ;
        RECT  5.485000 199.250000  5.685000 199.450000 ;
        RECT  5.485000 199.655000  5.685000 199.855000 ;
        RECT  5.880000  25.910000  6.080000  26.110000 ;
        RECT  5.880000  26.340000  6.080000  26.540000 ;
        RECT  5.880000  26.770000  6.080000  26.970000 ;
        RECT  5.880000  27.200000  6.080000  27.400000 ;
        RECT  5.880000  27.630000  6.080000  27.830000 ;
        RECT  5.880000  28.060000  6.080000  28.260000 ;
        RECT  5.880000  28.490000  6.080000  28.690000 ;
        RECT  5.880000  28.920000  6.080000  29.120000 ;
        RECT  5.880000  29.350000  6.080000  29.550000 ;
        RECT  5.880000  29.780000  6.080000  29.980000 ;
        RECT  5.880000  30.210000  6.080000  30.410000 ;
        RECT  5.885000 175.995000  6.085000 176.195000 ;
        RECT  5.885000 176.395000  6.085000 176.595000 ;
        RECT  5.885000 176.795000  6.085000 176.995000 ;
        RECT  5.885000 177.195000  6.085000 177.395000 ;
        RECT  5.885000 177.595000  6.085000 177.795000 ;
        RECT  5.885000 177.995000  6.085000 178.195000 ;
        RECT  5.885000 178.395000  6.085000 178.595000 ;
        RECT  5.885000 178.795000  6.085000 178.995000 ;
        RECT  5.885000 179.195000  6.085000 179.395000 ;
        RECT  5.885000 179.595000  6.085000 179.795000 ;
        RECT  5.885000 179.995000  6.085000 180.195000 ;
        RECT  5.885000 180.395000  6.085000 180.595000 ;
        RECT  5.885000 180.795000  6.085000 180.995000 ;
        RECT  5.885000 181.195000  6.085000 181.395000 ;
        RECT  5.885000 181.595000  6.085000 181.795000 ;
        RECT  5.885000 181.995000  6.085000 182.195000 ;
        RECT  5.885000 182.395000  6.085000 182.595000 ;
        RECT  5.885000 182.795000  6.085000 182.995000 ;
        RECT  5.885000 183.195000  6.085000 183.395000 ;
        RECT  5.885000 183.595000  6.085000 183.795000 ;
        RECT  5.885000 183.995000  6.085000 184.195000 ;
        RECT  5.885000 184.395000  6.085000 184.595000 ;
        RECT  5.885000 184.795000  6.085000 184.995000 ;
        RECT  5.885000 185.195000  6.085000 185.395000 ;
        RECT  5.885000 185.595000  6.085000 185.795000 ;
        RECT  5.885000 185.995000  6.085000 186.195000 ;
        RECT  5.885000 186.395000  6.085000 186.595000 ;
        RECT  5.885000 186.795000  6.085000 186.995000 ;
        RECT  5.885000 187.195000  6.085000 187.395000 ;
        RECT  5.885000 187.595000  6.085000 187.795000 ;
        RECT  5.885000 187.995000  6.085000 188.195000 ;
        RECT  5.885000 188.395000  6.085000 188.595000 ;
        RECT  5.885000 188.795000  6.085000 188.995000 ;
        RECT  5.885000 189.195000  6.085000 189.395000 ;
        RECT  5.885000 189.595000  6.085000 189.795000 ;
        RECT  5.885000 189.995000  6.085000 190.195000 ;
        RECT  5.885000 190.395000  6.085000 190.595000 ;
        RECT  5.885000 190.795000  6.085000 190.995000 ;
        RECT  5.885000 191.195000  6.085000 191.395000 ;
        RECT  5.885000 191.595000  6.085000 191.795000 ;
        RECT  5.885000 191.995000  6.085000 192.195000 ;
        RECT  5.885000 192.395000  6.085000 192.595000 ;
        RECT  5.885000 192.795000  6.085000 192.995000 ;
        RECT  5.885000 193.195000  6.085000 193.395000 ;
        RECT  5.885000 193.595000  6.085000 193.795000 ;
        RECT  5.885000 193.995000  6.085000 194.195000 ;
        RECT  5.885000 194.395000  6.085000 194.595000 ;
        RECT  5.885000 194.795000  6.085000 194.995000 ;
        RECT  5.885000 195.200000  6.085000 195.400000 ;
        RECT  5.885000 195.605000  6.085000 195.805000 ;
        RECT  5.885000 196.010000  6.085000 196.210000 ;
        RECT  5.885000 196.415000  6.085000 196.615000 ;
        RECT  5.885000 196.820000  6.085000 197.020000 ;
        RECT  5.885000 197.225000  6.085000 197.425000 ;
        RECT  5.885000 197.630000  6.085000 197.830000 ;
        RECT  5.885000 198.035000  6.085000 198.235000 ;
        RECT  5.885000 198.440000  6.085000 198.640000 ;
        RECT  5.885000 198.845000  6.085000 199.045000 ;
        RECT  5.885000 199.250000  6.085000 199.450000 ;
        RECT  5.885000 199.655000  6.085000 199.855000 ;
        RECT  6.285000  25.910000  6.485000  26.110000 ;
        RECT  6.285000  26.340000  6.485000  26.540000 ;
        RECT  6.285000  26.770000  6.485000  26.970000 ;
        RECT  6.285000  27.200000  6.485000  27.400000 ;
        RECT  6.285000  27.630000  6.485000  27.830000 ;
        RECT  6.285000  28.060000  6.485000  28.260000 ;
        RECT  6.285000  28.490000  6.485000  28.690000 ;
        RECT  6.285000  28.920000  6.485000  29.120000 ;
        RECT  6.285000  29.350000  6.485000  29.550000 ;
        RECT  6.285000  29.780000  6.485000  29.980000 ;
        RECT  6.285000  30.210000  6.485000  30.410000 ;
        RECT  6.285000 175.995000  6.485000 176.195000 ;
        RECT  6.285000 176.395000  6.485000 176.595000 ;
        RECT  6.285000 176.795000  6.485000 176.995000 ;
        RECT  6.285000 177.195000  6.485000 177.395000 ;
        RECT  6.285000 177.595000  6.485000 177.795000 ;
        RECT  6.285000 177.995000  6.485000 178.195000 ;
        RECT  6.285000 178.395000  6.485000 178.595000 ;
        RECT  6.285000 178.795000  6.485000 178.995000 ;
        RECT  6.285000 179.195000  6.485000 179.395000 ;
        RECT  6.285000 179.595000  6.485000 179.795000 ;
        RECT  6.285000 179.995000  6.485000 180.195000 ;
        RECT  6.285000 180.395000  6.485000 180.595000 ;
        RECT  6.285000 180.795000  6.485000 180.995000 ;
        RECT  6.285000 181.195000  6.485000 181.395000 ;
        RECT  6.285000 181.595000  6.485000 181.795000 ;
        RECT  6.285000 181.995000  6.485000 182.195000 ;
        RECT  6.285000 182.395000  6.485000 182.595000 ;
        RECT  6.285000 182.795000  6.485000 182.995000 ;
        RECT  6.285000 183.195000  6.485000 183.395000 ;
        RECT  6.285000 183.595000  6.485000 183.795000 ;
        RECT  6.285000 183.995000  6.485000 184.195000 ;
        RECT  6.285000 184.395000  6.485000 184.595000 ;
        RECT  6.285000 184.795000  6.485000 184.995000 ;
        RECT  6.285000 185.195000  6.485000 185.395000 ;
        RECT  6.285000 185.595000  6.485000 185.795000 ;
        RECT  6.285000 185.995000  6.485000 186.195000 ;
        RECT  6.285000 186.395000  6.485000 186.595000 ;
        RECT  6.285000 186.795000  6.485000 186.995000 ;
        RECT  6.285000 187.195000  6.485000 187.395000 ;
        RECT  6.285000 187.595000  6.485000 187.795000 ;
        RECT  6.285000 187.995000  6.485000 188.195000 ;
        RECT  6.285000 188.395000  6.485000 188.595000 ;
        RECT  6.285000 188.795000  6.485000 188.995000 ;
        RECT  6.285000 189.195000  6.485000 189.395000 ;
        RECT  6.285000 189.595000  6.485000 189.795000 ;
        RECT  6.285000 189.995000  6.485000 190.195000 ;
        RECT  6.285000 190.395000  6.485000 190.595000 ;
        RECT  6.285000 190.795000  6.485000 190.995000 ;
        RECT  6.285000 191.195000  6.485000 191.395000 ;
        RECT  6.285000 191.595000  6.485000 191.795000 ;
        RECT  6.285000 191.995000  6.485000 192.195000 ;
        RECT  6.285000 192.395000  6.485000 192.595000 ;
        RECT  6.285000 192.795000  6.485000 192.995000 ;
        RECT  6.285000 193.195000  6.485000 193.395000 ;
        RECT  6.285000 193.595000  6.485000 193.795000 ;
        RECT  6.285000 193.995000  6.485000 194.195000 ;
        RECT  6.285000 194.395000  6.485000 194.595000 ;
        RECT  6.285000 194.795000  6.485000 194.995000 ;
        RECT  6.285000 195.200000  6.485000 195.400000 ;
        RECT  6.285000 195.605000  6.485000 195.805000 ;
        RECT  6.285000 196.010000  6.485000 196.210000 ;
        RECT  6.285000 196.415000  6.485000 196.615000 ;
        RECT  6.285000 196.820000  6.485000 197.020000 ;
        RECT  6.285000 197.225000  6.485000 197.425000 ;
        RECT  6.285000 197.630000  6.485000 197.830000 ;
        RECT  6.285000 198.035000  6.485000 198.235000 ;
        RECT  6.285000 198.440000  6.485000 198.640000 ;
        RECT  6.285000 198.845000  6.485000 199.045000 ;
        RECT  6.285000 199.250000  6.485000 199.450000 ;
        RECT  6.285000 199.655000  6.485000 199.855000 ;
        RECT  6.685000 175.995000  6.885000 176.195000 ;
        RECT  6.685000 176.395000  6.885000 176.595000 ;
        RECT  6.685000 176.795000  6.885000 176.995000 ;
        RECT  6.685000 177.195000  6.885000 177.395000 ;
        RECT  6.685000 177.595000  6.885000 177.795000 ;
        RECT  6.685000 177.995000  6.885000 178.195000 ;
        RECT  6.685000 178.395000  6.885000 178.595000 ;
        RECT  6.685000 178.795000  6.885000 178.995000 ;
        RECT  6.685000 179.195000  6.885000 179.395000 ;
        RECT  6.685000 179.595000  6.885000 179.795000 ;
        RECT  6.685000 179.995000  6.885000 180.195000 ;
        RECT  6.685000 180.395000  6.885000 180.595000 ;
        RECT  6.685000 180.795000  6.885000 180.995000 ;
        RECT  6.685000 181.195000  6.885000 181.395000 ;
        RECT  6.685000 181.595000  6.885000 181.795000 ;
        RECT  6.685000 181.995000  6.885000 182.195000 ;
        RECT  6.685000 182.395000  6.885000 182.595000 ;
        RECT  6.685000 182.795000  6.885000 182.995000 ;
        RECT  6.685000 183.195000  6.885000 183.395000 ;
        RECT  6.685000 183.595000  6.885000 183.795000 ;
        RECT  6.685000 183.995000  6.885000 184.195000 ;
        RECT  6.685000 184.395000  6.885000 184.595000 ;
        RECT  6.685000 184.795000  6.885000 184.995000 ;
        RECT  6.685000 185.195000  6.885000 185.395000 ;
        RECT  6.685000 185.595000  6.885000 185.795000 ;
        RECT  6.685000 185.995000  6.885000 186.195000 ;
        RECT  6.685000 186.395000  6.885000 186.595000 ;
        RECT  6.685000 186.795000  6.885000 186.995000 ;
        RECT  6.685000 187.195000  6.885000 187.395000 ;
        RECT  6.685000 187.595000  6.885000 187.795000 ;
        RECT  6.685000 187.995000  6.885000 188.195000 ;
        RECT  6.685000 188.395000  6.885000 188.595000 ;
        RECT  6.685000 188.795000  6.885000 188.995000 ;
        RECT  6.685000 189.195000  6.885000 189.395000 ;
        RECT  6.685000 189.595000  6.885000 189.795000 ;
        RECT  6.685000 189.995000  6.885000 190.195000 ;
        RECT  6.685000 190.395000  6.885000 190.595000 ;
        RECT  6.685000 190.795000  6.885000 190.995000 ;
        RECT  6.685000 191.195000  6.885000 191.395000 ;
        RECT  6.685000 191.595000  6.885000 191.795000 ;
        RECT  6.685000 191.995000  6.885000 192.195000 ;
        RECT  6.685000 192.395000  6.885000 192.595000 ;
        RECT  6.685000 192.795000  6.885000 192.995000 ;
        RECT  6.685000 193.195000  6.885000 193.395000 ;
        RECT  6.685000 193.595000  6.885000 193.795000 ;
        RECT  6.685000 193.995000  6.885000 194.195000 ;
        RECT  6.685000 194.395000  6.885000 194.595000 ;
        RECT  6.685000 194.795000  6.885000 194.995000 ;
        RECT  6.685000 195.200000  6.885000 195.400000 ;
        RECT  6.685000 195.605000  6.885000 195.805000 ;
        RECT  6.685000 196.010000  6.885000 196.210000 ;
        RECT  6.685000 196.415000  6.885000 196.615000 ;
        RECT  6.685000 196.820000  6.885000 197.020000 ;
        RECT  6.685000 197.225000  6.885000 197.425000 ;
        RECT  6.685000 197.630000  6.885000 197.830000 ;
        RECT  6.685000 198.035000  6.885000 198.235000 ;
        RECT  6.685000 198.440000  6.885000 198.640000 ;
        RECT  6.685000 198.845000  6.885000 199.045000 ;
        RECT  6.685000 199.250000  6.885000 199.450000 ;
        RECT  6.685000 199.655000  6.885000 199.855000 ;
        RECT  6.690000  25.910000  6.890000  26.110000 ;
        RECT  6.690000  26.340000  6.890000  26.540000 ;
        RECT  6.690000  26.770000  6.890000  26.970000 ;
        RECT  6.690000  27.200000  6.890000  27.400000 ;
        RECT  6.690000  27.630000  6.890000  27.830000 ;
        RECT  6.690000  28.060000  6.890000  28.260000 ;
        RECT  6.690000  28.490000  6.890000  28.690000 ;
        RECT  6.690000  28.920000  6.890000  29.120000 ;
        RECT  6.690000  29.350000  6.890000  29.550000 ;
        RECT  6.690000  29.780000  6.890000  29.980000 ;
        RECT  6.690000  30.210000  6.890000  30.410000 ;
        RECT  7.085000 175.995000  7.285000 176.195000 ;
        RECT  7.085000 176.395000  7.285000 176.595000 ;
        RECT  7.085000 176.795000  7.285000 176.995000 ;
        RECT  7.085000 177.195000  7.285000 177.395000 ;
        RECT  7.085000 177.595000  7.285000 177.795000 ;
        RECT  7.085000 177.995000  7.285000 178.195000 ;
        RECT  7.085000 178.395000  7.285000 178.595000 ;
        RECT  7.085000 178.795000  7.285000 178.995000 ;
        RECT  7.085000 179.195000  7.285000 179.395000 ;
        RECT  7.085000 179.595000  7.285000 179.795000 ;
        RECT  7.085000 179.995000  7.285000 180.195000 ;
        RECT  7.085000 180.395000  7.285000 180.595000 ;
        RECT  7.085000 180.795000  7.285000 180.995000 ;
        RECT  7.085000 181.195000  7.285000 181.395000 ;
        RECT  7.085000 181.595000  7.285000 181.795000 ;
        RECT  7.085000 181.995000  7.285000 182.195000 ;
        RECT  7.085000 182.395000  7.285000 182.595000 ;
        RECT  7.085000 182.795000  7.285000 182.995000 ;
        RECT  7.085000 183.195000  7.285000 183.395000 ;
        RECT  7.085000 183.595000  7.285000 183.795000 ;
        RECT  7.085000 183.995000  7.285000 184.195000 ;
        RECT  7.085000 184.395000  7.285000 184.595000 ;
        RECT  7.085000 184.795000  7.285000 184.995000 ;
        RECT  7.085000 185.195000  7.285000 185.395000 ;
        RECT  7.085000 185.595000  7.285000 185.795000 ;
        RECT  7.085000 185.995000  7.285000 186.195000 ;
        RECT  7.085000 186.395000  7.285000 186.595000 ;
        RECT  7.085000 186.795000  7.285000 186.995000 ;
        RECT  7.085000 187.195000  7.285000 187.395000 ;
        RECT  7.085000 187.595000  7.285000 187.795000 ;
        RECT  7.085000 187.995000  7.285000 188.195000 ;
        RECT  7.085000 188.395000  7.285000 188.595000 ;
        RECT  7.085000 188.795000  7.285000 188.995000 ;
        RECT  7.085000 189.195000  7.285000 189.395000 ;
        RECT  7.085000 189.595000  7.285000 189.795000 ;
        RECT  7.085000 189.995000  7.285000 190.195000 ;
        RECT  7.085000 190.395000  7.285000 190.595000 ;
        RECT  7.085000 190.795000  7.285000 190.995000 ;
        RECT  7.085000 191.195000  7.285000 191.395000 ;
        RECT  7.085000 191.595000  7.285000 191.795000 ;
        RECT  7.085000 191.995000  7.285000 192.195000 ;
        RECT  7.085000 192.395000  7.285000 192.595000 ;
        RECT  7.085000 192.795000  7.285000 192.995000 ;
        RECT  7.085000 193.195000  7.285000 193.395000 ;
        RECT  7.085000 193.595000  7.285000 193.795000 ;
        RECT  7.085000 193.995000  7.285000 194.195000 ;
        RECT  7.085000 194.395000  7.285000 194.595000 ;
        RECT  7.085000 194.795000  7.285000 194.995000 ;
        RECT  7.085000 195.200000  7.285000 195.400000 ;
        RECT  7.085000 195.605000  7.285000 195.805000 ;
        RECT  7.085000 196.010000  7.285000 196.210000 ;
        RECT  7.085000 196.415000  7.285000 196.615000 ;
        RECT  7.085000 196.820000  7.285000 197.020000 ;
        RECT  7.085000 197.225000  7.285000 197.425000 ;
        RECT  7.085000 197.630000  7.285000 197.830000 ;
        RECT  7.085000 198.035000  7.285000 198.235000 ;
        RECT  7.085000 198.440000  7.285000 198.640000 ;
        RECT  7.085000 198.845000  7.285000 199.045000 ;
        RECT  7.085000 199.250000  7.285000 199.450000 ;
        RECT  7.085000 199.655000  7.285000 199.855000 ;
        RECT  7.095000  25.910000  7.295000  26.110000 ;
        RECT  7.095000  26.340000  7.295000  26.540000 ;
        RECT  7.095000  26.770000  7.295000  26.970000 ;
        RECT  7.095000  27.200000  7.295000  27.400000 ;
        RECT  7.095000  27.630000  7.295000  27.830000 ;
        RECT  7.095000  28.060000  7.295000  28.260000 ;
        RECT  7.095000  28.490000  7.295000  28.690000 ;
        RECT  7.095000  28.920000  7.295000  29.120000 ;
        RECT  7.095000  29.350000  7.295000  29.550000 ;
        RECT  7.095000  29.780000  7.295000  29.980000 ;
        RECT  7.095000  30.210000  7.295000  30.410000 ;
        RECT  7.485000 175.995000  7.685000 176.195000 ;
        RECT  7.485000 176.395000  7.685000 176.595000 ;
        RECT  7.485000 176.795000  7.685000 176.995000 ;
        RECT  7.485000 177.195000  7.685000 177.395000 ;
        RECT  7.485000 177.595000  7.685000 177.795000 ;
        RECT  7.485000 177.995000  7.685000 178.195000 ;
        RECT  7.485000 178.395000  7.685000 178.595000 ;
        RECT  7.485000 178.795000  7.685000 178.995000 ;
        RECT  7.485000 179.195000  7.685000 179.395000 ;
        RECT  7.485000 179.595000  7.685000 179.795000 ;
        RECT  7.485000 179.995000  7.685000 180.195000 ;
        RECT  7.485000 180.395000  7.685000 180.595000 ;
        RECT  7.485000 180.795000  7.685000 180.995000 ;
        RECT  7.485000 181.195000  7.685000 181.395000 ;
        RECT  7.485000 181.595000  7.685000 181.795000 ;
        RECT  7.485000 181.995000  7.685000 182.195000 ;
        RECT  7.485000 182.395000  7.685000 182.595000 ;
        RECT  7.485000 182.795000  7.685000 182.995000 ;
        RECT  7.485000 183.195000  7.685000 183.395000 ;
        RECT  7.485000 183.595000  7.685000 183.795000 ;
        RECT  7.485000 183.995000  7.685000 184.195000 ;
        RECT  7.485000 184.395000  7.685000 184.595000 ;
        RECT  7.485000 184.795000  7.685000 184.995000 ;
        RECT  7.485000 185.195000  7.685000 185.395000 ;
        RECT  7.485000 185.595000  7.685000 185.795000 ;
        RECT  7.485000 185.995000  7.685000 186.195000 ;
        RECT  7.485000 186.395000  7.685000 186.595000 ;
        RECT  7.485000 186.795000  7.685000 186.995000 ;
        RECT  7.485000 187.195000  7.685000 187.395000 ;
        RECT  7.485000 187.595000  7.685000 187.795000 ;
        RECT  7.485000 187.995000  7.685000 188.195000 ;
        RECT  7.485000 188.395000  7.685000 188.595000 ;
        RECT  7.485000 188.795000  7.685000 188.995000 ;
        RECT  7.485000 189.195000  7.685000 189.395000 ;
        RECT  7.485000 189.595000  7.685000 189.795000 ;
        RECT  7.485000 189.995000  7.685000 190.195000 ;
        RECT  7.485000 190.395000  7.685000 190.595000 ;
        RECT  7.485000 190.795000  7.685000 190.995000 ;
        RECT  7.485000 191.195000  7.685000 191.395000 ;
        RECT  7.485000 191.595000  7.685000 191.795000 ;
        RECT  7.485000 191.995000  7.685000 192.195000 ;
        RECT  7.485000 192.395000  7.685000 192.595000 ;
        RECT  7.485000 192.795000  7.685000 192.995000 ;
        RECT  7.485000 193.195000  7.685000 193.395000 ;
        RECT  7.485000 193.595000  7.685000 193.795000 ;
        RECT  7.485000 193.995000  7.685000 194.195000 ;
        RECT  7.485000 194.395000  7.685000 194.595000 ;
        RECT  7.485000 194.795000  7.685000 194.995000 ;
        RECT  7.485000 195.200000  7.685000 195.400000 ;
        RECT  7.485000 195.605000  7.685000 195.805000 ;
        RECT  7.485000 196.010000  7.685000 196.210000 ;
        RECT  7.485000 196.415000  7.685000 196.615000 ;
        RECT  7.485000 196.820000  7.685000 197.020000 ;
        RECT  7.485000 197.225000  7.685000 197.425000 ;
        RECT  7.485000 197.630000  7.685000 197.830000 ;
        RECT  7.485000 198.035000  7.685000 198.235000 ;
        RECT  7.485000 198.440000  7.685000 198.640000 ;
        RECT  7.485000 198.845000  7.685000 199.045000 ;
        RECT  7.485000 199.250000  7.685000 199.450000 ;
        RECT  7.485000 199.655000  7.685000 199.855000 ;
        RECT  7.500000  25.910000  7.700000  26.110000 ;
        RECT  7.500000  26.340000  7.700000  26.540000 ;
        RECT  7.500000  26.770000  7.700000  26.970000 ;
        RECT  7.500000  27.200000  7.700000  27.400000 ;
        RECT  7.500000  27.630000  7.700000  27.830000 ;
        RECT  7.500000  28.060000  7.700000  28.260000 ;
        RECT  7.500000  28.490000  7.700000  28.690000 ;
        RECT  7.500000  28.920000  7.700000  29.120000 ;
        RECT  7.500000  29.350000  7.700000  29.550000 ;
        RECT  7.500000  29.780000  7.700000  29.980000 ;
        RECT  7.500000  30.210000  7.700000  30.410000 ;
        RECT  7.885000 175.995000  8.085000 176.195000 ;
        RECT  7.885000 176.395000  8.085000 176.595000 ;
        RECT  7.885000 176.795000  8.085000 176.995000 ;
        RECT  7.885000 177.195000  8.085000 177.395000 ;
        RECT  7.885000 177.595000  8.085000 177.795000 ;
        RECT  7.885000 177.995000  8.085000 178.195000 ;
        RECT  7.885000 178.395000  8.085000 178.595000 ;
        RECT  7.885000 178.795000  8.085000 178.995000 ;
        RECT  7.885000 179.195000  8.085000 179.395000 ;
        RECT  7.885000 179.595000  8.085000 179.795000 ;
        RECT  7.885000 179.995000  8.085000 180.195000 ;
        RECT  7.885000 180.395000  8.085000 180.595000 ;
        RECT  7.885000 180.795000  8.085000 180.995000 ;
        RECT  7.885000 181.195000  8.085000 181.395000 ;
        RECT  7.885000 181.595000  8.085000 181.795000 ;
        RECT  7.885000 181.995000  8.085000 182.195000 ;
        RECT  7.885000 182.395000  8.085000 182.595000 ;
        RECT  7.885000 182.795000  8.085000 182.995000 ;
        RECT  7.885000 183.195000  8.085000 183.395000 ;
        RECT  7.885000 183.595000  8.085000 183.795000 ;
        RECT  7.885000 183.995000  8.085000 184.195000 ;
        RECT  7.885000 184.395000  8.085000 184.595000 ;
        RECT  7.885000 184.795000  8.085000 184.995000 ;
        RECT  7.885000 185.195000  8.085000 185.395000 ;
        RECT  7.885000 185.595000  8.085000 185.795000 ;
        RECT  7.885000 185.995000  8.085000 186.195000 ;
        RECT  7.885000 186.395000  8.085000 186.595000 ;
        RECT  7.885000 186.795000  8.085000 186.995000 ;
        RECT  7.885000 187.195000  8.085000 187.395000 ;
        RECT  7.885000 187.595000  8.085000 187.795000 ;
        RECT  7.885000 187.995000  8.085000 188.195000 ;
        RECT  7.885000 188.395000  8.085000 188.595000 ;
        RECT  7.885000 188.795000  8.085000 188.995000 ;
        RECT  7.885000 189.195000  8.085000 189.395000 ;
        RECT  7.885000 189.595000  8.085000 189.795000 ;
        RECT  7.885000 189.995000  8.085000 190.195000 ;
        RECT  7.885000 190.395000  8.085000 190.595000 ;
        RECT  7.885000 190.795000  8.085000 190.995000 ;
        RECT  7.885000 191.195000  8.085000 191.395000 ;
        RECT  7.885000 191.595000  8.085000 191.795000 ;
        RECT  7.885000 191.995000  8.085000 192.195000 ;
        RECT  7.885000 192.395000  8.085000 192.595000 ;
        RECT  7.885000 192.795000  8.085000 192.995000 ;
        RECT  7.885000 193.195000  8.085000 193.395000 ;
        RECT  7.885000 193.595000  8.085000 193.795000 ;
        RECT  7.885000 193.995000  8.085000 194.195000 ;
        RECT  7.885000 194.395000  8.085000 194.595000 ;
        RECT  7.885000 194.795000  8.085000 194.995000 ;
        RECT  7.885000 195.200000  8.085000 195.400000 ;
        RECT  7.885000 195.605000  8.085000 195.805000 ;
        RECT  7.885000 196.010000  8.085000 196.210000 ;
        RECT  7.885000 196.415000  8.085000 196.615000 ;
        RECT  7.885000 196.820000  8.085000 197.020000 ;
        RECT  7.885000 197.225000  8.085000 197.425000 ;
        RECT  7.885000 197.630000  8.085000 197.830000 ;
        RECT  7.885000 198.035000  8.085000 198.235000 ;
        RECT  7.885000 198.440000  8.085000 198.640000 ;
        RECT  7.885000 198.845000  8.085000 199.045000 ;
        RECT  7.885000 199.250000  8.085000 199.450000 ;
        RECT  7.885000 199.655000  8.085000 199.855000 ;
        RECT  7.905000  25.910000  8.105000  26.110000 ;
        RECT  7.905000  26.340000  8.105000  26.540000 ;
        RECT  7.905000  26.770000  8.105000  26.970000 ;
        RECT  7.905000  27.200000  8.105000  27.400000 ;
        RECT  7.905000  27.630000  8.105000  27.830000 ;
        RECT  7.905000  28.060000  8.105000  28.260000 ;
        RECT  7.905000  28.490000  8.105000  28.690000 ;
        RECT  7.905000  28.920000  8.105000  29.120000 ;
        RECT  7.905000  29.350000  8.105000  29.550000 ;
        RECT  7.905000  29.780000  8.105000  29.980000 ;
        RECT  7.905000  30.210000  8.105000  30.410000 ;
        RECT  8.285000 175.995000  8.485000 176.195000 ;
        RECT  8.285000 176.395000  8.485000 176.595000 ;
        RECT  8.285000 176.795000  8.485000 176.995000 ;
        RECT  8.285000 177.195000  8.485000 177.395000 ;
        RECT  8.285000 177.595000  8.485000 177.795000 ;
        RECT  8.285000 177.995000  8.485000 178.195000 ;
        RECT  8.285000 178.395000  8.485000 178.595000 ;
        RECT  8.285000 178.795000  8.485000 178.995000 ;
        RECT  8.285000 179.195000  8.485000 179.395000 ;
        RECT  8.285000 179.595000  8.485000 179.795000 ;
        RECT  8.285000 179.995000  8.485000 180.195000 ;
        RECT  8.285000 180.395000  8.485000 180.595000 ;
        RECT  8.285000 180.795000  8.485000 180.995000 ;
        RECT  8.285000 181.195000  8.485000 181.395000 ;
        RECT  8.285000 181.595000  8.485000 181.795000 ;
        RECT  8.285000 181.995000  8.485000 182.195000 ;
        RECT  8.285000 182.395000  8.485000 182.595000 ;
        RECT  8.285000 182.795000  8.485000 182.995000 ;
        RECT  8.285000 183.195000  8.485000 183.395000 ;
        RECT  8.285000 183.595000  8.485000 183.795000 ;
        RECT  8.285000 183.995000  8.485000 184.195000 ;
        RECT  8.285000 184.395000  8.485000 184.595000 ;
        RECT  8.285000 184.795000  8.485000 184.995000 ;
        RECT  8.285000 185.195000  8.485000 185.395000 ;
        RECT  8.285000 185.595000  8.485000 185.795000 ;
        RECT  8.285000 185.995000  8.485000 186.195000 ;
        RECT  8.285000 186.395000  8.485000 186.595000 ;
        RECT  8.285000 186.795000  8.485000 186.995000 ;
        RECT  8.285000 187.195000  8.485000 187.395000 ;
        RECT  8.285000 187.595000  8.485000 187.795000 ;
        RECT  8.285000 187.995000  8.485000 188.195000 ;
        RECT  8.285000 188.395000  8.485000 188.595000 ;
        RECT  8.285000 188.795000  8.485000 188.995000 ;
        RECT  8.285000 189.195000  8.485000 189.395000 ;
        RECT  8.285000 189.595000  8.485000 189.795000 ;
        RECT  8.285000 189.995000  8.485000 190.195000 ;
        RECT  8.285000 190.395000  8.485000 190.595000 ;
        RECT  8.285000 190.795000  8.485000 190.995000 ;
        RECT  8.285000 191.195000  8.485000 191.395000 ;
        RECT  8.285000 191.595000  8.485000 191.795000 ;
        RECT  8.285000 191.995000  8.485000 192.195000 ;
        RECT  8.285000 192.395000  8.485000 192.595000 ;
        RECT  8.285000 192.795000  8.485000 192.995000 ;
        RECT  8.285000 193.195000  8.485000 193.395000 ;
        RECT  8.285000 193.595000  8.485000 193.795000 ;
        RECT  8.285000 193.995000  8.485000 194.195000 ;
        RECT  8.285000 194.395000  8.485000 194.595000 ;
        RECT  8.285000 194.795000  8.485000 194.995000 ;
        RECT  8.285000 195.200000  8.485000 195.400000 ;
        RECT  8.285000 195.605000  8.485000 195.805000 ;
        RECT  8.285000 196.010000  8.485000 196.210000 ;
        RECT  8.285000 196.415000  8.485000 196.615000 ;
        RECT  8.285000 196.820000  8.485000 197.020000 ;
        RECT  8.285000 197.225000  8.485000 197.425000 ;
        RECT  8.285000 197.630000  8.485000 197.830000 ;
        RECT  8.285000 198.035000  8.485000 198.235000 ;
        RECT  8.285000 198.440000  8.485000 198.640000 ;
        RECT  8.285000 198.845000  8.485000 199.045000 ;
        RECT  8.285000 199.250000  8.485000 199.450000 ;
        RECT  8.285000 199.655000  8.485000 199.855000 ;
        RECT  8.310000  25.910000  8.510000  26.110000 ;
        RECT  8.310000  26.340000  8.510000  26.540000 ;
        RECT  8.310000  26.770000  8.510000  26.970000 ;
        RECT  8.310000  27.200000  8.510000  27.400000 ;
        RECT  8.310000  27.630000  8.510000  27.830000 ;
        RECT  8.310000  28.060000  8.510000  28.260000 ;
        RECT  8.310000  28.490000  8.510000  28.690000 ;
        RECT  8.310000  28.920000  8.510000  29.120000 ;
        RECT  8.310000  29.350000  8.510000  29.550000 ;
        RECT  8.310000  29.780000  8.510000  29.980000 ;
        RECT  8.310000  30.210000  8.510000  30.410000 ;
        RECT  8.685000 175.995000  8.885000 176.195000 ;
        RECT  8.685000 176.395000  8.885000 176.595000 ;
        RECT  8.685000 176.795000  8.885000 176.995000 ;
        RECT  8.685000 177.195000  8.885000 177.395000 ;
        RECT  8.685000 177.595000  8.885000 177.795000 ;
        RECT  8.685000 177.995000  8.885000 178.195000 ;
        RECT  8.685000 178.395000  8.885000 178.595000 ;
        RECT  8.685000 178.795000  8.885000 178.995000 ;
        RECT  8.685000 179.195000  8.885000 179.395000 ;
        RECT  8.685000 179.595000  8.885000 179.795000 ;
        RECT  8.685000 179.995000  8.885000 180.195000 ;
        RECT  8.685000 180.395000  8.885000 180.595000 ;
        RECT  8.685000 180.795000  8.885000 180.995000 ;
        RECT  8.685000 181.195000  8.885000 181.395000 ;
        RECT  8.685000 181.595000  8.885000 181.795000 ;
        RECT  8.685000 181.995000  8.885000 182.195000 ;
        RECT  8.685000 182.395000  8.885000 182.595000 ;
        RECT  8.685000 182.795000  8.885000 182.995000 ;
        RECT  8.685000 183.195000  8.885000 183.395000 ;
        RECT  8.685000 183.595000  8.885000 183.795000 ;
        RECT  8.685000 183.995000  8.885000 184.195000 ;
        RECT  8.685000 184.395000  8.885000 184.595000 ;
        RECT  8.685000 184.795000  8.885000 184.995000 ;
        RECT  8.685000 185.195000  8.885000 185.395000 ;
        RECT  8.685000 185.595000  8.885000 185.795000 ;
        RECT  8.685000 185.995000  8.885000 186.195000 ;
        RECT  8.685000 186.395000  8.885000 186.595000 ;
        RECT  8.685000 186.795000  8.885000 186.995000 ;
        RECT  8.685000 187.195000  8.885000 187.395000 ;
        RECT  8.685000 187.595000  8.885000 187.795000 ;
        RECT  8.685000 187.995000  8.885000 188.195000 ;
        RECT  8.685000 188.395000  8.885000 188.595000 ;
        RECT  8.685000 188.795000  8.885000 188.995000 ;
        RECT  8.685000 189.195000  8.885000 189.395000 ;
        RECT  8.685000 189.595000  8.885000 189.795000 ;
        RECT  8.685000 189.995000  8.885000 190.195000 ;
        RECT  8.685000 190.395000  8.885000 190.595000 ;
        RECT  8.685000 190.795000  8.885000 190.995000 ;
        RECT  8.685000 191.195000  8.885000 191.395000 ;
        RECT  8.685000 191.595000  8.885000 191.795000 ;
        RECT  8.685000 191.995000  8.885000 192.195000 ;
        RECT  8.685000 192.395000  8.885000 192.595000 ;
        RECT  8.685000 192.795000  8.885000 192.995000 ;
        RECT  8.685000 193.195000  8.885000 193.395000 ;
        RECT  8.685000 193.595000  8.885000 193.795000 ;
        RECT  8.685000 193.995000  8.885000 194.195000 ;
        RECT  8.685000 194.395000  8.885000 194.595000 ;
        RECT  8.685000 194.795000  8.885000 194.995000 ;
        RECT  8.685000 195.200000  8.885000 195.400000 ;
        RECT  8.685000 195.605000  8.885000 195.805000 ;
        RECT  8.685000 196.010000  8.885000 196.210000 ;
        RECT  8.685000 196.415000  8.885000 196.615000 ;
        RECT  8.685000 196.820000  8.885000 197.020000 ;
        RECT  8.685000 197.225000  8.885000 197.425000 ;
        RECT  8.685000 197.630000  8.885000 197.830000 ;
        RECT  8.685000 198.035000  8.885000 198.235000 ;
        RECT  8.685000 198.440000  8.885000 198.640000 ;
        RECT  8.685000 198.845000  8.885000 199.045000 ;
        RECT  8.685000 199.250000  8.885000 199.450000 ;
        RECT  8.685000 199.655000  8.885000 199.855000 ;
        RECT  8.715000  25.910000  8.915000  26.110000 ;
        RECT  8.715000  26.340000  8.915000  26.540000 ;
        RECT  8.715000  26.770000  8.915000  26.970000 ;
        RECT  8.715000  27.200000  8.915000  27.400000 ;
        RECT  8.715000  27.630000  8.915000  27.830000 ;
        RECT  8.715000  28.060000  8.915000  28.260000 ;
        RECT  8.715000  28.490000  8.915000  28.690000 ;
        RECT  8.715000  28.920000  8.915000  29.120000 ;
        RECT  8.715000  29.350000  8.915000  29.550000 ;
        RECT  8.715000  29.780000  8.915000  29.980000 ;
        RECT  8.715000  30.210000  8.915000  30.410000 ;
        RECT  9.085000 175.995000  9.285000 176.195000 ;
        RECT  9.085000 176.395000  9.285000 176.595000 ;
        RECT  9.085000 176.795000  9.285000 176.995000 ;
        RECT  9.085000 177.195000  9.285000 177.395000 ;
        RECT  9.085000 177.595000  9.285000 177.795000 ;
        RECT  9.085000 177.995000  9.285000 178.195000 ;
        RECT  9.085000 178.395000  9.285000 178.595000 ;
        RECT  9.085000 178.795000  9.285000 178.995000 ;
        RECT  9.085000 179.195000  9.285000 179.395000 ;
        RECT  9.085000 179.595000  9.285000 179.795000 ;
        RECT  9.085000 179.995000  9.285000 180.195000 ;
        RECT  9.085000 180.395000  9.285000 180.595000 ;
        RECT  9.085000 180.795000  9.285000 180.995000 ;
        RECT  9.085000 181.195000  9.285000 181.395000 ;
        RECT  9.085000 181.595000  9.285000 181.795000 ;
        RECT  9.085000 181.995000  9.285000 182.195000 ;
        RECT  9.085000 182.395000  9.285000 182.595000 ;
        RECT  9.085000 182.795000  9.285000 182.995000 ;
        RECT  9.085000 183.195000  9.285000 183.395000 ;
        RECT  9.085000 183.595000  9.285000 183.795000 ;
        RECT  9.085000 183.995000  9.285000 184.195000 ;
        RECT  9.085000 184.395000  9.285000 184.595000 ;
        RECT  9.085000 184.795000  9.285000 184.995000 ;
        RECT  9.085000 185.195000  9.285000 185.395000 ;
        RECT  9.085000 185.595000  9.285000 185.795000 ;
        RECT  9.085000 185.995000  9.285000 186.195000 ;
        RECT  9.085000 186.395000  9.285000 186.595000 ;
        RECT  9.085000 186.795000  9.285000 186.995000 ;
        RECT  9.085000 187.195000  9.285000 187.395000 ;
        RECT  9.085000 187.595000  9.285000 187.795000 ;
        RECT  9.085000 187.995000  9.285000 188.195000 ;
        RECT  9.085000 188.395000  9.285000 188.595000 ;
        RECT  9.085000 188.795000  9.285000 188.995000 ;
        RECT  9.085000 189.195000  9.285000 189.395000 ;
        RECT  9.085000 189.595000  9.285000 189.795000 ;
        RECT  9.085000 189.995000  9.285000 190.195000 ;
        RECT  9.085000 190.395000  9.285000 190.595000 ;
        RECT  9.085000 190.795000  9.285000 190.995000 ;
        RECT  9.085000 191.195000  9.285000 191.395000 ;
        RECT  9.085000 191.595000  9.285000 191.795000 ;
        RECT  9.085000 191.995000  9.285000 192.195000 ;
        RECT  9.085000 192.395000  9.285000 192.595000 ;
        RECT  9.085000 192.795000  9.285000 192.995000 ;
        RECT  9.085000 193.195000  9.285000 193.395000 ;
        RECT  9.085000 193.595000  9.285000 193.795000 ;
        RECT  9.085000 193.995000  9.285000 194.195000 ;
        RECT  9.085000 194.395000  9.285000 194.595000 ;
        RECT  9.085000 194.795000  9.285000 194.995000 ;
        RECT  9.085000 195.200000  9.285000 195.400000 ;
        RECT  9.085000 195.605000  9.285000 195.805000 ;
        RECT  9.085000 196.010000  9.285000 196.210000 ;
        RECT  9.085000 196.415000  9.285000 196.615000 ;
        RECT  9.085000 196.820000  9.285000 197.020000 ;
        RECT  9.085000 197.225000  9.285000 197.425000 ;
        RECT  9.085000 197.630000  9.285000 197.830000 ;
        RECT  9.085000 198.035000  9.285000 198.235000 ;
        RECT  9.085000 198.440000  9.285000 198.640000 ;
        RECT  9.085000 198.845000  9.285000 199.045000 ;
        RECT  9.085000 199.250000  9.285000 199.450000 ;
        RECT  9.085000 199.655000  9.285000 199.855000 ;
        RECT  9.120000  25.910000  9.320000  26.110000 ;
        RECT  9.120000  26.340000  9.320000  26.540000 ;
        RECT  9.120000  26.770000  9.320000  26.970000 ;
        RECT  9.120000  27.200000  9.320000  27.400000 ;
        RECT  9.120000  27.630000  9.320000  27.830000 ;
        RECT  9.120000  28.060000  9.320000  28.260000 ;
        RECT  9.120000  28.490000  9.320000  28.690000 ;
        RECT  9.120000  28.920000  9.320000  29.120000 ;
        RECT  9.120000  29.350000  9.320000  29.550000 ;
        RECT  9.120000  29.780000  9.320000  29.980000 ;
        RECT  9.120000  30.210000  9.320000  30.410000 ;
        RECT  9.485000 175.995000  9.685000 176.195000 ;
        RECT  9.485000 176.395000  9.685000 176.595000 ;
        RECT  9.485000 176.795000  9.685000 176.995000 ;
        RECT  9.485000 177.195000  9.685000 177.395000 ;
        RECT  9.485000 177.595000  9.685000 177.795000 ;
        RECT  9.485000 177.995000  9.685000 178.195000 ;
        RECT  9.485000 178.395000  9.685000 178.595000 ;
        RECT  9.485000 178.795000  9.685000 178.995000 ;
        RECT  9.485000 179.195000  9.685000 179.395000 ;
        RECT  9.485000 179.595000  9.685000 179.795000 ;
        RECT  9.485000 179.995000  9.685000 180.195000 ;
        RECT  9.485000 180.395000  9.685000 180.595000 ;
        RECT  9.485000 180.795000  9.685000 180.995000 ;
        RECT  9.485000 181.195000  9.685000 181.395000 ;
        RECT  9.485000 181.595000  9.685000 181.795000 ;
        RECT  9.485000 181.995000  9.685000 182.195000 ;
        RECT  9.485000 182.395000  9.685000 182.595000 ;
        RECT  9.485000 182.795000  9.685000 182.995000 ;
        RECT  9.485000 183.195000  9.685000 183.395000 ;
        RECT  9.485000 183.595000  9.685000 183.795000 ;
        RECT  9.485000 183.995000  9.685000 184.195000 ;
        RECT  9.485000 184.395000  9.685000 184.595000 ;
        RECT  9.485000 184.795000  9.685000 184.995000 ;
        RECT  9.485000 185.195000  9.685000 185.395000 ;
        RECT  9.485000 185.595000  9.685000 185.795000 ;
        RECT  9.485000 185.995000  9.685000 186.195000 ;
        RECT  9.485000 186.395000  9.685000 186.595000 ;
        RECT  9.485000 186.795000  9.685000 186.995000 ;
        RECT  9.485000 187.195000  9.685000 187.395000 ;
        RECT  9.485000 187.595000  9.685000 187.795000 ;
        RECT  9.485000 187.995000  9.685000 188.195000 ;
        RECT  9.485000 188.395000  9.685000 188.595000 ;
        RECT  9.485000 188.795000  9.685000 188.995000 ;
        RECT  9.485000 189.195000  9.685000 189.395000 ;
        RECT  9.485000 189.595000  9.685000 189.795000 ;
        RECT  9.485000 189.995000  9.685000 190.195000 ;
        RECT  9.485000 190.395000  9.685000 190.595000 ;
        RECT  9.485000 190.795000  9.685000 190.995000 ;
        RECT  9.485000 191.195000  9.685000 191.395000 ;
        RECT  9.485000 191.595000  9.685000 191.795000 ;
        RECT  9.485000 191.995000  9.685000 192.195000 ;
        RECT  9.485000 192.395000  9.685000 192.595000 ;
        RECT  9.485000 192.795000  9.685000 192.995000 ;
        RECT  9.485000 193.195000  9.685000 193.395000 ;
        RECT  9.485000 193.595000  9.685000 193.795000 ;
        RECT  9.485000 193.995000  9.685000 194.195000 ;
        RECT  9.485000 194.395000  9.685000 194.595000 ;
        RECT  9.485000 194.795000  9.685000 194.995000 ;
        RECT  9.485000 195.200000  9.685000 195.400000 ;
        RECT  9.485000 195.605000  9.685000 195.805000 ;
        RECT  9.485000 196.010000  9.685000 196.210000 ;
        RECT  9.485000 196.415000  9.685000 196.615000 ;
        RECT  9.485000 196.820000  9.685000 197.020000 ;
        RECT  9.485000 197.225000  9.685000 197.425000 ;
        RECT  9.485000 197.630000  9.685000 197.830000 ;
        RECT  9.485000 198.035000  9.685000 198.235000 ;
        RECT  9.485000 198.440000  9.685000 198.640000 ;
        RECT  9.485000 198.845000  9.685000 199.045000 ;
        RECT  9.485000 199.250000  9.685000 199.450000 ;
        RECT  9.485000 199.655000  9.685000 199.855000 ;
        RECT  9.525000  25.910000  9.725000  26.110000 ;
        RECT  9.525000  26.340000  9.725000  26.540000 ;
        RECT  9.525000  26.770000  9.725000  26.970000 ;
        RECT  9.525000  27.200000  9.725000  27.400000 ;
        RECT  9.525000  27.630000  9.725000  27.830000 ;
        RECT  9.525000  28.060000  9.725000  28.260000 ;
        RECT  9.525000  28.490000  9.725000  28.690000 ;
        RECT  9.525000  28.920000  9.725000  29.120000 ;
        RECT  9.525000  29.350000  9.725000  29.550000 ;
        RECT  9.525000  29.780000  9.725000  29.980000 ;
        RECT  9.525000  30.210000  9.725000  30.410000 ;
        RECT  9.885000 175.995000 10.085000 176.195000 ;
        RECT  9.885000 176.395000 10.085000 176.595000 ;
        RECT  9.885000 176.795000 10.085000 176.995000 ;
        RECT  9.885000 177.195000 10.085000 177.395000 ;
        RECT  9.885000 177.595000 10.085000 177.795000 ;
        RECT  9.885000 177.995000 10.085000 178.195000 ;
        RECT  9.885000 178.395000 10.085000 178.595000 ;
        RECT  9.885000 178.795000 10.085000 178.995000 ;
        RECT  9.885000 179.195000 10.085000 179.395000 ;
        RECT  9.885000 179.595000 10.085000 179.795000 ;
        RECT  9.885000 179.995000 10.085000 180.195000 ;
        RECT  9.885000 180.395000 10.085000 180.595000 ;
        RECT  9.885000 180.795000 10.085000 180.995000 ;
        RECT  9.885000 181.195000 10.085000 181.395000 ;
        RECT  9.885000 181.595000 10.085000 181.795000 ;
        RECT  9.885000 181.995000 10.085000 182.195000 ;
        RECT  9.885000 182.395000 10.085000 182.595000 ;
        RECT  9.885000 182.795000 10.085000 182.995000 ;
        RECT  9.885000 183.195000 10.085000 183.395000 ;
        RECT  9.885000 183.595000 10.085000 183.795000 ;
        RECT  9.885000 183.995000 10.085000 184.195000 ;
        RECT  9.885000 184.395000 10.085000 184.595000 ;
        RECT  9.885000 184.795000 10.085000 184.995000 ;
        RECT  9.885000 185.195000 10.085000 185.395000 ;
        RECT  9.885000 185.595000 10.085000 185.795000 ;
        RECT  9.885000 185.995000 10.085000 186.195000 ;
        RECT  9.885000 186.395000 10.085000 186.595000 ;
        RECT  9.885000 186.795000 10.085000 186.995000 ;
        RECT  9.885000 187.195000 10.085000 187.395000 ;
        RECT  9.885000 187.595000 10.085000 187.795000 ;
        RECT  9.885000 187.995000 10.085000 188.195000 ;
        RECT  9.885000 188.395000 10.085000 188.595000 ;
        RECT  9.885000 188.795000 10.085000 188.995000 ;
        RECT  9.885000 189.195000 10.085000 189.395000 ;
        RECT  9.885000 189.595000 10.085000 189.795000 ;
        RECT  9.885000 189.995000 10.085000 190.195000 ;
        RECT  9.885000 190.395000 10.085000 190.595000 ;
        RECT  9.885000 190.795000 10.085000 190.995000 ;
        RECT  9.885000 191.195000 10.085000 191.395000 ;
        RECT  9.885000 191.595000 10.085000 191.795000 ;
        RECT  9.885000 191.995000 10.085000 192.195000 ;
        RECT  9.885000 192.395000 10.085000 192.595000 ;
        RECT  9.885000 192.795000 10.085000 192.995000 ;
        RECT  9.885000 193.195000 10.085000 193.395000 ;
        RECT  9.885000 193.595000 10.085000 193.795000 ;
        RECT  9.885000 193.995000 10.085000 194.195000 ;
        RECT  9.885000 194.395000 10.085000 194.595000 ;
        RECT  9.885000 194.795000 10.085000 194.995000 ;
        RECT  9.885000 195.200000 10.085000 195.400000 ;
        RECT  9.885000 195.605000 10.085000 195.805000 ;
        RECT  9.885000 196.010000 10.085000 196.210000 ;
        RECT  9.885000 196.415000 10.085000 196.615000 ;
        RECT  9.885000 196.820000 10.085000 197.020000 ;
        RECT  9.885000 197.225000 10.085000 197.425000 ;
        RECT  9.885000 197.630000 10.085000 197.830000 ;
        RECT  9.885000 198.035000 10.085000 198.235000 ;
        RECT  9.885000 198.440000 10.085000 198.640000 ;
        RECT  9.885000 198.845000 10.085000 199.045000 ;
        RECT  9.885000 199.250000 10.085000 199.450000 ;
        RECT  9.885000 199.655000 10.085000 199.855000 ;
        RECT  9.930000  25.910000 10.130000  26.110000 ;
        RECT  9.930000  26.340000 10.130000  26.540000 ;
        RECT  9.930000  26.770000 10.130000  26.970000 ;
        RECT  9.930000  27.200000 10.130000  27.400000 ;
        RECT  9.930000  27.630000 10.130000  27.830000 ;
        RECT  9.930000  28.060000 10.130000  28.260000 ;
        RECT  9.930000  28.490000 10.130000  28.690000 ;
        RECT  9.930000  28.920000 10.130000  29.120000 ;
        RECT  9.930000  29.350000 10.130000  29.550000 ;
        RECT  9.930000  29.780000 10.130000  29.980000 ;
        RECT  9.930000  30.210000 10.130000  30.410000 ;
        RECT 10.285000 175.995000 10.485000 176.195000 ;
        RECT 10.285000 176.395000 10.485000 176.595000 ;
        RECT 10.285000 176.795000 10.485000 176.995000 ;
        RECT 10.285000 177.195000 10.485000 177.395000 ;
        RECT 10.285000 177.595000 10.485000 177.795000 ;
        RECT 10.285000 177.995000 10.485000 178.195000 ;
        RECT 10.285000 178.395000 10.485000 178.595000 ;
        RECT 10.285000 178.795000 10.485000 178.995000 ;
        RECT 10.285000 179.195000 10.485000 179.395000 ;
        RECT 10.285000 179.595000 10.485000 179.795000 ;
        RECT 10.285000 179.995000 10.485000 180.195000 ;
        RECT 10.285000 180.395000 10.485000 180.595000 ;
        RECT 10.285000 180.795000 10.485000 180.995000 ;
        RECT 10.285000 181.195000 10.485000 181.395000 ;
        RECT 10.285000 181.595000 10.485000 181.795000 ;
        RECT 10.285000 181.995000 10.485000 182.195000 ;
        RECT 10.285000 182.395000 10.485000 182.595000 ;
        RECT 10.285000 182.795000 10.485000 182.995000 ;
        RECT 10.285000 183.195000 10.485000 183.395000 ;
        RECT 10.285000 183.595000 10.485000 183.795000 ;
        RECT 10.285000 183.995000 10.485000 184.195000 ;
        RECT 10.285000 184.395000 10.485000 184.595000 ;
        RECT 10.285000 184.795000 10.485000 184.995000 ;
        RECT 10.285000 185.195000 10.485000 185.395000 ;
        RECT 10.285000 185.595000 10.485000 185.795000 ;
        RECT 10.285000 185.995000 10.485000 186.195000 ;
        RECT 10.285000 186.395000 10.485000 186.595000 ;
        RECT 10.285000 186.795000 10.485000 186.995000 ;
        RECT 10.285000 187.195000 10.485000 187.395000 ;
        RECT 10.285000 187.595000 10.485000 187.795000 ;
        RECT 10.285000 187.995000 10.485000 188.195000 ;
        RECT 10.285000 188.395000 10.485000 188.595000 ;
        RECT 10.285000 188.795000 10.485000 188.995000 ;
        RECT 10.285000 189.195000 10.485000 189.395000 ;
        RECT 10.285000 189.595000 10.485000 189.795000 ;
        RECT 10.285000 189.995000 10.485000 190.195000 ;
        RECT 10.285000 190.395000 10.485000 190.595000 ;
        RECT 10.285000 190.795000 10.485000 190.995000 ;
        RECT 10.285000 191.195000 10.485000 191.395000 ;
        RECT 10.285000 191.595000 10.485000 191.795000 ;
        RECT 10.285000 191.995000 10.485000 192.195000 ;
        RECT 10.285000 192.395000 10.485000 192.595000 ;
        RECT 10.285000 192.795000 10.485000 192.995000 ;
        RECT 10.285000 193.195000 10.485000 193.395000 ;
        RECT 10.285000 193.595000 10.485000 193.795000 ;
        RECT 10.285000 193.995000 10.485000 194.195000 ;
        RECT 10.285000 194.395000 10.485000 194.595000 ;
        RECT 10.285000 194.795000 10.485000 194.995000 ;
        RECT 10.285000 195.200000 10.485000 195.400000 ;
        RECT 10.285000 195.605000 10.485000 195.805000 ;
        RECT 10.285000 196.010000 10.485000 196.210000 ;
        RECT 10.285000 196.415000 10.485000 196.615000 ;
        RECT 10.285000 196.820000 10.485000 197.020000 ;
        RECT 10.285000 197.225000 10.485000 197.425000 ;
        RECT 10.285000 197.630000 10.485000 197.830000 ;
        RECT 10.285000 198.035000 10.485000 198.235000 ;
        RECT 10.285000 198.440000 10.485000 198.640000 ;
        RECT 10.285000 198.845000 10.485000 199.045000 ;
        RECT 10.285000 199.250000 10.485000 199.450000 ;
        RECT 10.285000 199.655000 10.485000 199.855000 ;
        RECT 10.335000  25.910000 10.535000  26.110000 ;
        RECT 10.335000  26.340000 10.535000  26.540000 ;
        RECT 10.335000  26.770000 10.535000  26.970000 ;
        RECT 10.335000  27.200000 10.535000  27.400000 ;
        RECT 10.335000  27.630000 10.535000  27.830000 ;
        RECT 10.335000  28.060000 10.535000  28.260000 ;
        RECT 10.335000  28.490000 10.535000  28.690000 ;
        RECT 10.335000  28.920000 10.535000  29.120000 ;
        RECT 10.335000  29.350000 10.535000  29.550000 ;
        RECT 10.335000  29.780000 10.535000  29.980000 ;
        RECT 10.335000  30.210000 10.535000  30.410000 ;
        RECT 10.685000 175.995000 10.885000 176.195000 ;
        RECT 10.685000 176.395000 10.885000 176.595000 ;
        RECT 10.685000 176.795000 10.885000 176.995000 ;
        RECT 10.685000 177.195000 10.885000 177.395000 ;
        RECT 10.685000 177.595000 10.885000 177.795000 ;
        RECT 10.685000 177.995000 10.885000 178.195000 ;
        RECT 10.685000 178.395000 10.885000 178.595000 ;
        RECT 10.685000 178.795000 10.885000 178.995000 ;
        RECT 10.685000 179.195000 10.885000 179.395000 ;
        RECT 10.685000 179.595000 10.885000 179.795000 ;
        RECT 10.685000 179.995000 10.885000 180.195000 ;
        RECT 10.685000 180.395000 10.885000 180.595000 ;
        RECT 10.685000 180.795000 10.885000 180.995000 ;
        RECT 10.685000 181.195000 10.885000 181.395000 ;
        RECT 10.685000 181.595000 10.885000 181.795000 ;
        RECT 10.685000 181.995000 10.885000 182.195000 ;
        RECT 10.685000 182.395000 10.885000 182.595000 ;
        RECT 10.685000 182.795000 10.885000 182.995000 ;
        RECT 10.685000 183.195000 10.885000 183.395000 ;
        RECT 10.685000 183.595000 10.885000 183.795000 ;
        RECT 10.685000 183.995000 10.885000 184.195000 ;
        RECT 10.685000 184.395000 10.885000 184.595000 ;
        RECT 10.685000 184.795000 10.885000 184.995000 ;
        RECT 10.685000 185.195000 10.885000 185.395000 ;
        RECT 10.685000 185.595000 10.885000 185.795000 ;
        RECT 10.685000 185.995000 10.885000 186.195000 ;
        RECT 10.685000 186.395000 10.885000 186.595000 ;
        RECT 10.685000 186.795000 10.885000 186.995000 ;
        RECT 10.685000 187.195000 10.885000 187.395000 ;
        RECT 10.685000 187.595000 10.885000 187.795000 ;
        RECT 10.685000 187.995000 10.885000 188.195000 ;
        RECT 10.685000 188.395000 10.885000 188.595000 ;
        RECT 10.685000 188.795000 10.885000 188.995000 ;
        RECT 10.685000 189.195000 10.885000 189.395000 ;
        RECT 10.685000 189.595000 10.885000 189.795000 ;
        RECT 10.685000 189.995000 10.885000 190.195000 ;
        RECT 10.685000 190.395000 10.885000 190.595000 ;
        RECT 10.685000 190.795000 10.885000 190.995000 ;
        RECT 10.685000 191.195000 10.885000 191.395000 ;
        RECT 10.685000 191.595000 10.885000 191.795000 ;
        RECT 10.685000 191.995000 10.885000 192.195000 ;
        RECT 10.685000 192.395000 10.885000 192.595000 ;
        RECT 10.685000 192.795000 10.885000 192.995000 ;
        RECT 10.685000 193.195000 10.885000 193.395000 ;
        RECT 10.685000 193.595000 10.885000 193.795000 ;
        RECT 10.685000 193.995000 10.885000 194.195000 ;
        RECT 10.685000 194.395000 10.885000 194.595000 ;
        RECT 10.685000 194.795000 10.885000 194.995000 ;
        RECT 10.685000 195.200000 10.885000 195.400000 ;
        RECT 10.685000 195.605000 10.885000 195.805000 ;
        RECT 10.685000 196.010000 10.885000 196.210000 ;
        RECT 10.685000 196.415000 10.885000 196.615000 ;
        RECT 10.685000 196.820000 10.885000 197.020000 ;
        RECT 10.685000 197.225000 10.885000 197.425000 ;
        RECT 10.685000 197.630000 10.885000 197.830000 ;
        RECT 10.685000 198.035000 10.885000 198.235000 ;
        RECT 10.685000 198.440000 10.885000 198.640000 ;
        RECT 10.685000 198.845000 10.885000 199.045000 ;
        RECT 10.685000 199.250000 10.885000 199.450000 ;
        RECT 10.685000 199.655000 10.885000 199.855000 ;
        RECT 10.740000  25.910000 10.940000  26.110000 ;
        RECT 10.740000  26.340000 10.940000  26.540000 ;
        RECT 10.740000  26.770000 10.940000  26.970000 ;
        RECT 10.740000  27.200000 10.940000  27.400000 ;
        RECT 10.740000  27.630000 10.940000  27.830000 ;
        RECT 10.740000  28.060000 10.940000  28.260000 ;
        RECT 10.740000  28.490000 10.940000  28.690000 ;
        RECT 10.740000  28.920000 10.940000  29.120000 ;
        RECT 10.740000  29.350000 10.940000  29.550000 ;
        RECT 10.740000  29.780000 10.940000  29.980000 ;
        RECT 10.740000  30.210000 10.940000  30.410000 ;
        RECT 11.085000 175.995000 11.285000 176.195000 ;
        RECT 11.085000 176.395000 11.285000 176.595000 ;
        RECT 11.085000 176.795000 11.285000 176.995000 ;
        RECT 11.085000 177.195000 11.285000 177.395000 ;
        RECT 11.085000 177.595000 11.285000 177.795000 ;
        RECT 11.085000 177.995000 11.285000 178.195000 ;
        RECT 11.085000 178.395000 11.285000 178.595000 ;
        RECT 11.085000 178.795000 11.285000 178.995000 ;
        RECT 11.085000 179.195000 11.285000 179.395000 ;
        RECT 11.085000 179.595000 11.285000 179.795000 ;
        RECT 11.085000 179.995000 11.285000 180.195000 ;
        RECT 11.085000 180.395000 11.285000 180.595000 ;
        RECT 11.085000 180.795000 11.285000 180.995000 ;
        RECT 11.085000 181.195000 11.285000 181.395000 ;
        RECT 11.085000 181.595000 11.285000 181.795000 ;
        RECT 11.085000 181.995000 11.285000 182.195000 ;
        RECT 11.085000 182.395000 11.285000 182.595000 ;
        RECT 11.085000 182.795000 11.285000 182.995000 ;
        RECT 11.085000 183.195000 11.285000 183.395000 ;
        RECT 11.085000 183.595000 11.285000 183.795000 ;
        RECT 11.085000 183.995000 11.285000 184.195000 ;
        RECT 11.085000 184.395000 11.285000 184.595000 ;
        RECT 11.085000 184.795000 11.285000 184.995000 ;
        RECT 11.085000 185.195000 11.285000 185.395000 ;
        RECT 11.085000 185.595000 11.285000 185.795000 ;
        RECT 11.085000 185.995000 11.285000 186.195000 ;
        RECT 11.085000 186.395000 11.285000 186.595000 ;
        RECT 11.085000 186.795000 11.285000 186.995000 ;
        RECT 11.085000 187.195000 11.285000 187.395000 ;
        RECT 11.085000 187.595000 11.285000 187.795000 ;
        RECT 11.085000 187.995000 11.285000 188.195000 ;
        RECT 11.085000 188.395000 11.285000 188.595000 ;
        RECT 11.085000 188.795000 11.285000 188.995000 ;
        RECT 11.085000 189.195000 11.285000 189.395000 ;
        RECT 11.085000 189.595000 11.285000 189.795000 ;
        RECT 11.085000 189.995000 11.285000 190.195000 ;
        RECT 11.085000 190.395000 11.285000 190.595000 ;
        RECT 11.085000 190.795000 11.285000 190.995000 ;
        RECT 11.085000 191.195000 11.285000 191.395000 ;
        RECT 11.085000 191.595000 11.285000 191.795000 ;
        RECT 11.085000 191.995000 11.285000 192.195000 ;
        RECT 11.085000 192.395000 11.285000 192.595000 ;
        RECT 11.085000 192.795000 11.285000 192.995000 ;
        RECT 11.085000 193.195000 11.285000 193.395000 ;
        RECT 11.085000 193.595000 11.285000 193.795000 ;
        RECT 11.085000 193.995000 11.285000 194.195000 ;
        RECT 11.085000 194.395000 11.285000 194.595000 ;
        RECT 11.085000 194.795000 11.285000 194.995000 ;
        RECT 11.085000 195.200000 11.285000 195.400000 ;
        RECT 11.085000 195.605000 11.285000 195.805000 ;
        RECT 11.085000 196.010000 11.285000 196.210000 ;
        RECT 11.085000 196.415000 11.285000 196.615000 ;
        RECT 11.085000 196.820000 11.285000 197.020000 ;
        RECT 11.085000 197.225000 11.285000 197.425000 ;
        RECT 11.085000 197.630000 11.285000 197.830000 ;
        RECT 11.085000 198.035000 11.285000 198.235000 ;
        RECT 11.085000 198.440000 11.285000 198.640000 ;
        RECT 11.085000 198.845000 11.285000 199.045000 ;
        RECT 11.085000 199.250000 11.285000 199.450000 ;
        RECT 11.085000 199.655000 11.285000 199.855000 ;
        RECT 11.145000  25.910000 11.345000  26.110000 ;
        RECT 11.145000  26.340000 11.345000  26.540000 ;
        RECT 11.145000  26.770000 11.345000  26.970000 ;
        RECT 11.145000  27.200000 11.345000  27.400000 ;
        RECT 11.145000  27.630000 11.345000  27.830000 ;
        RECT 11.145000  28.060000 11.345000  28.260000 ;
        RECT 11.145000  28.490000 11.345000  28.690000 ;
        RECT 11.145000  28.920000 11.345000  29.120000 ;
        RECT 11.145000  29.350000 11.345000  29.550000 ;
        RECT 11.145000  29.780000 11.345000  29.980000 ;
        RECT 11.145000  30.210000 11.345000  30.410000 ;
        RECT 11.485000 175.995000 11.685000 176.195000 ;
        RECT 11.485000 176.395000 11.685000 176.595000 ;
        RECT 11.485000 176.795000 11.685000 176.995000 ;
        RECT 11.485000 177.195000 11.685000 177.395000 ;
        RECT 11.485000 177.595000 11.685000 177.795000 ;
        RECT 11.485000 177.995000 11.685000 178.195000 ;
        RECT 11.485000 178.395000 11.685000 178.595000 ;
        RECT 11.485000 178.795000 11.685000 178.995000 ;
        RECT 11.485000 179.195000 11.685000 179.395000 ;
        RECT 11.485000 179.595000 11.685000 179.795000 ;
        RECT 11.485000 179.995000 11.685000 180.195000 ;
        RECT 11.485000 180.395000 11.685000 180.595000 ;
        RECT 11.485000 180.795000 11.685000 180.995000 ;
        RECT 11.485000 181.195000 11.685000 181.395000 ;
        RECT 11.485000 181.595000 11.685000 181.795000 ;
        RECT 11.485000 181.995000 11.685000 182.195000 ;
        RECT 11.485000 182.395000 11.685000 182.595000 ;
        RECT 11.485000 182.795000 11.685000 182.995000 ;
        RECT 11.485000 183.195000 11.685000 183.395000 ;
        RECT 11.485000 183.595000 11.685000 183.795000 ;
        RECT 11.485000 183.995000 11.685000 184.195000 ;
        RECT 11.485000 184.395000 11.685000 184.595000 ;
        RECT 11.485000 184.795000 11.685000 184.995000 ;
        RECT 11.485000 185.195000 11.685000 185.395000 ;
        RECT 11.485000 185.595000 11.685000 185.795000 ;
        RECT 11.485000 185.995000 11.685000 186.195000 ;
        RECT 11.485000 186.395000 11.685000 186.595000 ;
        RECT 11.485000 186.795000 11.685000 186.995000 ;
        RECT 11.485000 187.195000 11.685000 187.395000 ;
        RECT 11.485000 187.595000 11.685000 187.795000 ;
        RECT 11.485000 187.995000 11.685000 188.195000 ;
        RECT 11.485000 188.395000 11.685000 188.595000 ;
        RECT 11.485000 188.795000 11.685000 188.995000 ;
        RECT 11.485000 189.195000 11.685000 189.395000 ;
        RECT 11.485000 189.595000 11.685000 189.795000 ;
        RECT 11.485000 189.995000 11.685000 190.195000 ;
        RECT 11.485000 190.395000 11.685000 190.595000 ;
        RECT 11.485000 190.795000 11.685000 190.995000 ;
        RECT 11.485000 191.195000 11.685000 191.395000 ;
        RECT 11.485000 191.595000 11.685000 191.795000 ;
        RECT 11.485000 191.995000 11.685000 192.195000 ;
        RECT 11.485000 192.395000 11.685000 192.595000 ;
        RECT 11.485000 192.795000 11.685000 192.995000 ;
        RECT 11.485000 193.195000 11.685000 193.395000 ;
        RECT 11.485000 193.595000 11.685000 193.795000 ;
        RECT 11.485000 193.995000 11.685000 194.195000 ;
        RECT 11.485000 194.395000 11.685000 194.595000 ;
        RECT 11.485000 194.795000 11.685000 194.995000 ;
        RECT 11.485000 195.200000 11.685000 195.400000 ;
        RECT 11.485000 195.605000 11.685000 195.805000 ;
        RECT 11.485000 196.010000 11.685000 196.210000 ;
        RECT 11.485000 196.415000 11.685000 196.615000 ;
        RECT 11.485000 196.820000 11.685000 197.020000 ;
        RECT 11.485000 197.225000 11.685000 197.425000 ;
        RECT 11.485000 197.630000 11.685000 197.830000 ;
        RECT 11.485000 198.035000 11.685000 198.235000 ;
        RECT 11.485000 198.440000 11.685000 198.640000 ;
        RECT 11.485000 198.845000 11.685000 199.045000 ;
        RECT 11.485000 199.250000 11.685000 199.450000 ;
        RECT 11.485000 199.655000 11.685000 199.855000 ;
        RECT 11.550000  25.910000 11.750000  26.110000 ;
        RECT 11.550000  26.340000 11.750000  26.540000 ;
        RECT 11.550000  26.770000 11.750000  26.970000 ;
        RECT 11.550000  27.200000 11.750000  27.400000 ;
        RECT 11.550000  27.630000 11.750000  27.830000 ;
        RECT 11.550000  28.060000 11.750000  28.260000 ;
        RECT 11.550000  28.490000 11.750000  28.690000 ;
        RECT 11.550000  28.920000 11.750000  29.120000 ;
        RECT 11.550000  29.350000 11.750000  29.550000 ;
        RECT 11.550000  29.780000 11.750000  29.980000 ;
        RECT 11.550000  30.210000 11.750000  30.410000 ;
        RECT 11.885000 175.995000 12.085000 176.195000 ;
        RECT 11.885000 176.395000 12.085000 176.595000 ;
        RECT 11.885000 176.795000 12.085000 176.995000 ;
        RECT 11.885000 177.195000 12.085000 177.395000 ;
        RECT 11.885000 177.595000 12.085000 177.795000 ;
        RECT 11.885000 177.995000 12.085000 178.195000 ;
        RECT 11.885000 178.395000 12.085000 178.595000 ;
        RECT 11.885000 178.795000 12.085000 178.995000 ;
        RECT 11.885000 179.195000 12.085000 179.395000 ;
        RECT 11.885000 179.595000 12.085000 179.795000 ;
        RECT 11.885000 179.995000 12.085000 180.195000 ;
        RECT 11.885000 180.395000 12.085000 180.595000 ;
        RECT 11.885000 180.795000 12.085000 180.995000 ;
        RECT 11.885000 181.195000 12.085000 181.395000 ;
        RECT 11.885000 181.595000 12.085000 181.795000 ;
        RECT 11.885000 181.995000 12.085000 182.195000 ;
        RECT 11.885000 182.395000 12.085000 182.595000 ;
        RECT 11.885000 182.795000 12.085000 182.995000 ;
        RECT 11.885000 183.195000 12.085000 183.395000 ;
        RECT 11.885000 183.595000 12.085000 183.795000 ;
        RECT 11.885000 183.995000 12.085000 184.195000 ;
        RECT 11.885000 184.395000 12.085000 184.595000 ;
        RECT 11.885000 184.795000 12.085000 184.995000 ;
        RECT 11.885000 185.195000 12.085000 185.395000 ;
        RECT 11.885000 185.595000 12.085000 185.795000 ;
        RECT 11.885000 185.995000 12.085000 186.195000 ;
        RECT 11.885000 186.395000 12.085000 186.595000 ;
        RECT 11.885000 186.795000 12.085000 186.995000 ;
        RECT 11.885000 187.195000 12.085000 187.395000 ;
        RECT 11.885000 187.595000 12.085000 187.795000 ;
        RECT 11.885000 187.995000 12.085000 188.195000 ;
        RECT 11.885000 188.395000 12.085000 188.595000 ;
        RECT 11.885000 188.795000 12.085000 188.995000 ;
        RECT 11.885000 189.195000 12.085000 189.395000 ;
        RECT 11.885000 189.595000 12.085000 189.795000 ;
        RECT 11.885000 189.995000 12.085000 190.195000 ;
        RECT 11.885000 190.395000 12.085000 190.595000 ;
        RECT 11.885000 190.795000 12.085000 190.995000 ;
        RECT 11.885000 191.195000 12.085000 191.395000 ;
        RECT 11.885000 191.595000 12.085000 191.795000 ;
        RECT 11.885000 191.995000 12.085000 192.195000 ;
        RECT 11.885000 192.395000 12.085000 192.595000 ;
        RECT 11.885000 192.795000 12.085000 192.995000 ;
        RECT 11.885000 193.195000 12.085000 193.395000 ;
        RECT 11.885000 193.595000 12.085000 193.795000 ;
        RECT 11.885000 193.995000 12.085000 194.195000 ;
        RECT 11.885000 194.395000 12.085000 194.595000 ;
        RECT 11.885000 194.795000 12.085000 194.995000 ;
        RECT 11.885000 195.200000 12.085000 195.400000 ;
        RECT 11.885000 195.605000 12.085000 195.805000 ;
        RECT 11.885000 196.010000 12.085000 196.210000 ;
        RECT 11.885000 196.415000 12.085000 196.615000 ;
        RECT 11.885000 196.820000 12.085000 197.020000 ;
        RECT 11.885000 197.225000 12.085000 197.425000 ;
        RECT 11.885000 197.630000 12.085000 197.830000 ;
        RECT 11.885000 198.035000 12.085000 198.235000 ;
        RECT 11.885000 198.440000 12.085000 198.640000 ;
        RECT 11.885000 198.845000 12.085000 199.045000 ;
        RECT 11.885000 199.250000 12.085000 199.450000 ;
        RECT 11.885000 199.655000 12.085000 199.855000 ;
        RECT 11.955000  25.910000 12.155000  26.110000 ;
        RECT 11.955000  26.340000 12.155000  26.540000 ;
        RECT 11.955000  26.770000 12.155000  26.970000 ;
        RECT 11.955000  27.200000 12.155000  27.400000 ;
        RECT 11.955000  27.630000 12.155000  27.830000 ;
        RECT 11.955000  28.060000 12.155000  28.260000 ;
        RECT 11.955000  28.490000 12.155000  28.690000 ;
        RECT 11.955000  28.920000 12.155000  29.120000 ;
        RECT 11.955000  29.350000 12.155000  29.550000 ;
        RECT 11.955000  29.780000 12.155000  29.980000 ;
        RECT 11.955000  30.210000 12.155000  30.410000 ;
        RECT 12.285000 175.995000 12.485000 176.195000 ;
        RECT 12.285000 176.395000 12.485000 176.595000 ;
        RECT 12.285000 176.795000 12.485000 176.995000 ;
        RECT 12.285000 177.195000 12.485000 177.395000 ;
        RECT 12.285000 177.595000 12.485000 177.795000 ;
        RECT 12.285000 177.995000 12.485000 178.195000 ;
        RECT 12.285000 178.395000 12.485000 178.595000 ;
        RECT 12.285000 178.795000 12.485000 178.995000 ;
        RECT 12.285000 179.195000 12.485000 179.395000 ;
        RECT 12.285000 179.595000 12.485000 179.795000 ;
        RECT 12.285000 179.995000 12.485000 180.195000 ;
        RECT 12.285000 180.395000 12.485000 180.595000 ;
        RECT 12.285000 180.795000 12.485000 180.995000 ;
        RECT 12.285000 181.195000 12.485000 181.395000 ;
        RECT 12.285000 181.595000 12.485000 181.795000 ;
        RECT 12.285000 181.995000 12.485000 182.195000 ;
        RECT 12.285000 182.395000 12.485000 182.595000 ;
        RECT 12.285000 182.795000 12.485000 182.995000 ;
        RECT 12.285000 183.195000 12.485000 183.395000 ;
        RECT 12.285000 183.595000 12.485000 183.795000 ;
        RECT 12.285000 183.995000 12.485000 184.195000 ;
        RECT 12.285000 184.395000 12.485000 184.595000 ;
        RECT 12.285000 184.795000 12.485000 184.995000 ;
        RECT 12.285000 185.195000 12.485000 185.395000 ;
        RECT 12.285000 185.595000 12.485000 185.795000 ;
        RECT 12.285000 185.995000 12.485000 186.195000 ;
        RECT 12.285000 186.395000 12.485000 186.595000 ;
        RECT 12.285000 186.795000 12.485000 186.995000 ;
        RECT 12.285000 187.195000 12.485000 187.395000 ;
        RECT 12.285000 187.595000 12.485000 187.795000 ;
        RECT 12.285000 187.995000 12.485000 188.195000 ;
        RECT 12.285000 188.395000 12.485000 188.595000 ;
        RECT 12.285000 188.795000 12.485000 188.995000 ;
        RECT 12.285000 189.195000 12.485000 189.395000 ;
        RECT 12.285000 189.595000 12.485000 189.795000 ;
        RECT 12.285000 189.995000 12.485000 190.195000 ;
        RECT 12.285000 190.395000 12.485000 190.595000 ;
        RECT 12.285000 190.795000 12.485000 190.995000 ;
        RECT 12.285000 191.195000 12.485000 191.395000 ;
        RECT 12.285000 191.595000 12.485000 191.795000 ;
        RECT 12.285000 191.995000 12.485000 192.195000 ;
        RECT 12.285000 192.395000 12.485000 192.595000 ;
        RECT 12.285000 192.795000 12.485000 192.995000 ;
        RECT 12.285000 193.195000 12.485000 193.395000 ;
        RECT 12.285000 193.595000 12.485000 193.795000 ;
        RECT 12.285000 193.995000 12.485000 194.195000 ;
        RECT 12.285000 194.395000 12.485000 194.595000 ;
        RECT 12.285000 194.795000 12.485000 194.995000 ;
        RECT 12.285000 195.200000 12.485000 195.400000 ;
        RECT 12.285000 195.605000 12.485000 195.805000 ;
        RECT 12.285000 196.010000 12.485000 196.210000 ;
        RECT 12.285000 196.415000 12.485000 196.615000 ;
        RECT 12.285000 196.820000 12.485000 197.020000 ;
        RECT 12.285000 197.225000 12.485000 197.425000 ;
        RECT 12.285000 197.630000 12.485000 197.830000 ;
        RECT 12.285000 198.035000 12.485000 198.235000 ;
        RECT 12.285000 198.440000 12.485000 198.640000 ;
        RECT 12.285000 198.845000 12.485000 199.045000 ;
        RECT 12.285000 199.250000 12.485000 199.450000 ;
        RECT 12.285000 199.655000 12.485000 199.855000 ;
        RECT 12.360000  25.910000 12.560000  26.110000 ;
        RECT 12.360000  26.340000 12.560000  26.540000 ;
        RECT 12.360000  26.770000 12.560000  26.970000 ;
        RECT 12.360000  27.200000 12.560000  27.400000 ;
        RECT 12.360000  27.630000 12.560000  27.830000 ;
        RECT 12.360000  28.060000 12.560000  28.260000 ;
        RECT 12.360000  28.490000 12.560000  28.690000 ;
        RECT 12.360000  28.920000 12.560000  29.120000 ;
        RECT 12.360000  29.350000 12.560000  29.550000 ;
        RECT 12.360000  29.780000 12.560000  29.980000 ;
        RECT 12.360000  30.210000 12.560000  30.410000 ;
        RECT 12.685000 175.995000 12.885000 176.195000 ;
        RECT 12.685000 176.395000 12.885000 176.595000 ;
        RECT 12.685000 176.795000 12.885000 176.995000 ;
        RECT 12.685000 177.195000 12.885000 177.395000 ;
        RECT 12.685000 177.595000 12.885000 177.795000 ;
        RECT 12.685000 177.995000 12.885000 178.195000 ;
        RECT 12.685000 178.395000 12.885000 178.595000 ;
        RECT 12.685000 178.795000 12.885000 178.995000 ;
        RECT 12.685000 179.195000 12.885000 179.395000 ;
        RECT 12.685000 179.595000 12.885000 179.795000 ;
        RECT 12.685000 179.995000 12.885000 180.195000 ;
        RECT 12.685000 180.395000 12.885000 180.595000 ;
        RECT 12.685000 180.795000 12.885000 180.995000 ;
        RECT 12.685000 181.195000 12.885000 181.395000 ;
        RECT 12.685000 181.595000 12.885000 181.795000 ;
        RECT 12.685000 181.995000 12.885000 182.195000 ;
        RECT 12.685000 182.395000 12.885000 182.595000 ;
        RECT 12.685000 182.795000 12.885000 182.995000 ;
        RECT 12.685000 183.195000 12.885000 183.395000 ;
        RECT 12.685000 183.595000 12.885000 183.795000 ;
        RECT 12.685000 183.995000 12.885000 184.195000 ;
        RECT 12.685000 184.395000 12.885000 184.595000 ;
        RECT 12.685000 184.795000 12.885000 184.995000 ;
        RECT 12.685000 185.195000 12.885000 185.395000 ;
        RECT 12.685000 185.595000 12.885000 185.795000 ;
        RECT 12.685000 185.995000 12.885000 186.195000 ;
        RECT 12.685000 186.395000 12.885000 186.595000 ;
        RECT 12.685000 186.795000 12.885000 186.995000 ;
        RECT 12.685000 187.195000 12.885000 187.395000 ;
        RECT 12.685000 187.595000 12.885000 187.795000 ;
        RECT 12.685000 187.995000 12.885000 188.195000 ;
        RECT 12.685000 188.395000 12.885000 188.595000 ;
        RECT 12.685000 188.795000 12.885000 188.995000 ;
        RECT 12.685000 189.195000 12.885000 189.395000 ;
        RECT 12.685000 189.595000 12.885000 189.795000 ;
        RECT 12.685000 189.995000 12.885000 190.195000 ;
        RECT 12.685000 190.395000 12.885000 190.595000 ;
        RECT 12.685000 190.795000 12.885000 190.995000 ;
        RECT 12.685000 191.195000 12.885000 191.395000 ;
        RECT 12.685000 191.595000 12.885000 191.795000 ;
        RECT 12.685000 191.995000 12.885000 192.195000 ;
        RECT 12.685000 192.395000 12.885000 192.595000 ;
        RECT 12.685000 192.795000 12.885000 192.995000 ;
        RECT 12.685000 193.195000 12.885000 193.395000 ;
        RECT 12.685000 193.595000 12.885000 193.795000 ;
        RECT 12.685000 193.995000 12.885000 194.195000 ;
        RECT 12.685000 194.395000 12.885000 194.595000 ;
        RECT 12.685000 194.795000 12.885000 194.995000 ;
        RECT 12.685000 195.200000 12.885000 195.400000 ;
        RECT 12.685000 195.605000 12.885000 195.805000 ;
        RECT 12.685000 196.010000 12.885000 196.210000 ;
        RECT 12.685000 196.415000 12.885000 196.615000 ;
        RECT 12.685000 196.820000 12.885000 197.020000 ;
        RECT 12.685000 197.225000 12.885000 197.425000 ;
        RECT 12.685000 197.630000 12.885000 197.830000 ;
        RECT 12.685000 198.035000 12.885000 198.235000 ;
        RECT 12.685000 198.440000 12.885000 198.640000 ;
        RECT 12.685000 198.845000 12.885000 199.045000 ;
        RECT 12.685000 199.250000 12.885000 199.450000 ;
        RECT 12.685000 199.655000 12.885000 199.855000 ;
        RECT 12.765000  25.910000 12.965000  26.110000 ;
        RECT 12.765000  26.340000 12.965000  26.540000 ;
        RECT 12.765000  26.770000 12.965000  26.970000 ;
        RECT 12.765000  27.200000 12.965000  27.400000 ;
        RECT 12.765000  27.630000 12.965000  27.830000 ;
        RECT 12.765000  28.060000 12.965000  28.260000 ;
        RECT 12.765000  28.490000 12.965000  28.690000 ;
        RECT 12.765000  28.920000 12.965000  29.120000 ;
        RECT 12.765000  29.350000 12.965000  29.550000 ;
        RECT 12.765000  29.780000 12.965000  29.980000 ;
        RECT 12.765000  30.210000 12.965000  30.410000 ;
        RECT 13.085000 175.995000 13.285000 176.195000 ;
        RECT 13.085000 176.395000 13.285000 176.595000 ;
        RECT 13.085000 176.795000 13.285000 176.995000 ;
        RECT 13.085000 177.195000 13.285000 177.395000 ;
        RECT 13.085000 177.595000 13.285000 177.795000 ;
        RECT 13.085000 177.995000 13.285000 178.195000 ;
        RECT 13.085000 178.395000 13.285000 178.595000 ;
        RECT 13.085000 178.795000 13.285000 178.995000 ;
        RECT 13.085000 179.195000 13.285000 179.395000 ;
        RECT 13.085000 179.595000 13.285000 179.795000 ;
        RECT 13.085000 179.995000 13.285000 180.195000 ;
        RECT 13.085000 180.395000 13.285000 180.595000 ;
        RECT 13.085000 180.795000 13.285000 180.995000 ;
        RECT 13.085000 181.195000 13.285000 181.395000 ;
        RECT 13.085000 181.595000 13.285000 181.795000 ;
        RECT 13.085000 181.995000 13.285000 182.195000 ;
        RECT 13.085000 182.395000 13.285000 182.595000 ;
        RECT 13.085000 182.795000 13.285000 182.995000 ;
        RECT 13.085000 183.195000 13.285000 183.395000 ;
        RECT 13.085000 183.595000 13.285000 183.795000 ;
        RECT 13.085000 183.995000 13.285000 184.195000 ;
        RECT 13.085000 184.395000 13.285000 184.595000 ;
        RECT 13.085000 184.795000 13.285000 184.995000 ;
        RECT 13.085000 185.195000 13.285000 185.395000 ;
        RECT 13.085000 185.595000 13.285000 185.795000 ;
        RECT 13.085000 185.995000 13.285000 186.195000 ;
        RECT 13.085000 186.395000 13.285000 186.595000 ;
        RECT 13.085000 186.795000 13.285000 186.995000 ;
        RECT 13.085000 187.195000 13.285000 187.395000 ;
        RECT 13.085000 187.595000 13.285000 187.795000 ;
        RECT 13.085000 187.995000 13.285000 188.195000 ;
        RECT 13.085000 188.395000 13.285000 188.595000 ;
        RECT 13.085000 188.795000 13.285000 188.995000 ;
        RECT 13.085000 189.195000 13.285000 189.395000 ;
        RECT 13.085000 189.595000 13.285000 189.795000 ;
        RECT 13.085000 189.995000 13.285000 190.195000 ;
        RECT 13.085000 190.395000 13.285000 190.595000 ;
        RECT 13.085000 190.795000 13.285000 190.995000 ;
        RECT 13.085000 191.195000 13.285000 191.395000 ;
        RECT 13.085000 191.595000 13.285000 191.795000 ;
        RECT 13.085000 191.995000 13.285000 192.195000 ;
        RECT 13.085000 192.395000 13.285000 192.595000 ;
        RECT 13.085000 192.795000 13.285000 192.995000 ;
        RECT 13.085000 193.195000 13.285000 193.395000 ;
        RECT 13.085000 193.595000 13.285000 193.795000 ;
        RECT 13.085000 193.995000 13.285000 194.195000 ;
        RECT 13.085000 194.395000 13.285000 194.595000 ;
        RECT 13.085000 194.795000 13.285000 194.995000 ;
        RECT 13.085000 195.200000 13.285000 195.400000 ;
        RECT 13.085000 195.605000 13.285000 195.805000 ;
        RECT 13.085000 196.010000 13.285000 196.210000 ;
        RECT 13.085000 196.415000 13.285000 196.615000 ;
        RECT 13.085000 196.820000 13.285000 197.020000 ;
        RECT 13.085000 197.225000 13.285000 197.425000 ;
        RECT 13.085000 197.630000 13.285000 197.830000 ;
        RECT 13.085000 198.035000 13.285000 198.235000 ;
        RECT 13.085000 198.440000 13.285000 198.640000 ;
        RECT 13.085000 198.845000 13.285000 199.045000 ;
        RECT 13.085000 199.250000 13.285000 199.450000 ;
        RECT 13.085000 199.655000 13.285000 199.855000 ;
        RECT 13.170000  25.910000 13.370000  26.110000 ;
        RECT 13.170000  26.340000 13.370000  26.540000 ;
        RECT 13.170000  26.770000 13.370000  26.970000 ;
        RECT 13.170000  27.200000 13.370000  27.400000 ;
        RECT 13.170000  27.630000 13.370000  27.830000 ;
        RECT 13.170000  28.060000 13.370000  28.260000 ;
        RECT 13.170000  28.490000 13.370000  28.690000 ;
        RECT 13.170000  28.920000 13.370000  29.120000 ;
        RECT 13.170000  29.350000 13.370000  29.550000 ;
        RECT 13.170000  29.780000 13.370000  29.980000 ;
        RECT 13.170000  30.210000 13.370000  30.410000 ;
        RECT 13.575000  25.910000 13.775000  26.110000 ;
        RECT 13.575000  26.340000 13.775000  26.540000 ;
        RECT 13.575000  26.770000 13.775000  26.970000 ;
        RECT 13.575000  27.200000 13.775000  27.400000 ;
        RECT 13.575000  27.630000 13.775000  27.830000 ;
        RECT 13.575000  28.060000 13.775000  28.260000 ;
        RECT 13.575000  28.490000 13.775000  28.690000 ;
        RECT 13.575000  28.920000 13.775000  29.120000 ;
        RECT 13.575000  29.350000 13.775000  29.550000 ;
        RECT 13.575000  29.780000 13.775000  29.980000 ;
        RECT 13.575000  30.210000 13.775000  30.410000 ;
        RECT 13.695000 197.250000 13.895000 197.450000 ;
        RECT 13.695000 197.650000 13.895000 197.850000 ;
        RECT 13.695000 198.050000 13.895000 198.250000 ;
        RECT 13.695000 198.450000 13.895000 198.650000 ;
        RECT 13.695000 198.850000 13.895000 199.050000 ;
        RECT 13.695000 199.250000 13.895000 199.450000 ;
        RECT 13.695000 199.650000 13.895000 199.850000 ;
        RECT 13.825000 196.295000 14.025000 196.495000 ;
        RECT 13.825000 196.705000 14.025000 196.905000 ;
        RECT 13.980000  25.910000 14.180000  26.110000 ;
        RECT 13.980000  26.340000 14.180000  26.540000 ;
        RECT 13.980000  26.770000 14.180000  26.970000 ;
        RECT 13.980000  27.200000 14.180000  27.400000 ;
        RECT 13.980000  27.630000 14.180000  27.830000 ;
        RECT 13.980000  28.060000 14.180000  28.260000 ;
        RECT 13.980000  28.490000 14.180000  28.690000 ;
        RECT 13.980000  28.920000 14.180000  29.120000 ;
        RECT 13.980000  29.350000 14.180000  29.550000 ;
        RECT 13.980000  29.780000 14.180000  29.980000 ;
        RECT 13.980000  30.210000 14.180000  30.410000 ;
        RECT 14.100000 197.250000 14.300000 197.450000 ;
        RECT 14.100000 197.650000 14.300000 197.850000 ;
        RECT 14.100000 198.050000 14.300000 198.250000 ;
        RECT 14.100000 198.450000 14.300000 198.650000 ;
        RECT 14.100000 198.850000 14.300000 199.050000 ;
        RECT 14.100000 199.250000 14.300000 199.450000 ;
        RECT 14.100000 199.650000 14.300000 199.850000 ;
        RECT 14.385000  25.910000 14.585000  26.110000 ;
        RECT 14.385000  26.340000 14.585000  26.540000 ;
        RECT 14.385000  26.770000 14.585000  26.970000 ;
        RECT 14.385000  27.200000 14.585000  27.400000 ;
        RECT 14.385000  27.630000 14.585000  27.830000 ;
        RECT 14.385000  28.060000 14.585000  28.260000 ;
        RECT 14.385000  28.490000 14.585000  28.690000 ;
        RECT 14.385000  28.920000 14.585000  29.120000 ;
        RECT 14.385000  29.350000 14.585000  29.550000 ;
        RECT 14.385000  29.780000 14.585000  29.980000 ;
        RECT 14.385000  30.210000 14.585000  30.410000 ;
        RECT 14.505000 197.250000 14.705000 197.450000 ;
        RECT 14.505000 197.650000 14.705000 197.850000 ;
        RECT 14.505000 198.050000 14.705000 198.250000 ;
        RECT 14.505000 198.450000 14.705000 198.650000 ;
        RECT 14.505000 198.850000 14.705000 199.050000 ;
        RECT 14.505000 199.250000 14.705000 199.450000 ;
        RECT 14.505000 199.650000 14.705000 199.850000 ;
        RECT 14.790000  25.910000 14.990000  26.110000 ;
        RECT 14.790000  26.340000 14.990000  26.540000 ;
        RECT 14.790000  26.770000 14.990000  26.970000 ;
        RECT 14.790000  27.200000 14.990000  27.400000 ;
        RECT 14.790000  27.630000 14.990000  27.830000 ;
        RECT 14.790000  28.060000 14.990000  28.260000 ;
        RECT 14.790000  28.490000 14.990000  28.690000 ;
        RECT 14.790000  28.920000 14.990000  29.120000 ;
        RECT 14.790000  29.350000 14.990000  29.550000 ;
        RECT 14.790000  29.780000 14.990000  29.980000 ;
        RECT 14.790000  30.210000 14.990000  30.410000 ;
        RECT 14.910000 197.250000 15.110000 197.450000 ;
        RECT 14.910000 197.650000 15.110000 197.850000 ;
        RECT 14.910000 198.050000 15.110000 198.250000 ;
        RECT 14.910000 198.450000 15.110000 198.650000 ;
        RECT 14.910000 198.850000 15.110000 199.050000 ;
        RECT 14.910000 199.250000 15.110000 199.450000 ;
        RECT 14.910000 199.650000 15.110000 199.850000 ;
        RECT 15.195000  25.910000 15.395000  26.110000 ;
        RECT 15.195000  26.340000 15.395000  26.540000 ;
        RECT 15.195000  26.770000 15.395000  26.970000 ;
        RECT 15.195000  27.200000 15.395000  27.400000 ;
        RECT 15.195000  27.630000 15.395000  27.830000 ;
        RECT 15.195000  28.060000 15.395000  28.260000 ;
        RECT 15.195000  28.490000 15.395000  28.690000 ;
        RECT 15.195000  28.920000 15.395000  29.120000 ;
        RECT 15.195000  29.350000 15.395000  29.550000 ;
        RECT 15.195000  29.780000 15.395000  29.980000 ;
        RECT 15.195000  30.210000 15.395000  30.410000 ;
        RECT 15.315000 197.250000 15.515000 197.450000 ;
        RECT 15.315000 197.650000 15.515000 197.850000 ;
        RECT 15.315000 198.050000 15.515000 198.250000 ;
        RECT 15.315000 198.450000 15.515000 198.650000 ;
        RECT 15.315000 198.850000 15.515000 199.050000 ;
        RECT 15.315000 199.250000 15.515000 199.450000 ;
        RECT 15.315000 199.650000 15.515000 199.850000 ;
        RECT 15.600000  25.910000 15.800000  26.110000 ;
        RECT 15.600000  26.340000 15.800000  26.540000 ;
        RECT 15.600000  26.770000 15.800000  26.970000 ;
        RECT 15.600000  27.200000 15.800000  27.400000 ;
        RECT 15.600000  27.630000 15.800000  27.830000 ;
        RECT 15.600000  28.060000 15.800000  28.260000 ;
        RECT 15.600000  28.490000 15.800000  28.690000 ;
        RECT 15.600000  28.920000 15.800000  29.120000 ;
        RECT 15.600000  29.350000 15.800000  29.550000 ;
        RECT 15.600000  29.780000 15.800000  29.980000 ;
        RECT 15.600000  30.210000 15.800000  30.410000 ;
        RECT 15.720000 197.250000 15.920000 197.450000 ;
        RECT 15.720000 197.650000 15.920000 197.850000 ;
        RECT 15.720000 198.050000 15.920000 198.250000 ;
        RECT 15.720000 198.450000 15.920000 198.650000 ;
        RECT 15.720000 198.850000 15.920000 199.050000 ;
        RECT 15.720000 199.250000 15.920000 199.450000 ;
        RECT 15.720000 199.650000 15.920000 199.850000 ;
        RECT 16.005000  25.910000 16.205000  26.110000 ;
        RECT 16.005000  26.340000 16.205000  26.540000 ;
        RECT 16.005000  26.770000 16.205000  26.970000 ;
        RECT 16.005000  27.200000 16.205000  27.400000 ;
        RECT 16.005000  27.630000 16.205000  27.830000 ;
        RECT 16.005000  28.060000 16.205000  28.260000 ;
        RECT 16.005000  28.490000 16.205000  28.690000 ;
        RECT 16.005000  28.920000 16.205000  29.120000 ;
        RECT 16.005000  29.350000 16.205000  29.550000 ;
        RECT 16.005000  29.780000 16.205000  29.980000 ;
        RECT 16.005000  30.210000 16.205000  30.410000 ;
        RECT 16.125000 197.250000 16.325000 197.450000 ;
        RECT 16.125000 197.650000 16.325000 197.850000 ;
        RECT 16.125000 198.050000 16.325000 198.250000 ;
        RECT 16.125000 198.450000 16.325000 198.650000 ;
        RECT 16.125000 198.850000 16.325000 199.050000 ;
        RECT 16.125000 199.250000 16.325000 199.450000 ;
        RECT 16.125000 199.650000 16.325000 199.850000 ;
        RECT 16.410000  25.910000 16.610000  26.110000 ;
        RECT 16.410000  26.340000 16.610000  26.540000 ;
        RECT 16.410000  26.770000 16.610000  26.970000 ;
        RECT 16.410000  27.200000 16.610000  27.400000 ;
        RECT 16.410000  27.630000 16.610000  27.830000 ;
        RECT 16.410000  28.060000 16.610000  28.260000 ;
        RECT 16.410000  28.490000 16.610000  28.690000 ;
        RECT 16.410000  28.920000 16.610000  29.120000 ;
        RECT 16.410000  29.350000 16.610000  29.550000 ;
        RECT 16.410000  29.780000 16.610000  29.980000 ;
        RECT 16.410000  30.210000 16.610000  30.410000 ;
        RECT 16.530000 197.250000 16.730000 197.450000 ;
        RECT 16.530000 197.650000 16.730000 197.850000 ;
        RECT 16.530000 198.050000 16.730000 198.250000 ;
        RECT 16.530000 198.450000 16.730000 198.650000 ;
        RECT 16.530000 198.850000 16.730000 199.050000 ;
        RECT 16.530000 199.250000 16.730000 199.450000 ;
        RECT 16.530000 199.650000 16.730000 199.850000 ;
        RECT 16.815000  25.910000 17.015000  26.110000 ;
        RECT 16.815000  26.340000 17.015000  26.540000 ;
        RECT 16.815000  26.770000 17.015000  26.970000 ;
        RECT 16.815000  27.200000 17.015000  27.400000 ;
        RECT 16.815000  27.630000 17.015000  27.830000 ;
        RECT 16.815000  28.060000 17.015000  28.260000 ;
        RECT 16.815000  28.490000 17.015000  28.690000 ;
        RECT 16.815000  28.920000 17.015000  29.120000 ;
        RECT 16.815000  29.350000 17.015000  29.550000 ;
        RECT 16.815000  29.780000 17.015000  29.980000 ;
        RECT 16.815000  30.210000 17.015000  30.410000 ;
        RECT 16.935000 197.250000 17.135000 197.450000 ;
        RECT 16.935000 197.650000 17.135000 197.850000 ;
        RECT 16.935000 198.050000 17.135000 198.250000 ;
        RECT 16.935000 198.450000 17.135000 198.650000 ;
        RECT 16.935000 198.850000 17.135000 199.050000 ;
        RECT 16.935000 199.250000 17.135000 199.450000 ;
        RECT 16.935000 199.650000 17.135000 199.850000 ;
        RECT 17.220000  25.910000 17.420000  26.110000 ;
        RECT 17.220000  26.340000 17.420000  26.540000 ;
        RECT 17.220000  26.770000 17.420000  26.970000 ;
        RECT 17.220000  27.200000 17.420000  27.400000 ;
        RECT 17.220000  27.630000 17.420000  27.830000 ;
        RECT 17.220000  28.060000 17.420000  28.260000 ;
        RECT 17.220000  28.490000 17.420000  28.690000 ;
        RECT 17.220000  28.920000 17.420000  29.120000 ;
        RECT 17.220000  29.350000 17.420000  29.550000 ;
        RECT 17.220000  29.780000 17.420000  29.980000 ;
        RECT 17.220000  30.210000 17.420000  30.410000 ;
        RECT 17.340000 197.250000 17.540000 197.450000 ;
        RECT 17.340000 197.650000 17.540000 197.850000 ;
        RECT 17.340000 198.050000 17.540000 198.250000 ;
        RECT 17.340000 198.450000 17.540000 198.650000 ;
        RECT 17.340000 198.850000 17.540000 199.050000 ;
        RECT 17.340000 199.250000 17.540000 199.450000 ;
        RECT 17.340000 199.650000 17.540000 199.850000 ;
        RECT 17.625000  25.910000 17.825000  26.110000 ;
        RECT 17.625000  26.340000 17.825000  26.540000 ;
        RECT 17.625000  26.770000 17.825000  26.970000 ;
        RECT 17.625000  27.200000 17.825000  27.400000 ;
        RECT 17.625000  27.630000 17.825000  27.830000 ;
        RECT 17.625000  28.060000 17.825000  28.260000 ;
        RECT 17.625000  28.490000 17.825000  28.690000 ;
        RECT 17.625000  28.920000 17.825000  29.120000 ;
        RECT 17.625000  29.350000 17.825000  29.550000 ;
        RECT 17.625000  29.780000 17.825000  29.980000 ;
        RECT 17.625000  30.210000 17.825000  30.410000 ;
        RECT 17.745000 197.250000 17.945000 197.450000 ;
        RECT 17.745000 197.650000 17.945000 197.850000 ;
        RECT 17.745000 198.050000 17.945000 198.250000 ;
        RECT 17.745000 198.450000 17.945000 198.650000 ;
        RECT 17.745000 198.850000 17.945000 199.050000 ;
        RECT 17.745000 199.250000 17.945000 199.450000 ;
        RECT 17.745000 199.650000 17.945000 199.850000 ;
        RECT 18.030000  25.910000 18.230000  26.110000 ;
        RECT 18.030000  26.340000 18.230000  26.540000 ;
        RECT 18.030000  26.770000 18.230000  26.970000 ;
        RECT 18.030000  27.200000 18.230000  27.400000 ;
        RECT 18.030000  27.630000 18.230000  27.830000 ;
        RECT 18.030000  28.060000 18.230000  28.260000 ;
        RECT 18.030000  28.490000 18.230000  28.690000 ;
        RECT 18.030000  28.920000 18.230000  29.120000 ;
        RECT 18.030000  29.350000 18.230000  29.550000 ;
        RECT 18.030000  29.780000 18.230000  29.980000 ;
        RECT 18.030000  30.210000 18.230000  30.410000 ;
        RECT 18.150000 197.250000 18.350000 197.450000 ;
        RECT 18.150000 197.650000 18.350000 197.850000 ;
        RECT 18.150000 198.050000 18.350000 198.250000 ;
        RECT 18.150000 198.450000 18.350000 198.650000 ;
        RECT 18.150000 198.850000 18.350000 199.050000 ;
        RECT 18.150000 199.250000 18.350000 199.450000 ;
        RECT 18.150000 199.650000 18.350000 199.850000 ;
        RECT 18.435000  25.910000 18.635000  26.110000 ;
        RECT 18.435000  26.340000 18.635000  26.540000 ;
        RECT 18.435000  26.770000 18.635000  26.970000 ;
        RECT 18.435000  27.200000 18.635000  27.400000 ;
        RECT 18.435000  27.630000 18.635000  27.830000 ;
        RECT 18.435000  28.060000 18.635000  28.260000 ;
        RECT 18.435000  28.490000 18.635000  28.690000 ;
        RECT 18.435000  28.920000 18.635000  29.120000 ;
        RECT 18.435000  29.350000 18.635000  29.550000 ;
        RECT 18.435000  29.780000 18.635000  29.980000 ;
        RECT 18.435000  30.210000 18.635000  30.410000 ;
        RECT 18.555000 197.250000 18.755000 197.450000 ;
        RECT 18.555000 197.650000 18.755000 197.850000 ;
        RECT 18.555000 198.050000 18.755000 198.250000 ;
        RECT 18.555000 198.450000 18.755000 198.650000 ;
        RECT 18.555000 198.850000 18.755000 199.050000 ;
        RECT 18.555000 199.250000 18.755000 199.450000 ;
        RECT 18.555000 199.650000 18.755000 199.850000 ;
        RECT 18.840000  25.910000 19.040000  26.110000 ;
        RECT 18.840000  26.340000 19.040000  26.540000 ;
        RECT 18.840000  26.770000 19.040000  26.970000 ;
        RECT 18.840000  27.200000 19.040000  27.400000 ;
        RECT 18.840000  27.630000 19.040000  27.830000 ;
        RECT 18.840000  28.060000 19.040000  28.260000 ;
        RECT 18.840000  28.490000 19.040000  28.690000 ;
        RECT 18.840000  28.920000 19.040000  29.120000 ;
        RECT 18.840000  29.350000 19.040000  29.550000 ;
        RECT 18.840000  29.780000 19.040000  29.980000 ;
        RECT 18.840000  30.210000 19.040000  30.410000 ;
        RECT 18.960000 197.250000 19.160000 197.450000 ;
        RECT 18.960000 197.650000 19.160000 197.850000 ;
        RECT 18.960000 198.050000 19.160000 198.250000 ;
        RECT 18.960000 198.450000 19.160000 198.650000 ;
        RECT 18.960000 198.850000 19.160000 199.050000 ;
        RECT 18.960000 199.250000 19.160000 199.450000 ;
        RECT 18.960000 199.650000 19.160000 199.850000 ;
        RECT 19.245000  25.910000 19.445000  26.110000 ;
        RECT 19.245000  26.340000 19.445000  26.540000 ;
        RECT 19.245000  26.770000 19.445000  26.970000 ;
        RECT 19.245000  27.200000 19.445000  27.400000 ;
        RECT 19.245000  27.630000 19.445000  27.830000 ;
        RECT 19.245000  28.060000 19.445000  28.260000 ;
        RECT 19.245000  28.490000 19.445000  28.690000 ;
        RECT 19.245000  28.920000 19.445000  29.120000 ;
        RECT 19.245000  29.350000 19.445000  29.550000 ;
        RECT 19.245000  29.780000 19.445000  29.980000 ;
        RECT 19.245000  30.210000 19.445000  30.410000 ;
        RECT 19.365000 197.250000 19.565000 197.450000 ;
        RECT 19.365000 197.650000 19.565000 197.850000 ;
        RECT 19.365000 198.050000 19.565000 198.250000 ;
        RECT 19.365000 198.450000 19.565000 198.650000 ;
        RECT 19.365000 198.850000 19.565000 199.050000 ;
        RECT 19.365000 199.250000 19.565000 199.450000 ;
        RECT 19.365000 199.650000 19.565000 199.850000 ;
        RECT 19.650000  25.910000 19.850000  26.110000 ;
        RECT 19.650000  26.340000 19.850000  26.540000 ;
        RECT 19.650000  26.770000 19.850000  26.970000 ;
        RECT 19.650000  27.200000 19.850000  27.400000 ;
        RECT 19.650000  27.630000 19.850000  27.830000 ;
        RECT 19.650000  28.060000 19.850000  28.260000 ;
        RECT 19.650000  28.490000 19.850000  28.690000 ;
        RECT 19.650000  28.920000 19.850000  29.120000 ;
        RECT 19.650000  29.350000 19.850000  29.550000 ;
        RECT 19.650000  29.780000 19.850000  29.980000 ;
        RECT 19.650000  30.210000 19.850000  30.410000 ;
        RECT 19.770000 197.250000 19.970000 197.450000 ;
        RECT 19.770000 197.650000 19.970000 197.850000 ;
        RECT 19.770000 198.050000 19.970000 198.250000 ;
        RECT 19.770000 198.450000 19.970000 198.650000 ;
        RECT 19.770000 198.850000 19.970000 199.050000 ;
        RECT 19.770000 199.250000 19.970000 199.450000 ;
        RECT 19.770000 199.650000 19.970000 199.850000 ;
        RECT 20.055000  25.910000 20.255000  26.110000 ;
        RECT 20.055000  26.340000 20.255000  26.540000 ;
        RECT 20.055000  26.770000 20.255000  26.970000 ;
        RECT 20.055000  27.200000 20.255000  27.400000 ;
        RECT 20.055000  27.630000 20.255000  27.830000 ;
        RECT 20.055000  28.060000 20.255000  28.260000 ;
        RECT 20.055000  28.490000 20.255000  28.690000 ;
        RECT 20.055000  28.920000 20.255000  29.120000 ;
        RECT 20.055000  29.350000 20.255000  29.550000 ;
        RECT 20.055000  29.780000 20.255000  29.980000 ;
        RECT 20.055000  30.210000 20.255000  30.410000 ;
        RECT 20.175000 197.250000 20.375000 197.450000 ;
        RECT 20.175000 197.650000 20.375000 197.850000 ;
        RECT 20.175000 198.050000 20.375000 198.250000 ;
        RECT 20.175000 198.450000 20.375000 198.650000 ;
        RECT 20.175000 198.850000 20.375000 199.050000 ;
        RECT 20.175000 199.250000 20.375000 199.450000 ;
        RECT 20.175000 199.650000 20.375000 199.850000 ;
        RECT 20.460000  25.910000 20.660000  26.110000 ;
        RECT 20.460000  26.340000 20.660000  26.540000 ;
        RECT 20.460000  26.770000 20.660000  26.970000 ;
        RECT 20.460000  27.200000 20.660000  27.400000 ;
        RECT 20.460000  27.630000 20.660000  27.830000 ;
        RECT 20.460000  28.060000 20.660000  28.260000 ;
        RECT 20.460000  28.490000 20.660000  28.690000 ;
        RECT 20.460000  28.920000 20.660000  29.120000 ;
        RECT 20.460000  29.350000 20.660000  29.550000 ;
        RECT 20.460000  29.780000 20.660000  29.980000 ;
        RECT 20.460000  30.210000 20.660000  30.410000 ;
        RECT 20.580000 197.250000 20.780000 197.450000 ;
        RECT 20.580000 197.650000 20.780000 197.850000 ;
        RECT 20.580000 198.050000 20.780000 198.250000 ;
        RECT 20.580000 198.450000 20.780000 198.650000 ;
        RECT 20.580000 198.850000 20.780000 199.050000 ;
        RECT 20.580000 199.250000 20.780000 199.450000 ;
        RECT 20.580000 199.650000 20.780000 199.850000 ;
        RECT 20.865000  25.910000 21.065000  26.110000 ;
        RECT 20.865000  26.340000 21.065000  26.540000 ;
        RECT 20.865000  26.770000 21.065000  26.970000 ;
        RECT 20.865000  27.200000 21.065000  27.400000 ;
        RECT 20.865000  27.630000 21.065000  27.830000 ;
        RECT 20.865000  28.060000 21.065000  28.260000 ;
        RECT 20.865000  28.490000 21.065000  28.690000 ;
        RECT 20.865000  28.920000 21.065000  29.120000 ;
        RECT 20.865000  29.350000 21.065000  29.550000 ;
        RECT 20.865000  29.780000 21.065000  29.980000 ;
        RECT 20.865000  30.210000 21.065000  30.410000 ;
        RECT 20.985000 197.250000 21.185000 197.450000 ;
        RECT 20.985000 197.650000 21.185000 197.850000 ;
        RECT 20.985000 198.050000 21.185000 198.250000 ;
        RECT 20.985000 198.450000 21.185000 198.650000 ;
        RECT 20.985000 198.850000 21.185000 199.050000 ;
        RECT 20.985000 199.250000 21.185000 199.450000 ;
        RECT 20.985000 199.650000 21.185000 199.850000 ;
        RECT 21.270000  25.910000 21.470000  26.110000 ;
        RECT 21.270000  26.340000 21.470000  26.540000 ;
        RECT 21.270000  26.770000 21.470000  26.970000 ;
        RECT 21.270000  27.200000 21.470000  27.400000 ;
        RECT 21.270000  27.630000 21.470000  27.830000 ;
        RECT 21.270000  28.060000 21.470000  28.260000 ;
        RECT 21.270000  28.490000 21.470000  28.690000 ;
        RECT 21.270000  28.920000 21.470000  29.120000 ;
        RECT 21.270000  29.350000 21.470000  29.550000 ;
        RECT 21.270000  29.780000 21.470000  29.980000 ;
        RECT 21.270000  30.210000 21.470000  30.410000 ;
        RECT 21.390000 197.250000 21.590000 197.450000 ;
        RECT 21.390000 197.650000 21.590000 197.850000 ;
        RECT 21.390000 198.050000 21.590000 198.250000 ;
        RECT 21.390000 198.450000 21.590000 198.650000 ;
        RECT 21.390000 198.850000 21.590000 199.050000 ;
        RECT 21.390000 199.250000 21.590000 199.450000 ;
        RECT 21.390000 199.650000 21.590000 199.850000 ;
        RECT 21.675000  25.910000 21.875000  26.110000 ;
        RECT 21.675000  26.340000 21.875000  26.540000 ;
        RECT 21.675000  26.770000 21.875000  26.970000 ;
        RECT 21.675000  27.200000 21.875000  27.400000 ;
        RECT 21.675000  27.630000 21.875000  27.830000 ;
        RECT 21.675000  28.060000 21.875000  28.260000 ;
        RECT 21.675000  28.490000 21.875000  28.690000 ;
        RECT 21.675000  28.920000 21.875000  29.120000 ;
        RECT 21.675000  29.350000 21.875000  29.550000 ;
        RECT 21.675000  29.780000 21.875000  29.980000 ;
        RECT 21.675000  30.210000 21.875000  30.410000 ;
        RECT 21.795000 197.250000 21.995000 197.450000 ;
        RECT 21.795000 197.650000 21.995000 197.850000 ;
        RECT 21.795000 198.050000 21.995000 198.250000 ;
        RECT 21.795000 198.450000 21.995000 198.650000 ;
        RECT 21.795000 198.850000 21.995000 199.050000 ;
        RECT 21.795000 199.250000 21.995000 199.450000 ;
        RECT 21.795000 199.650000 21.995000 199.850000 ;
        RECT 22.080000  25.910000 22.280000  26.110000 ;
        RECT 22.080000  26.340000 22.280000  26.540000 ;
        RECT 22.080000  26.770000 22.280000  26.970000 ;
        RECT 22.080000  27.200000 22.280000  27.400000 ;
        RECT 22.080000  27.630000 22.280000  27.830000 ;
        RECT 22.080000  28.060000 22.280000  28.260000 ;
        RECT 22.080000  28.490000 22.280000  28.690000 ;
        RECT 22.080000  28.920000 22.280000  29.120000 ;
        RECT 22.080000  29.350000 22.280000  29.550000 ;
        RECT 22.080000  29.780000 22.280000  29.980000 ;
        RECT 22.080000  30.210000 22.280000  30.410000 ;
        RECT 22.200000 197.250000 22.400000 197.450000 ;
        RECT 22.200000 197.650000 22.400000 197.850000 ;
        RECT 22.200000 198.050000 22.400000 198.250000 ;
        RECT 22.200000 198.450000 22.400000 198.650000 ;
        RECT 22.200000 198.850000 22.400000 199.050000 ;
        RECT 22.200000 199.250000 22.400000 199.450000 ;
        RECT 22.200000 199.650000 22.400000 199.850000 ;
        RECT 22.485000  25.910000 22.685000  26.110000 ;
        RECT 22.485000  26.340000 22.685000  26.540000 ;
        RECT 22.485000  26.770000 22.685000  26.970000 ;
        RECT 22.485000  27.200000 22.685000  27.400000 ;
        RECT 22.485000  27.630000 22.685000  27.830000 ;
        RECT 22.485000  28.060000 22.685000  28.260000 ;
        RECT 22.485000  28.490000 22.685000  28.690000 ;
        RECT 22.485000  28.920000 22.685000  29.120000 ;
        RECT 22.485000  29.350000 22.685000  29.550000 ;
        RECT 22.485000  29.780000 22.685000  29.980000 ;
        RECT 22.485000  30.210000 22.685000  30.410000 ;
        RECT 22.605000 197.250000 22.805000 197.450000 ;
        RECT 22.605000 197.650000 22.805000 197.850000 ;
        RECT 22.605000 198.050000 22.805000 198.250000 ;
        RECT 22.605000 198.450000 22.805000 198.650000 ;
        RECT 22.605000 198.850000 22.805000 199.050000 ;
        RECT 22.605000 199.250000 22.805000 199.450000 ;
        RECT 22.605000 199.650000 22.805000 199.850000 ;
        RECT 22.890000  25.910000 23.090000  26.110000 ;
        RECT 22.890000  26.340000 23.090000  26.540000 ;
        RECT 22.890000  26.770000 23.090000  26.970000 ;
        RECT 22.890000  27.200000 23.090000  27.400000 ;
        RECT 22.890000  27.630000 23.090000  27.830000 ;
        RECT 22.890000  28.060000 23.090000  28.260000 ;
        RECT 22.890000  28.490000 23.090000  28.690000 ;
        RECT 22.890000  28.920000 23.090000  29.120000 ;
        RECT 22.890000  29.350000 23.090000  29.550000 ;
        RECT 22.890000  29.780000 23.090000  29.980000 ;
        RECT 22.890000  30.210000 23.090000  30.410000 ;
        RECT 23.010000 197.250000 23.210000 197.450000 ;
        RECT 23.010000 197.650000 23.210000 197.850000 ;
        RECT 23.010000 198.050000 23.210000 198.250000 ;
        RECT 23.010000 198.450000 23.210000 198.650000 ;
        RECT 23.010000 198.850000 23.210000 199.050000 ;
        RECT 23.010000 199.250000 23.210000 199.450000 ;
        RECT 23.010000 199.650000 23.210000 199.850000 ;
        RECT 23.295000  25.910000 23.495000  26.110000 ;
        RECT 23.295000  26.340000 23.495000  26.540000 ;
        RECT 23.295000  26.770000 23.495000  26.970000 ;
        RECT 23.295000  27.200000 23.495000  27.400000 ;
        RECT 23.295000  27.630000 23.495000  27.830000 ;
        RECT 23.295000  28.060000 23.495000  28.260000 ;
        RECT 23.295000  28.490000 23.495000  28.690000 ;
        RECT 23.295000  28.920000 23.495000  29.120000 ;
        RECT 23.295000  29.350000 23.495000  29.550000 ;
        RECT 23.295000  29.780000 23.495000  29.980000 ;
        RECT 23.295000  30.210000 23.495000  30.410000 ;
        RECT 23.415000 197.250000 23.615000 197.450000 ;
        RECT 23.415000 197.650000 23.615000 197.850000 ;
        RECT 23.415000 198.050000 23.615000 198.250000 ;
        RECT 23.415000 198.450000 23.615000 198.650000 ;
        RECT 23.415000 198.850000 23.615000 199.050000 ;
        RECT 23.415000 199.250000 23.615000 199.450000 ;
        RECT 23.415000 199.650000 23.615000 199.850000 ;
        RECT 23.700000  25.910000 23.900000  26.110000 ;
        RECT 23.700000  26.340000 23.900000  26.540000 ;
        RECT 23.700000  26.770000 23.900000  26.970000 ;
        RECT 23.700000  27.200000 23.900000  27.400000 ;
        RECT 23.700000  27.630000 23.900000  27.830000 ;
        RECT 23.700000  28.060000 23.900000  28.260000 ;
        RECT 23.700000  28.490000 23.900000  28.690000 ;
        RECT 23.700000  28.920000 23.900000  29.120000 ;
        RECT 23.700000  29.350000 23.900000  29.550000 ;
        RECT 23.700000  29.780000 23.900000  29.980000 ;
        RECT 23.700000  30.210000 23.900000  30.410000 ;
        RECT 23.820000 197.250000 24.020000 197.450000 ;
        RECT 23.820000 197.650000 24.020000 197.850000 ;
        RECT 23.820000 198.050000 24.020000 198.250000 ;
        RECT 23.820000 198.450000 24.020000 198.650000 ;
        RECT 23.820000 198.850000 24.020000 199.050000 ;
        RECT 23.820000 199.250000 24.020000 199.450000 ;
        RECT 23.820000 199.650000 24.020000 199.850000 ;
        RECT 24.105000  25.910000 24.305000  26.110000 ;
        RECT 24.105000  26.340000 24.305000  26.540000 ;
        RECT 24.105000  26.770000 24.305000  26.970000 ;
        RECT 24.105000  27.200000 24.305000  27.400000 ;
        RECT 24.105000  27.630000 24.305000  27.830000 ;
        RECT 24.105000  28.060000 24.305000  28.260000 ;
        RECT 24.105000  28.490000 24.305000  28.690000 ;
        RECT 24.105000  28.920000 24.305000  29.120000 ;
        RECT 24.105000  29.350000 24.305000  29.550000 ;
        RECT 24.105000  29.780000 24.305000  29.980000 ;
        RECT 24.105000  30.210000 24.305000  30.410000 ;
        RECT 24.225000 197.250000 24.425000 197.450000 ;
        RECT 24.225000 197.650000 24.425000 197.850000 ;
        RECT 24.225000 198.050000 24.425000 198.250000 ;
        RECT 24.225000 198.450000 24.425000 198.650000 ;
        RECT 24.225000 198.850000 24.425000 199.050000 ;
        RECT 24.225000 199.250000 24.425000 199.450000 ;
        RECT 24.225000 199.650000 24.425000 199.850000 ;
        RECT 24.630000 197.250000 24.830000 197.450000 ;
        RECT 24.630000 197.650000 24.830000 197.850000 ;
        RECT 24.630000 198.050000 24.830000 198.250000 ;
        RECT 24.630000 198.450000 24.830000 198.650000 ;
        RECT 24.630000 198.850000 24.830000 199.050000 ;
        RECT 24.630000 199.250000 24.830000 199.450000 ;
        RECT 24.630000 199.650000 24.830000 199.850000 ;
        RECT 25.035000 197.250000 25.235000 197.450000 ;
        RECT 25.035000 197.650000 25.235000 197.850000 ;
        RECT 25.035000 198.050000 25.235000 198.250000 ;
        RECT 25.035000 198.450000 25.235000 198.650000 ;
        RECT 25.035000 198.850000 25.235000 199.050000 ;
        RECT 25.035000 199.250000 25.235000 199.450000 ;
        RECT 25.035000 199.650000 25.235000 199.850000 ;
        RECT 25.440000 197.250000 25.640000 197.450000 ;
        RECT 25.440000 197.650000 25.640000 197.850000 ;
        RECT 25.440000 198.050000 25.640000 198.250000 ;
        RECT 25.440000 198.450000 25.640000 198.650000 ;
        RECT 25.440000 198.850000 25.640000 199.050000 ;
        RECT 25.440000 199.250000 25.640000 199.450000 ;
        RECT 25.440000 199.650000 25.640000 199.850000 ;
        RECT 25.845000 197.250000 26.045000 197.450000 ;
        RECT 25.845000 197.650000 26.045000 197.850000 ;
        RECT 25.845000 198.050000 26.045000 198.250000 ;
        RECT 25.845000 198.450000 26.045000 198.650000 ;
        RECT 25.845000 198.850000 26.045000 199.050000 ;
        RECT 25.845000 199.250000 26.045000 199.450000 ;
        RECT 25.845000 199.650000 26.045000 199.850000 ;
        RECT 26.250000 197.250000 26.450000 197.450000 ;
        RECT 26.250000 197.650000 26.450000 197.850000 ;
        RECT 26.250000 198.050000 26.450000 198.250000 ;
        RECT 26.250000 198.450000 26.450000 198.650000 ;
        RECT 26.250000 198.850000 26.450000 199.050000 ;
        RECT 26.250000 199.250000 26.450000 199.450000 ;
        RECT 26.250000 199.650000 26.450000 199.850000 ;
        RECT 26.655000 197.250000 26.855000 197.450000 ;
        RECT 26.655000 197.650000 26.855000 197.850000 ;
        RECT 26.655000 198.050000 26.855000 198.250000 ;
        RECT 26.655000 198.450000 26.855000 198.650000 ;
        RECT 26.655000 198.850000 26.855000 199.050000 ;
        RECT 26.655000 199.250000 26.855000 199.450000 ;
        RECT 26.655000 199.650000 26.855000 199.850000 ;
        RECT 27.060000 197.250000 27.260000 197.450000 ;
        RECT 27.060000 197.650000 27.260000 197.850000 ;
        RECT 27.060000 198.050000 27.260000 198.250000 ;
        RECT 27.060000 198.450000 27.260000 198.650000 ;
        RECT 27.060000 198.850000 27.260000 199.050000 ;
        RECT 27.060000 199.250000 27.260000 199.450000 ;
        RECT 27.060000 199.650000 27.260000 199.850000 ;
        RECT 27.460000 197.250000 27.660000 197.450000 ;
        RECT 27.460000 197.650000 27.660000 197.850000 ;
        RECT 27.460000 198.050000 27.660000 198.250000 ;
        RECT 27.460000 198.450000 27.660000 198.650000 ;
        RECT 27.460000 198.850000 27.660000 199.050000 ;
        RECT 27.460000 199.250000 27.660000 199.450000 ;
        RECT 27.460000 199.650000 27.660000 199.850000 ;
        RECT 27.860000 197.250000 28.060000 197.450000 ;
        RECT 27.860000 197.650000 28.060000 197.850000 ;
        RECT 27.860000 198.050000 28.060000 198.250000 ;
        RECT 27.860000 198.450000 28.060000 198.650000 ;
        RECT 27.860000 198.850000 28.060000 199.050000 ;
        RECT 27.860000 199.250000 28.060000 199.450000 ;
        RECT 27.860000 199.650000 28.060000 199.850000 ;
        RECT 28.260000 197.250000 28.460000 197.450000 ;
        RECT 28.260000 197.650000 28.460000 197.850000 ;
        RECT 28.260000 198.050000 28.460000 198.250000 ;
        RECT 28.260000 198.450000 28.460000 198.650000 ;
        RECT 28.260000 198.850000 28.460000 199.050000 ;
        RECT 28.260000 199.250000 28.460000 199.450000 ;
        RECT 28.260000 199.650000 28.460000 199.850000 ;
        RECT 28.660000 197.250000 28.860000 197.450000 ;
        RECT 28.660000 197.650000 28.860000 197.850000 ;
        RECT 28.660000 198.050000 28.860000 198.250000 ;
        RECT 28.660000 198.450000 28.860000 198.650000 ;
        RECT 28.660000 198.850000 28.860000 199.050000 ;
        RECT 28.660000 199.250000 28.860000 199.450000 ;
        RECT 28.660000 199.650000 28.860000 199.850000 ;
        RECT 29.060000 197.250000 29.260000 197.450000 ;
        RECT 29.060000 197.650000 29.260000 197.850000 ;
        RECT 29.060000 198.050000 29.260000 198.250000 ;
        RECT 29.060000 198.450000 29.260000 198.650000 ;
        RECT 29.060000 198.850000 29.260000 199.050000 ;
        RECT 29.060000 199.250000 29.260000 199.450000 ;
        RECT 29.060000 199.650000 29.260000 199.850000 ;
        RECT 29.460000 197.250000 29.660000 197.450000 ;
        RECT 29.460000 197.650000 29.660000 197.850000 ;
        RECT 29.460000 198.050000 29.660000 198.250000 ;
        RECT 29.460000 198.450000 29.660000 198.650000 ;
        RECT 29.460000 198.850000 29.660000 199.050000 ;
        RECT 29.460000 199.250000 29.660000 199.450000 ;
        RECT 29.460000 199.650000 29.660000 199.850000 ;
        RECT 29.860000 197.250000 30.060000 197.450000 ;
        RECT 29.860000 197.650000 30.060000 197.850000 ;
        RECT 29.860000 198.050000 30.060000 198.250000 ;
        RECT 29.860000 198.450000 30.060000 198.650000 ;
        RECT 29.860000 198.850000 30.060000 199.050000 ;
        RECT 29.860000 199.250000 30.060000 199.450000 ;
        RECT 29.860000 199.650000 30.060000 199.850000 ;
        RECT 30.260000 197.250000 30.460000 197.450000 ;
        RECT 30.260000 197.650000 30.460000 197.850000 ;
        RECT 30.260000 198.050000 30.460000 198.250000 ;
        RECT 30.260000 198.450000 30.460000 198.650000 ;
        RECT 30.260000 198.850000 30.460000 199.050000 ;
        RECT 30.260000 199.250000 30.460000 199.450000 ;
        RECT 30.260000 199.650000 30.460000 199.850000 ;
        RECT 30.660000 197.250000 30.860000 197.450000 ;
        RECT 30.660000 197.650000 30.860000 197.850000 ;
        RECT 30.660000 198.050000 30.860000 198.250000 ;
        RECT 30.660000 198.450000 30.860000 198.650000 ;
        RECT 30.660000 198.850000 30.860000 199.050000 ;
        RECT 30.660000 199.250000 30.860000 199.450000 ;
        RECT 30.660000 199.650000 30.860000 199.850000 ;
        RECT 31.060000 197.250000 31.260000 197.450000 ;
        RECT 31.060000 197.650000 31.260000 197.850000 ;
        RECT 31.060000 198.050000 31.260000 198.250000 ;
        RECT 31.060000 198.450000 31.260000 198.650000 ;
        RECT 31.060000 198.850000 31.260000 199.050000 ;
        RECT 31.060000 199.250000 31.260000 199.450000 ;
        RECT 31.060000 199.650000 31.260000 199.850000 ;
        RECT 31.460000 197.250000 31.660000 197.450000 ;
        RECT 31.460000 197.650000 31.660000 197.850000 ;
        RECT 31.460000 198.050000 31.660000 198.250000 ;
        RECT 31.460000 198.450000 31.660000 198.650000 ;
        RECT 31.460000 198.850000 31.660000 199.050000 ;
        RECT 31.460000 199.250000 31.660000 199.450000 ;
        RECT 31.460000 199.650000 31.660000 199.850000 ;
        RECT 31.860000 197.250000 32.060000 197.450000 ;
        RECT 31.860000 197.650000 32.060000 197.850000 ;
        RECT 31.860000 198.050000 32.060000 198.250000 ;
        RECT 31.860000 198.450000 32.060000 198.650000 ;
        RECT 31.860000 198.850000 32.060000 199.050000 ;
        RECT 31.860000 199.250000 32.060000 199.450000 ;
        RECT 31.860000 199.650000 32.060000 199.850000 ;
        RECT 32.260000 197.250000 32.460000 197.450000 ;
        RECT 32.260000 197.650000 32.460000 197.850000 ;
        RECT 32.260000 198.050000 32.460000 198.250000 ;
        RECT 32.260000 198.450000 32.460000 198.650000 ;
        RECT 32.260000 198.850000 32.460000 199.050000 ;
        RECT 32.260000 199.250000 32.460000 199.450000 ;
        RECT 32.260000 199.650000 32.460000 199.850000 ;
        RECT 32.660000 197.250000 32.860000 197.450000 ;
        RECT 32.660000 197.650000 32.860000 197.850000 ;
        RECT 32.660000 198.050000 32.860000 198.250000 ;
        RECT 32.660000 198.450000 32.860000 198.650000 ;
        RECT 32.660000 198.850000 32.860000 199.050000 ;
        RECT 32.660000 199.250000 32.860000 199.450000 ;
        RECT 32.660000 199.650000 32.860000 199.850000 ;
        RECT 33.060000 197.250000 33.260000 197.450000 ;
        RECT 33.060000 197.650000 33.260000 197.850000 ;
        RECT 33.060000 198.050000 33.260000 198.250000 ;
        RECT 33.060000 198.450000 33.260000 198.650000 ;
        RECT 33.060000 198.850000 33.260000 199.050000 ;
        RECT 33.060000 199.250000 33.260000 199.450000 ;
        RECT 33.060000 199.650000 33.260000 199.850000 ;
        RECT 33.460000 197.250000 33.660000 197.450000 ;
        RECT 33.460000 197.650000 33.660000 197.850000 ;
        RECT 33.460000 198.050000 33.660000 198.250000 ;
        RECT 33.460000 198.450000 33.660000 198.650000 ;
        RECT 33.460000 198.850000 33.660000 199.050000 ;
        RECT 33.460000 199.250000 33.660000 199.450000 ;
        RECT 33.460000 199.650000 33.660000 199.850000 ;
        RECT 33.860000 197.250000 34.060000 197.450000 ;
        RECT 33.860000 197.650000 34.060000 197.850000 ;
        RECT 33.860000 198.050000 34.060000 198.250000 ;
        RECT 33.860000 198.450000 34.060000 198.650000 ;
        RECT 33.860000 198.850000 34.060000 199.050000 ;
        RECT 33.860000 199.250000 34.060000 199.450000 ;
        RECT 33.860000 199.650000 34.060000 199.850000 ;
        RECT 34.260000 197.250000 34.460000 197.450000 ;
        RECT 34.260000 197.650000 34.460000 197.850000 ;
        RECT 34.260000 198.050000 34.460000 198.250000 ;
        RECT 34.260000 198.450000 34.460000 198.650000 ;
        RECT 34.260000 198.850000 34.460000 199.050000 ;
        RECT 34.260000 199.250000 34.460000 199.450000 ;
        RECT 34.260000 199.650000 34.460000 199.850000 ;
        RECT 34.660000 197.250000 34.860000 197.450000 ;
        RECT 34.660000 197.650000 34.860000 197.850000 ;
        RECT 34.660000 198.050000 34.860000 198.250000 ;
        RECT 34.660000 198.450000 34.860000 198.650000 ;
        RECT 34.660000 198.850000 34.860000 199.050000 ;
        RECT 34.660000 199.250000 34.860000 199.450000 ;
        RECT 34.660000 199.650000 34.860000 199.850000 ;
        RECT 35.060000 197.250000 35.260000 197.450000 ;
        RECT 35.060000 197.650000 35.260000 197.850000 ;
        RECT 35.060000 198.050000 35.260000 198.250000 ;
        RECT 35.060000 198.450000 35.260000 198.650000 ;
        RECT 35.060000 198.850000 35.260000 199.050000 ;
        RECT 35.060000 199.250000 35.260000 199.450000 ;
        RECT 35.060000 199.650000 35.260000 199.850000 ;
        RECT 35.460000 197.250000 35.660000 197.450000 ;
        RECT 35.460000 197.650000 35.660000 197.850000 ;
        RECT 35.460000 198.050000 35.660000 198.250000 ;
        RECT 35.460000 198.450000 35.660000 198.650000 ;
        RECT 35.460000 198.850000 35.660000 199.050000 ;
        RECT 35.460000 199.250000 35.660000 199.450000 ;
        RECT 35.460000 199.650000 35.660000 199.850000 ;
        RECT 35.860000 197.250000 36.060000 197.450000 ;
        RECT 35.860000 197.650000 36.060000 197.850000 ;
        RECT 35.860000 198.050000 36.060000 198.250000 ;
        RECT 35.860000 198.450000 36.060000 198.650000 ;
        RECT 35.860000 198.850000 36.060000 199.050000 ;
        RECT 35.860000 199.250000 36.060000 199.450000 ;
        RECT 35.860000 199.650000 36.060000 199.850000 ;
        RECT 36.260000 197.250000 36.460000 197.450000 ;
        RECT 36.260000 197.650000 36.460000 197.850000 ;
        RECT 36.260000 198.050000 36.460000 198.250000 ;
        RECT 36.260000 198.450000 36.460000 198.650000 ;
        RECT 36.260000 198.850000 36.460000 199.050000 ;
        RECT 36.260000 199.250000 36.460000 199.450000 ;
        RECT 36.260000 199.650000 36.460000 199.850000 ;
        RECT 36.660000 197.250000 36.860000 197.450000 ;
        RECT 36.660000 197.650000 36.860000 197.850000 ;
        RECT 36.660000 198.050000 36.860000 198.250000 ;
        RECT 36.660000 198.450000 36.860000 198.650000 ;
        RECT 36.660000 198.850000 36.860000 199.050000 ;
        RECT 36.660000 199.250000 36.860000 199.450000 ;
        RECT 36.660000 199.650000 36.860000 199.850000 ;
        RECT 37.060000 197.250000 37.260000 197.450000 ;
        RECT 37.060000 197.650000 37.260000 197.850000 ;
        RECT 37.060000 198.050000 37.260000 198.250000 ;
        RECT 37.060000 198.450000 37.260000 198.650000 ;
        RECT 37.060000 198.850000 37.260000 199.050000 ;
        RECT 37.060000 199.250000 37.260000 199.450000 ;
        RECT 37.060000 199.650000 37.260000 199.850000 ;
        RECT 37.460000 197.250000 37.660000 197.450000 ;
        RECT 37.460000 197.650000 37.660000 197.850000 ;
        RECT 37.460000 198.050000 37.660000 198.250000 ;
        RECT 37.460000 198.450000 37.660000 198.650000 ;
        RECT 37.460000 198.850000 37.660000 199.050000 ;
        RECT 37.460000 199.250000 37.660000 199.450000 ;
        RECT 37.460000 199.650000 37.660000 199.850000 ;
        RECT 37.860000 197.250000 38.060000 197.450000 ;
        RECT 37.860000 197.650000 38.060000 197.850000 ;
        RECT 37.860000 198.050000 38.060000 198.250000 ;
        RECT 37.860000 198.450000 38.060000 198.650000 ;
        RECT 37.860000 198.850000 38.060000 199.050000 ;
        RECT 37.860000 199.250000 38.060000 199.450000 ;
        RECT 37.860000 199.650000 38.060000 199.850000 ;
        RECT 38.260000 197.250000 38.460000 197.450000 ;
        RECT 38.260000 197.650000 38.460000 197.850000 ;
        RECT 38.260000 198.050000 38.460000 198.250000 ;
        RECT 38.260000 198.450000 38.460000 198.650000 ;
        RECT 38.260000 198.850000 38.460000 199.050000 ;
        RECT 38.260000 199.250000 38.460000 199.450000 ;
        RECT 38.260000 199.650000 38.460000 199.850000 ;
        RECT 38.660000 197.250000 38.860000 197.450000 ;
        RECT 38.660000 197.650000 38.860000 197.850000 ;
        RECT 38.660000 198.050000 38.860000 198.250000 ;
        RECT 38.660000 198.450000 38.860000 198.650000 ;
        RECT 38.660000 198.850000 38.860000 199.050000 ;
        RECT 38.660000 199.250000 38.860000 199.450000 ;
        RECT 38.660000 199.650000 38.860000 199.850000 ;
        RECT 39.060000 197.250000 39.260000 197.450000 ;
        RECT 39.060000 197.650000 39.260000 197.850000 ;
        RECT 39.060000 198.050000 39.260000 198.250000 ;
        RECT 39.060000 198.450000 39.260000 198.650000 ;
        RECT 39.060000 198.850000 39.260000 199.050000 ;
        RECT 39.060000 199.250000 39.260000 199.450000 ;
        RECT 39.060000 199.650000 39.260000 199.850000 ;
        RECT 39.460000 197.250000 39.660000 197.450000 ;
        RECT 39.460000 197.650000 39.660000 197.850000 ;
        RECT 39.460000 198.050000 39.660000 198.250000 ;
        RECT 39.460000 198.450000 39.660000 198.650000 ;
        RECT 39.460000 198.850000 39.660000 199.050000 ;
        RECT 39.460000 199.250000 39.660000 199.450000 ;
        RECT 39.460000 199.650000 39.660000 199.850000 ;
        RECT 39.860000 197.250000 40.060000 197.450000 ;
        RECT 39.860000 197.650000 40.060000 197.850000 ;
        RECT 39.860000 198.050000 40.060000 198.250000 ;
        RECT 39.860000 198.450000 40.060000 198.650000 ;
        RECT 39.860000 198.850000 40.060000 199.050000 ;
        RECT 39.860000 199.250000 40.060000 199.450000 ;
        RECT 39.860000 199.650000 40.060000 199.850000 ;
        RECT 40.260000 197.250000 40.460000 197.450000 ;
        RECT 40.260000 197.650000 40.460000 197.850000 ;
        RECT 40.260000 198.050000 40.460000 198.250000 ;
        RECT 40.260000 198.450000 40.460000 198.650000 ;
        RECT 40.260000 198.850000 40.460000 199.050000 ;
        RECT 40.260000 199.250000 40.460000 199.450000 ;
        RECT 40.260000 199.650000 40.460000 199.850000 ;
        RECT 40.660000 197.250000 40.860000 197.450000 ;
        RECT 40.660000 197.650000 40.860000 197.850000 ;
        RECT 40.660000 198.050000 40.860000 198.250000 ;
        RECT 40.660000 198.450000 40.860000 198.650000 ;
        RECT 40.660000 198.850000 40.860000 199.050000 ;
        RECT 40.660000 199.250000 40.860000 199.450000 ;
        RECT 40.660000 199.650000 40.860000 199.850000 ;
        RECT 41.060000 197.250000 41.260000 197.450000 ;
        RECT 41.060000 197.650000 41.260000 197.850000 ;
        RECT 41.060000 198.050000 41.260000 198.250000 ;
        RECT 41.060000 198.450000 41.260000 198.650000 ;
        RECT 41.060000 198.850000 41.260000 199.050000 ;
        RECT 41.060000 199.250000 41.260000 199.450000 ;
        RECT 41.060000 199.650000 41.260000 199.850000 ;
        RECT 41.460000 197.250000 41.660000 197.450000 ;
        RECT 41.460000 197.650000 41.660000 197.850000 ;
        RECT 41.460000 198.050000 41.660000 198.250000 ;
        RECT 41.460000 198.450000 41.660000 198.650000 ;
        RECT 41.460000 198.850000 41.660000 199.050000 ;
        RECT 41.460000 199.250000 41.660000 199.450000 ;
        RECT 41.460000 199.650000 41.660000 199.850000 ;
        RECT 41.860000 197.250000 42.060000 197.450000 ;
        RECT 41.860000 197.650000 42.060000 197.850000 ;
        RECT 41.860000 198.050000 42.060000 198.250000 ;
        RECT 41.860000 198.450000 42.060000 198.650000 ;
        RECT 41.860000 198.850000 42.060000 199.050000 ;
        RECT 41.860000 199.250000 42.060000 199.450000 ;
        RECT 41.860000 199.650000 42.060000 199.850000 ;
        RECT 42.260000 197.250000 42.460000 197.450000 ;
        RECT 42.260000 197.650000 42.460000 197.850000 ;
        RECT 42.260000 198.050000 42.460000 198.250000 ;
        RECT 42.260000 198.450000 42.460000 198.650000 ;
        RECT 42.260000 198.850000 42.460000 199.050000 ;
        RECT 42.260000 199.250000 42.460000 199.450000 ;
        RECT 42.260000 199.650000 42.460000 199.850000 ;
        RECT 42.660000 197.250000 42.860000 197.450000 ;
        RECT 42.660000 197.650000 42.860000 197.850000 ;
        RECT 42.660000 198.050000 42.860000 198.250000 ;
        RECT 42.660000 198.450000 42.860000 198.650000 ;
        RECT 42.660000 198.850000 42.860000 199.050000 ;
        RECT 42.660000 199.250000 42.860000 199.450000 ;
        RECT 42.660000 199.650000 42.860000 199.850000 ;
        RECT 43.060000 197.250000 43.260000 197.450000 ;
        RECT 43.060000 197.650000 43.260000 197.850000 ;
        RECT 43.060000 198.050000 43.260000 198.250000 ;
        RECT 43.060000 198.450000 43.260000 198.650000 ;
        RECT 43.060000 198.850000 43.260000 199.050000 ;
        RECT 43.060000 199.250000 43.260000 199.450000 ;
        RECT 43.060000 199.650000 43.260000 199.850000 ;
        RECT 43.460000 197.250000 43.660000 197.450000 ;
        RECT 43.460000 197.650000 43.660000 197.850000 ;
        RECT 43.460000 198.050000 43.660000 198.250000 ;
        RECT 43.460000 198.450000 43.660000 198.650000 ;
        RECT 43.460000 198.850000 43.660000 199.050000 ;
        RECT 43.460000 199.250000 43.660000 199.450000 ;
        RECT 43.460000 199.650000 43.660000 199.850000 ;
        RECT 43.860000 197.250000 44.060000 197.450000 ;
        RECT 43.860000 197.650000 44.060000 197.850000 ;
        RECT 43.860000 198.050000 44.060000 198.250000 ;
        RECT 43.860000 198.450000 44.060000 198.650000 ;
        RECT 43.860000 198.850000 44.060000 199.050000 ;
        RECT 43.860000 199.250000 44.060000 199.450000 ;
        RECT 43.860000 199.650000 44.060000 199.850000 ;
        RECT 44.260000 197.250000 44.460000 197.450000 ;
        RECT 44.260000 197.650000 44.460000 197.850000 ;
        RECT 44.260000 198.050000 44.460000 198.250000 ;
        RECT 44.260000 198.450000 44.460000 198.650000 ;
        RECT 44.260000 198.850000 44.460000 199.050000 ;
        RECT 44.260000 199.250000 44.460000 199.450000 ;
        RECT 44.260000 199.650000 44.460000 199.850000 ;
        RECT 44.660000 197.250000 44.860000 197.450000 ;
        RECT 44.660000 197.650000 44.860000 197.850000 ;
        RECT 44.660000 198.050000 44.860000 198.250000 ;
        RECT 44.660000 198.450000 44.860000 198.650000 ;
        RECT 44.660000 198.850000 44.860000 199.050000 ;
        RECT 44.660000 199.250000 44.860000 199.450000 ;
        RECT 44.660000 199.650000 44.860000 199.850000 ;
        RECT 45.060000 197.250000 45.260000 197.450000 ;
        RECT 45.060000 197.650000 45.260000 197.850000 ;
        RECT 45.060000 198.050000 45.260000 198.250000 ;
        RECT 45.060000 198.450000 45.260000 198.650000 ;
        RECT 45.060000 198.850000 45.260000 199.050000 ;
        RECT 45.060000 199.250000 45.260000 199.450000 ;
        RECT 45.060000 199.650000 45.260000 199.850000 ;
        RECT 45.460000 197.250000 45.660000 197.450000 ;
        RECT 45.460000 197.650000 45.660000 197.850000 ;
        RECT 45.460000 198.050000 45.660000 198.250000 ;
        RECT 45.460000 198.450000 45.660000 198.650000 ;
        RECT 45.460000 198.850000 45.660000 199.050000 ;
        RECT 45.460000 199.250000 45.660000 199.450000 ;
        RECT 45.460000 199.650000 45.660000 199.850000 ;
        RECT 45.860000 197.250000 46.060000 197.450000 ;
        RECT 45.860000 197.650000 46.060000 197.850000 ;
        RECT 45.860000 198.050000 46.060000 198.250000 ;
        RECT 45.860000 198.450000 46.060000 198.650000 ;
        RECT 45.860000 198.850000 46.060000 199.050000 ;
        RECT 45.860000 199.250000 46.060000 199.450000 ;
        RECT 45.860000 199.650000 46.060000 199.850000 ;
        RECT 46.260000 197.250000 46.460000 197.450000 ;
        RECT 46.260000 197.650000 46.460000 197.850000 ;
        RECT 46.260000 198.050000 46.460000 198.250000 ;
        RECT 46.260000 198.450000 46.460000 198.650000 ;
        RECT 46.260000 198.850000 46.460000 199.050000 ;
        RECT 46.260000 199.250000 46.460000 199.450000 ;
        RECT 46.260000 199.650000 46.460000 199.850000 ;
        RECT 46.660000 197.250000 46.860000 197.450000 ;
        RECT 46.660000 197.650000 46.860000 197.850000 ;
        RECT 46.660000 198.050000 46.860000 198.250000 ;
        RECT 46.660000 198.450000 46.860000 198.650000 ;
        RECT 46.660000 198.850000 46.860000 199.050000 ;
        RECT 46.660000 199.250000 46.860000 199.450000 ;
        RECT 46.660000 199.650000 46.860000 199.850000 ;
        RECT 47.060000 197.250000 47.260000 197.450000 ;
        RECT 47.060000 197.650000 47.260000 197.850000 ;
        RECT 47.060000 198.050000 47.260000 198.250000 ;
        RECT 47.060000 198.450000 47.260000 198.650000 ;
        RECT 47.060000 198.850000 47.260000 199.050000 ;
        RECT 47.060000 199.250000 47.260000 199.450000 ;
        RECT 47.060000 199.650000 47.260000 199.850000 ;
        RECT 47.460000 197.250000 47.660000 197.450000 ;
        RECT 47.460000 197.650000 47.660000 197.850000 ;
        RECT 47.460000 198.050000 47.660000 198.250000 ;
        RECT 47.460000 198.450000 47.660000 198.650000 ;
        RECT 47.460000 198.850000 47.660000 199.050000 ;
        RECT 47.460000 199.250000 47.660000 199.450000 ;
        RECT 47.460000 199.650000 47.660000 199.850000 ;
        RECT 47.860000 197.250000 48.060000 197.450000 ;
        RECT 47.860000 197.650000 48.060000 197.850000 ;
        RECT 47.860000 198.050000 48.060000 198.250000 ;
        RECT 47.860000 198.450000 48.060000 198.650000 ;
        RECT 47.860000 198.850000 48.060000 199.050000 ;
        RECT 47.860000 199.250000 48.060000 199.450000 ;
        RECT 47.860000 199.650000 48.060000 199.850000 ;
        RECT 48.260000 197.250000 48.460000 197.450000 ;
        RECT 48.260000 197.650000 48.460000 197.850000 ;
        RECT 48.260000 198.050000 48.460000 198.250000 ;
        RECT 48.260000 198.450000 48.460000 198.650000 ;
        RECT 48.260000 198.850000 48.460000 199.050000 ;
        RECT 48.260000 199.250000 48.460000 199.450000 ;
        RECT 48.260000 199.650000 48.460000 199.850000 ;
        RECT 48.660000 197.250000 48.860000 197.450000 ;
        RECT 48.660000 197.650000 48.860000 197.850000 ;
        RECT 48.660000 198.050000 48.860000 198.250000 ;
        RECT 48.660000 198.450000 48.860000 198.650000 ;
        RECT 48.660000 198.850000 48.860000 199.050000 ;
        RECT 48.660000 199.250000 48.860000 199.450000 ;
        RECT 48.660000 199.650000 48.860000 199.850000 ;
        RECT 49.060000 197.250000 49.260000 197.450000 ;
        RECT 49.060000 197.650000 49.260000 197.850000 ;
        RECT 49.060000 198.050000 49.260000 198.250000 ;
        RECT 49.060000 198.450000 49.260000 198.650000 ;
        RECT 49.060000 198.850000 49.260000 199.050000 ;
        RECT 49.060000 199.250000 49.260000 199.450000 ;
        RECT 49.060000 199.650000 49.260000 199.850000 ;
        RECT 49.460000 197.250000 49.660000 197.450000 ;
        RECT 49.460000 197.650000 49.660000 197.850000 ;
        RECT 49.460000 198.050000 49.660000 198.250000 ;
        RECT 49.460000 198.450000 49.660000 198.650000 ;
        RECT 49.460000 198.850000 49.660000 199.050000 ;
        RECT 49.460000 199.250000 49.660000 199.450000 ;
        RECT 49.460000 199.650000 49.660000 199.850000 ;
        RECT 49.860000 197.250000 50.060000 197.450000 ;
        RECT 49.860000 197.650000 50.060000 197.850000 ;
        RECT 49.860000 198.050000 50.060000 198.250000 ;
        RECT 49.860000 198.450000 50.060000 198.650000 ;
        RECT 49.860000 198.850000 50.060000 199.050000 ;
        RECT 49.860000 199.250000 50.060000 199.450000 ;
        RECT 49.860000 199.650000 50.060000 199.850000 ;
        RECT 50.260000 197.250000 50.460000 197.450000 ;
        RECT 50.260000 197.650000 50.460000 197.850000 ;
        RECT 50.260000 198.050000 50.460000 198.250000 ;
        RECT 50.260000 198.450000 50.460000 198.650000 ;
        RECT 50.260000 198.850000 50.460000 199.050000 ;
        RECT 50.260000 199.250000 50.460000 199.450000 ;
        RECT 50.260000 199.650000 50.460000 199.850000 ;
        RECT 50.480000  25.910000 50.680000  26.110000 ;
        RECT 50.480000  26.340000 50.680000  26.540000 ;
        RECT 50.480000  26.770000 50.680000  26.970000 ;
        RECT 50.480000  27.200000 50.680000  27.400000 ;
        RECT 50.480000  27.630000 50.680000  27.830000 ;
        RECT 50.480000  28.060000 50.680000  28.260000 ;
        RECT 50.480000  28.490000 50.680000  28.690000 ;
        RECT 50.480000  28.920000 50.680000  29.120000 ;
        RECT 50.480000  29.350000 50.680000  29.550000 ;
        RECT 50.480000  29.780000 50.680000  29.980000 ;
        RECT 50.480000  30.210000 50.680000  30.410000 ;
        RECT 50.660000 197.250000 50.860000 197.450000 ;
        RECT 50.660000 197.650000 50.860000 197.850000 ;
        RECT 50.660000 198.050000 50.860000 198.250000 ;
        RECT 50.660000 198.450000 50.860000 198.650000 ;
        RECT 50.660000 198.850000 50.860000 199.050000 ;
        RECT 50.660000 199.250000 50.860000 199.450000 ;
        RECT 50.660000 199.650000 50.860000 199.850000 ;
        RECT 50.890000  25.910000 51.090000  26.110000 ;
        RECT 50.890000  26.340000 51.090000  26.540000 ;
        RECT 50.890000  26.770000 51.090000  26.970000 ;
        RECT 50.890000  27.200000 51.090000  27.400000 ;
        RECT 50.890000  27.630000 51.090000  27.830000 ;
        RECT 50.890000  28.060000 51.090000  28.260000 ;
        RECT 50.890000  28.490000 51.090000  28.690000 ;
        RECT 50.890000  28.920000 51.090000  29.120000 ;
        RECT 50.890000  29.350000 51.090000  29.550000 ;
        RECT 50.890000  29.780000 51.090000  29.980000 ;
        RECT 50.890000  30.210000 51.090000  30.410000 ;
        RECT 51.060000 197.250000 51.260000 197.450000 ;
        RECT 51.060000 197.650000 51.260000 197.850000 ;
        RECT 51.060000 198.050000 51.260000 198.250000 ;
        RECT 51.060000 198.450000 51.260000 198.650000 ;
        RECT 51.060000 198.850000 51.260000 199.050000 ;
        RECT 51.060000 199.250000 51.260000 199.450000 ;
        RECT 51.060000 199.650000 51.260000 199.850000 ;
        RECT 51.300000  25.910000 51.500000  26.110000 ;
        RECT 51.300000  26.340000 51.500000  26.540000 ;
        RECT 51.300000  26.770000 51.500000  26.970000 ;
        RECT 51.300000  27.200000 51.500000  27.400000 ;
        RECT 51.300000  27.630000 51.500000  27.830000 ;
        RECT 51.300000  28.060000 51.500000  28.260000 ;
        RECT 51.300000  28.490000 51.500000  28.690000 ;
        RECT 51.300000  28.920000 51.500000  29.120000 ;
        RECT 51.300000  29.350000 51.500000  29.550000 ;
        RECT 51.300000  29.780000 51.500000  29.980000 ;
        RECT 51.300000  30.210000 51.500000  30.410000 ;
        RECT 51.460000 197.250000 51.660000 197.450000 ;
        RECT 51.460000 197.650000 51.660000 197.850000 ;
        RECT 51.460000 198.050000 51.660000 198.250000 ;
        RECT 51.460000 198.450000 51.660000 198.650000 ;
        RECT 51.460000 198.850000 51.660000 199.050000 ;
        RECT 51.460000 199.250000 51.660000 199.450000 ;
        RECT 51.460000 199.650000 51.660000 199.850000 ;
        RECT 51.710000  25.910000 51.910000  26.110000 ;
        RECT 51.710000  26.340000 51.910000  26.540000 ;
        RECT 51.710000  26.770000 51.910000  26.970000 ;
        RECT 51.710000  27.200000 51.910000  27.400000 ;
        RECT 51.710000  27.630000 51.910000  27.830000 ;
        RECT 51.710000  28.060000 51.910000  28.260000 ;
        RECT 51.710000  28.490000 51.910000  28.690000 ;
        RECT 51.710000  28.920000 51.910000  29.120000 ;
        RECT 51.710000  29.350000 51.910000  29.550000 ;
        RECT 51.710000  29.780000 51.910000  29.980000 ;
        RECT 51.710000  30.210000 51.910000  30.410000 ;
        RECT 51.860000 197.250000 52.060000 197.450000 ;
        RECT 51.860000 197.650000 52.060000 197.850000 ;
        RECT 51.860000 198.050000 52.060000 198.250000 ;
        RECT 51.860000 198.450000 52.060000 198.650000 ;
        RECT 51.860000 198.850000 52.060000 199.050000 ;
        RECT 51.860000 199.250000 52.060000 199.450000 ;
        RECT 51.860000 199.650000 52.060000 199.850000 ;
        RECT 52.120000  25.910000 52.320000  26.110000 ;
        RECT 52.120000  26.340000 52.320000  26.540000 ;
        RECT 52.120000  26.770000 52.320000  26.970000 ;
        RECT 52.120000  27.200000 52.320000  27.400000 ;
        RECT 52.120000  27.630000 52.320000  27.830000 ;
        RECT 52.120000  28.060000 52.320000  28.260000 ;
        RECT 52.120000  28.490000 52.320000  28.690000 ;
        RECT 52.120000  28.920000 52.320000  29.120000 ;
        RECT 52.120000  29.350000 52.320000  29.550000 ;
        RECT 52.120000  29.780000 52.320000  29.980000 ;
        RECT 52.120000  30.210000 52.320000  30.410000 ;
        RECT 52.260000 197.250000 52.460000 197.450000 ;
        RECT 52.260000 197.650000 52.460000 197.850000 ;
        RECT 52.260000 198.050000 52.460000 198.250000 ;
        RECT 52.260000 198.450000 52.460000 198.650000 ;
        RECT 52.260000 198.850000 52.460000 199.050000 ;
        RECT 52.260000 199.250000 52.460000 199.450000 ;
        RECT 52.260000 199.650000 52.460000 199.850000 ;
        RECT 52.530000  25.910000 52.730000  26.110000 ;
        RECT 52.530000  26.340000 52.730000  26.540000 ;
        RECT 52.530000  26.770000 52.730000  26.970000 ;
        RECT 52.530000  27.200000 52.730000  27.400000 ;
        RECT 52.530000  27.630000 52.730000  27.830000 ;
        RECT 52.530000  28.060000 52.730000  28.260000 ;
        RECT 52.530000  28.490000 52.730000  28.690000 ;
        RECT 52.530000  28.920000 52.730000  29.120000 ;
        RECT 52.530000  29.350000 52.730000  29.550000 ;
        RECT 52.530000  29.780000 52.730000  29.980000 ;
        RECT 52.530000  30.210000 52.730000  30.410000 ;
        RECT 52.660000 197.250000 52.860000 197.450000 ;
        RECT 52.660000 197.650000 52.860000 197.850000 ;
        RECT 52.660000 198.050000 52.860000 198.250000 ;
        RECT 52.660000 198.450000 52.860000 198.650000 ;
        RECT 52.660000 198.850000 52.860000 199.050000 ;
        RECT 52.660000 199.250000 52.860000 199.450000 ;
        RECT 52.660000 199.650000 52.860000 199.850000 ;
        RECT 52.940000  25.910000 53.140000  26.110000 ;
        RECT 52.940000  26.340000 53.140000  26.540000 ;
        RECT 52.940000  26.770000 53.140000  26.970000 ;
        RECT 52.940000  27.200000 53.140000  27.400000 ;
        RECT 52.940000  27.630000 53.140000  27.830000 ;
        RECT 52.940000  28.060000 53.140000  28.260000 ;
        RECT 52.940000  28.490000 53.140000  28.690000 ;
        RECT 52.940000  28.920000 53.140000  29.120000 ;
        RECT 52.940000  29.350000 53.140000  29.550000 ;
        RECT 52.940000  29.780000 53.140000  29.980000 ;
        RECT 52.940000  30.210000 53.140000  30.410000 ;
        RECT 53.060000 197.250000 53.260000 197.450000 ;
        RECT 53.060000 197.650000 53.260000 197.850000 ;
        RECT 53.060000 198.050000 53.260000 198.250000 ;
        RECT 53.060000 198.450000 53.260000 198.650000 ;
        RECT 53.060000 198.850000 53.260000 199.050000 ;
        RECT 53.060000 199.250000 53.260000 199.450000 ;
        RECT 53.060000 199.650000 53.260000 199.850000 ;
        RECT 53.345000  25.910000 53.545000  26.110000 ;
        RECT 53.345000  26.340000 53.545000  26.540000 ;
        RECT 53.345000  26.770000 53.545000  26.970000 ;
        RECT 53.345000  27.200000 53.545000  27.400000 ;
        RECT 53.345000  27.630000 53.545000  27.830000 ;
        RECT 53.345000  28.060000 53.545000  28.260000 ;
        RECT 53.345000  28.490000 53.545000  28.690000 ;
        RECT 53.345000  28.920000 53.545000  29.120000 ;
        RECT 53.345000  29.350000 53.545000  29.550000 ;
        RECT 53.345000  29.780000 53.545000  29.980000 ;
        RECT 53.345000  30.210000 53.545000  30.410000 ;
        RECT 53.460000 197.250000 53.660000 197.450000 ;
        RECT 53.460000 197.650000 53.660000 197.850000 ;
        RECT 53.460000 198.050000 53.660000 198.250000 ;
        RECT 53.460000 198.450000 53.660000 198.650000 ;
        RECT 53.460000 198.850000 53.660000 199.050000 ;
        RECT 53.460000 199.250000 53.660000 199.450000 ;
        RECT 53.460000 199.650000 53.660000 199.850000 ;
        RECT 53.750000  25.910000 53.950000  26.110000 ;
        RECT 53.750000  26.340000 53.950000  26.540000 ;
        RECT 53.750000  26.770000 53.950000  26.970000 ;
        RECT 53.750000  27.200000 53.950000  27.400000 ;
        RECT 53.750000  27.630000 53.950000  27.830000 ;
        RECT 53.750000  28.060000 53.950000  28.260000 ;
        RECT 53.750000  28.490000 53.950000  28.690000 ;
        RECT 53.750000  28.920000 53.950000  29.120000 ;
        RECT 53.750000  29.350000 53.950000  29.550000 ;
        RECT 53.750000  29.780000 53.950000  29.980000 ;
        RECT 53.750000  30.210000 53.950000  30.410000 ;
        RECT 53.860000 197.250000 54.060000 197.450000 ;
        RECT 53.860000 197.650000 54.060000 197.850000 ;
        RECT 53.860000 198.050000 54.060000 198.250000 ;
        RECT 53.860000 198.450000 54.060000 198.650000 ;
        RECT 53.860000 198.850000 54.060000 199.050000 ;
        RECT 53.860000 199.250000 54.060000 199.450000 ;
        RECT 53.860000 199.650000 54.060000 199.850000 ;
        RECT 54.155000  25.910000 54.355000  26.110000 ;
        RECT 54.155000  26.340000 54.355000  26.540000 ;
        RECT 54.155000  26.770000 54.355000  26.970000 ;
        RECT 54.155000  27.200000 54.355000  27.400000 ;
        RECT 54.155000  27.630000 54.355000  27.830000 ;
        RECT 54.155000  28.060000 54.355000  28.260000 ;
        RECT 54.155000  28.490000 54.355000  28.690000 ;
        RECT 54.155000  28.920000 54.355000  29.120000 ;
        RECT 54.155000  29.350000 54.355000  29.550000 ;
        RECT 54.155000  29.780000 54.355000  29.980000 ;
        RECT 54.155000  30.210000 54.355000  30.410000 ;
        RECT 54.260000 197.250000 54.460000 197.450000 ;
        RECT 54.260000 197.650000 54.460000 197.850000 ;
        RECT 54.260000 198.050000 54.460000 198.250000 ;
        RECT 54.260000 198.450000 54.460000 198.650000 ;
        RECT 54.260000 198.850000 54.460000 199.050000 ;
        RECT 54.260000 199.250000 54.460000 199.450000 ;
        RECT 54.260000 199.650000 54.460000 199.850000 ;
        RECT 54.560000  25.910000 54.760000  26.110000 ;
        RECT 54.560000  26.340000 54.760000  26.540000 ;
        RECT 54.560000  26.770000 54.760000  26.970000 ;
        RECT 54.560000  27.200000 54.760000  27.400000 ;
        RECT 54.560000  27.630000 54.760000  27.830000 ;
        RECT 54.560000  28.060000 54.760000  28.260000 ;
        RECT 54.560000  28.490000 54.760000  28.690000 ;
        RECT 54.560000  28.920000 54.760000  29.120000 ;
        RECT 54.560000  29.350000 54.760000  29.550000 ;
        RECT 54.560000  29.780000 54.760000  29.980000 ;
        RECT 54.560000  30.210000 54.760000  30.410000 ;
        RECT 54.660000 197.250000 54.860000 197.450000 ;
        RECT 54.660000 197.650000 54.860000 197.850000 ;
        RECT 54.660000 198.050000 54.860000 198.250000 ;
        RECT 54.660000 198.450000 54.860000 198.650000 ;
        RECT 54.660000 198.850000 54.860000 199.050000 ;
        RECT 54.660000 199.250000 54.860000 199.450000 ;
        RECT 54.660000 199.650000 54.860000 199.850000 ;
        RECT 54.965000  25.910000 55.165000  26.110000 ;
        RECT 54.965000  26.340000 55.165000  26.540000 ;
        RECT 54.965000  26.770000 55.165000  26.970000 ;
        RECT 54.965000  27.200000 55.165000  27.400000 ;
        RECT 54.965000  27.630000 55.165000  27.830000 ;
        RECT 54.965000  28.060000 55.165000  28.260000 ;
        RECT 54.965000  28.490000 55.165000  28.690000 ;
        RECT 54.965000  28.920000 55.165000  29.120000 ;
        RECT 54.965000  29.350000 55.165000  29.550000 ;
        RECT 54.965000  29.780000 55.165000  29.980000 ;
        RECT 54.965000  30.210000 55.165000  30.410000 ;
        RECT 55.060000 197.250000 55.260000 197.450000 ;
        RECT 55.060000 197.650000 55.260000 197.850000 ;
        RECT 55.060000 198.050000 55.260000 198.250000 ;
        RECT 55.060000 198.450000 55.260000 198.650000 ;
        RECT 55.060000 198.850000 55.260000 199.050000 ;
        RECT 55.060000 199.250000 55.260000 199.450000 ;
        RECT 55.060000 199.650000 55.260000 199.850000 ;
        RECT 55.370000  25.910000 55.570000  26.110000 ;
        RECT 55.370000  26.340000 55.570000  26.540000 ;
        RECT 55.370000  26.770000 55.570000  26.970000 ;
        RECT 55.370000  27.200000 55.570000  27.400000 ;
        RECT 55.370000  27.630000 55.570000  27.830000 ;
        RECT 55.370000  28.060000 55.570000  28.260000 ;
        RECT 55.370000  28.490000 55.570000  28.690000 ;
        RECT 55.370000  28.920000 55.570000  29.120000 ;
        RECT 55.370000  29.350000 55.570000  29.550000 ;
        RECT 55.370000  29.780000 55.570000  29.980000 ;
        RECT 55.370000  30.210000 55.570000  30.410000 ;
        RECT 55.460000 197.250000 55.660000 197.450000 ;
        RECT 55.460000 197.650000 55.660000 197.850000 ;
        RECT 55.460000 198.050000 55.660000 198.250000 ;
        RECT 55.460000 198.450000 55.660000 198.650000 ;
        RECT 55.460000 198.850000 55.660000 199.050000 ;
        RECT 55.460000 199.250000 55.660000 199.450000 ;
        RECT 55.460000 199.650000 55.660000 199.850000 ;
        RECT 55.775000  25.910000 55.975000  26.110000 ;
        RECT 55.775000  26.340000 55.975000  26.540000 ;
        RECT 55.775000  26.770000 55.975000  26.970000 ;
        RECT 55.775000  27.200000 55.975000  27.400000 ;
        RECT 55.775000  27.630000 55.975000  27.830000 ;
        RECT 55.775000  28.060000 55.975000  28.260000 ;
        RECT 55.775000  28.490000 55.975000  28.690000 ;
        RECT 55.775000  28.920000 55.975000  29.120000 ;
        RECT 55.775000  29.350000 55.975000  29.550000 ;
        RECT 55.775000  29.780000 55.975000  29.980000 ;
        RECT 55.775000  30.210000 55.975000  30.410000 ;
        RECT 55.860000 197.250000 56.060000 197.450000 ;
        RECT 55.860000 197.650000 56.060000 197.850000 ;
        RECT 55.860000 198.050000 56.060000 198.250000 ;
        RECT 55.860000 198.450000 56.060000 198.650000 ;
        RECT 55.860000 198.850000 56.060000 199.050000 ;
        RECT 55.860000 199.250000 56.060000 199.450000 ;
        RECT 55.860000 199.650000 56.060000 199.850000 ;
        RECT 56.180000  25.910000 56.380000  26.110000 ;
        RECT 56.180000  26.340000 56.380000  26.540000 ;
        RECT 56.180000  26.770000 56.380000  26.970000 ;
        RECT 56.180000  27.200000 56.380000  27.400000 ;
        RECT 56.180000  27.630000 56.380000  27.830000 ;
        RECT 56.180000  28.060000 56.380000  28.260000 ;
        RECT 56.180000  28.490000 56.380000  28.690000 ;
        RECT 56.180000  28.920000 56.380000  29.120000 ;
        RECT 56.180000  29.350000 56.380000  29.550000 ;
        RECT 56.180000  29.780000 56.380000  29.980000 ;
        RECT 56.180000  30.210000 56.380000  30.410000 ;
        RECT 56.260000 197.250000 56.460000 197.450000 ;
        RECT 56.260000 197.650000 56.460000 197.850000 ;
        RECT 56.260000 198.050000 56.460000 198.250000 ;
        RECT 56.260000 198.450000 56.460000 198.650000 ;
        RECT 56.260000 198.850000 56.460000 199.050000 ;
        RECT 56.260000 199.250000 56.460000 199.450000 ;
        RECT 56.260000 199.650000 56.460000 199.850000 ;
        RECT 56.585000  25.910000 56.785000  26.110000 ;
        RECT 56.585000  26.340000 56.785000  26.540000 ;
        RECT 56.585000  26.770000 56.785000  26.970000 ;
        RECT 56.585000  27.200000 56.785000  27.400000 ;
        RECT 56.585000  27.630000 56.785000  27.830000 ;
        RECT 56.585000  28.060000 56.785000  28.260000 ;
        RECT 56.585000  28.490000 56.785000  28.690000 ;
        RECT 56.585000  28.920000 56.785000  29.120000 ;
        RECT 56.585000  29.350000 56.785000  29.550000 ;
        RECT 56.585000  29.780000 56.785000  29.980000 ;
        RECT 56.585000  30.210000 56.785000  30.410000 ;
        RECT 56.660000 197.250000 56.860000 197.450000 ;
        RECT 56.660000 197.650000 56.860000 197.850000 ;
        RECT 56.660000 198.050000 56.860000 198.250000 ;
        RECT 56.660000 198.450000 56.860000 198.650000 ;
        RECT 56.660000 198.850000 56.860000 199.050000 ;
        RECT 56.660000 199.250000 56.860000 199.450000 ;
        RECT 56.660000 199.650000 56.860000 199.850000 ;
        RECT 56.990000  25.910000 57.190000  26.110000 ;
        RECT 56.990000  26.340000 57.190000  26.540000 ;
        RECT 56.990000  26.770000 57.190000  26.970000 ;
        RECT 56.990000  27.200000 57.190000  27.400000 ;
        RECT 56.990000  27.630000 57.190000  27.830000 ;
        RECT 56.990000  28.060000 57.190000  28.260000 ;
        RECT 56.990000  28.490000 57.190000  28.690000 ;
        RECT 56.990000  28.920000 57.190000  29.120000 ;
        RECT 56.990000  29.350000 57.190000  29.550000 ;
        RECT 56.990000  29.780000 57.190000  29.980000 ;
        RECT 56.990000  30.210000 57.190000  30.410000 ;
        RECT 57.060000 197.250000 57.260000 197.450000 ;
        RECT 57.060000 197.650000 57.260000 197.850000 ;
        RECT 57.060000 198.050000 57.260000 198.250000 ;
        RECT 57.060000 198.450000 57.260000 198.650000 ;
        RECT 57.060000 198.850000 57.260000 199.050000 ;
        RECT 57.060000 199.250000 57.260000 199.450000 ;
        RECT 57.060000 199.650000 57.260000 199.850000 ;
        RECT 57.395000  25.910000 57.595000  26.110000 ;
        RECT 57.395000  26.340000 57.595000  26.540000 ;
        RECT 57.395000  26.770000 57.595000  26.970000 ;
        RECT 57.395000  27.200000 57.595000  27.400000 ;
        RECT 57.395000  27.630000 57.595000  27.830000 ;
        RECT 57.395000  28.060000 57.595000  28.260000 ;
        RECT 57.395000  28.490000 57.595000  28.690000 ;
        RECT 57.395000  28.920000 57.595000  29.120000 ;
        RECT 57.395000  29.350000 57.595000  29.550000 ;
        RECT 57.395000  29.780000 57.595000  29.980000 ;
        RECT 57.395000  30.210000 57.595000  30.410000 ;
        RECT 57.460000 197.250000 57.660000 197.450000 ;
        RECT 57.460000 197.650000 57.660000 197.850000 ;
        RECT 57.460000 198.050000 57.660000 198.250000 ;
        RECT 57.460000 198.450000 57.660000 198.650000 ;
        RECT 57.460000 198.850000 57.660000 199.050000 ;
        RECT 57.460000 199.250000 57.660000 199.450000 ;
        RECT 57.460000 199.650000 57.660000 199.850000 ;
        RECT 57.800000  25.910000 58.000000  26.110000 ;
        RECT 57.800000  26.340000 58.000000  26.540000 ;
        RECT 57.800000  26.770000 58.000000  26.970000 ;
        RECT 57.800000  27.200000 58.000000  27.400000 ;
        RECT 57.800000  27.630000 58.000000  27.830000 ;
        RECT 57.800000  28.060000 58.000000  28.260000 ;
        RECT 57.800000  28.490000 58.000000  28.690000 ;
        RECT 57.800000  28.920000 58.000000  29.120000 ;
        RECT 57.800000  29.350000 58.000000  29.550000 ;
        RECT 57.800000  29.780000 58.000000  29.980000 ;
        RECT 57.800000  30.210000 58.000000  30.410000 ;
        RECT 57.860000 197.250000 58.060000 197.450000 ;
        RECT 57.860000 197.650000 58.060000 197.850000 ;
        RECT 57.860000 198.050000 58.060000 198.250000 ;
        RECT 57.860000 198.450000 58.060000 198.650000 ;
        RECT 57.860000 198.850000 58.060000 199.050000 ;
        RECT 57.860000 199.250000 58.060000 199.450000 ;
        RECT 57.860000 199.650000 58.060000 199.850000 ;
        RECT 58.205000  25.910000 58.405000  26.110000 ;
        RECT 58.205000  26.340000 58.405000  26.540000 ;
        RECT 58.205000  26.770000 58.405000  26.970000 ;
        RECT 58.205000  27.200000 58.405000  27.400000 ;
        RECT 58.205000  27.630000 58.405000  27.830000 ;
        RECT 58.205000  28.060000 58.405000  28.260000 ;
        RECT 58.205000  28.490000 58.405000  28.690000 ;
        RECT 58.205000  28.920000 58.405000  29.120000 ;
        RECT 58.205000  29.350000 58.405000  29.550000 ;
        RECT 58.205000  29.780000 58.405000  29.980000 ;
        RECT 58.205000  30.210000 58.405000  30.410000 ;
        RECT 58.260000 197.250000 58.460000 197.450000 ;
        RECT 58.260000 197.650000 58.460000 197.850000 ;
        RECT 58.260000 198.050000 58.460000 198.250000 ;
        RECT 58.260000 198.450000 58.460000 198.650000 ;
        RECT 58.260000 198.850000 58.460000 199.050000 ;
        RECT 58.260000 199.250000 58.460000 199.450000 ;
        RECT 58.260000 199.650000 58.460000 199.850000 ;
        RECT 58.610000  25.910000 58.810000  26.110000 ;
        RECT 58.610000  26.340000 58.810000  26.540000 ;
        RECT 58.610000  26.770000 58.810000  26.970000 ;
        RECT 58.610000  27.200000 58.810000  27.400000 ;
        RECT 58.610000  27.630000 58.810000  27.830000 ;
        RECT 58.610000  28.060000 58.810000  28.260000 ;
        RECT 58.610000  28.490000 58.810000  28.690000 ;
        RECT 58.610000  28.920000 58.810000  29.120000 ;
        RECT 58.610000  29.350000 58.810000  29.550000 ;
        RECT 58.610000  29.780000 58.810000  29.980000 ;
        RECT 58.610000  30.210000 58.810000  30.410000 ;
        RECT 58.660000 197.250000 58.860000 197.450000 ;
        RECT 58.660000 197.650000 58.860000 197.850000 ;
        RECT 58.660000 198.050000 58.860000 198.250000 ;
        RECT 58.660000 198.450000 58.860000 198.650000 ;
        RECT 58.660000 198.850000 58.860000 199.050000 ;
        RECT 58.660000 199.250000 58.860000 199.450000 ;
        RECT 58.660000 199.650000 58.860000 199.850000 ;
        RECT 59.015000  25.910000 59.215000  26.110000 ;
        RECT 59.015000  26.340000 59.215000  26.540000 ;
        RECT 59.015000  26.770000 59.215000  26.970000 ;
        RECT 59.015000  27.200000 59.215000  27.400000 ;
        RECT 59.015000  27.630000 59.215000  27.830000 ;
        RECT 59.015000  28.060000 59.215000  28.260000 ;
        RECT 59.015000  28.490000 59.215000  28.690000 ;
        RECT 59.015000  28.920000 59.215000  29.120000 ;
        RECT 59.015000  29.350000 59.215000  29.550000 ;
        RECT 59.015000  29.780000 59.215000  29.980000 ;
        RECT 59.015000  30.210000 59.215000  30.410000 ;
        RECT 59.060000 197.250000 59.260000 197.450000 ;
        RECT 59.060000 197.650000 59.260000 197.850000 ;
        RECT 59.060000 198.050000 59.260000 198.250000 ;
        RECT 59.060000 198.450000 59.260000 198.650000 ;
        RECT 59.060000 198.850000 59.260000 199.050000 ;
        RECT 59.060000 199.250000 59.260000 199.450000 ;
        RECT 59.060000 199.650000 59.260000 199.850000 ;
        RECT 59.420000  25.910000 59.620000  26.110000 ;
        RECT 59.420000  26.340000 59.620000  26.540000 ;
        RECT 59.420000  26.770000 59.620000  26.970000 ;
        RECT 59.420000  27.200000 59.620000  27.400000 ;
        RECT 59.420000  27.630000 59.620000  27.830000 ;
        RECT 59.420000  28.060000 59.620000  28.260000 ;
        RECT 59.420000  28.490000 59.620000  28.690000 ;
        RECT 59.420000  28.920000 59.620000  29.120000 ;
        RECT 59.420000  29.350000 59.620000  29.550000 ;
        RECT 59.420000  29.780000 59.620000  29.980000 ;
        RECT 59.420000  30.210000 59.620000  30.410000 ;
        RECT 59.460000 197.250000 59.660000 197.450000 ;
        RECT 59.460000 197.650000 59.660000 197.850000 ;
        RECT 59.460000 198.050000 59.660000 198.250000 ;
        RECT 59.460000 198.450000 59.660000 198.650000 ;
        RECT 59.460000 198.850000 59.660000 199.050000 ;
        RECT 59.460000 199.250000 59.660000 199.450000 ;
        RECT 59.460000 199.650000 59.660000 199.850000 ;
        RECT 59.825000  25.910000 60.025000  26.110000 ;
        RECT 59.825000  26.340000 60.025000  26.540000 ;
        RECT 59.825000  26.770000 60.025000  26.970000 ;
        RECT 59.825000  27.200000 60.025000  27.400000 ;
        RECT 59.825000  27.630000 60.025000  27.830000 ;
        RECT 59.825000  28.060000 60.025000  28.260000 ;
        RECT 59.825000  28.490000 60.025000  28.690000 ;
        RECT 59.825000  28.920000 60.025000  29.120000 ;
        RECT 59.825000  29.350000 60.025000  29.550000 ;
        RECT 59.825000  29.780000 60.025000  29.980000 ;
        RECT 59.825000  30.210000 60.025000  30.410000 ;
        RECT 59.860000 197.250000 60.060000 197.450000 ;
        RECT 59.860000 197.650000 60.060000 197.850000 ;
        RECT 59.860000 198.050000 60.060000 198.250000 ;
        RECT 59.860000 198.450000 60.060000 198.650000 ;
        RECT 59.860000 198.850000 60.060000 199.050000 ;
        RECT 59.860000 199.250000 60.060000 199.450000 ;
        RECT 59.860000 199.650000 60.060000 199.850000 ;
        RECT 60.230000  25.910000 60.430000  26.110000 ;
        RECT 60.230000  26.340000 60.430000  26.540000 ;
        RECT 60.230000  26.770000 60.430000  26.970000 ;
        RECT 60.230000  27.200000 60.430000  27.400000 ;
        RECT 60.230000  27.630000 60.430000  27.830000 ;
        RECT 60.230000  28.060000 60.430000  28.260000 ;
        RECT 60.230000  28.490000 60.430000  28.690000 ;
        RECT 60.230000  28.920000 60.430000  29.120000 ;
        RECT 60.230000  29.350000 60.430000  29.550000 ;
        RECT 60.230000  29.780000 60.430000  29.980000 ;
        RECT 60.230000  30.210000 60.430000  30.410000 ;
        RECT 60.260000 197.250000 60.460000 197.450000 ;
        RECT 60.260000 197.650000 60.460000 197.850000 ;
        RECT 60.260000 198.050000 60.460000 198.250000 ;
        RECT 60.260000 198.450000 60.460000 198.650000 ;
        RECT 60.260000 198.850000 60.460000 199.050000 ;
        RECT 60.260000 199.250000 60.460000 199.450000 ;
        RECT 60.260000 199.650000 60.460000 199.850000 ;
        RECT 60.635000  25.910000 60.835000  26.110000 ;
        RECT 60.635000  26.340000 60.835000  26.540000 ;
        RECT 60.635000  26.770000 60.835000  26.970000 ;
        RECT 60.635000  27.200000 60.835000  27.400000 ;
        RECT 60.635000  27.630000 60.835000  27.830000 ;
        RECT 60.635000  28.060000 60.835000  28.260000 ;
        RECT 60.635000  28.490000 60.835000  28.690000 ;
        RECT 60.635000  28.920000 60.835000  29.120000 ;
        RECT 60.635000  29.350000 60.835000  29.550000 ;
        RECT 60.635000  29.780000 60.835000  29.980000 ;
        RECT 60.635000  30.210000 60.835000  30.410000 ;
        RECT 60.660000 197.250000 60.860000 197.450000 ;
        RECT 60.660000 197.650000 60.860000 197.850000 ;
        RECT 60.660000 198.050000 60.860000 198.250000 ;
        RECT 60.660000 198.450000 60.860000 198.650000 ;
        RECT 60.660000 198.850000 60.860000 199.050000 ;
        RECT 60.660000 199.250000 60.860000 199.450000 ;
        RECT 60.660000 199.650000 60.860000 199.850000 ;
        RECT 60.910000 196.295000 61.110000 196.495000 ;
        RECT 60.910000 196.705000 61.110000 196.905000 ;
        RECT 61.040000  25.910000 61.240000  26.110000 ;
        RECT 61.040000  26.340000 61.240000  26.540000 ;
        RECT 61.040000  26.770000 61.240000  26.970000 ;
        RECT 61.040000  27.200000 61.240000  27.400000 ;
        RECT 61.040000  27.630000 61.240000  27.830000 ;
        RECT 61.040000  28.060000 61.240000  28.260000 ;
        RECT 61.040000  28.490000 61.240000  28.690000 ;
        RECT 61.040000  28.920000 61.240000  29.120000 ;
        RECT 61.040000  29.350000 61.240000  29.550000 ;
        RECT 61.040000  29.780000 61.240000  29.980000 ;
        RECT 61.040000  30.210000 61.240000  30.410000 ;
        RECT 61.060000 197.250000 61.260000 197.450000 ;
        RECT 61.060000 197.650000 61.260000 197.850000 ;
        RECT 61.060000 198.050000 61.260000 198.250000 ;
        RECT 61.060000 198.450000 61.260000 198.650000 ;
        RECT 61.060000 198.850000 61.260000 199.050000 ;
        RECT 61.060000 199.250000 61.260000 199.450000 ;
        RECT 61.060000 199.650000 61.260000 199.850000 ;
        RECT 61.445000  25.910000 61.645000  26.110000 ;
        RECT 61.445000  26.340000 61.645000  26.540000 ;
        RECT 61.445000  26.770000 61.645000  26.970000 ;
        RECT 61.445000  27.200000 61.645000  27.400000 ;
        RECT 61.445000  27.630000 61.645000  27.830000 ;
        RECT 61.445000  28.060000 61.645000  28.260000 ;
        RECT 61.445000  28.490000 61.645000  28.690000 ;
        RECT 61.445000  28.920000 61.645000  29.120000 ;
        RECT 61.445000  29.350000 61.645000  29.550000 ;
        RECT 61.445000  29.780000 61.645000  29.980000 ;
        RECT 61.445000  30.210000 61.645000  30.410000 ;
        RECT 61.590000 175.995000 61.790000 176.195000 ;
        RECT 61.590000 176.395000 61.790000 176.595000 ;
        RECT 61.590000 176.795000 61.790000 176.995000 ;
        RECT 61.590000 177.195000 61.790000 177.395000 ;
        RECT 61.590000 177.595000 61.790000 177.795000 ;
        RECT 61.590000 177.995000 61.790000 178.195000 ;
        RECT 61.590000 178.395000 61.790000 178.595000 ;
        RECT 61.590000 178.795000 61.790000 178.995000 ;
        RECT 61.590000 179.195000 61.790000 179.395000 ;
        RECT 61.590000 179.595000 61.790000 179.795000 ;
        RECT 61.590000 179.995000 61.790000 180.195000 ;
        RECT 61.590000 180.395000 61.790000 180.595000 ;
        RECT 61.590000 180.795000 61.790000 180.995000 ;
        RECT 61.590000 181.195000 61.790000 181.395000 ;
        RECT 61.590000 181.595000 61.790000 181.795000 ;
        RECT 61.590000 181.995000 61.790000 182.195000 ;
        RECT 61.590000 182.395000 61.790000 182.595000 ;
        RECT 61.590000 182.795000 61.790000 182.995000 ;
        RECT 61.590000 183.195000 61.790000 183.395000 ;
        RECT 61.590000 183.595000 61.790000 183.795000 ;
        RECT 61.590000 183.995000 61.790000 184.195000 ;
        RECT 61.590000 184.395000 61.790000 184.595000 ;
        RECT 61.590000 184.795000 61.790000 184.995000 ;
        RECT 61.590000 185.195000 61.790000 185.395000 ;
        RECT 61.590000 185.595000 61.790000 185.795000 ;
        RECT 61.590000 185.995000 61.790000 186.195000 ;
        RECT 61.590000 186.395000 61.790000 186.595000 ;
        RECT 61.590000 186.795000 61.790000 186.995000 ;
        RECT 61.590000 187.195000 61.790000 187.395000 ;
        RECT 61.590000 187.595000 61.790000 187.795000 ;
        RECT 61.590000 187.995000 61.790000 188.195000 ;
        RECT 61.590000 188.395000 61.790000 188.595000 ;
        RECT 61.590000 188.795000 61.790000 188.995000 ;
        RECT 61.590000 189.195000 61.790000 189.395000 ;
        RECT 61.590000 189.595000 61.790000 189.795000 ;
        RECT 61.590000 189.995000 61.790000 190.195000 ;
        RECT 61.590000 190.395000 61.790000 190.595000 ;
        RECT 61.590000 190.795000 61.790000 190.995000 ;
        RECT 61.590000 191.195000 61.790000 191.395000 ;
        RECT 61.590000 191.595000 61.790000 191.795000 ;
        RECT 61.590000 191.995000 61.790000 192.195000 ;
        RECT 61.590000 192.395000 61.790000 192.595000 ;
        RECT 61.590000 192.795000 61.790000 192.995000 ;
        RECT 61.590000 193.195000 61.790000 193.395000 ;
        RECT 61.590000 193.595000 61.790000 193.795000 ;
        RECT 61.590000 193.995000 61.790000 194.195000 ;
        RECT 61.590000 194.395000 61.790000 194.595000 ;
        RECT 61.590000 194.795000 61.790000 194.995000 ;
        RECT 61.590000 195.200000 61.790000 195.400000 ;
        RECT 61.590000 195.605000 61.790000 195.805000 ;
        RECT 61.590000 196.010000 61.790000 196.210000 ;
        RECT 61.590000 196.415000 61.790000 196.615000 ;
        RECT 61.590000 196.820000 61.790000 197.020000 ;
        RECT 61.590000 197.225000 61.790000 197.425000 ;
        RECT 61.590000 197.630000 61.790000 197.830000 ;
        RECT 61.590000 198.035000 61.790000 198.235000 ;
        RECT 61.590000 198.440000 61.790000 198.640000 ;
        RECT 61.590000 198.845000 61.790000 199.045000 ;
        RECT 61.590000 199.250000 61.790000 199.450000 ;
        RECT 61.590000 199.655000 61.790000 199.855000 ;
        RECT 61.850000  25.910000 62.050000  26.110000 ;
        RECT 61.850000  26.340000 62.050000  26.540000 ;
        RECT 61.850000  26.770000 62.050000  26.970000 ;
        RECT 61.850000  27.200000 62.050000  27.400000 ;
        RECT 61.850000  27.630000 62.050000  27.830000 ;
        RECT 61.850000  28.060000 62.050000  28.260000 ;
        RECT 61.850000  28.490000 62.050000  28.690000 ;
        RECT 61.850000  28.920000 62.050000  29.120000 ;
        RECT 61.850000  29.350000 62.050000  29.550000 ;
        RECT 61.850000  29.780000 62.050000  29.980000 ;
        RECT 61.850000  30.210000 62.050000  30.410000 ;
        RECT 61.990000 175.995000 62.190000 176.195000 ;
        RECT 61.990000 176.395000 62.190000 176.595000 ;
        RECT 61.990000 176.795000 62.190000 176.995000 ;
        RECT 61.990000 177.195000 62.190000 177.395000 ;
        RECT 61.990000 177.595000 62.190000 177.795000 ;
        RECT 61.990000 177.995000 62.190000 178.195000 ;
        RECT 61.990000 178.395000 62.190000 178.595000 ;
        RECT 61.990000 178.795000 62.190000 178.995000 ;
        RECT 61.990000 179.195000 62.190000 179.395000 ;
        RECT 61.990000 179.595000 62.190000 179.795000 ;
        RECT 61.990000 179.995000 62.190000 180.195000 ;
        RECT 61.990000 180.395000 62.190000 180.595000 ;
        RECT 61.990000 180.795000 62.190000 180.995000 ;
        RECT 61.990000 181.195000 62.190000 181.395000 ;
        RECT 61.990000 181.595000 62.190000 181.795000 ;
        RECT 61.990000 181.995000 62.190000 182.195000 ;
        RECT 61.990000 182.395000 62.190000 182.595000 ;
        RECT 61.990000 182.795000 62.190000 182.995000 ;
        RECT 61.990000 183.195000 62.190000 183.395000 ;
        RECT 61.990000 183.595000 62.190000 183.795000 ;
        RECT 61.990000 183.995000 62.190000 184.195000 ;
        RECT 61.990000 184.395000 62.190000 184.595000 ;
        RECT 61.990000 184.795000 62.190000 184.995000 ;
        RECT 61.990000 185.195000 62.190000 185.395000 ;
        RECT 61.990000 185.595000 62.190000 185.795000 ;
        RECT 61.990000 185.995000 62.190000 186.195000 ;
        RECT 61.990000 186.395000 62.190000 186.595000 ;
        RECT 61.990000 186.795000 62.190000 186.995000 ;
        RECT 61.990000 187.195000 62.190000 187.395000 ;
        RECT 61.990000 187.595000 62.190000 187.795000 ;
        RECT 61.990000 187.995000 62.190000 188.195000 ;
        RECT 61.990000 188.395000 62.190000 188.595000 ;
        RECT 61.990000 188.795000 62.190000 188.995000 ;
        RECT 61.990000 189.195000 62.190000 189.395000 ;
        RECT 61.990000 189.595000 62.190000 189.795000 ;
        RECT 61.990000 189.995000 62.190000 190.195000 ;
        RECT 61.990000 190.395000 62.190000 190.595000 ;
        RECT 61.990000 190.795000 62.190000 190.995000 ;
        RECT 61.990000 191.195000 62.190000 191.395000 ;
        RECT 61.990000 191.595000 62.190000 191.795000 ;
        RECT 61.990000 191.995000 62.190000 192.195000 ;
        RECT 61.990000 192.395000 62.190000 192.595000 ;
        RECT 61.990000 192.795000 62.190000 192.995000 ;
        RECT 61.990000 193.195000 62.190000 193.395000 ;
        RECT 61.990000 193.595000 62.190000 193.795000 ;
        RECT 61.990000 193.995000 62.190000 194.195000 ;
        RECT 61.990000 194.395000 62.190000 194.595000 ;
        RECT 61.990000 194.795000 62.190000 194.995000 ;
        RECT 61.990000 195.200000 62.190000 195.400000 ;
        RECT 61.990000 195.605000 62.190000 195.805000 ;
        RECT 61.990000 196.010000 62.190000 196.210000 ;
        RECT 61.990000 196.415000 62.190000 196.615000 ;
        RECT 61.990000 196.820000 62.190000 197.020000 ;
        RECT 61.990000 197.225000 62.190000 197.425000 ;
        RECT 61.990000 197.630000 62.190000 197.830000 ;
        RECT 61.990000 198.035000 62.190000 198.235000 ;
        RECT 61.990000 198.440000 62.190000 198.640000 ;
        RECT 61.990000 198.845000 62.190000 199.045000 ;
        RECT 61.990000 199.250000 62.190000 199.450000 ;
        RECT 61.990000 199.655000 62.190000 199.855000 ;
        RECT 62.255000  25.910000 62.455000  26.110000 ;
        RECT 62.255000  26.340000 62.455000  26.540000 ;
        RECT 62.255000  26.770000 62.455000  26.970000 ;
        RECT 62.255000  27.200000 62.455000  27.400000 ;
        RECT 62.255000  27.630000 62.455000  27.830000 ;
        RECT 62.255000  28.060000 62.455000  28.260000 ;
        RECT 62.255000  28.490000 62.455000  28.690000 ;
        RECT 62.255000  28.920000 62.455000  29.120000 ;
        RECT 62.255000  29.350000 62.455000  29.550000 ;
        RECT 62.255000  29.780000 62.455000  29.980000 ;
        RECT 62.255000  30.210000 62.455000  30.410000 ;
        RECT 62.390000 175.995000 62.590000 176.195000 ;
        RECT 62.390000 176.395000 62.590000 176.595000 ;
        RECT 62.390000 176.795000 62.590000 176.995000 ;
        RECT 62.390000 177.195000 62.590000 177.395000 ;
        RECT 62.390000 177.595000 62.590000 177.795000 ;
        RECT 62.390000 177.995000 62.590000 178.195000 ;
        RECT 62.390000 178.395000 62.590000 178.595000 ;
        RECT 62.390000 178.795000 62.590000 178.995000 ;
        RECT 62.390000 179.195000 62.590000 179.395000 ;
        RECT 62.390000 179.595000 62.590000 179.795000 ;
        RECT 62.390000 179.995000 62.590000 180.195000 ;
        RECT 62.390000 180.395000 62.590000 180.595000 ;
        RECT 62.390000 180.795000 62.590000 180.995000 ;
        RECT 62.390000 181.195000 62.590000 181.395000 ;
        RECT 62.390000 181.595000 62.590000 181.795000 ;
        RECT 62.390000 181.995000 62.590000 182.195000 ;
        RECT 62.390000 182.395000 62.590000 182.595000 ;
        RECT 62.390000 182.795000 62.590000 182.995000 ;
        RECT 62.390000 183.195000 62.590000 183.395000 ;
        RECT 62.390000 183.595000 62.590000 183.795000 ;
        RECT 62.390000 183.995000 62.590000 184.195000 ;
        RECT 62.390000 184.395000 62.590000 184.595000 ;
        RECT 62.390000 184.795000 62.590000 184.995000 ;
        RECT 62.390000 185.195000 62.590000 185.395000 ;
        RECT 62.390000 185.595000 62.590000 185.795000 ;
        RECT 62.390000 185.995000 62.590000 186.195000 ;
        RECT 62.390000 186.395000 62.590000 186.595000 ;
        RECT 62.390000 186.795000 62.590000 186.995000 ;
        RECT 62.390000 187.195000 62.590000 187.395000 ;
        RECT 62.390000 187.595000 62.590000 187.795000 ;
        RECT 62.390000 187.995000 62.590000 188.195000 ;
        RECT 62.390000 188.395000 62.590000 188.595000 ;
        RECT 62.390000 188.795000 62.590000 188.995000 ;
        RECT 62.390000 189.195000 62.590000 189.395000 ;
        RECT 62.390000 189.595000 62.590000 189.795000 ;
        RECT 62.390000 189.995000 62.590000 190.195000 ;
        RECT 62.390000 190.395000 62.590000 190.595000 ;
        RECT 62.390000 190.795000 62.590000 190.995000 ;
        RECT 62.390000 191.195000 62.590000 191.395000 ;
        RECT 62.390000 191.595000 62.590000 191.795000 ;
        RECT 62.390000 191.995000 62.590000 192.195000 ;
        RECT 62.390000 192.395000 62.590000 192.595000 ;
        RECT 62.390000 192.795000 62.590000 192.995000 ;
        RECT 62.390000 193.195000 62.590000 193.395000 ;
        RECT 62.390000 193.595000 62.590000 193.795000 ;
        RECT 62.390000 193.995000 62.590000 194.195000 ;
        RECT 62.390000 194.395000 62.590000 194.595000 ;
        RECT 62.390000 194.795000 62.590000 194.995000 ;
        RECT 62.390000 195.200000 62.590000 195.400000 ;
        RECT 62.390000 195.605000 62.590000 195.805000 ;
        RECT 62.390000 196.010000 62.590000 196.210000 ;
        RECT 62.390000 196.415000 62.590000 196.615000 ;
        RECT 62.390000 196.820000 62.590000 197.020000 ;
        RECT 62.390000 197.225000 62.590000 197.425000 ;
        RECT 62.390000 197.630000 62.590000 197.830000 ;
        RECT 62.390000 198.035000 62.590000 198.235000 ;
        RECT 62.390000 198.440000 62.590000 198.640000 ;
        RECT 62.390000 198.845000 62.590000 199.045000 ;
        RECT 62.390000 199.250000 62.590000 199.450000 ;
        RECT 62.390000 199.655000 62.590000 199.855000 ;
        RECT 62.660000  25.910000 62.860000  26.110000 ;
        RECT 62.660000  26.340000 62.860000  26.540000 ;
        RECT 62.660000  26.770000 62.860000  26.970000 ;
        RECT 62.660000  27.200000 62.860000  27.400000 ;
        RECT 62.660000  27.630000 62.860000  27.830000 ;
        RECT 62.660000  28.060000 62.860000  28.260000 ;
        RECT 62.660000  28.490000 62.860000  28.690000 ;
        RECT 62.660000  28.920000 62.860000  29.120000 ;
        RECT 62.660000  29.350000 62.860000  29.550000 ;
        RECT 62.660000  29.780000 62.860000  29.980000 ;
        RECT 62.660000  30.210000 62.860000  30.410000 ;
        RECT 62.790000 175.995000 62.990000 176.195000 ;
        RECT 62.790000 176.395000 62.990000 176.595000 ;
        RECT 62.790000 176.795000 62.990000 176.995000 ;
        RECT 62.790000 177.195000 62.990000 177.395000 ;
        RECT 62.790000 177.595000 62.990000 177.795000 ;
        RECT 62.790000 177.995000 62.990000 178.195000 ;
        RECT 62.790000 178.395000 62.990000 178.595000 ;
        RECT 62.790000 178.795000 62.990000 178.995000 ;
        RECT 62.790000 179.195000 62.990000 179.395000 ;
        RECT 62.790000 179.595000 62.990000 179.795000 ;
        RECT 62.790000 179.995000 62.990000 180.195000 ;
        RECT 62.790000 180.395000 62.990000 180.595000 ;
        RECT 62.790000 180.795000 62.990000 180.995000 ;
        RECT 62.790000 181.195000 62.990000 181.395000 ;
        RECT 62.790000 181.595000 62.990000 181.795000 ;
        RECT 62.790000 181.995000 62.990000 182.195000 ;
        RECT 62.790000 182.395000 62.990000 182.595000 ;
        RECT 62.790000 182.795000 62.990000 182.995000 ;
        RECT 62.790000 183.195000 62.990000 183.395000 ;
        RECT 62.790000 183.595000 62.990000 183.795000 ;
        RECT 62.790000 183.995000 62.990000 184.195000 ;
        RECT 62.790000 184.395000 62.990000 184.595000 ;
        RECT 62.790000 184.795000 62.990000 184.995000 ;
        RECT 62.790000 185.195000 62.990000 185.395000 ;
        RECT 62.790000 185.595000 62.990000 185.795000 ;
        RECT 62.790000 185.995000 62.990000 186.195000 ;
        RECT 62.790000 186.395000 62.990000 186.595000 ;
        RECT 62.790000 186.795000 62.990000 186.995000 ;
        RECT 62.790000 187.195000 62.990000 187.395000 ;
        RECT 62.790000 187.595000 62.990000 187.795000 ;
        RECT 62.790000 187.995000 62.990000 188.195000 ;
        RECT 62.790000 188.395000 62.990000 188.595000 ;
        RECT 62.790000 188.795000 62.990000 188.995000 ;
        RECT 62.790000 189.195000 62.990000 189.395000 ;
        RECT 62.790000 189.595000 62.990000 189.795000 ;
        RECT 62.790000 189.995000 62.990000 190.195000 ;
        RECT 62.790000 190.395000 62.990000 190.595000 ;
        RECT 62.790000 190.795000 62.990000 190.995000 ;
        RECT 62.790000 191.195000 62.990000 191.395000 ;
        RECT 62.790000 191.595000 62.990000 191.795000 ;
        RECT 62.790000 191.995000 62.990000 192.195000 ;
        RECT 62.790000 192.395000 62.990000 192.595000 ;
        RECT 62.790000 192.795000 62.990000 192.995000 ;
        RECT 62.790000 193.195000 62.990000 193.395000 ;
        RECT 62.790000 193.595000 62.990000 193.795000 ;
        RECT 62.790000 193.995000 62.990000 194.195000 ;
        RECT 62.790000 194.395000 62.990000 194.595000 ;
        RECT 62.790000 194.795000 62.990000 194.995000 ;
        RECT 62.790000 195.200000 62.990000 195.400000 ;
        RECT 62.790000 195.605000 62.990000 195.805000 ;
        RECT 62.790000 196.010000 62.990000 196.210000 ;
        RECT 62.790000 196.415000 62.990000 196.615000 ;
        RECT 62.790000 196.820000 62.990000 197.020000 ;
        RECT 62.790000 197.225000 62.990000 197.425000 ;
        RECT 62.790000 197.630000 62.990000 197.830000 ;
        RECT 62.790000 198.035000 62.990000 198.235000 ;
        RECT 62.790000 198.440000 62.990000 198.640000 ;
        RECT 62.790000 198.845000 62.990000 199.045000 ;
        RECT 62.790000 199.250000 62.990000 199.450000 ;
        RECT 62.790000 199.655000 62.990000 199.855000 ;
        RECT 63.065000  25.910000 63.265000  26.110000 ;
        RECT 63.065000  26.340000 63.265000  26.540000 ;
        RECT 63.065000  26.770000 63.265000  26.970000 ;
        RECT 63.065000  27.200000 63.265000  27.400000 ;
        RECT 63.065000  27.630000 63.265000  27.830000 ;
        RECT 63.065000  28.060000 63.265000  28.260000 ;
        RECT 63.065000  28.490000 63.265000  28.690000 ;
        RECT 63.065000  28.920000 63.265000  29.120000 ;
        RECT 63.065000  29.350000 63.265000  29.550000 ;
        RECT 63.065000  29.780000 63.265000  29.980000 ;
        RECT 63.065000  30.210000 63.265000  30.410000 ;
        RECT 63.190000 175.995000 63.390000 176.195000 ;
        RECT 63.190000 176.395000 63.390000 176.595000 ;
        RECT 63.190000 176.795000 63.390000 176.995000 ;
        RECT 63.190000 177.195000 63.390000 177.395000 ;
        RECT 63.190000 177.595000 63.390000 177.795000 ;
        RECT 63.190000 177.995000 63.390000 178.195000 ;
        RECT 63.190000 178.395000 63.390000 178.595000 ;
        RECT 63.190000 178.795000 63.390000 178.995000 ;
        RECT 63.190000 179.195000 63.390000 179.395000 ;
        RECT 63.190000 179.595000 63.390000 179.795000 ;
        RECT 63.190000 179.995000 63.390000 180.195000 ;
        RECT 63.190000 180.395000 63.390000 180.595000 ;
        RECT 63.190000 180.795000 63.390000 180.995000 ;
        RECT 63.190000 181.195000 63.390000 181.395000 ;
        RECT 63.190000 181.595000 63.390000 181.795000 ;
        RECT 63.190000 181.995000 63.390000 182.195000 ;
        RECT 63.190000 182.395000 63.390000 182.595000 ;
        RECT 63.190000 182.795000 63.390000 182.995000 ;
        RECT 63.190000 183.195000 63.390000 183.395000 ;
        RECT 63.190000 183.595000 63.390000 183.795000 ;
        RECT 63.190000 183.995000 63.390000 184.195000 ;
        RECT 63.190000 184.395000 63.390000 184.595000 ;
        RECT 63.190000 184.795000 63.390000 184.995000 ;
        RECT 63.190000 185.195000 63.390000 185.395000 ;
        RECT 63.190000 185.595000 63.390000 185.795000 ;
        RECT 63.190000 185.995000 63.390000 186.195000 ;
        RECT 63.190000 186.395000 63.390000 186.595000 ;
        RECT 63.190000 186.795000 63.390000 186.995000 ;
        RECT 63.190000 187.195000 63.390000 187.395000 ;
        RECT 63.190000 187.595000 63.390000 187.795000 ;
        RECT 63.190000 187.995000 63.390000 188.195000 ;
        RECT 63.190000 188.395000 63.390000 188.595000 ;
        RECT 63.190000 188.795000 63.390000 188.995000 ;
        RECT 63.190000 189.195000 63.390000 189.395000 ;
        RECT 63.190000 189.595000 63.390000 189.795000 ;
        RECT 63.190000 189.995000 63.390000 190.195000 ;
        RECT 63.190000 190.395000 63.390000 190.595000 ;
        RECT 63.190000 190.795000 63.390000 190.995000 ;
        RECT 63.190000 191.195000 63.390000 191.395000 ;
        RECT 63.190000 191.595000 63.390000 191.795000 ;
        RECT 63.190000 191.995000 63.390000 192.195000 ;
        RECT 63.190000 192.395000 63.390000 192.595000 ;
        RECT 63.190000 192.795000 63.390000 192.995000 ;
        RECT 63.190000 193.195000 63.390000 193.395000 ;
        RECT 63.190000 193.595000 63.390000 193.795000 ;
        RECT 63.190000 193.995000 63.390000 194.195000 ;
        RECT 63.190000 194.395000 63.390000 194.595000 ;
        RECT 63.190000 194.795000 63.390000 194.995000 ;
        RECT 63.190000 195.200000 63.390000 195.400000 ;
        RECT 63.190000 195.605000 63.390000 195.805000 ;
        RECT 63.190000 196.010000 63.390000 196.210000 ;
        RECT 63.190000 196.415000 63.390000 196.615000 ;
        RECT 63.190000 196.820000 63.390000 197.020000 ;
        RECT 63.190000 197.225000 63.390000 197.425000 ;
        RECT 63.190000 197.630000 63.390000 197.830000 ;
        RECT 63.190000 198.035000 63.390000 198.235000 ;
        RECT 63.190000 198.440000 63.390000 198.640000 ;
        RECT 63.190000 198.845000 63.390000 199.045000 ;
        RECT 63.190000 199.250000 63.390000 199.450000 ;
        RECT 63.190000 199.655000 63.390000 199.855000 ;
        RECT 63.470000  25.910000 63.670000  26.110000 ;
        RECT 63.470000  26.340000 63.670000  26.540000 ;
        RECT 63.470000  26.770000 63.670000  26.970000 ;
        RECT 63.470000  27.200000 63.670000  27.400000 ;
        RECT 63.470000  27.630000 63.670000  27.830000 ;
        RECT 63.470000  28.060000 63.670000  28.260000 ;
        RECT 63.470000  28.490000 63.670000  28.690000 ;
        RECT 63.470000  28.920000 63.670000  29.120000 ;
        RECT 63.470000  29.350000 63.670000  29.550000 ;
        RECT 63.470000  29.780000 63.670000  29.980000 ;
        RECT 63.470000  30.210000 63.670000  30.410000 ;
        RECT 63.590000 175.995000 63.790000 176.195000 ;
        RECT 63.590000 176.395000 63.790000 176.595000 ;
        RECT 63.590000 176.795000 63.790000 176.995000 ;
        RECT 63.590000 177.195000 63.790000 177.395000 ;
        RECT 63.590000 177.595000 63.790000 177.795000 ;
        RECT 63.590000 177.995000 63.790000 178.195000 ;
        RECT 63.590000 178.395000 63.790000 178.595000 ;
        RECT 63.590000 178.795000 63.790000 178.995000 ;
        RECT 63.590000 179.195000 63.790000 179.395000 ;
        RECT 63.590000 179.595000 63.790000 179.795000 ;
        RECT 63.590000 179.995000 63.790000 180.195000 ;
        RECT 63.590000 180.395000 63.790000 180.595000 ;
        RECT 63.590000 180.795000 63.790000 180.995000 ;
        RECT 63.590000 181.195000 63.790000 181.395000 ;
        RECT 63.590000 181.595000 63.790000 181.795000 ;
        RECT 63.590000 181.995000 63.790000 182.195000 ;
        RECT 63.590000 182.395000 63.790000 182.595000 ;
        RECT 63.590000 182.795000 63.790000 182.995000 ;
        RECT 63.590000 183.195000 63.790000 183.395000 ;
        RECT 63.590000 183.595000 63.790000 183.795000 ;
        RECT 63.590000 183.995000 63.790000 184.195000 ;
        RECT 63.590000 184.395000 63.790000 184.595000 ;
        RECT 63.590000 184.795000 63.790000 184.995000 ;
        RECT 63.590000 185.195000 63.790000 185.395000 ;
        RECT 63.590000 185.595000 63.790000 185.795000 ;
        RECT 63.590000 185.995000 63.790000 186.195000 ;
        RECT 63.590000 186.395000 63.790000 186.595000 ;
        RECT 63.590000 186.795000 63.790000 186.995000 ;
        RECT 63.590000 187.195000 63.790000 187.395000 ;
        RECT 63.590000 187.595000 63.790000 187.795000 ;
        RECT 63.590000 187.995000 63.790000 188.195000 ;
        RECT 63.590000 188.395000 63.790000 188.595000 ;
        RECT 63.590000 188.795000 63.790000 188.995000 ;
        RECT 63.590000 189.195000 63.790000 189.395000 ;
        RECT 63.590000 189.595000 63.790000 189.795000 ;
        RECT 63.590000 189.995000 63.790000 190.195000 ;
        RECT 63.590000 190.395000 63.790000 190.595000 ;
        RECT 63.590000 190.795000 63.790000 190.995000 ;
        RECT 63.590000 191.195000 63.790000 191.395000 ;
        RECT 63.590000 191.595000 63.790000 191.795000 ;
        RECT 63.590000 191.995000 63.790000 192.195000 ;
        RECT 63.590000 192.395000 63.790000 192.595000 ;
        RECT 63.590000 192.795000 63.790000 192.995000 ;
        RECT 63.590000 193.195000 63.790000 193.395000 ;
        RECT 63.590000 193.595000 63.790000 193.795000 ;
        RECT 63.590000 193.995000 63.790000 194.195000 ;
        RECT 63.590000 194.395000 63.790000 194.595000 ;
        RECT 63.590000 194.795000 63.790000 194.995000 ;
        RECT 63.590000 195.200000 63.790000 195.400000 ;
        RECT 63.590000 195.605000 63.790000 195.805000 ;
        RECT 63.590000 196.010000 63.790000 196.210000 ;
        RECT 63.590000 196.415000 63.790000 196.615000 ;
        RECT 63.590000 196.820000 63.790000 197.020000 ;
        RECT 63.590000 197.225000 63.790000 197.425000 ;
        RECT 63.590000 197.630000 63.790000 197.830000 ;
        RECT 63.590000 198.035000 63.790000 198.235000 ;
        RECT 63.590000 198.440000 63.790000 198.640000 ;
        RECT 63.590000 198.845000 63.790000 199.045000 ;
        RECT 63.590000 199.250000 63.790000 199.450000 ;
        RECT 63.590000 199.655000 63.790000 199.855000 ;
        RECT 63.875000  25.910000 64.075000  26.110000 ;
        RECT 63.875000  26.340000 64.075000  26.540000 ;
        RECT 63.875000  26.770000 64.075000  26.970000 ;
        RECT 63.875000  27.200000 64.075000  27.400000 ;
        RECT 63.875000  27.630000 64.075000  27.830000 ;
        RECT 63.875000  28.060000 64.075000  28.260000 ;
        RECT 63.875000  28.490000 64.075000  28.690000 ;
        RECT 63.875000  28.920000 64.075000  29.120000 ;
        RECT 63.875000  29.350000 64.075000  29.550000 ;
        RECT 63.875000  29.780000 64.075000  29.980000 ;
        RECT 63.875000  30.210000 64.075000  30.410000 ;
        RECT 63.990000 175.995000 64.190000 176.195000 ;
        RECT 63.990000 176.395000 64.190000 176.595000 ;
        RECT 63.990000 176.795000 64.190000 176.995000 ;
        RECT 63.990000 177.195000 64.190000 177.395000 ;
        RECT 63.990000 177.595000 64.190000 177.795000 ;
        RECT 63.990000 177.995000 64.190000 178.195000 ;
        RECT 63.990000 178.395000 64.190000 178.595000 ;
        RECT 63.990000 178.795000 64.190000 178.995000 ;
        RECT 63.990000 179.195000 64.190000 179.395000 ;
        RECT 63.990000 179.595000 64.190000 179.795000 ;
        RECT 63.990000 179.995000 64.190000 180.195000 ;
        RECT 63.990000 180.395000 64.190000 180.595000 ;
        RECT 63.990000 180.795000 64.190000 180.995000 ;
        RECT 63.990000 181.195000 64.190000 181.395000 ;
        RECT 63.990000 181.595000 64.190000 181.795000 ;
        RECT 63.990000 181.995000 64.190000 182.195000 ;
        RECT 63.990000 182.395000 64.190000 182.595000 ;
        RECT 63.990000 182.795000 64.190000 182.995000 ;
        RECT 63.990000 183.195000 64.190000 183.395000 ;
        RECT 63.990000 183.595000 64.190000 183.795000 ;
        RECT 63.990000 183.995000 64.190000 184.195000 ;
        RECT 63.990000 184.395000 64.190000 184.595000 ;
        RECT 63.990000 184.795000 64.190000 184.995000 ;
        RECT 63.990000 185.195000 64.190000 185.395000 ;
        RECT 63.990000 185.595000 64.190000 185.795000 ;
        RECT 63.990000 185.995000 64.190000 186.195000 ;
        RECT 63.990000 186.395000 64.190000 186.595000 ;
        RECT 63.990000 186.795000 64.190000 186.995000 ;
        RECT 63.990000 187.195000 64.190000 187.395000 ;
        RECT 63.990000 187.595000 64.190000 187.795000 ;
        RECT 63.990000 187.995000 64.190000 188.195000 ;
        RECT 63.990000 188.395000 64.190000 188.595000 ;
        RECT 63.990000 188.795000 64.190000 188.995000 ;
        RECT 63.990000 189.195000 64.190000 189.395000 ;
        RECT 63.990000 189.595000 64.190000 189.795000 ;
        RECT 63.990000 189.995000 64.190000 190.195000 ;
        RECT 63.990000 190.395000 64.190000 190.595000 ;
        RECT 63.990000 190.795000 64.190000 190.995000 ;
        RECT 63.990000 191.195000 64.190000 191.395000 ;
        RECT 63.990000 191.595000 64.190000 191.795000 ;
        RECT 63.990000 191.995000 64.190000 192.195000 ;
        RECT 63.990000 192.395000 64.190000 192.595000 ;
        RECT 63.990000 192.795000 64.190000 192.995000 ;
        RECT 63.990000 193.195000 64.190000 193.395000 ;
        RECT 63.990000 193.595000 64.190000 193.795000 ;
        RECT 63.990000 193.995000 64.190000 194.195000 ;
        RECT 63.990000 194.395000 64.190000 194.595000 ;
        RECT 63.990000 194.795000 64.190000 194.995000 ;
        RECT 63.990000 195.200000 64.190000 195.400000 ;
        RECT 63.990000 195.605000 64.190000 195.805000 ;
        RECT 63.990000 196.010000 64.190000 196.210000 ;
        RECT 63.990000 196.415000 64.190000 196.615000 ;
        RECT 63.990000 196.820000 64.190000 197.020000 ;
        RECT 63.990000 197.225000 64.190000 197.425000 ;
        RECT 63.990000 197.630000 64.190000 197.830000 ;
        RECT 63.990000 198.035000 64.190000 198.235000 ;
        RECT 63.990000 198.440000 64.190000 198.640000 ;
        RECT 63.990000 198.845000 64.190000 199.045000 ;
        RECT 63.990000 199.250000 64.190000 199.450000 ;
        RECT 63.990000 199.655000 64.190000 199.855000 ;
        RECT 64.280000  25.910000 64.480000  26.110000 ;
        RECT 64.280000  26.340000 64.480000  26.540000 ;
        RECT 64.280000  26.770000 64.480000  26.970000 ;
        RECT 64.280000  27.200000 64.480000  27.400000 ;
        RECT 64.280000  27.630000 64.480000  27.830000 ;
        RECT 64.280000  28.060000 64.480000  28.260000 ;
        RECT 64.280000  28.490000 64.480000  28.690000 ;
        RECT 64.280000  28.920000 64.480000  29.120000 ;
        RECT 64.280000  29.350000 64.480000  29.550000 ;
        RECT 64.280000  29.780000 64.480000  29.980000 ;
        RECT 64.280000  30.210000 64.480000  30.410000 ;
        RECT 64.390000 175.995000 64.590000 176.195000 ;
        RECT 64.390000 176.395000 64.590000 176.595000 ;
        RECT 64.390000 176.795000 64.590000 176.995000 ;
        RECT 64.390000 177.195000 64.590000 177.395000 ;
        RECT 64.390000 177.595000 64.590000 177.795000 ;
        RECT 64.390000 177.995000 64.590000 178.195000 ;
        RECT 64.390000 178.395000 64.590000 178.595000 ;
        RECT 64.390000 178.795000 64.590000 178.995000 ;
        RECT 64.390000 179.195000 64.590000 179.395000 ;
        RECT 64.390000 179.595000 64.590000 179.795000 ;
        RECT 64.390000 179.995000 64.590000 180.195000 ;
        RECT 64.390000 180.395000 64.590000 180.595000 ;
        RECT 64.390000 180.795000 64.590000 180.995000 ;
        RECT 64.390000 181.195000 64.590000 181.395000 ;
        RECT 64.390000 181.595000 64.590000 181.795000 ;
        RECT 64.390000 181.995000 64.590000 182.195000 ;
        RECT 64.390000 182.395000 64.590000 182.595000 ;
        RECT 64.390000 182.795000 64.590000 182.995000 ;
        RECT 64.390000 183.195000 64.590000 183.395000 ;
        RECT 64.390000 183.595000 64.590000 183.795000 ;
        RECT 64.390000 183.995000 64.590000 184.195000 ;
        RECT 64.390000 184.395000 64.590000 184.595000 ;
        RECT 64.390000 184.795000 64.590000 184.995000 ;
        RECT 64.390000 185.195000 64.590000 185.395000 ;
        RECT 64.390000 185.595000 64.590000 185.795000 ;
        RECT 64.390000 185.995000 64.590000 186.195000 ;
        RECT 64.390000 186.395000 64.590000 186.595000 ;
        RECT 64.390000 186.795000 64.590000 186.995000 ;
        RECT 64.390000 187.195000 64.590000 187.395000 ;
        RECT 64.390000 187.595000 64.590000 187.795000 ;
        RECT 64.390000 187.995000 64.590000 188.195000 ;
        RECT 64.390000 188.395000 64.590000 188.595000 ;
        RECT 64.390000 188.795000 64.590000 188.995000 ;
        RECT 64.390000 189.195000 64.590000 189.395000 ;
        RECT 64.390000 189.595000 64.590000 189.795000 ;
        RECT 64.390000 189.995000 64.590000 190.195000 ;
        RECT 64.390000 190.395000 64.590000 190.595000 ;
        RECT 64.390000 190.795000 64.590000 190.995000 ;
        RECT 64.390000 191.195000 64.590000 191.395000 ;
        RECT 64.390000 191.595000 64.590000 191.795000 ;
        RECT 64.390000 191.995000 64.590000 192.195000 ;
        RECT 64.390000 192.395000 64.590000 192.595000 ;
        RECT 64.390000 192.795000 64.590000 192.995000 ;
        RECT 64.390000 193.195000 64.590000 193.395000 ;
        RECT 64.390000 193.595000 64.590000 193.795000 ;
        RECT 64.390000 193.995000 64.590000 194.195000 ;
        RECT 64.390000 194.395000 64.590000 194.595000 ;
        RECT 64.390000 194.795000 64.590000 194.995000 ;
        RECT 64.390000 195.200000 64.590000 195.400000 ;
        RECT 64.390000 195.605000 64.590000 195.805000 ;
        RECT 64.390000 196.010000 64.590000 196.210000 ;
        RECT 64.390000 196.415000 64.590000 196.615000 ;
        RECT 64.390000 196.820000 64.590000 197.020000 ;
        RECT 64.390000 197.225000 64.590000 197.425000 ;
        RECT 64.390000 197.630000 64.590000 197.830000 ;
        RECT 64.390000 198.035000 64.590000 198.235000 ;
        RECT 64.390000 198.440000 64.590000 198.640000 ;
        RECT 64.390000 198.845000 64.590000 199.045000 ;
        RECT 64.390000 199.250000 64.590000 199.450000 ;
        RECT 64.390000 199.655000 64.590000 199.855000 ;
        RECT 64.685000  25.910000 64.885000  26.110000 ;
        RECT 64.685000  26.340000 64.885000  26.540000 ;
        RECT 64.685000  26.770000 64.885000  26.970000 ;
        RECT 64.685000  27.200000 64.885000  27.400000 ;
        RECT 64.685000  27.630000 64.885000  27.830000 ;
        RECT 64.685000  28.060000 64.885000  28.260000 ;
        RECT 64.685000  28.490000 64.885000  28.690000 ;
        RECT 64.685000  28.920000 64.885000  29.120000 ;
        RECT 64.685000  29.350000 64.885000  29.550000 ;
        RECT 64.685000  29.780000 64.885000  29.980000 ;
        RECT 64.685000  30.210000 64.885000  30.410000 ;
        RECT 64.790000 175.995000 64.990000 176.195000 ;
        RECT 64.790000 176.395000 64.990000 176.595000 ;
        RECT 64.790000 176.795000 64.990000 176.995000 ;
        RECT 64.790000 177.195000 64.990000 177.395000 ;
        RECT 64.790000 177.595000 64.990000 177.795000 ;
        RECT 64.790000 177.995000 64.990000 178.195000 ;
        RECT 64.790000 178.395000 64.990000 178.595000 ;
        RECT 64.790000 178.795000 64.990000 178.995000 ;
        RECT 64.790000 179.195000 64.990000 179.395000 ;
        RECT 64.790000 179.595000 64.990000 179.795000 ;
        RECT 64.790000 179.995000 64.990000 180.195000 ;
        RECT 64.790000 180.395000 64.990000 180.595000 ;
        RECT 64.790000 180.795000 64.990000 180.995000 ;
        RECT 64.790000 181.195000 64.990000 181.395000 ;
        RECT 64.790000 181.595000 64.990000 181.795000 ;
        RECT 64.790000 181.995000 64.990000 182.195000 ;
        RECT 64.790000 182.395000 64.990000 182.595000 ;
        RECT 64.790000 182.795000 64.990000 182.995000 ;
        RECT 64.790000 183.195000 64.990000 183.395000 ;
        RECT 64.790000 183.595000 64.990000 183.795000 ;
        RECT 64.790000 183.995000 64.990000 184.195000 ;
        RECT 64.790000 184.395000 64.990000 184.595000 ;
        RECT 64.790000 184.795000 64.990000 184.995000 ;
        RECT 64.790000 185.195000 64.990000 185.395000 ;
        RECT 64.790000 185.595000 64.990000 185.795000 ;
        RECT 64.790000 185.995000 64.990000 186.195000 ;
        RECT 64.790000 186.395000 64.990000 186.595000 ;
        RECT 64.790000 186.795000 64.990000 186.995000 ;
        RECT 64.790000 187.195000 64.990000 187.395000 ;
        RECT 64.790000 187.595000 64.990000 187.795000 ;
        RECT 64.790000 187.995000 64.990000 188.195000 ;
        RECT 64.790000 188.395000 64.990000 188.595000 ;
        RECT 64.790000 188.795000 64.990000 188.995000 ;
        RECT 64.790000 189.195000 64.990000 189.395000 ;
        RECT 64.790000 189.595000 64.990000 189.795000 ;
        RECT 64.790000 189.995000 64.990000 190.195000 ;
        RECT 64.790000 190.395000 64.990000 190.595000 ;
        RECT 64.790000 190.795000 64.990000 190.995000 ;
        RECT 64.790000 191.195000 64.990000 191.395000 ;
        RECT 64.790000 191.595000 64.990000 191.795000 ;
        RECT 64.790000 191.995000 64.990000 192.195000 ;
        RECT 64.790000 192.395000 64.990000 192.595000 ;
        RECT 64.790000 192.795000 64.990000 192.995000 ;
        RECT 64.790000 193.195000 64.990000 193.395000 ;
        RECT 64.790000 193.595000 64.990000 193.795000 ;
        RECT 64.790000 193.995000 64.990000 194.195000 ;
        RECT 64.790000 194.395000 64.990000 194.595000 ;
        RECT 64.790000 194.795000 64.990000 194.995000 ;
        RECT 64.790000 195.200000 64.990000 195.400000 ;
        RECT 64.790000 195.605000 64.990000 195.805000 ;
        RECT 64.790000 196.010000 64.990000 196.210000 ;
        RECT 64.790000 196.415000 64.990000 196.615000 ;
        RECT 64.790000 196.820000 64.990000 197.020000 ;
        RECT 64.790000 197.225000 64.990000 197.425000 ;
        RECT 64.790000 197.630000 64.990000 197.830000 ;
        RECT 64.790000 198.035000 64.990000 198.235000 ;
        RECT 64.790000 198.440000 64.990000 198.640000 ;
        RECT 64.790000 198.845000 64.990000 199.045000 ;
        RECT 64.790000 199.250000 64.990000 199.450000 ;
        RECT 64.790000 199.655000 64.990000 199.855000 ;
        RECT 65.090000  25.910000 65.290000  26.110000 ;
        RECT 65.090000  26.340000 65.290000  26.540000 ;
        RECT 65.090000  26.770000 65.290000  26.970000 ;
        RECT 65.090000  27.200000 65.290000  27.400000 ;
        RECT 65.090000  27.630000 65.290000  27.830000 ;
        RECT 65.090000  28.060000 65.290000  28.260000 ;
        RECT 65.090000  28.490000 65.290000  28.690000 ;
        RECT 65.090000  28.920000 65.290000  29.120000 ;
        RECT 65.090000  29.350000 65.290000  29.550000 ;
        RECT 65.090000  29.780000 65.290000  29.980000 ;
        RECT 65.090000  30.210000 65.290000  30.410000 ;
        RECT 65.190000 175.995000 65.390000 176.195000 ;
        RECT 65.190000 176.395000 65.390000 176.595000 ;
        RECT 65.190000 176.795000 65.390000 176.995000 ;
        RECT 65.190000 177.195000 65.390000 177.395000 ;
        RECT 65.190000 177.595000 65.390000 177.795000 ;
        RECT 65.190000 177.995000 65.390000 178.195000 ;
        RECT 65.190000 178.395000 65.390000 178.595000 ;
        RECT 65.190000 178.795000 65.390000 178.995000 ;
        RECT 65.190000 179.195000 65.390000 179.395000 ;
        RECT 65.190000 179.595000 65.390000 179.795000 ;
        RECT 65.190000 179.995000 65.390000 180.195000 ;
        RECT 65.190000 180.395000 65.390000 180.595000 ;
        RECT 65.190000 180.795000 65.390000 180.995000 ;
        RECT 65.190000 181.195000 65.390000 181.395000 ;
        RECT 65.190000 181.595000 65.390000 181.795000 ;
        RECT 65.190000 181.995000 65.390000 182.195000 ;
        RECT 65.190000 182.395000 65.390000 182.595000 ;
        RECT 65.190000 182.795000 65.390000 182.995000 ;
        RECT 65.190000 183.195000 65.390000 183.395000 ;
        RECT 65.190000 183.595000 65.390000 183.795000 ;
        RECT 65.190000 183.995000 65.390000 184.195000 ;
        RECT 65.190000 184.395000 65.390000 184.595000 ;
        RECT 65.190000 184.795000 65.390000 184.995000 ;
        RECT 65.190000 185.195000 65.390000 185.395000 ;
        RECT 65.190000 185.595000 65.390000 185.795000 ;
        RECT 65.190000 185.995000 65.390000 186.195000 ;
        RECT 65.190000 186.395000 65.390000 186.595000 ;
        RECT 65.190000 186.795000 65.390000 186.995000 ;
        RECT 65.190000 187.195000 65.390000 187.395000 ;
        RECT 65.190000 187.595000 65.390000 187.795000 ;
        RECT 65.190000 187.995000 65.390000 188.195000 ;
        RECT 65.190000 188.395000 65.390000 188.595000 ;
        RECT 65.190000 188.795000 65.390000 188.995000 ;
        RECT 65.190000 189.195000 65.390000 189.395000 ;
        RECT 65.190000 189.595000 65.390000 189.795000 ;
        RECT 65.190000 189.995000 65.390000 190.195000 ;
        RECT 65.190000 190.395000 65.390000 190.595000 ;
        RECT 65.190000 190.795000 65.390000 190.995000 ;
        RECT 65.190000 191.195000 65.390000 191.395000 ;
        RECT 65.190000 191.595000 65.390000 191.795000 ;
        RECT 65.190000 191.995000 65.390000 192.195000 ;
        RECT 65.190000 192.395000 65.390000 192.595000 ;
        RECT 65.190000 192.795000 65.390000 192.995000 ;
        RECT 65.190000 193.195000 65.390000 193.395000 ;
        RECT 65.190000 193.595000 65.390000 193.795000 ;
        RECT 65.190000 193.995000 65.390000 194.195000 ;
        RECT 65.190000 194.395000 65.390000 194.595000 ;
        RECT 65.190000 194.795000 65.390000 194.995000 ;
        RECT 65.190000 195.200000 65.390000 195.400000 ;
        RECT 65.190000 195.605000 65.390000 195.805000 ;
        RECT 65.190000 196.010000 65.390000 196.210000 ;
        RECT 65.190000 196.415000 65.390000 196.615000 ;
        RECT 65.190000 196.820000 65.390000 197.020000 ;
        RECT 65.190000 197.225000 65.390000 197.425000 ;
        RECT 65.190000 197.630000 65.390000 197.830000 ;
        RECT 65.190000 198.035000 65.390000 198.235000 ;
        RECT 65.190000 198.440000 65.390000 198.640000 ;
        RECT 65.190000 198.845000 65.390000 199.045000 ;
        RECT 65.190000 199.250000 65.390000 199.450000 ;
        RECT 65.190000 199.655000 65.390000 199.855000 ;
        RECT 65.495000  25.910000 65.695000  26.110000 ;
        RECT 65.495000  26.340000 65.695000  26.540000 ;
        RECT 65.495000  26.770000 65.695000  26.970000 ;
        RECT 65.495000  27.200000 65.695000  27.400000 ;
        RECT 65.495000  27.630000 65.695000  27.830000 ;
        RECT 65.495000  28.060000 65.695000  28.260000 ;
        RECT 65.495000  28.490000 65.695000  28.690000 ;
        RECT 65.495000  28.920000 65.695000  29.120000 ;
        RECT 65.495000  29.350000 65.695000  29.550000 ;
        RECT 65.495000  29.780000 65.695000  29.980000 ;
        RECT 65.495000  30.210000 65.695000  30.410000 ;
        RECT 65.590000 175.995000 65.790000 176.195000 ;
        RECT 65.590000 176.395000 65.790000 176.595000 ;
        RECT 65.590000 176.795000 65.790000 176.995000 ;
        RECT 65.590000 177.195000 65.790000 177.395000 ;
        RECT 65.590000 177.595000 65.790000 177.795000 ;
        RECT 65.590000 177.995000 65.790000 178.195000 ;
        RECT 65.590000 178.395000 65.790000 178.595000 ;
        RECT 65.590000 178.795000 65.790000 178.995000 ;
        RECT 65.590000 179.195000 65.790000 179.395000 ;
        RECT 65.590000 179.595000 65.790000 179.795000 ;
        RECT 65.590000 179.995000 65.790000 180.195000 ;
        RECT 65.590000 180.395000 65.790000 180.595000 ;
        RECT 65.590000 180.795000 65.790000 180.995000 ;
        RECT 65.590000 181.195000 65.790000 181.395000 ;
        RECT 65.590000 181.595000 65.790000 181.795000 ;
        RECT 65.590000 181.995000 65.790000 182.195000 ;
        RECT 65.590000 182.395000 65.790000 182.595000 ;
        RECT 65.590000 182.795000 65.790000 182.995000 ;
        RECT 65.590000 183.195000 65.790000 183.395000 ;
        RECT 65.590000 183.595000 65.790000 183.795000 ;
        RECT 65.590000 183.995000 65.790000 184.195000 ;
        RECT 65.590000 184.395000 65.790000 184.595000 ;
        RECT 65.590000 184.795000 65.790000 184.995000 ;
        RECT 65.590000 185.195000 65.790000 185.395000 ;
        RECT 65.590000 185.595000 65.790000 185.795000 ;
        RECT 65.590000 185.995000 65.790000 186.195000 ;
        RECT 65.590000 186.395000 65.790000 186.595000 ;
        RECT 65.590000 186.795000 65.790000 186.995000 ;
        RECT 65.590000 187.195000 65.790000 187.395000 ;
        RECT 65.590000 187.595000 65.790000 187.795000 ;
        RECT 65.590000 187.995000 65.790000 188.195000 ;
        RECT 65.590000 188.395000 65.790000 188.595000 ;
        RECT 65.590000 188.795000 65.790000 188.995000 ;
        RECT 65.590000 189.195000 65.790000 189.395000 ;
        RECT 65.590000 189.595000 65.790000 189.795000 ;
        RECT 65.590000 189.995000 65.790000 190.195000 ;
        RECT 65.590000 190.395000 65.790000 190.595000 ;
        RECT 65.590000 190.795000 65.790000 190.995000 ;
        RECT 65.590000 191.195000 65.790000 191.395000 ;
        RECT 65.590000 191.595000 65.790000 191.795000 ;
        RECT 65.590000 191.995000 65.790000 192.195000 ;
        RECT 65.590000 192.395000 65.790000 192.595000 ;
        RECT 65.590000 192.795000 65.790000 192.995000 ;
        RECT 65.590000 193.195000 65.790000 193.395000 ;
        RECT 65.590000 193.595000 65.790000 193.795000 ;
        RECT 65.590000 193.995000 65.790000 194.195000 ;
        RECT 65.590000 194.395000 65.790000 194.595000 ;
        RECT 65.590000 194.795000 65.790000 194.995000 ;
        RECT 65.590000 195.200000 65.790000 195.400000 ;
        RECT 65.590000 195.605000 65.790000 195.805000 ;
        RECT 65.590000 196.010000 65.790000 196.210000 ;
        RECT 65.590000 196.415000 65.790000 196.615000 ;
        RECT 65.590000 196.820000 65.790000 197.020000 ;
        RECT 65.590000 197.225000 65.790000 197.425000 ;
        RECT 65.590000 197.630000 65.790000 197.830000 ;
        RECT 65.590000 198.035000 65.790000 198.235000 ;
        RECT 65.590000 198.440000 65.790000 198.640000 ;
        RECT 65.590000 198.845000 65.790000 199.045000 ;
        RECT 65.590000 199.250000 65.790000 199.450000 ;
        RECT 65.590000 199.655000 65.790000 199.855000 ;
        RECT 65.900000  25.910000 66.100000  26.110000 ;
        RECT 65.900000  26.340000 66.100000  26.540000 ;
        RECT 65.900000  26.770000 66.100000  26.970000 ;
        RECT 65.900000  27.200000 66.100000  27.400000 ;
        RECT 65.900000  27.630000 66.100000  27.830000 ;
        RECT 65.900000  28.060000 66.100000  28.260000 ;
        RECT 65.900000  28.490000 66.100000  28.690000 ;
        RECT 65.900000  28.920000 66.100000  29.120000 ;
        RECT 65.900000  29.350000 66.100000  29.550000 ;
        RECT 65.900000  29.780000 66.100000  29.980000 ;
        RECT 65.900000  30.210000 66.100000  30.410000 ;
        RECT 65.990000 175.995000 66.190000 176.195000 ;
        RECT 65.990000 176.395000 66.190000 176.595000 ;
        RECT 65.990000 176.795000 66.190000 176.995000 ;
        RECT 65.990000 177.195000 66.190000 177.395000 ;
        RECT 65.990000 177.595000 66.190000 177.795000 ;
        RECT 65.990000 177.995000 66.190000 178.195000 ;
        RECT 65.990000 178.395000 66.190000 178.595000 ;
        RECT 65.990000 178.795000 66.190000 178.995000 ;
        RECT 65.990000 179.195000 66.190000 179.395000 ;
        RECT 65.990000 179.595000 66.190000 179.795000 ;
        RECT 65.990000 179.995000 66.190000 180.195000 ;
        RECT 65.990000 180.395000 66.190000 180.595000 ;
        RECT 65.990000 180.795000 66.190000 180.995000 ;
        RECT 65.990000 181.195000 66.190000 181.395000 ;
        RECT 65.990000 181.595000 66.190000 181.795000 ;
        RECT 65.990000 181.995000 66.190000 182.195000 ;
        RECT 65.990000 182.395000 66.190000 182.595000 ;
        RECT 65.990000 182.795000 66.190000 182.995000 ;
        RECT 65.990000 183.195000 66.190000 183.395000 ;
        RECT 65.990000 183.595000 66.190000 183.795000 ;
        RECT 65.990000 183.995000 66.190000 184.195000 ;
        RECT 65.990000 184.395000 66.190000 184.595000 ;
        RECT 65.990000 184.795000 66.190000 184.995000 ;
        RECT 65.990000 185.195000 66.190000 185.395000 ;
        RECT 65.990000 185.595000 66.190000 185.795000 ;
        RECT 65.990000 185.995000 66.190000 186.195000 ;
        RECT 65.990000 186.395000 66.190000 186.595000 ;
        RECT 65.990000 186.795000 66.190000 186.995000 ;
        RECT 65.990000 187.195000 66.190000 187.395000 ;
        RECT 65.990000 187.595000 66.190000 187.795000 ;
        RECT 65.990000 187.995000 66.190000 188.195000 ;
        RECT 65.990000 188.395000 66.190000 188.595000 ;
        RECT 65.990000 188.795000 66.190000 188.995000 ;
        RECT 65.990000 189.195000 66.190000 189.395000 ;
        RECT 65.990000 189.595000 66.190000 189.795000 ;
        RECT 65.990000 189.995000 66.190000 190.195000 ;
        RECT 65.990000 190.395000 66.190000 190.595000 ;
        RECT 65.990000 190.795000 66.190000 190.995000 ;
        RECT 65.990000 191.195000 66.190000 191.395000 ;
        RECT 65.990000 191.595000 66.190000 191.795000 ;
        RECT 65.990000 191.995000 66.190000 192.195000 ;
        RECT 65.990000 192.395000 66.190000 192.595000 ;
        RECT 65.990000 192.795000 66.190000 192.995000 ;
        RECT 65.990000 193.195000 66.190000 193.395000 ;
        RECT 65.990000 193.595000 66.190000 193.795000 ;
        RECT 65.990000 193.995000 66.190000 194.195000 ;
        RECT 65.990000 194.395000 66.190000 194.595000 ;
        RECT 65.990000 194.795000 66.190000 194.995000 ;
        RECT 65.990000 195.200000 66.190000 195.400000 ;
        RECT 65.990000 195.605000 66.190000 195.805000 ;
        RECT 65.990000 196.010000 66.190000 196.210000 ;
        RECT 65.990000 196.415000 66.190000 196.615000 ;
        RECT 65.990000 196.820000 66.190000 197.020000 ;
        RECT 65.990000 197.225000 66.190000 197.425000 ;
        RECT 65.990000 197.630000 66.190000 197.830000 ;
        RECT 65.990000 198.035000 66.190000 198.235000 ;
        RECT 65.990000 198.440000 66.190000 198.640000 ;
        RECT 65.990000 198.845000 66.190000 199.045000 ;
        RECT 65.990000 199.250000 66.190000 199.450000 ;
        RECT 65.990000 199.655000 66.190000 199.855000 ;
        RECT 66.305000  25.910000 66.505000  26.110000 ;
        RECT 66.305000  26.340000 66.505000  26.540000 ;
        RECT 66.305000  26.770000 66.505000  26.970000 ;
        RECT 66.305000  27.200000 66.505000  27.400000 ;
        RECT 66.305000  27.630000 66.505000  27.830000 ;
        RECT 66.305000  28.060000 66.505000  28.260000 ;
        RECT 66.305000  28.490000 66.505000  28.690000 ;
        RECT 66.305000  28.920000 66.505000  29.120000 ;
        RECT 66.305000  29.350000 66.505000  29.550000 ;
        RECT 66.305000  29.780000 66.505000  29.980000 ;
        RECT 66.305000  30.210000 66.505000  30.410000 ;
        RECT 66.390000 175.995000 66.590000 176.195000 ;
        RECT 66.390000 176.395000 66.590000 176.595000 ;
        RECT 66.390000 176.795000 66.590000 176.995000 ;
        RECT 66.390000 177.195000 66.590000 177.395000 ;
        RECT 66.390000 177.595000 66.590000 177.795000 ;
        RECT 66.390000 177.995000 66.590000 178.195000 ;
        RECT 66.390000 178.395000 66.590000 178.595000 ;
        RECT 66.390000 178.795000 66.590000 178.995000 ;
        RECT 66.390000 179.195000 66.590000 179.395000 ;
        RECT 66.390000 179.595000 66.590000 179.795000 ;
        RECT 66.390000 179.995000 66.590000 180.195000 ;
        RECT 66.390000 180.395000 66.590000 180.595000 ;
        RECT 66.390000 180.795000 66.590000 180.995000 ;
        RECT 66.390000 181.195000 66.590000 181.395000 ;
        RECT 66.390000 181.595000 66.590000 181.795000 ;
        RECT 66.390000 181.995000 66.590000 182.195000 ;
        RECT 66.390000 182.395000 66.590000 182.595000 ;
        RECT 66.390000 182.795000 66.590000 182.995000 ;
        RECT 66.390000 183.195000 66.590000 183.395000 ;
        RECT 66.390000 183.595000 66.590000 183.795000 ;
        RECT 66.390000 183.995000 66.590000 184.195000 ;
        RECT 66.390000 184.395000 66.590000 184.595000 ;
        RECT 66.390000 184.795000 66.590000 184.995000 ;
        RECT 66.390000 185.195000 66.590000 185.395000 ;
        RECT 66.390000 185.595000 66.590000 185.795000 ;
        RECT 66.390000 185.995000 66.590000 186.195000 ;
        RECT 66.390000 186.395000 66.590000 186.595000 ;
        RECT 66.390000 186.795000 66.590000 186.995000 ;
        RECT 66.390000 187.195000 66.590000 187.395000 ;
        RECT 66.390000 187.595000 66.590000 187.795000 ;
        RECT 66.390000 187.995000 66.590000 188.195000 ;
        RECT 66.390000 188.395000 66.590000 188.595000 ;
        RECT 66.390000 188.795000 66.590000 188.995000 ;
        RECT 66.390000 189.195000 66.590000 189.395000 ;
        RECT 66.390000 189.595000 66.590000 189.795000 ;
        RECT 66.390000 189.995000 66.590000 190.195000 ;
        RECT 66.390000 190.395000 66.590000 190.595000 ;
        RECT 66.390000 190.795000 66.590000 190.995000 ;
        RECT 66.390000 191.195000 66.590000 191.395000 ;
        RECT 66.390000 191.595000 66.590000 191.795000 ;
        RECT 66.390000 191.995000 66.590000 192.195000 ;
        RECT 66.390000 192.395000 66.590000 192.595000 ;
        RECT 66.390000 192.795000 66.590000 192.995000 ;
        RECT 66.390000 193.195000 66.590000 193.395000 ;
        RECT 66.390000 193.595000 66.590000 193.795000 ;
        RECT 66.390000 193.995000 66.590000 194.195000 ;
        RECT 66.390000 194.395000 66.590000 194.595000 ;
        RECT 66.390000 194.795000 66.590000 194.995000 ;
        RECT 66.390000 195.200000 66.590000 195.400000 ;
        RECT 66.390000 195.605000 66.590000 195.805000 ;
        RECT 66.390000 196.010000 66.590000 196.210000 ;
        RECT 66.390000 196.415000 66.590000 196.615000 ;
        RECT 66.390000 196.820000 66.590000 197.020000 ;
        RECT 66.390000 197.225000 66.590000 197.425000 ;
        RECT 66.390000 197.630000 66.590000 197.830000 ;
        RECT 66.390000 198.035000 66.590000 198.235000 ;
        RECT 66.390000 198.440000 66.590000 198.640000 ;
        RECT 66.390000 198.845000 66.590000 199.045000 ;
        RECT 66.390000 199.250000 66.590000 199.450000 ;
        RECT 66.390000 199.655000 66.590000 199.855000 ;
        RECT 66.710000  25.910000 66.910000  26.110000 ;
        RECT 66.710000  26.340000 66.910000  26.540000 ;
        RECT 66.710000  26.770000 66.910000  26.970000 ;
        RECT 66.710000  27.200000 66.910000  27.400000 ;
        RECT 66.710000  27.630000 66.910000  27.830000 ;
        RECT 66.710000  28.060000 66.910000  28.260000 ;
        RECT 66.710000  28.490000 66.910000  28.690000 ;
        RECT 66.710000  28.920000 66.910000  29.120000 ;
        RECT 66.710000  29.350000 66.910000  29.550000 ;
        RECT 66.710000  29.780000 66.910000  29.980000 ;
        RECT 66.710000  30.210000 66.910000  30.410000 ;
        RECT 66.790000 175.995000 66.990000 176.195000 ;
        RECT 66.790000 176.395000 66.990000 176.595000 ;
        RECT 66.790000 176.795000 66.990000 176.995000 ;
        RECT 66.790000 177.195000 66.990000 177.395000 ;
        RECT 66.790000 177.595000 66.990000 177.795000 ;
        RECT 66.790000 177.995000 66.990000 178.195000 ;
        RECT 66.790000 178.395000 66.990000 178.595000 ;
        RECT 66.790000 178.795000 66.990000 178.995000 ;
        RECT 66.790000 179.195000 66.990000 179.395000 ;
        RECT 66.790000 179.595000 66.990000 179.795000 ;
        RECT 66.790000 179.995000 66.990000 180.195000 ;
        RECT 66.790000 180.395000 66.990000 180.595000 ;
        RECT 66.790000 180.795000 66.990000 180.995000 ;
        RECT 66.790000 181.195000 66.990000 181.395000 ;
        RECT 66.790000 181.595000 66.990000 181.795000 ;
        RECT 66.790000 181.995000 66.990000 182.195000 ;
        RECT 66.790000 182.395000 66.990000 182.595000 ;
        RECT 66.790000 182.795000 66.990000 182.995000 ;
        RECT 66.790000 183.195000 66.990000 183.395000 ;
        RECT 66.790000 183.595000 66.990000 183.795000 ;
        RECT 66.790000 183.995000 66.990000 184.195000 ;
        RECT 66.790000 184.395000 66.990000 184.595000 ;
        RECT 66.790000 184.795000 66.990000 184.995000 ;
        RECT 66.790000 185.195000 66.990000 185.395000 ;
        RECT 66.790000 185.595000 66.990000 185.795000 ;
        RECT 66.790000 185.995000 66.990000 186.195000 ;
        RECT 66.790000 186.395000 66.990000 186.595000 ;
        RECT 66.790000 186.795000 66.990000 186.995000 ;
        RECT 66.790000 187.195000 66.990000 187.395000 ;
        RECT 66.790000 187.595000 66.990000 187.795000 ;
        RECT 66.790000 187.995000 66.990000 188.195000 ;
        RECT 66.790000 188.395000 66.990000 188.595000 ;
        RECT 66.790000 188.795000 66.990000 188.995000 ;
        RECT 66.790000 189.195000 66.990000 189.395000 ;
        RECT 66.790000 189.595000 66.990000 189.795000 ;
        RECT 66.790000 189.995000 66.990000 190.195000 ;
        RECT 66.790000 190.395000 66.990000 190.595000 ;
        RECT 66.790000 190.795000 66.990000 190.995000 ;
        RECT 66.790000 191.195000 66.990000 191.395000 ;
        RECT 66.790000 191.595000 66.990000 191.795000 ;
        RECT 66.790000 191.995000 66.990000 192.195000 ;
        RECT 66.790000 192.395000 66.990000 192.595000 ;
        RECT 66.790000 192.795000 66.990000 192.995000 ;
        RECT 66.790000 193.195000 66.990000 193.395000 ;
        RECT 66.790000 193.595000 66.990000 193.795000 ;
        RECT 66.790000 193.995000 66.990000 194.195000 ;
        RECT 66.790000 194.395000 66.990000 194.595000 ;
        RECT 66.790000 194.795000 66.990000 194.995000 ;
        RECT 66.790000 195.200000 66.990000 195.400000 ;
        RECT 66.790000 195.605000 66.990000 195.805000 ;
        RECT 66.790000 196.010000 66.990000 196.210000 ;
        RECT 66.790000 196.415000 66.990000 196.615000 ;
        RECT 66.790000 196.820000 66.990000 197.020000 ;
        RECT 66.790000 197.225000 66.990000 197.425000 ;
        RECT 66.790000 197.630000 66.990000 197.830000 ;
        RECT 66.790000 198.035000 66.990000 198.235000 ;
        RECT 66.790000 198.440000 66.990000 198.640000 ;
        RECT 66.790000 198.845000 66.990000 199.045000 ;
        RECT 66.790000 199.250000 66.990000 199.450000 ;
        RECT 66.790000 199.655000 66.990000 199.855000 ;
        RECT 67.115000  25.910000 67.315000  26.110000 ;
        RECT 67.115000  26.340000 67.315000  26.540000 ;
        RECT 67.115000  26.770000 67.315000  26.970000 ;
        RECT 67.115000  27.200000 67.315000  27.400000 ;
        RECT 67.115000  27.630000 67.315000  27.830000 ;
        RECT 67.115000  28.060000 67.315000  28.260000 ;
        RECT 67.115000  28.490000 67.315000  28.690000 ;
        RECT 67.115000  28.920000 67.315000  29.120000 ;
        RECT 67.115000  29.350000 67.315000  29.550000 ;
        RECT 67.115000  29.780000 67.315000  29.980000 ;
        RECT 67.115000  30.210000 67.315000  30.410000 ;
        RECT 67.190000 175.995000 67.390000 176.195000 ;
        RECT 67.190000 176.395000 67.390000 176.595000 ;
        RECT 67.190000 176.795000 67.390000 176.995000 ;
        RECT 67.190000 177.195000 67.390000 177.395000 ;
        RECT 67.190000 177.595000 67.390000 177.795000 ;
        RECT 67.190000 177.995000 67.390000 178.195000 ;
        RECT 67.190000 178.395000 67.390000 178.595000 ;
        RECT 67.190000 178.795000 67.390000 178.995000 ;
        RECT 67.190000 179.195000 67.390000 179.395000 ;
        RECT 67.190000 179.595000 67.390000 179.795000 ;
        RECT 67.190000 179.995000 67.390000 180.195000 ;
        RECT 67.190000 180.395000 67.390000 180.595000 ;
        RECT 67.190000 180.795000 67.390000 180.995000 ;
        RECT 67.190000 181.195000 67.390000 181.395000 ;
        RECT 67.190000 181.595000 67.390000 181.795000 ;
        RECT 67.190000 181.995000 67.390000 182.195000 ;
        RECT 67.190000 182.395000 67.390000 182.595000 ;
        RECT 67.190000 182.795000 67.390000 182.995000 ;
        RECT 67.190000 183.195000 67.390000 183.395000 ;
        RECT 67.190000 183.595000 67.390000 183.795000 ;
        RECT 67.190000 183.995000 67.390000 184.195000 ;
        RECT 67.190000 184.395000 67.390000 184.595000 ;
        RECT 67.190000 184.795000 67.390000 184.995000 ;
        RECT 67.190000 185.195000 67.390000 185.395000 ;
        RECT 67.190000 185.595000 67.390000 185.795000 ;
        RECT 67.190000 185.995000 67.390000 186.195000 ;
        RECT 67.190000 186.395000 67.390000 186.595000 ;
        RECT 67.190000 186.795000 67.390000 186.995000 ;
        RECT 67.190000 187.195000 67.390000 187.395000 ;
        RECT 67.190000 187.595000 67.390000 187.795000 ;
        RECT 67.190000 187.995000 67.390000 188.195000 ;
        RECT 67.190000 188.395000 67.390000 188.595000 ;
        RECT 67.190000 188.795000 67.390000 188.995000 ;
        RECT 67.190000 189.195000 67.390000 189.395000 ;
        RECT 67.190000 189.595000 67.390000 189.795000 ;
        RECT 67.190000 189.995000 67.390000 190.195000 ;
        RECT 67.190000 190.395000 67.390000 190.595000 ;
        RECT 67.190000 190.795000 67.390000 190.995000 ;
        RECT 67.190000 191.195000 67.390000 191.395000 ;
        RECT 67.190000 191.595000 67.390000 191.795000 ;
        RECT 67.190000 191.995000 67.390000 192.195000 ;
        RECT 67.190000 192.395000 67.390000 192.595000 ;
        RECT 67.190000 192.795000 67.390000 192.995000 ;
        RECT 67.190000 193.195000 67.390000 193.395000 ;
        RECT 67.190000 193.595000 67.390000 193.795000 ;
        RECT 67.190000 193.995000 67.390000 194.195000 ;
        RECT 67.190000 194.395000 67.390000 194.595000 ;
        RECT 67.190000 194.795000 67.390000 194.995000 ;
        RECT 67.190000 195.200000 67.390000 195.400000 ;
        RECT 67.190000 195.605000 67.390000 195.805000 ;
        RECT 67.190000 196.010000 67.390000 196.210000 ;
        RECT 67.190000 196.415000 67.390000 196.615000 ;
        RECT 67.190000 196.820000 67.390000 197.020000 ;
        RECT 67.190000 197.225000 67.390000 197.425000 ;
        RECT 67.190000 197.630000 67.390000 197.830000 ;
        RECT 67.190000 198.035000 67.390000 198.235000 ;
        RECT 67.190000 198.440000 67.390000 198.640000 ;
        RECT 67.190000 198.845000 67.390000 199.045000 ;
        RECT 67.190000 199.250000 67.390000 199.450000 ;
        RECT 67.190000 199.655000 67.390000 199.855000 ;
        RECT 67.520000  25.910000 67.720000  26.110000 ;
        RECT 67.520000  26.340000 67.720000  26.540000 ;
        RECT 67.520000  26.770000 67.720000  26.970000 ;
        RECT 67.520000  27.200000 67.720000  27.400000 ;
        RECT 67.520000  27.630000 67.720000  27.830000 ;
        RECT 67.520000  28.060000 67.720000  28.260000 ;
        RECT 67.520000  28.490000 67.720000  28.690000 ;
        RECT 67.520000  28.920000 67.720000  29.120000 ;
        RECT 67.520000  29.350000 67.720000  29.550000 ;
        RECT 67.520000  29.780000 67.720000  29.980000 ;
        RECT 67.520000  30.210000 67.720000  30.410000 ;
        RECT 67.590000 175.995000 67.790000 176.195000 ;
        RECT 67.590000 176.395000 67.790000 176.595000 ;
        RECT 67.590000 176.795000 67.790000 176.995000 ;
        RECT 67.590000 177.195000 67.790000 177.395000 ;
        RECT 67.590000 177.595000 67.790000 177.795000 ;
        RECT 67.590000 177.995000 67.790000 178.195000 ;
        RECT 67.590000 178.395000 67.790000 178.595000 ;
        RECT 67.590000 178.795000 67.790000 178.995000 ;
        RECT 67.590000 179.195000 67.790000 179.395000 ;
        RECT 67.590000 179.595000 67.790000 179.795000 ;
        RECT 67.590000 179.995000 67.790000 180.195000 ;
        RECT 67.590000 180.395000 67.790000 180.595000 ;
        RECT 67.590000 180.795000 67.790000 180.995000 ;
        RECT 67.590000 181.195000 67.790000 181.395000 ;
        RECT 67.590000 181.595000 67.790000 181.795000 ;
        RECT 67.590000 181.995000 67.790000 182.195000 ;
        RECT 67.590000 182.395000 67.790000 182.595000 ;
        RECT 67.590000 182.795000 67.790000 182.995000 ;
        RECT 67.590000 183.195000 67.790000 183.395000 ;
        RECT 67.590000 183.595000 67.790000 183.795000 ;
        RECT 67.590000 183.995000 67.790000 184.195000 ;
        RECT 67.590000 184.395000 67.790000 184.595000 ;
        RECT 67.590000 184.795000 67.790000 184.995000 ;
        RECT 67.590000 185.195000 67.790000 185.395000 ;
        RECT 67.590000 185.595000 67.790000 185.795000 ;
        RECT 67.590000 185.995000 67.790000 186.195000 ;
        RECT 67.590000 186.395000 67.790000 186.595000 ;
        RECT 67.590000 186.795000 67.790000 186.995000 ;
        RECT 67.590000 187.195000 67.790000 187.395000 ;
        RECT 67.590000 187.595000 67.790000 187.795000 ;
        RECT 67.590000 187.995000 67.790000 188.195000 ;
        RECT 67.590000 188.395000 67.790000 188.595000 ;
        RECT 67.590000 188.795000 67.790000 188.995000 ;
        RECT 67.590000 189.195000 67.790000 189.395000 ;
        RECT 67.590000 189.595000 67.790000 189.795000 ;
        RECT 67.590000 189.995000 67.790000 190.195000 ;
        RECT 67.590000 190.395000 67.790000 190.595000 ;
        RECT 67.590000 190.795000 67.790000 190.995000 ;
        RECT 67.590000 191.195000 67.790000 191.395000 ;
        RECT 67.590000 191.595000 67.790000 191.795000 ;
        RECT 67.590000 191.995000 67.790000 192.195000 ;
        RECT 67.590000 192.395000 67.790000 192.595000 ;
        RECT 67.590000 192.795000 67.790000 192.995000 ;
        RECT 67.590000 193.195000 67.790000 193.395000 ;
        RECT 67.590000 193.595000 67.790000 193.795000 ;
        RECT 67.590000 193.995000 67.790000 194.195000 ;
        RECT 67.590000 194.395000 67.790000 194.595000 ;
        RECT 67.590000 194.795000 67.790000 194.995000 ;
        RECT 67.590000 195.200000 67.790000 195.400000 ;
        RECT 67.590000 195.605000 67.790000 195.805000 ;
        RECT 67.590000 196.010000 67.790000 196.210000 ;
        RECT 67.590000 196.415000 67.790000 196.615000 ;
        RECT 67.590000 196.820000 67.790000 197.020000 ;
        RECT 67.590000 197.225000 67.790000 197.425000 ;
        RECT 67.590000 197.630000 67.790000 197.830000 ;
        RECT 67.590000 198.035000 67.790000 198.235000 ;
        RECT 67.590000 198.440000 67.790000 198.640000 ;
        RECT 67.590000 198.845000 67.790000 199.045000 ;
        RECT 67.590000 199.250000 67.790000 199.450000 ;
        RECT 67.590000 199.655000 67.790000 199.855000 ;
        RECT 67.925000  25.910000 68.125000  26.110000 ;
        RECT 67.925000  26.340000 68.125000  26.540000 ;
        RECT 67.925000  26.770000 68.125000  26.970000 ;
        RECT 67.925000  27.200000 68.125000  27.400000 ;
        RECT 67.925000  27.630000 68.125000  27.830000 ;
        RECT 67.925000  28.060000 68.125000  28.260000 ;
        RECT 67.925000  28.490000 68.125000  28.690000 ;
        RECT 67.925000  28.920000 68.125000  29.120000 ;
        RECT 67.925000  29.350000 68.125000  29.550000 ;
        RECT 67.925000  29.780000 68.125000  29.980000 ;
        RECT 67.925000  30.210000 68.125000  30.410000 ;
        RECT 67.990000 175.995000 68.190000 176.195000 ;
        RECT 67.990000 176.395000 68.190000 176.595000 ;
        RECT 67.990000 176.795000 68.190000 176.995000 ;
        RECT 67.990000 177.195000 68.190000 177.395000 ;
        RECT 67.990000 177.595000 68.190000 177.795000 ;
        RECT 67.990000 177.995000 68.190000 178.195000 ;
        RECT 67.990000 178.395000 68.190000 178.595000 ;
        RECT 67.990000 178.795000 68.190000 178.995000 ;
        RECT 67.990000 179.195000 68.190000 179.395000 ;
        RECT 67.990000 179.595000 68.190000 179.795000 ;
        RECT 67.990000 179.995000 68.190000 180.195000 ;
        RECT 67.990000 180.395000 68.190000 180.595000 ;
        RECT 67.990000 180.795000 68.190000 180.995000 ;
        RECT 67.990000 181.195000 68.190000 181.395000 ;
        RECT 67.990000 181.595000 68.190000 181.795000 ;
        RECT 67.990000 181.995000 68.190000 182.195000 ;
        RECT 67.990000 182.395000 68.190000 182.595000 ;
        RECT 67.990000 182.795000 68.190000 182.995000 ;
        RECT 67.990000 183.195000 68.190000 183.395000 ;
        RECT 67.990000 183.595000 68.190000 183.795000 ;
        RECT 67.990000 183.995000 68.190000 184.195000 ;
        RECT 67.990000 184.395000 68.190000 184.595000 ;
        RECT 67.990000 184.795000 68.190000 184.995000 ;
        RECT 67.990000 185.195000 68.190000 185.395000 ;
        RECT 67.990000 185.595000 68.190000 185.795000 ;
        RECT 67.990000 185.995000 68.190000 186.195000 ;
        RECT 67.990000 186.395000 68.190000 186.595000 ;
        RECT 67.990000 186.795000 68.190000 186.995000 ;
        RECT 67.990000 187.195000 68.190000 187.395000 ;
        RECT 67.990000 187.595000 68.190000 187.795000 ;
        RECT 67.990000 187.995000 68.190000 188.195000 ;
        RECT 67.990000 188.395000 68.190000 188.595000 ;
        RECT 67.990000 188.795000 68.190000 188.995000 ;
        RECT 67.990000 189.195000 68.190000 189.395000 ;
        RECT 67.990000 189.595000 68.190000 189.795000 ;
        RECT 67.990000 189.995000 68.190000 190.195000 ;
        RECT 67.990000 190.395000 68.190000 190.595000 ;
        RECT 67.990000 190.795000 68.190000 190.995000 ;
        RECT 67.990000 191.195000 68.190000 191.395000 ;
        RECT 67.990000 191.595000 68.190000 191.795000 ;
        RECT 67.990000 191.995000 68.190000 192.195000 ;
        RECT 67.990000 192.395000 68.190000 192.595000 ;
        RECT 67.990000 192.795000 68.190000 192.995000 ;
        RECT 67.990000 193.195000 68.190000 193.395000 ;
        RECT 67.990000 193.595000 68.190000 193.795000 ;
        RECT 67.990000 193.995000 68.190000 194.195000 ;
        RECT 67.990000 194.395000 68.190000 194.595000 ;
        RECT 67.990000 194.795000 68.190000 194.995000 ;
        RECT 67.990000 195.200000 68.190000 195.400000 ;
        RECT 67.990000 195.605000 68.190000 195.805000 ;
        RECT 67.990000 196.010000 68.190000 196.210000 ;
        RECT 67.990000 196.415000 68.190000 196.615000 ;
        RECT 67.990000 196.820000 68.190000 197.020000 ;
        RECT 67.990000 197.225000 68.190000 197.425000 ;
        RECT 67.990000 197.630000 68.190000 197.830000 ;
        RECT 67.990000 198.035000 68.190000 198.235000 ;
        RECT 67.990000 198.440000 68.190000 198.640000 ;
        RECT 67.990000 198.845000 68.190000 199.045000 ;
        RECT 67.990000 199.250000 68.190000 199.450000 ;
        RECT 67.990000 199.655000 68.190000 199.855000 ;
        RECT 68.330000  25.910000 68.530000  26.110000 ;
        RECT 68.330000  26.340000 68.530000  26.540000 ;
        RECT 68.330000  26.770000 68.530000  26.970000 ;
        RECT 68.330000  27.200000 68.530000  27.400000 ;
        RECT 68.330000  27.630000 68.530000  27.830000 ;
        RECT 68.330000  28.060000 68.530000  28.260000 ;
        RECT 68.330000  28.490000 68.530000  28.690000 ;
        RECT 68.330000  28.920000 68.530000  29.120000 ;
        RECT 68.330000  29.350000 68.530000  29.550000 ;
        RECT 68.330000  29.780000 68.530000  29.980000 ;
        RECT 68.330000  30.210000 68.530000  30.410000 ;
        RECT 68.390000 175.995000 68.590000 176.195000 ;
        RECT 68.390000 176.395000 68.590000 176.595000 ;
        RECT 68.390000 176.795000 68.590000 176.995000 ;
        RECT 68.390000 177.195000 68.590000 177.395000 ;
        RECT 68.390000 177.595000 68.590000 177.795000 ;
        RECT 68.390000 177.995000 68.590000 178.195000 ;
        RECT 68.390000 178.395000 68.590000 178.595000 ;
        RECT 68.390000 178.795000 68.590000 178.995000 ;
        RECT 68.390000 179.195000 68.590000 179.395000 ;
        RECT 68.390000 179.595000 68.590000 179.795000 ;
        RECT 68.390000 179.995000 68.590000 180.195000 ;
        RECT 68.390000 180.395000 68.590000 180.595000 ;
        RECT 68.390000 180.795000 68.590000 180.995000 ;
        RECT 68.390000 181.195000 68.590000 181.395000 ;
        RECT 68.390000 181.595000 68.590000 181.795000 ;
        RECT 68.390000 181.995000 68.590000 182.195000 ;
        RECT 68.390000 182.395000 68.590000 182.595000 ;
        RECT 68.390000 182.795000 68.590000 182.995000 ;
        RECT 68.390000 183.195000 68.590000 183.395000 ;
        RECT 68.390000 183.595000 68.590000 183.795000 ;
        RECT 68.390000 183.995000 68.590000 184.195000 ;
        RECT 68.390000 184.395000 68.590000 184.595000 ;
        RECT 68.390000 184.795000 68.590000 184.995000 ;
        RECT 68.390000 185.195000 68.590000 185.395000 ;
        RECT 68.390000 185.595000 68.590000 185.795000 ;
        RECT 68.390000 185.995000 68.590000 186.195000 ;
        RECT 68.390000 186.395000 68.590000 186.595000 ;
        RECT 68.390000 186.795000 68.590000 186.995000 ;
        RECT 68.390000 187.195000 68.590000 187.395000 ;
        RECT 68.390000 187.595000 68.590000 187.795000 ;
        RECT 68.390000 187.995000 68.590000 188.195000 ;
        RECT 68.390000 188.395000 68.590000 188.595000 ;
        RECT 68.390000 188.795000 68.590000 188.995000 ;
        RECT 68.390000 189.195000 68.590000 189.395000 ;
        RECT 68.390000 189.595000 68.590000 189.795000 ;
        RECT 68.390000 189.995000 68.590000 190.195000 ;
        RECT 68.390000 190.395000 68.590000 190.595000 ;
        RECT 68.390000 190.795000 68.590000 190.995000 ;
        RECT 68.390000 191.195000 68.590000 191.395000 ;
        RECT 68.390000 191.595000 68.590000 191.795000 ;
        RECT 68.390000 191.995000 68.590000 192.195000 ;
        RECT 68.390000 192.395000 68.590000 192.595000 ;
        RECT 68.390000 192.795000 68.590000 192.995000 ;
        RECT 68.390000 193.195000 68.590000 193.395000 ;
        RECT 68.390000 193.595000 68.590000 193.795000 ;
        RECT 68.390000 193.995000 68.590000 194.195000 ;
        RECT 68.390000 194.395000 68.590000 194.595000 ;
        RECT 68.390000 194.795000 68.590000 194.995000 ;
        RECT 68.390000 195.200000 68.590000 195.400000 ;
        RECT 68.390000 195.605000 68.590000 195.805000 ;
        RECT 68.390000 196.010000 68.590000 196.210000 ;
        RECT 68.390000 196.415000 68.590000 196.615000 ;
        RECT 68.390000 196.820000 68.590000 197.020000 ;
        RECT 68.390000 197.225000 68.590000 197.425000 ;
        RECT 68.390000 197.630000 68.590000 197.830000 ;
        RECT 68.390000 198.035000 68.590000 198.235000 ;
        RECT 68.390000 198.440000 68.590000 198.640000 ;
        RECT 68.390000 198.845000 68.590000 199.045000 ;
        RECT 68.390000 199.250000 68.590000 199.450000 ;
        RECT 68.390000 199.655000 68.590000 199.855000 ;
        RECT 68.735000  25.910000 68.935000  26.110000 ;
        RECT 68.735000  26.340000 68.935000  26.540000 ;
        RECT 68.735000  26.770000 68.935000  26.970000 ;
        RECT 68.735000  27.200000 68.935000  27.400000 ;
        RECT 68.735000  27.630000 68.935000  27.830000 ;
        RECT 68.735000  28.060000 68.935000  28.260000 ;
        RECT 68.735000  28.490000 68.935000  28.690000 ;
        RECT 68.735000  28.920000 68.935000  29.120000 ;
        RECT 68.735000  29.350000 68.935000  29.550000 ;
        RECT 68.735000  29.780000 68.935000  29.980000 ;
        RECT 68.735000  30.210000 68.935000  30.410000 ;
        RECT 68.790000 175.995000 68.990000 176.195000 ;
        RECT 68.790000 176.395000 68.990000 176.595000 ;
        RECT 68.790000 176.795000 68.990000 176.995000 ;
        RECT 68.790000 177.195000 68.990000 177.395000 ;
        RECT 68.790000 177.595000 68.990000 177.795000 ;
        RECT 68.790000 177.995000 68.990000 178.195000 ;
        RECT 68.790000 178.395000 68.990000 178.595000 ;
        RECT 68.790000 178.795000 68.990000 178.995000 ;
        RECT 68.790000 179.195000 68.990000 179.395000 ;
        RECT 68.790000 179.595000 68.990000 179.795000 ;
        RECT 68.790000 179.995000 68.990000 180.195000 ;
        RECT 68.790000 180.395000 68.990000 180.595000 ;
        RECT 68.790000 180.795000 68.990000 180.995000 ;
        RECT 68.790000 181.195000 68.990000 181.395000 ;
        RECT 68.790000 181.595000 68.990000 181.795000 ;
        RECT 68.790000 181.995000 68.990000 182.195000 ;
        RECT 68.790000 182.395000 68.990000 182.595000 ;
        RECT 68.790000 182.795000 68.990000 182.995000 ;
        RECT 68.790000 183.195000 68.990000 183.395000 ;
        RECT 68.790000 183.595000 68.990000 183.795000 ;
        RECT 68.790000 183.995000 68.990000 184.195000 ;
        RECT 68.790000 184.395000 68.990000 184.595000 ;
        RECT 68.790000 184.795000 68.990000 184.995000 ;
        RECT 68.790000 185.195000 68.990000 185.395000 ;
        RECT 68.790000 185.595000 68.990000 185.795000 ;
        RECT 68.790000 185.995000 68.990000 186.195000 ;
        RECT 68.790000 186.395000 68.990000 186.595000 ;
        RECT 68.790000 186.795000 68.990000 186.995000 ;
        RECT 68.790000 187.195000 68.990000 187.395000 ;
        RECT 68.790000 187.595000 68.990000 187.795000 ;
        RECT 68.790000 187.995000 68.990000 188.195000 ;
        RECT 68.790000 188.395000 68.990000 188.595000 ;
        RECT 68.790000 188.795000 68.990000 188.995000 ;
        RECT 68.790000 189.195000 68.990000 189.395000 ;
        RECT 68.790000 189.595000 68.990000 189.795000 ;
        RECT 68.790000 189.995000 68.990000 190.195000 ;
        RECT 68.790000 190.395000 68.990000 190.595000 ;
        RECT 68.790000 190.795000 68.990000 190.995000 ;
        RECT 68.790000 191.195000 68.990000 191.395000 ;
        RECT 68.790000 191.595000 68.990000 191.795000 ;
        RECT 68.790000 191.995000 68.990000 192.195000 ;
        RECT 68.790000 192.395000 68.990000 192.595000 ;
        RECT 68.790000 192.795000 68.990000 192.995000 ;
        RECT 68.790000 193.195000 68.990000 193.395000 ;
        RECT 68.790000 193.595000 68.990000 193.795000 ;
        RECT 68.790000 193.995000 68.990000 194.195000 ;
        RECT 68.790000 194.395000 68.990000 194.595000 ;
        RECT 68.790000 194.795000 68.990000 194.995000 ;
        RECT 68.790000 195.200000 68.990000 195.400000 ;
        RECT 68.790000 195.605000 68.990000 195.805000 ;
        RECT 68.790000 196.010000 68.990000 196.210000 ;
        RECT 68.790000 196.415000 68.990000 196.615000 ;
        RECT 68.790000 196.820000 68.990000 197.020000 ;
        RECT 68.790000 197.225000 68.990000 197.425000 ;
        RECT 68.790000 197.630000 68.990000 197.830000 ;
        RECT 68.790000 198.035000 68.990000 198.235000 ;
        RECT 68.790000 198.440000 68.990000 198.640000 ;
        RECT 68.790000 198.845000 68.990000 199.045000 ;
        RECT 68.790000 199.250000 68.990000 199.450000 ;
        RECT 68.790000 199.655000 68.990000 199.855000 ;
        RECT 69.140000  25.910000 69.340000  26.110000 ;
        RECT 69.140000  26.340000 69.340000  26.540000 ;
        RECT 69.140000  26.770000 69.340000  26.970000 ;
        RECT 69.140000  27.200000 69.340000  27.400000 ;
        RECT 69.140000  27.630000 69.340000  27.830000 ;
        RECT 69.140000  28.060000 69.340000  28.260000 ;
        RECT 69.140000  28.490000 69.340000  28.690000 ;
        RECT 69.140000  28.920000 69.340000  29.120000 ;
        RECT 69.140000  29.350000 69.340000  29.550000 ;
        RECT 69.140000  29.780000 69.340000  29.980000 ;
        RECT 69.140000  30.210000 69.340000  30.410000 ;
        RECT 69.190000 175.995000 69.390000 176.195000 ;
        RECT 69.190000 176.395000 69.390000 176.595000 ;
        RECT 69.190000 176.795000 69.390000 176.995000 ;
        RECT 69.190000 177.195000 69.390000 177.395000 ;
        RECT 69.190000 177.595000 69.390000 177.795000 ;
        RECT 69.190000 177.995000 69.390000 178.195000 ;
        RECT 69.190000 178.395000 69.390000 178.595000 ;
        RECT 69.190000 178.795000 69.390000 178.995000 ;
        RECT 69.190000 179.195000 69.390000 179.395000 ;
        RECT 69.190000 179.595000 69.390000 179.795000 ;
        RECT 69.190000 179.995000 69.390000 180.195000 ;
        RECT 69.190000 180.395000 69.390000 180.595000 ;
        RECT 69.190000 180.795000 69.390000 180.995000 ;
        RECT 69.190000 181.195000 69.390000 181.395000 ;
        RECT 69.190000 181.595000 69.390000 181.795000 ;
        RECT 69.190000 181.995000 69.390000 182.195000 ;
        RECT 69.190000 182.395000 69.390000 182.595000 ;
        RECT 69.190000 182.795000 69.390000 182.995000 ;
        RECT 69.190000 183.195000 69.390000 183.395000 ;
        RECT 69.190000 183.595000 69.390000 183.795000 ;
        RECT 69.190000 183.995000 69.390000 184.195000 ;
        RECT 69.190000 184.395000 69.390000 184.595000 ;
        RECT 69.190000 184.795000 69.390000 184.995000 ;
        RECT 69.190000 185.195000 69.390000 185.395000 ;
        RECT 69.190000 185.595000 69.390000 185.795000 ;
        RECT 69.190000 185.995000 69.390000 186.195000 ;
        RECT 69.190000 186.395000 69.390000 186.595000 ;
        RECT 69.190000 186.795000 69.390000 186.995000 ;
        RECT 69.190000 187.195000 69.390000 187.395000 ;
        RECT 69.190000 187.595000 69.390000 187.795000 ;
        RECT 69.190000 187.995000 69.390000 188.195000 ;
        RECT 69.190000 188.395000 69.390000 188.595000 ;
        RECT 69.190000 188.795000 69.390000 188.995000 ;
        RECT 69.190000 189.195000 69.390000 189.395000 ;
        RECT 69.190000 189.595000 69.390000 189.795000 ;
        RECT 69.190000 189.995000 69.390000 190.195000 ;
        RECT 69.190000 190.395000 69.390000 190.595000 ;
        RECT 69.190000 190.795000 69.390000 190.995000 ;
        RECT 69.190000 191.195000 69.390000 191.395000 ;
        RECT 69.190000 191.595000 69.390000 191.795000 ;
        RECT 69.190000 191.995000 69.390000 192.195000 ;
        RECT 69.190000 192.395000 69.390000 192.595000 ;
        RECT 69.190000 192.795000 69.390000 192.995000 ;
        RECT 69.190000 193.195000 69.390000 193.395000 ;
        RECT 69.190000 193.595000 69.390000 193.795000 ;
        RECT 69.190000 193.995000 69.390000 194.195000 ;
        RECT 69.190000 194.395000 69.390000 194.595000 ;
        RECT 69.190000 194.795000 69.390000 194.995000 ;
        RECT 69.190000 195.200000 69.390000 195.400000 ;
        RECT 69.190000 195.605000 69.390000 195.805000 ;
        RECT 69.190000 196.010000 69.390000 196.210000 ;
        RECT 69.190000 196.415000 69.390000 196.615000 ;
        RECT 69.190000 196.820000 69.390000 197.020000 ;
        RECT 69.190000 197.225000 69.390000 197.425000 ;
        RECT 69.190000 197.630000 69.390000 197.830000 ;
        RECT 69.190000 198.035000 69.390000 198.235000 ;
        RECT 69.190000 198.440000 69.390000 198.640000 ;
        RECT 69.190000 198.845000 69.390000 199.045000 ;
        RECT 69.190000 199.250000 69.390000 199.450000 ;
        RECT 69.190000 199.655000 69.390000 199.855000 ;
        RECT 69.545000  25.910000 69.745000  26.110000 ;
        RECT 69.545000  26.340000 69.745000  26.540000 ;
        RECT 69.545000  26.770000 69.745000  26.970000 ;
        RECT 69.545000  27.200000 69.745000  27.400000 ;
        RECT 69.545000  27.630000 69.745000  27.830000 ;
        RECT 69.545000  28.060000 69.745000  28.260000 ;
        RECT 69.545000  28.490000 69.745000  28.690000 ;
        RECT 69.545000  28.920000 69.745000  29.120000 ;
        RECT 69.545000  29.350000 69.745000  29.550000 ;
        RECT 69.545000  29.780000 69.745000  29.980000 ;
        RECT 69.545000  30.210000 69.745000  30.410000 ;
        RECT 69.590000 175.995000 69.790000 176.195000 ;
        RECT 69.590000 176.395000 69.790000 176.595000 ;
        RECT 69.590000 176.795000 69.790000 176.995000 ;
        RECT 69.590000 177.195000 69.790000 177.395000 ;
        RECT 69.590000 177.595000 69.790000 177.795000 ;
        RECT 69.590000 177.995000 69.790000 178.195000 ;
        RECT 69.590000 178.395000 69.790000 178.595000 ;
        RECT 69.590000 178.795000 69.790000 178.995000 ;
        RECT 69.590000 179.195000 69.790000 179.395000 ;
        RECT 69.590000 179.595000 69.790000 179.795000 ;
        RECT 69.590000 179.995000 69.790000 180.195000 ;
        RECT 69.590000 180.395000 69.790000 180.595000 ;
        RECT 69.590000 180.795000 69.790000 180.995000 ;
        RECT 69.590000 181.195000 69.790000 181.395000 ;
        RECT 69.590000 181.595000 69.790000 181.795000 ;
        RECT 69.590000 181.995000 69.790000 182.195000 ;
        RECT 69.590000 182.395000 69.790000 182.595000 ;
        RECT 69.590000 182.795000 69.790000 182.995000 ;
        RECT 69.590000 183.195000 69.790000 183.395000 ;
        RECT 69.590000 183.595000 69.790000 183.795000 ;
        RECT 69.590000 183.995000 69.790000 184.195000 ;
        RECT 69.590000 184.395000 69.790000 184.595000 ;
        RECT 69.590000 184.795000 69.790000 184.995000 ;
        RECT 69.590000 185.195000 69.790000 185.395000 ;
        RECT 69.590000 185.595000 69.790000 185.795000 ;
        RECT 69.590000 185.995000 69.790000 186.195000 ;
        RECT 69.590000 186.395000 69.790000 186.595000 ;
        RECT 69.590000 186.795000 69.790000 186.995000 ;
        RECT 69.590000 187.195000 69.790000 187.395000 ;
        RECT 69.590000 187.595000 69.790000 187.795000 ;
        RECT 69.590000 187.995000 69.790000 188.195000 ;
        RECT 69.590000 188.395000 69.790000 188.595000 ;
        RECT 69.590000 188.795000 69.790000 188.995000 ;
        RECT 69.590000 189.195000 69.790000 189.395000 ;
        RECT 69.590000 189.595000 69.790000 189.795000 ;
        RECT 69.590000 189.995000 69.790000 190.195000 ;
        RECT 69.590000 190.395000 69.790000 190.595000 ;
        RECT 69.590000 190.795000 69.790000 190.995000 ;
        RECT 69.590000 191.195000 69.790000 191.395000 ;
        RECT 69.590000 191.595000 69.790000 191.795000 ;
        RECT 69.590000 191.995000 69.790000 192.195000 ;
        RECT 69.590000 192.395000 69.790000 192.595000 ;
        RECT 69.590000 192.795000 69.790000 192.995000 ;
        RECT 69.590000 193.195000 69.790000 193.395000 ;
        RECT 69.590000 193.595000 69.790000 193.795000 ;
        RECT 69.590000 193.995000 69.790000 194.195000 ;
        RECT 69.590000 194.395000 69.790000 194.595000 ;
        RECT 69.590000 194.795000 69.790000 194.995000 ;
        RECT 69.590000 195.200000 69.790000 195.400000 ;
        RECT 69.590000 195.605000 69.790000 195.805000 ;
        RECT 69.590000 196.010000 69.790000 196.210000 ;
        RECT 69.590000 196.415000 69.790000 196.615000 ;
        RECT 69.590000 196.820000 69.790000 197.020000 ;
        RECT 69.590000 197.225000 69.790000 197.425000 ;
        RECT 69.590000 197.630000 69.790000 197.830000 ;
        RECT 69.590000 198.035000 69.790000 198.235000 ;
        RECT 69.590000 198.440000 69.790000 198.640000 ;
        RECT 69.590000 198.845000 69.790000 199.045000 ;
        RECT 69.590000 199.250000 69.790000 199.450000 ;
        RECT 69.590000 199.655000 69.790000 199.855000 ;
        RECT 69.950000  25.910000 70.150000  26.110000 ;
        RECT 69.950000  26.340000 70.150000  26.540000 ;
        RECT 69.950000  26.770000 70.150000  26.970000 ;
        RECT 69.950000  27.200000 70.150000  27.400000 ;
        RECT 69.950000  27.630000 70.150000  27.830000 ;
        RECT 69.950000  28.060000 70.150000  28.260000 ;
        RECT 69.950000  28.490000 70.150000  28.690000 ;
        RECT 69.950000  28.920000 70.150000  29.120000 ;
        RECT 69.950000  29.350000 70.150000  29.550000 ;
        RECT 69.950000  29.780000 70.150000  29.980000 ;
        RECT 69.950000  30.210000 70.150000  30.410000 ;
        RECT 69.990000 175.995000 70.190000 176.195000 ;
        RECT 69.990000 176.395000 70.190000 176.595000 ;
        RECT 69.990000 176.795000 70.190000 176.995000 ;
        RECT 69.990000 177.195000 70.190000 177.395000 ;
        RECT 69.990000 177.595000 70.190000 177.795000 ;
        RECT 69.990000 177.995000 70.190000 178.195000 ;
        RECT 69.990000 178.395000 70.190000 178.595000 ;
        RECT 69.990000 178.795000 70.190000 178.995000 ;
        RECT 69.990000 179.195000 70.190000 179.395000 ;
        RECT 69.990000 179.595000 70.190000 179.795000 ;
        RECT 69.990000 179.995000 70.190000 180.195000 ;
        RECT 69.990000 180.395000 70.190000 180.595000 ;
        RECT 69.990000 180.795000 70.190000 180.995000 ;
        RECT 69.990000 181.195000 70.190000 181.395000 ;
        RECT 69.990000 181.595000 70.190000 181.795000 ;
        RECT 69.990000 181.995000 70.190000 182.195000 ;
        RECT 69.990000 182.395000 70.190000 182.595000 ;
        RECT 69.990000 182.795000 70.190000 182.995000 ;
        RECT 69.990000 183.195000 70.190000 183.395000 ;
        RECT 69.990000 183.595000 70.190000 183.795000 ;
        RECT 69.990000 183.995000 70.190000 184.195000 ;
        RECT 69.990000 184.395000 70.190000 184.595000 ;
        RECT 69.990000 184.795000 70.190000 184.995000 ;
        RECT 69.990000 185.195000 70.190000 185.395000 ;
        RECT 69.990000 185.595000 70.190000 185.795000 ;
        RECT 69.990000 185.995000 70.190000 186.195000 ;
        RECT 69.990000 186.395000 70.190000 186.595000 ;
        RECT 69.990000 186.795000 70.190000 186.995000 ;
        RECT 69.990000 187.195000 70.190000 187.395000 ;
        RECT 69.990000 187.595000 70.190000 187.795000 ;
        RECT 69.990000 187.995000 70.190000 188.195000 ;
        RECT 69.990000 188.395000 70.190000 188.595000 ;
        RECT 69.990000 188.795000 70.190000 188.995000 ;
        RECT 69.990000 189.195000 70.190000 189.395000 ;
        RECT 69.990000 189.595000 70.190000 189.795000 ;
        RECT 69.990000 189.995000 70.190000 190.195000 ;
        RECT 69.990000 190.395000 70.190000 190.595000 ;
        RECT 69.990000 190.795000 70.190000 190.995000 ;
        RECT 69.990000 191.195000 70.190000 191.395000 ;
        RECT 69.990000 191.595000 70.190000 191.795000 ;
        RECT 69.990000 191.995000 70.190000 192.195000 ;
        RECT 69.990000 192.395000 70.190000 192.595000 ;
        RECT 69.990000 192.795000 70.190000 192.995000 ;
        RECT 69.990000 193.195000 70.190000 193.395000 ;
        RECT 69.990000 193.595000 70.190000 193.795000 ;
        RECT 69.990000 193.995000 70.190000 194.195000 ;
        RECT 69.990000 194.395000 70.190000 194.595000 ;
        RECT 69.990000 194.795000 70.190000 194.995000 ;
        RECT 69.990000 195.200000 70.190000 195.400000 ;
        RECT 69.990000 195.605000 70.190000 195.805000 ;
        RECT 69.990000 196.010000 70.190000 196.210000 ;
        RECT 69.990000 196.415000 70.190000 196.615000 ;
        RECT 69.990000 196.820000 70.190000 197.020000 ;
        RECT 69.990000 197.225000 70.190000 197.425000 ;
        RECT 69.990000 197.630000 70.190000 197.830000 ;
        RECT 69.990000 198.035000 70.190000 198.235000 ;
        RECT 69.990000 198.440000 70.190000 198.640000 ;
        RECT 69.990000 198.845000 70.190000 199.045000 ;
        RECT 69.990000 199.250000 70.190000 199.450000 ;
        RECT 69.990000 199.655000 70.190000 199.855000 ;
        RECT 70.355000  25.910000 70.555000  26.110000 ;
        RECT 70.355000  26.340000 70.555000  26.540000 ;
        RECT 70.355000  26.770000 70.555000  26.970000 ;
        RECT 70.355000  27.200000 70.555000  27.400000 ;
        RECT 70.355000  27.630000 70.555000  27.830000 ;
        RECT 70.355000  28.060000 70.555000  28.260000 ;
        RECT 70.355000  28.490000 70.555000  28.690000 ;
        RECT 70.355000  28.920000 70.555000  29.120000 ;
        RECT 70.355000  29.350000 70.555000  29.550000 ;
        RECT 70.355000  29.780000 70.555000  29.980000 ;
        RECT 70.355000  30.210000 70.555000  30.410000 ;
        RECT 70.390000 175.995000 70.590000 176.195000 ;
        RECT 70.390000 176.395000 70.590000 176.595000 ;
        RECT 70.390000 176.795000 70.590000 176.995000 ;
        RECT 70.390000 177.195000 70.590000 177.395000 ;
        RECT 70.390000 177.595000 70.590000 177.795000 ;
        RECT 70.390000 177.995000 70.590000 178.195000 ;
        RECT 70.390000 178.395000 70.590000 178.595000 ;
        RECT 70.390000 178.795000 70.590000 178.995000 ;
        RECT 70.390000 179.195000 70.590000 179.395000 ;
        RECT 70.390000 179.595000 70.590000 179.795000 ;
        RECT 70.390000 179.995000 70.590000 180.195000 ;
        RECT 70.390000 180.395000 70.590000 180.595000 ;
        RECT 70.390000 180.795000 70.590000 180.995000 ;
        RECT 70.390000 181.195000 70.590000 181.395000 ;
        RECT 70.390000 181.595000 70.590000 181.795000 ;
        RECT 70.390000 181.995000 70.590000 182.195000 ;
        RECT 70.390000 182.395000 70.590000 182.595000 ;
        RECT 70.390000 182.795000 70.590000 182.995000 ;
        RECT 70.390000 183.195000 70.590000 183.395000 ;
        RECT 70.390000 183.595000 70.590000 183.795000 ;
        RECT 70.390000 183.995000 70.590000 184.195000 ;
        RECT 70.390000 184.395000 70.590000 184.595000 ;
        RECT 70.390000 184.795000 70.590000 184.995000 ;
        RECT 70.390000 185.195000 70.590000 185.395000 ;
        RECT 70.390000 185.595000 70.590000 185.795000 ;
        RECT 70.390000 185.995000 70.590000 186.195000 ;
        RECT 70.390000 186.395000 70.590000 186.595000 ;
        RECT 70.390000 186.795000 70.590000 186.995000 ;
        RECT 70.390000 187.195000 70.590000 187.395000 ;
        RECT 70.390000 187.595000 70.590000 187.795000 ;
        RECT 70.390000 187.995000 70.590000 188.195000 ;
        RECT 70.390000 188.395000 70.590000 188.595000 ;
        RECT 70.390000 188.795000 70.590000 188.995000 ;
        RECT 70.390000 189.195000 70.590000 189.395000 ;
        RECT 70.390000 189.595000 70.590000 189.795000 ;
        RECT 70.390000 189.995000 70.590000 190.195000 ;
        RECT 70.390000 190.395000 70.590000 190.595000 ;
        RECT 70.390000 190.795000 70.590000 190.995000 ;
        RECT 70.390000 191.195000 70.590000 191.395000 ;
        RECT 70.390000 191.595000 70.590000 191.795000 ;
        RECT 70.390000 191.995000 70.590000 192.195000 ;
        RECT 70.390000 192.395000 70.590000 192.595000 ;
        RECT 70.390000 192.795000 70.590000 192.995000 ;
        RECT 70.390000 193.195000 70.590000 193.395000 ;
        RECT 70.390000 193.595000 70.590000 193.795000 ;
        RECT 70.390000 193.995000 70.590000 194.195000 ;
        RECT 70.390000 194.395000 70.590000 194.595000 ;
        RECT 70.390000 194.795000 70.590000 194.995000 ;
        RECT 70.390000 195.200000 70.590000 195.400000 ;
        RECT 70.390000 195.605000 70.590000 195.805000 ;
        RECT 70.390000 196.010000 70.590000 196.210000 ;
        RECT 70.390000 196.415000 70.590000 196.615000 ;
        RECT 70.390000 196.820000 70.590000 197.020000 ;
        RECT 70.390000 197.225000 70.590000 197.425000 ;
        RECT 70.390000 197.630000 70.590000 197.830000 ;
        RECT 70.390000 198.035000 70.590000 198.235000 ;
        RECT 70.390000 198.440000 70.590000 198.640000 ;
        RECT 70.390000 198.845000 70.590000 199.045000 ;
        RECT 70.390000 199.250000 70.590000 199.450000 ;
        RECT 70.390000 199.655000 70.590000 199.855000 ;
        RECT 70.760000  25.910000 70.960000  26.110000 ;
        RECT 70.760000  26.340000 70.960000  26.540000 ;
        RECT 70.760000  26.770000 70.960000  26.970000 ;
        RECT 70.760000  27.200000 70.960000  27.400000 ;
        RECT 70.760000  27.630000 70.960000  27.830000 ;
        RECT 70.760000  28.060000 70.960000  28.260000 ;
        RECT 70.760000  28.490000 70.960000  28.690000 ;
        RECT 70.760000  28.920000 70.960000  29.120000 ;
        RECT 70.760000  29.350000 70.960000  29.550000 ;
        RECT 70.760000  29.780000 70.960000  29.980000 ;
        RECT 70.760000  30.210000 70.960000  30.410000 ;
        RECT 70.790000 175.995000 70.990000 176.195000 ;
        RECT 70.790000 176.395000 70.990000 176.595000 ;
        RECT 70.790000 176.795000 70.990000 176.995000 ;
        RECT 70.790000 177.195000 70.990000 177.395000 ;
        RECT 70.790000 177.595000 70.990000 177.795000 ;
        RECT 70.790000 177.995000 70.990000 178.195000 ;
        RECT 70.790000 178.395000 70.990000 178.595000 ;
        RECT 70.790000 178.795000 70.990000 178.995000 ;
        RECT 70.790000 179.195000 70.990000 179.395000 ;
        RECT 70.790000 179.595000 70.990000 179.795000 ;
        RECT 70.790000 179.995000 70.990000 180.195000 ;
        RECT 70.790000 180.395000 70.990000 180.595000 ;
        RECT 70.790000 180.795000 70.990000 180.995000 ;
        RECT 70.790000 181.195000 70.990000 181.395000 ;
        RECT 70.790000 181.595000 70.990000 181.795000 ;
        RECT 70.790000 181.995000 70.990000 182.195000 ;
        RECT 70.790000 182.395000 70.990000 182.595000 ;
        RECT 70.790000 182.795000 70.990000 182.995000 ;
        RECT 70.790000 183.195000 70.990000 183.395000 ;
        RECT 70.790000 183.595000 70.990000 183.795000 ;
        RECT 70.790000 183.995000 70.990000 184.195000 ;
        RECT 70.790000 184.395000 70.990000 184.595000 ;
        RECT 70.790000 184.795000 70.990000 184.995000 ;
        RECT 70.790000 185.195000 70.990000 185.395000 ;
        RECT 70.790000 185.595000 70.990000 185.795000 ;
        RECT 70.790000 185.995000 70.990000 186.195000 ;
        RECT 70.790000 186.395000 70.990000 186.595000 ;
        RECT 70.790000 186.795000 70.990000 186.995000 ;
        RECT 70.790000 187.195000 70.990000 187.395000 ;
        RECT 70.790000 187.595000 70.990000 187.795000 ;
        RECT 70.790000 187.995000 70.990000 188.195000 ;
        RECT 70.790000 188.395000 70.990000 188.595000 ;
        RECT 70.790000 188.795000 70.990000 188.995000 ;
        RECT 70.790000 189.195000 70.990000 189.395000 ;
        RECT 70.790000 189.595000 70.990000 189.795000 ;
        RECT 70.790000 189.995000 70.990000 190.195000 ;
        RECT 70.790000 190.395000 70.990000 190.595000 ;
        RECT 70.790000 190.795000 70.990000 190.995000 ;
        RECT 70.790000 191.195000 70.990000 191.395000 ;
        RECT 70.790000 191.595000 70.990000 191.795000 ;
        RECT 70.790000 191.995000 70.990000 192.195000 ;
        RECT 70.790000 192.395000 70.990000 192.595000 ;
        RECT 70.790000 192.795000 70.990000 192.995000 ;
        RECT 70.790000 193.195000 70.990000 193.395000 ;
        RECT 70.790000 193.595000 70.990000 193.795000 ;
        RECT 70.790000 193.995000 70.990000 194.195000 ;
        RECT 70.790000 194.395000 70.990000 194.595000 ;
        RECT 70.790000 194.795000 70.990000 194.995000 ;
        RECT 70.790000 195.200000 70.990000 195.400000 ;
        RECT 70.790000 195.605000 70.990000 195.805000 ;
        RECT 70.790000 196.010000 70.990000 196.210000 ;
        RECT 70.790000 196.415000 70.990000 196.615000 ;
        RECT 70.790000 196.820000 70.990000 197.020000 ;
        RECT 70.790000 197.225000 70.990000 197.425000 ;
        RECT 70.790000 197.630000 70.990000 197.830000 ;
        RECT 70.790000 198.035000 70.990000 198.235000 ;
        RECT 70.790000 198.440000 70.990000 198.640000 ;
        RECT 70.790000 198.845000 70.990000 199.045000 ;
        RECT 70.790000 199.250000 70.990000 199.450000 ;
        RECT 70.790000 199.655000 70.990000 199.855000 ;
        RECT 71.165000  25.910000 71.365000  26.110000 ;
        RECT 71.165000  26.340000 71.365000  26.540000 ;
        RECT 71.165000  26.770000 71.365000  26.970000 ;
        RECT 71.165000  27.200000 71.365000  27.400000 ;
        RECT 71.165000  27.630000 71.365000  27.830000 ;
        RECT 71.165000  28.060000 71.365000  28.260000 ;
        RECT 71.165000  28.490000 71.365000  28.690000 ;
        RECT 71.165000  28.920000 71.365000  29.120000 ;
        RECT 71.165000  29.350000 71.365000  29.550000 ;
        RECT 71.165000  29.780000 71.365000  29.980000 ;
        RECT 71.165000  30.210000 71.365000  30.410000 ;
        RECT 71.190000 175.995000 71.390000 176.195000 ;
        RECT 71.190000 176.395000 71.390000 176.595000 ;
        RECT 71.190000 176.795000 71.390000 176.995000 ;
        RECT 71.190000 177.195000 71.390000 177.395000 ;
        RECT 71.190000 177.595000 71.390000 177.795000 ;
        RECT 71.190000 177.995000 71.390000 178.195000 ;
        RECT 71.190000 178.395000 71.390000 178.595000 ;
        RECT 71.190000 178.795000 71.390000 178.995000 ;
        RECT 71.190000 179.195000 71.390000 179.395000 ;
        RECT 71.190000 179.595000 71.390000 179.795000 ;
        RECT 71.190000 179.995000 71.390000 180.195000 ;
        RECT 71.190000 180.395000 71.390000 180.595000 ;
        RECT 71.190000 180.795000 71.390000 180.995000 ;
        RECT 71.190000 181.195000 71.390000 181.395000 ;
        RECT 71.190000 181.595000 71.390000 181.795000 ;
        RECT 71.190000 181.995000 71.390000 182.195000 ;
        RECT 71.190000 182.395000 71.390000 182.595000 ;
        RECT 71.190000 182.795000 71.390000 182.995000 ;
        RECT 71.190000 183.195000 71.390000 183.395000 ;
        RECT 71.190000 183.595000 71.390000 183.795000 ;
        RECT 71.190000 183.995000 71.390000 184.195000 ;
        RECT 71.190000 184.395000 71.390000 184.595000 ;
        RECT 71.190000 184.795000 71.390000 184.995000 ;
        RECT 71.190000 185.195000 71.390000 185.395000 ;
        RECT 71.190000 185.595000 71.390000 185.795000 ;
        RECT 71.190000 185.995000 71.390000 186.195000 ;
        RECT 71.190000 186.395000 71.390000 186.595000 ;
        RECT 71.190000 186.795000 71.390000 186.995000 ;
        RECT 71.190000 187.195000 71.390000 187.395000 ;
        RECT 71.190000 187.595000 71.390000 187.795000 ;
        RECT 71.190000 187.995000 71.390000 188.195000 ;
        RECT 71.190000 188.395000 71.390000 188.595000 ;
        RECT 71.190000 188.795000 71.390000 188.995000 ;
        RECT 71.190000 189.195000 71.390000 189.395000 ;
        RECT 71.190000 189.595000 71.390000 189.795000 ;
        RECT 71.190000 189.995000 71.390000 190.195000 ;
        RECT 71.190000 190.395000 71.390000 190.595000 ;
        RECT 71.190000 190.795000 71.390000 190.995000 ;
        RECT 71.190000 191.195000 71.390000 191.395000 ;
        RECT 71.190000 191.595000 71.390000 191.795000 ;
        RECT 71.190000 191.995000 71.390000 192.195000 ;
        RECT 71.190000 192.395000 71.390000 192.595000 ;
        RECT 71.190000 192.795000 71.390000 192.995000 ;
        RECT 71.190000 193.195000 71.390000 193.395000 ;
        RECT 71.190000 193.595000 71.390000 193.795000 ;
        RECT 71.190000 193.995000 71.390000 194.195000 ;
        RECT 71.190000 194.395000 71.390000 194.595000 ;
        RECT 71.190000 194.795000 71.390000 194.995000 ;
        RECT 71.190000 195.200000 71.390000 195.400000 ;
        RECT 71.190000 195.605000 71.390000 195.805000 ;
        RECT 71.190000 196.010000 71.390000 196.210000 ;
        RECT 71.190000 196.415000 71.390000 196.615000 ;
        RECT 71.190000 196.820000 71.390000 197.020000 ;
        RECT 71.190000 197.225000 71.390000 197.425000 ;
        RECT 71.190000 197.630000 71.390000 197.830000 ;
        RECT 71.190000 198.035000 71.390000 198.235000 ;
        RECT 71.190000 198.440000 71.390000 198.640000 ;
        RECT 71.190000 198.845000 71.390000 199.045000 ;
        RECT 71.190000 199.250000 71.390000 199.450000 ;
        RECT 71.190000 199.655000 71.390000 199.855000 ;
        RECT 71.570000  25.910000 71.770000  26.110000 ;
        RECT 71.570000  26.340000 71.770000  26.540000 ;
        RECT 71.570000  26.770000 71.770000  26.970000 ;
        RECT 71.570000  27.200000 71.770000  27.400000 ;
        RECT 71.570000  27.630000 71.770000  27.830000 ;
        RECT 71.570000  28.060000 71.770000  28.260000 ;
        RECT 71.570000  28.490000 71.770000  28.690000 ;
        RECT 71.570000  28.920000 71.770000  29.120000 ;
        RECT 71.570000  29.350000 71.770000  29.550000 ;
        RECT 71.570000  29.780000 71.770000  29.980000 ;
        RECT 71.570000  30.210000 71.770000  30.410000 ;
        RECT 71.590000 175.995000 71.790000 176.195000 ;
        RECT 71.590000 176.395000 71.790000 176.595000 ;
        RECT 71.590000 176.795000 71.790000 176.995000 ;
        RECT 71.590000 177.195000 71.790000 177.395000 ;
        RECT 71.590000 177.595000 71.790000 177.795000 ;
        RECT 71.590000 177.995000 71.790000 178.195000 ;
        RECT 71.590000 178.395000 71.790000 178.595000 ;
        RECT 71.590000 178.795000 71.790000 178.995000 ;
        RECT 71.590000 179.195000 71.790000 179.395000 ;
        RECT 71.590000 179.595000 71.790000 179.795000 ;
        RECT 71.590000 179.995000 71.790000 180.195000 ;
        RECT 71.590000 180.395000 71.790000 180.595000 ;
        RECT 71.590000 180.795000 71.790000 180.995000 ;
        RECT 71.590000 181.195000 71.790000 181.395000 ;
        RECT 71.590000 181.595000 71.790000 181.795000 ;
        RECT 71.590000 181.995000 71.790000 182.195000 ;
        RECT 71.590000 182.395000 71.790000 182.595000 ;
        RECT 71.590000 182.795000 71.790000 182.995000 ;
        RECT 71.590000 183.195000 71.790000 183.395000 ;
        RECT 71.590000 183.595000 71.790000 183.795000 ;
        RECT 71.590000 183.995000 71.790000 184.195000 ;
        RECT 71.590000 184.395000 71.790000 184.595000 ;
        RECT 71.590000 184.795000 71.790000 184.995000 ;
        RECT 71.590000 185.195000 71.790000 185.395000 ;
        RECT 71.590000 185.595000 71.790000 185.795000 ;
        RECT 71.590000 185.995000 71.790000 186.195000 ;
        RECT 71.590000 186.395000 71.790000 186.595000 ;
        RECT 71.590000 186.795000 71.790000 186.995000 ;
        RECT 71.590000 187.195000 71.790000 187.395000 ;
        RECT 71.590000 187.595000 71.790000 187.795000 ;
        RECT 71.590000 187.995000 71.790000 188.195000 ;
        RECT 71.590000 188.395000 71.790000 188.595000 ;
        RECT 71.590000 188.795000 71.790000 188.995000 ;
        RECT 71.590000 189.195000 71.790000 189.395000 ;
        RECT 71.590000 189.595000 71.790000 189.795000 ;
        RECT 71.590000 189.995000 71.790000 190.195000 ;
        RECT 71.590000 190.395000 71.790000 190.595000 ;
        RECT 71.590000 190.795000 71.790000 190.995000 ;
        RECT 71.590000 191.195000 71.790000 191.395000 ;
        RECT 71.590000 191.595000 71.790000 191.795000 ;
        RECT 71.590000 191.995000 71.790000 192.195000 ;
        RECT 71.590000 192.395000 71.790000 192.595000 ;
        RECT 71.590000 192.795000 71.790000 192.995000 ;
        RECT 71.590000 193.195000 71.790000 193.395000 ;
        RECT 71.590000 193.595000 71.790000 193.795000 ;
        RECT 71.590000 193.995000 71.790000 194.195000 ;
        RECT 71.590000 194.395000 71.790000 194.595000 ;
        RECT 71.590000 194.795000 71.790000 194.995000 ;
        RECT 71.590000 195.200000 71.790000 195.400000 ;
        RECT 71.590000 195.605000 71.790000 195.805000 ;
        RECT 71.590000 196.010000 71.790000 196.210000 ;
        RECT 71.590000 196.415000 71.790000 196.615000 ;
        RECT 71.590000 196.820000 71.790000 197.020000 ;
        RECT 71.590000 197.225000 71.790000 197.425000 ;
        RECT 71.590000 197.630000 71.790000 197.830000 ;
        RECT 71.590000 198.035000 71.790000 198.235000 ;
        RECT 71.590000 198.440000 71.790000 198.640000 ;
        RECT 71.590000 198.845000 71.790000 199.045000 ;
        RECT 71.590000 199.250000 71.790000 199.450000 ;
        RECT 71.590000 199.655000 71.790000 199.855000 ;
        RECT 71.975000  25.910000 72.175000  26.110000 ;
        RECT 71.975000  26.340000 72.175000  26.540000 ;
        RECT 71.975000  26.770000 72.175000  26.970000 ;
        RECT 71.975000  27.200000 72.175000  27.400000 ;
        RECT 71.975000  27.630000 72.175000  27.830000 ;
        RECT 71.975000  28.060000 72.175000  28.260000 ;
        RECT 71.975000  28.490000 72.175000  28.690000 ;
        RECT 71.975000  28.920000 72.175000  29.120000 ;
        RECT 71.975000  29.350000 72.175000  29.550000 ;
        RECT 71.975000  29.780000 72.175000  29.980000 ;
        RECT 71.975000  30.210000 72.175000  30.410000 ;
        RECT 71.990000 175.995000 72.190000 176.195000 ;
        RECT 71.990000 176.395000 72.190000 176.595000 ;
        RECT 71.990000 176.795000 72.190000 176.995000 ;
        RECT 71.990000 177.195000 72.190000 177.395000 ;
        RECT 71.990000 177.595000 72.190000 177.795000 ;
        RECT 71.990000 177.995000 72.190000 178.195000 ;
        RECT 71.990000 178.395000 72.190000 178.595000 ;
        RECT 71.990000 178.795000 72.190000 178.995000 ;
        RECT 71.990000 179.195000 72.190000 179.395000 ;
        RECT 71.990000 179.595000 72.190000 179.795000 ;
        RECT 71.990000 179.995000 72.190000 180.195000 ;
        RECT 71.990000 180.395000 72.190000 180.595000 ;
        RECT 71.990000 180.795000 72.190000 180.995000 ;
        RECT 71.990000 181.195000 72.190000 181.395000 ;
        RECT 71.990000 181.595000 72.190000 181.795000 ;
        RECT 71.990000 181.995000 72.190000 182.195000 ;
        RECT 71.990000 182.395000 72.190000 182.595000 ;
        RECT 71.990000 182.795000 72.190000 182.995000 ;
        RECT 71.990000 183.195000 72.190000 183.395000 ;
        RECT 71.990000 183.595000 72.190000 183.795000 ;
        RECT 71.990000 183.995000 72.190000 184.195000 ;
        RECT 71.990000 184.395000 72.190000 184.595000 ;
        RECT 71.990000 184.795000 72.190000 184.995000 ;
        RECT 71.990000 185.195000 72.190000 185.395000 ;
        RECT 71.990000 185.595000 72.190000 185.795000 ;
        RECT 71.990000 185.995000 72.190000 186.195000 ;
        RECT 71.990000 186.395000 72.190000 186.595000 ;
        RECT 71.990000 186.795000 72.190000 186.995000 ;
        RECT 71.990000 187.195000 72.190000 187.395000 ;
        RECT 71.990000 187.595000 72.190000 187.795000 ;
        RECT 71.990000 187.995000 72.190000 188.195000 ;
        RECT 71.990000 188.395000 72.190000 188.595000 ;
        RECT 71.990000 188.795000 72.190000 188.995000 ;
        RECT 71.990000 189.195000 72.190000 189.395000 ;
        RECT 71.990000 189.595000 72.190000 189.795000 ;
        RECT 71.990000 189.995000 72.190000 190.195000 ;
        RECT 71.990000 190.395000 72.190000 190.595000 ;
        RECT 71.990000 190.795000 72.190000 190.995000 ;
        RECT 71.990000 191.195000 72.190000 191.395000 ;
        RECT 71.990000 191.595000 72.190000 191.795000 ;
        RECT 71.990000 191.995000 72.190000 192.195000 ;
        RECT 71.990000 192.395000 72.190000 192.595000 ;
        RECT 71.990000 192.795000 72.190000 192.995000 ;
        RECT 71.990000 193.195000 72.190000 193.395000 ;
        RECT 71.990000 193.595000 72.190000 193.795000 ;
        RECT 71.990000 193.995000 72.190000 194.195000 ;
        RECT 71.990000 194.395000 72.190000 194.595000 ;
        RECT 71.990000 194.795000 72.190000 194.995000 ;
        RECT 71.990000 195.200000 72.190000 195.400000 ;
        RECT 71.990000 195.605000 72.190000 195.805000 ;
        RECT 71.990000 196.010000 72.190000 196.210000 ;
        RECT 71.990000 196.415000 72.190000 196.615000 ;
        RECT 71.990000 196.820000 72.190000 197.020000 ;
        RECT 71.990000 197.225000 72.190000 197.425000 ;
        RECT 71.990000 197.630000 72.190000 197.830000 ;
        RECT 71.990000 198.035000 72.190000 198.235000 ;
        RECT 71.990000 198.440000 72.190000 198.640000 ;
        RECT 71.990000 198.845000 72.190000 199.045000 ;
        RECT 71.990000 199.250000 72.190000 199.450000 ;
        RECT 71.990000 199.655000 72.190000 199.855000 ;
        RECT 72.380000  25.910000 72.580000  26.110000 ;
        RECT 72.380000  26.340000 72.580000  26.540000 ;
        RECT 72.380000  26.770000 72.580000  26.970000 ;
        RECT 72.380000  27.200000 72.580000  27.400000 ;
        RECT 72.380000  27.630000 72.580000  27.830000 ;
        RECT 72.380000  28.060000 72.580000  28.260000 ;
        RECT 72.380000  28.490000 72.580000  28.690000 ;
        RECT 72.380000  28.920000 72.580000  29.120000 ;
        RECT 72.380000  29.350000 72.580000  29.550000 ;
        RECT 72.380000  29.780000 72.580000  29.980000 ;
        RECT 72.380000  30.210000 72.580000  30.410000 ;
        RECT 72.390000 175.995000 72.590000 176.195000 ;
        RECT 72.390000 176.395000 72.590000 176.595000 ;
        RECT 72.390000 176.795000 72.590000 176.995000 ;
        RECT 72.390000 177.195000 72.590000 177.395000 ;
        RECT 72.390000 177.595000 72.590000 177.795000 ;
        RECT 72.390000 177.995000 72.590000 178.195000 ;
        RECT 72.390000 178.395000 72.590000 178.595000 ;
        RECT 72.390000 178.795000 72.590000 178.995000 ;
        RECT 72.390000 179.195000 72.590000 179.395000 ;
        RECT 72.390000 179.595000 72.590000 179.795000 ;
        RECT 72.390000 179.995000 72.590000 180.195000 ;
        RECT 72.390000 180.395000 72.590000 180.595000 ;
        RECT 72.390000 180.795000 72.590000 180.995000 ;
        RECT 72.390000 181.195000 72.590000 181.395000 ;
        RECT 72.390000 181.595000 72.590000 181.795000 ;
        RECT 72.390000 181.995000 72.590000 182.195000 ;
        RECT 72.390000 182.395000 72.590000 182.595000 ;
        RECT 72.390000 182.795000 72.590000 182.995000 ;
        RECT 72.390000 183.195000 72.590000 183.395000 ;
        RECT 72.390000 183.595000 72.590000 183.795000 ;
        RECT 72.390000 183.995000 72.590000 184.195000 ;
        RECT 72.390000 184.395000 72.590000 184.595000 ;
        RECT 72.390000 184.795000 72.590000 184.995000 ;
        RECT 72.390000 185.195000 72.590000 185.395000 ;
        RECT 72.390000 185.595000 72.590000 185.795000 ;
        RECT 72.390000 185.995000 72.590000 186.195000 ;
        RECT 72.390000 186.395000 72.590000 186.595000 ;
        RECT 72.390000 186.795000 72.590000 186.995000 ;
        RECT 72.390000 187.195000 72.590000 187.395000 ;
        RECT 72.390000 187.595000 72.590000 187.795000 ;
        RECT 72.390000 187.995000 72.590000 188.195000 ;
        RECT 72.390000 188.395000 72.590000 188.595000 ;
        RECT 72.390000 188.795000 72.590000 188.995000 ;
        RECT 72.390000 189.195000 72.590000 189.395000 ;
        RECT 72.390000 189.595000 72.590000 189.795000 ;
        RECT 72.390000 189.995000 72.590000 190.195000 ;
        RECT 72.390000 190.395000 72.590000 190.595000 ;
        RECT 72.390000 190.795000 72.590000 190.995000 ;
        RECT 72.390000 191.195000 72.590000 191.395000 ;
        RECT 72.390000 191.595000 72.590000 191.795000 ;
        RECT 72.390000 191.995000 72.590000 192.195000 ;
        RECT 72.390000 192.395000 72.590000 192.595000 ;
        RECT 72.390000 192.795000 72.590000 192.995000 ;
        RECT 72.390000 193.195000 72.590000 193.395000 ;
        RECT 72.390000 193.595000 72.590000 193.795000 ;
        RECT 72.390000 193.995000 72.590000 194.195000 ;
        RECT 72.390000 194.395000 72.590000 194.595000 ;
        RECT 72.390000 194.795000 72.590000 194.995000 ;
        RECT 72.390000 195.200000 72.590000 195.400000 ;
        RECT 72.390000 195.605000 72.590000 195.805000 ;
        RECT 72.390000 196.010000 72.590000 196.210000 ;
        RECT 72.390000 196.415000 72.590000 196.615000 ;
        RECT 72.390000 196.820000 72.590000 197.020000 ;
        RECT 72.390000 197.225000 72.590000 197.425000 ;
        RECT 72.390000 197.630000 72.590000 197.830000 ;
        RECT 72.390000 198.035000 72.590000 198.235000 ;
        RECT 72.390000 198.440000 72.590000 198.640000 ;
        RECT 72.390000 198.845000 72.590000 199.045000 ;
        RECT 72.390000 199.250000 72.590000 199.450000 ;
        RECT 72.390000 199.655000 72.590000 199.855000 ;
        RECT 72.785000  25.910000 72.985000  26.110000 ;
        RECT 72.785000  26.340000 72.985000  26.540000 ;
        RECT 72.785000  26.770000 72.985000  26.970000 ;
        RECT 72.785000  27.200000 72.985000  27.400000 ;
        RECT 72.785000  27.630000 72.985000  27.830000 ;
        RECT 72.785000  28.060000 72.985000  28.260000 ;
        RECT 72.785000  28.490000 72.985000  28.690000 ;
        RECT 72.785000  28.920000 72.985000  29.120000 ;
        RECT 72.785000  29.350000 72.985000  29.550000 ;
        RECT 72.785000  29.780000 72.985000  29.980000 ;
        RECT 72.785000  30.210000 72.985000  30.410000 ;
        RECT 72.790000 175.995000 72.990000 176.195000 ;
        RECT 72.790000 176.395000 72.990000 176.595000 ;
        RECT 72.790000 176.795000 72.990000 176.995000 ;
        RECT 72.790000 177.195000 72.990000 177.395000 ;
        RECT 72.790000 177.595000 72.990000 177.795000 ;
        RECT 72.790000 177.995000 72.990000 178.195000 ;
        RECT 72.790000 178.395000 72.990000 178.595000 ;
        RECT 72.790000 178.795000 72.990000 178.995000 ;
        RECT 72.790000 179.195000 72.990000 179.395000 ;
        RECT 72.790000 179.595000 72.990000 179.795000 ;
        RECT 72.790000 179.995000 72.990000 180.195000 ;
        RECT 72.790000 180.395000 72.990000 180.595000 ;
        RECT 72.790000 180.795000 72.990000 180.995000 ;
        RECT 72.790000 181.195000 72.990000 181.395000 ;
        RECT 72.790000 181.595000 72.990000 181.795000 ;
        RECT 72.790000 181.995000 72.990000 182.195000 ;
        RECT 72.790000 182.395000 72.990000 182.595000 ;
        RECT 72.790000 182.795000 72.990000 182.995000 ;
        RECT 72.790000 183.195000 72.990000 183.395000 ;
        RECT 72.790000 183.595000 72.990000 183.795000 ;
        RECT 72.790000 183.995000 72.990000 184.195000 ;
        RECT 72.790000 184.395000 72.990000 184.595000 ;
        RECT 72.790000 184.795000 72.990000 184.995000 ;
        RECT 72.790000 185.195000 72.990000 185.395000 ;
        RECT 72.790000 185.595000 72.990000 185.795000 ;
        RECT 72.790000 185.995000 72.990000 186.195000 ;
        RECT 72.790000 186.395000 72.990000 186.595000 ;
        RECT 72.790000 186.795000 72.990000 186.995000 ;
        RECT 72.790000 187.195000 72.990000 187.395000 ;
        RECT 72.790000 187.595000 72.990000 187.795000 ;
        RECT 72.790000 187.995000 72.990000 188.195000 ;
        RECT 72.790000 188.395000 72.990000 188.595000 ;
        RECT 72.790000 188.795000 72.990000 188.995000 ;
        RECT 72.790000 189.195000 72.990000 189.395000 ;
        RECT 72.790000 189.595000 72.990000 189.795000 ;
        RECT 72.790000 189.995000 72.990000 190.195000 ;
        RECT 72.790000 190.395000 72.990000 190.595000 ;
        RECT 72.790000 190.795000 72.990000 190.995000 ;
        RECT 72.790000 191.195000 72.990000 191.395000 ;
        RECT 72.790000 191.595000 72.990000 191.795000 ;
        RECT 72.790000 191.995000 72.990000 192.195000 ;
        RECT 72.790000 192.395000 72.990000 192.595000 ;
        RECT 72.790000 192.795000 72.990000 192.995000 ;
        RECT 72.790000 193.195000 72.990000 193.395000 ;
        RECT 72.790000 193.595000 72.990000 193.795000 ;
        RECT 72.790000 193.995000 72.990000 194.195000 ;
        RECT 72.790000 194.395000 72.990000 194.595000 ;
        RECT 72.790000 194.795000 72.990000 194.995000 ;
        RECT 72.790000 195.200000 72.990000 195.400000 ;
        RECT 72.790000 195.605000 72.990000 195.805000 ;
        RECT 72.790000 196.010000 72.990000 196.210000 ;
        RECT 72.790000 196.415000 72.990000 196.615000 ;
        RECT 72.790000 196.820000 72.990000 197.020000 ;
        RECT 72.790000 197.225000 72.990000 197.425000 ;
        RECT 72.790000 197.630000 72.990000 197.830000 ;
        RECT 72.790000 198.035000 72.990000 198.235000 ;
        RECT 72.790000 198.440000 72.990000 198.640000 ;
        RECT 72.790000 198.845000 72.990000 199.045000 ;
        RECT 72.790000 199.250000 72.990000 199.450000 ;
        RECT 72.790000 199.655000 72.990000 199.855000 ;
        RECT 73.190000  25.910000 73.390000  26.110000 ;
        RECT 73.190000  26.340000 73.390000  26.540000 ;
        RECT 73.190000  26.770000 73.390000  26.970000 ;
        RECT 73.190000  27.200000 73.390000  27.400000 ;
        RECT 73.190000  27.630000 73.390000  27.830000 ;
        RECT 73.190000  28.060000 73.390000  28.260000 ;
        RECT 73.190000  28.490000 73.390000  28.690000 ;
        RECT 73.190000  28.920000 73.390000  29.120000 ;
        RECT 73.190000  29.350000 73.390000  29.550000 ;
        RECT 73.190000  29.780000 73.390000  29.980000 ;
        RECT 73.190000  30.210000 73.390000  30.410000 ;
        RECT 73.190000 175.995000 73.390000 176.195000 ;
        RECT 73.190000 176.395000 73.390000 176.595000 ;
        RECT 73.190000 176.795000 73.390000 176.995000 ;
        RECT 73.190000 177.195000 73.390000 177.395000 ;
        RECT 73.190000 177.595000 73.390000 177.795000 ;
        RECT 73.190000 177.995000 73.390000 178.195000 ;
        RECT 73.190000 178.395000 73.390000 178.595000 ;
        RECT 73.190000 178.795000 73.390000 178.995000 ;
        RECT 73.190000 179.195000 73.390000 179.395000 ;
        RECT 73.190000 179.595000 73.390000 179.795000 ;
        RECT 73.190000 179.995000 73.390000 180.195000 ;
        RECT 73.190000 180.395000 73.390000 180.595000 ;
        RECT 73.190000 180.795000 73.390000 180.995000 ;
        RECT 73.190000 181.195000 73.390000 181.395000 ;
        RECT 73.190000 181.595000 73.390000 181.795000 ;
        RECT 73.190000 181.995000 73.390000 182.195000 ;
        RECT 73.190000 182.395000 73.390000 182.595000 ;
        RECT 73.190000 182.795000 73.390000 182.995000 ;
        RECT 73.190000 183.195000 73.390000 183.395000 ;
        RECT 73.190000 183.595000 73.390000 183.795000 ;
        RECT 73.190000 183.995000 73.390000 184.195000 ;
        RECT 73.190000 184.395000 73.390000 184.595000 ;
        RECT 73.190000 184.795000 73.390000 184.995000 ;
        RECT 73.190000 185.195000 73.390000 185.395000 ;
        RECT 73.190000 185.595000 73.390000 185.795000 ;
        RECT 73.190000 185.995000 73.390000 186.195000 ;
        RECT 73.190000 186.395000 73.390000 186.595000 ;
        RECT 73.190000 186.795000 73.390000 186.995000 ;
        RECT 73.190000 187.195000 73.390000 187.395000 ;
        RECT 73.190000 187.595000 73.390000 187.795000 ;
        RECT 73.190000 187.995000 73.390000 188.195000 ;
        RECT 73.190000 188.395000 73.390000 188.595000 ;
        RECT 73.190000 188.795000 73.390000 188.995000 ;
        RECT 73.190000 189.195000 73.390000 189.395000 ;
        RECT 73.190000 189.595000 73.390000 189.795000 ;
        RECT 73.190000 189.995000 73.390000 190.195000 ;
        RECT 73.190000 190.395000 73.390000 190.595000 ;
        RECT 73.190000 190.795000 73.390000 190.995000 ;
        RECT 73.190000 191.195000 73.390000 191.395000 ;
        RECT 73.190000 191.595000 73.390000 191.795000 ;
        RECT 73.190000 191.995000 73.390000 192.195000 ;
        RECT 73.190000 192.395000 73.390000 192.595000 ;
        RECT 73.190000 192.795000 73.390000 192.995000 ;
        RECT 73.190000 193.195000 73.390000 193.395000 ;
        RECT 73.190000 193.595000 73.390000 193.795000 ;
        RECT 73.190000 193.995000 73.390000 194.195000 ;
        RECT 73.190000 194.395000 73.390000 194.595000 ;
        RECT 73.190000 194.795000 73.390000 194.995000 ;
        RECT 73.190000 195.200000 73.390000 195.400000 ;
        RECT 73.190000 195.605000 73.390000 195.805000 ;
        RECT 73.190000 196.010000 73.390000 196.210000 ;
        RECT 73.190000 196.415000 73.390000 196.615000 ;
        RECT 73.190000 196.820000 73.390000 197.020000 ;
        RECT 73.190000 197.225000 73.390000 197.425000 ;
        RECT 73.190000 197.630000 73.390000 197.830000 ;
        RECT 73.190000 198.035000 73.390000 198.235000 ;
        RECT 73.190000 198.440000 73.390000 198.640000 ;
        RECT 73.190000 198.845000 73.390000 199.045000 ;
        RECT 73.190000 199.250000 73.390000 199.450000 ;
        RECT 73.190000 199.655000 73.390000 199.855000 ;
        RECT 73.590000 175.995000 73.790000 176.195000 ;
        RECT 73.590000 176.395000 73.790000 176.595000 ;
        RECT 73.590000 176.795000 73.790000 176.995000 ;
        RECT 73.590000 177.195000 73.790000 177.395000 ;
        RECT 73.590000 177.595000 73.790000 177.795000 ;
        RECT 73.590000 177.995000 73.790000 178.195000 ;
        RECT 73.590000 178.395000 73.790000 178.595000 ;
        RECT 73.590000 178.795000 73.790000 178.995000 ;
        RECT 73.590000 179.195000 73.790000 179.395000 ;
        RECT 73.590000 179.595000 73.790000 179.795000 ;
        RECT 73.590000 179.995000 73.790000 180.195000 ;
        RECT 73.590000 180.395000 73.790000 180.595000 ;
        RECT 73.590000 180.795000 73.790000 180.995000 ;
        RECT 73.590000 181.195000 73.790000 181.395000 ;
        RECT 73.590000 181.595000 73.790000 181.795000 ;
        RECT 73.590000 181.995000 73.790000 182.195000 ;
        RECT 73.590000 182.395000 73.790000 182.595000 ;
        RECT 73.590000 182.795000 73.790000 182.995000 ;
        RECT 73.590000 183.195000 73.790000 183.395000 ;
        RECT 73.590000 183.595000 73.790000 183.795000 ;
        RECT 73.590000 183.995000 73.790000 184.195000 ;
        RECT 73.590000 184.395000 73.790000 184.595000 ;
        RECT 73.590000 184.795000 73.790000 184.995000 ;
        RECT 73.590000 185.195000 73.790000 185.395000 ;
        RECT 73.590000 185.595000 73.790000 185.795000 ;
        RECT 73.590000 185.995000 73.790000 186.195000 ;
        RECT 73.590000 186.395000 73.790000 186.595000 ;
        RECT 73.590000 186.795000 73.790000 186.995000 ;
        RECT 73.590000 187.195000 73.790000 187.395000 ;
        RECT 73.590000 187.595000 73.790000 187.795000 ;
        RECT 73.590000 187.995000 73.790000 188.195000 ;
        RECT 73.590000 188.395000 73.790000 188.595000 ;
        RECT 73.590000 188.795000 73.790000 188.995000 ;
        RECT 73.590000 189.195000 73.790000 189.395000 ;
        RECT 73.590000 189.595000 73.790000 189.795000 ;
        RECT 73.590000 189.995000 73.790000 190.195000 ;
        RECT 73.590000 190.395000 73.790000 190.595000 ;
        RECT 73.590000 190.795000 73.790000 190.995000 ;
        RECT 73.590000 191.195000 73.790000 191.395000 ;
        RECT 73.590000 191.595000 73.790000 191.795000 ;
        RECT 73.590000 191.995000 73.790000 192.195000 ;
        RECT 73.590000 192.395000 73.790000 192.595000 ;
        RECT 73.590000 192.795000 73.790000 192.995000 ;
        RECT 73.590000 193.195000 73.790000 193.395000 ;
        RECT 73.590000 193.595000 73.790000 193.795000 ;
        RECT 73.590000 193.995000 73.790000 194.195000 ;
        RECT 73.590000 194.395000 73.790000 194.595000 ;
        RECT 73.590000 194.795000 73.790000 194.995000 ;
        RECT 73.590000 195.200000 73.790000 195.400000 ;
        RECT 73.590000 195.605000 73.790000 195.805000 ;
        RECT 73.590000 196.010000 73.790000 196.210000 ;
        RECT 73.590000 196.415000 73.790000 196.615000 ;
        RECT 73.590000 196.820000 73.790000 197.020000 ;
        RECT 73.590000 197.225000 73.790000 197.425000 ;
        RECT 73.590000 197.630000 73.790000 197.830000 ;
        RECT 73.590000 198.035000 73.790000 198.235000 ;
        RECT 73.590000 198.440000 73.790000 198.640000 ;
        RECT 73.590000 198.845000 73.790000 199.045000 ;
        RECT 73.590000 199.250000 73.790000 199.450000 ;
        RECT 73.590000 199.655000 73.790000 199.855000 ;
        RECT 73.595000  25.910000 73.795000  26.110000 ;
        RECT 73.595000  26.340000 73.795000  26.540000 ;
        RECT 73.595000  26.770000 73.795000  26.970000 ;
        RECT 73.595000  27.200000 73.795000  27.400000 ;
        RECT 73.595000  27.630000 73.795000  27.830000 ;
        RECT 73.595000  28.060000 73.795000  28.260000 ;
        RECT 73.595000  28.490000 73.795000  28.690000 ;
        RECT 73.595000  28.920000 73.795000  29.120000 ;
        RECT 73.595000  29.350000 73.795000  29.550000 ;
        RECT 73.595000  29.780000 73.795000  29.980000 ;
        RECT 73.595000  30.210000 73.795000  30.410000 ;
        RECT 73.990000 175.995000 74.190000 176.195000 ;
        RECT 73.990000 176.395000 74.190000 176.595000 ;
        RECT 73.990000 176.795000 74.190000 176.995000 ;
        RECT 73.990000 177.195000 74.190000 177.395000 ;
        RECT 73.990000 177.595000 74.190000 177.795000 ;
        RECT 73.990000 177.995000 74.190000 178.195000 ;
        RECT 73.990000 178.395000 74.190000 178.595000 ;
        RECT 73.990000 178.795000 74.190000 178.995000 ;
        RECT 73.990000 179.195000 74.190000 179.395000 ;
        RECT 73.990000 179.595000 74.190000 179.795000 ;
        RECT 73.990000 179.995000 74.190000 180.195000 ;
        RECT 73.990000 180.395000 74.190000 180.595000 ;
        RECT 73.990000 180.795000 74.190000 180.995000 ;
        RECT 73.990000 181.195000 74.190000 181.395000 ;
        RECT 73.990000 181.595000 74.190000 181.795000 ;
        RECT 73.990000 181.995000 74.190000 182.195000 ;
        RECT 73.990000 182.395000 74.190000 182.595000 ;
        RECT 73.990000 182.795000 74.190000 182.995000 ;
        RECT 73.990000 183.195000 74.190000 183.395000 ;
        RECT 73.990000 183.595000 74.190000 183.795000 ;
        RECT 73.990000 183.995000 74.190000 184.195000 ;
        RECT 73.990000 184.395000 74.190000 184.595000 ;
        RECT 73.990000 184.795000 74.190000 184.995000 ;
        RECT 73.990000 185.195000 74.190000 185.395000 ;
        RECT 73.990000 185.595000 74.190000 185.795000 ;
        RECT 73.990000 185.995000 74.190000 186.195000 ;
        RECT 73.990000 186.395000 74.190000 186.595000 ;
        RECT 73.990000 186.795000 74.190000 186.995000 ;
        RECT 73.990000 187.195000 74.190000 187.395000 ;
        RECT 73.990000 187.595000 74.190000 187.795000 ;
        RECT 73.990000 187.995000 74.190000 188.195000 ;
        RECT 73.990000 188.395000 74.190000 188.595000 ;
        RECT 73.990000 188.795000 74.190000 188.995000 ;
        RECT 73.990000 189.195000 74.190000 189.395000 ;
        RECT 73.990000 189.595000 74.190000 189.795000 ;
        RECT 73.990000 189.995000 74.190000 190.195000 ;
        RECT 73.990000 190.395000 74.190000 190.595000 ;
        RECT 73.990000 190.795000 74.190000 190.995000 ;
        RECT 73.990000 191.195000 74.190000 191.395000 ;
        RECT 73.990000 191.595000 74.190000 191.795000 ;
        RECT 73.990000 191.995000 74.190000 192.195000 ;
        RECT 73.990000 192.395000 74.190000 192.595000 ;
        RECT 73.990000 192.795000 74.190000 192.995000 ;
        RECT 73.990000 193.195000 74.190000 193.395000 ;
        RECT 73.990000 193.595000 74.190000 193.795000 ;
        RECT 73.990000 193.995000 74.190000 194.195000 ;
        RECT 73.990000 194.395000 74.190000 194.595000 ;
        RECT 73.990000 194.795000 74.190000 194.995000 ;
        RECT 73.990000 195.200000 74.190000 195.400000 ;
        RECT 73.990000 195.605000 74.190000 195.805000 ;
        RECT 73.990000 196.010000 74.190000 196.210000 ;
        RECT 73.990000 196.415000 74.190000 196.615000 ;
        RECT 73.990000 196.820000 74.190000 197.020000 ;
        RECT 73.990000 197.225000 74.190000 197.425000 ;
        RECT 73.990000 197.630000 74.190000 197.830000 ;
        RECT 73.990000 198.035000 74.190000 198.235000 ;
        RECT 73.990000 198.440000 74.190000 198.640000 ;
        RECT 73.990000 198.845000 74.190000 199.045000 ;
        RECT 73.990000 199.250000 74.190000 199.450000 ;
        RECT 73.990000 199.655000 74.190000 199.855000 ;
        RECT 74.000000  25.910000 74.200000  26.110000 ;
        RECT 74.000000  26.340000 74.200000  26.540000 ;
        RECT 74.000000  26.770000 74.200000  26.970000 ;
        RECT 74.000000  27.200000 74.200000  27.400000 ;
        RECT 74.000000  27.630000 74.200000  27.830000 ;
        RECT 74.000000  28.060000 74.200000  28.260000 ;
        RECT 74.000000  28.490000 74.200000  28.690000 ;
        RECT 74.000000  28.920000 74.200000  29.120000 ;
        RECT 74.000000  29.350000 74.200000  29.550000 ;
        RECT 74.000000  29.780000 74.200000  29.980000 ;
        RECT 74.000000  30.210000 74.200000  30.410000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.495000 58.240000 24.395000 62.680000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390000 58.240000 74.290000 62.680000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 24.370000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.415000 58.235000 75.000000 62.685000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 58.335000 1.270000 62.585000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
    PORT
      LAYER via3 ;
        RECT  0.585000 58.310000  0.785000 58.510000 ;
        RECT  0.585000 58.720000  0.785000 58.920000 ;
        RECT  0.585000 59.130000  0.785000 59.330000 ;
        RECT  0.585000 59.540000  0.785000 59.740000 ;
        RECT  0.585000 59.950000  0.785000 60.150000 ;
        RECT  0.585000 60.360000  0.785000 60.560000 ;
        RECT  0.585000 60.770000  0.785000 60.970000 ;
        RECT  0.585000 61.180000  0.785000 61.380000 ;
        RECT  0.585000 61.590000  0.785000 61.790000 ;
        RECT  0.585000 62.000000  0.785000 62.200000 ;
        RECT  0.585000 62.410000  0.785000 62.610000 ;
        RECT  0.995000 58.310000  1.195000 58.510000 ;
        RECT  0.995000 58.720000  1.195000 58.920000 ;
        RECT  0.995000 59.130000  1.195000 59.330000 ;
        RECT  0.995000 59.540000  1.195000 59.740000 ;
        RECT  0.995000 59.950000  1.195000 60.150000 ;
        RECT  0.995000 60.360000  1.195000 60.560000 ;
        RECT  0.995000 60.770000  1.195000 60.970000 ;
        RECT  0.995000 61.180000  1.195000 61.380000 ;
        RECT  0.995000 61.590000  1.195000 61.790000 ;
        RECT  0.995000 62.000000  1.195000 62.200000 ;
        RECT  0.995000 62.410000  1.195000 62.610000 ;
        RECT  1.405000 58.310000  1.605000 58.510000 ;
        RECT  1.405000 58.720000  1.605000 58.920000 ;
        RECT  1.405000 59.130000  1.605000 59.330000 ;
        RECT  1.405000 59.540000  1.605000 59.740000 ;
        RECT  1.405000 59.950000  1.605000 60.150000 ;
        RECT  1.405000 60.360000  1.605000 60.560000 ;
        RECT  1.405000 60.770000  1.605000 60.970000 ;
        RECT  1.405000 61.180000  1.605000 61.380000 ;
        RECT  1.405000 61.590000  1.605000 61.790000 ;
        RECT  1.405000 62.000000  1.605000 62.200000 ;
        RECT  1.405000 62.410000  1.605000 62.610000 ;
        RECT  1.815000 58.310000  2.015000 58.510000 ;
        RECT  1.815000 58.720000  2.015000 58.920000 ;
        RECT  1.815000 59.130000  2.015000 59.330000 ;
        RECT  1.815000 59.540000  2.015000 59.740000 ;
        RECT  1.815000 59.950000  2.015000 60.150000 ;
        RECT  1.815000 60.360000  2.015000 60.560000 ;
        RECT  1.815000 60.770000  2.015000 60.970000 ;
        RECT  1.815000 61.180000  2.015000 61.380000 ;
        RECT  1.815000 61.590000  2.015000 61.790000 ;
        RECT  1.815000 62.000000  2.015000 62.200000 ;
        RECT  1.815000 62.410000  2.015000 62.610000 ;
        RECT  2.225000 58.310000  2.425000 58.510000 ;
        RECT  2.225000 58.720000  2.425000 58.920000 ;
        RECT  2.225000 59.130000  2.425000 59.330000 ;
        RECT  2.225000 59.540000  2.425000 59.740000 ;
        RECT  2.225000 59.950000  2.425000 60.150000 ;
        RECT  2.225000 60.360000  2.425000 60.560000 ;
        RECT  2.225000 60.770000  2.425000 60.970000 ;
        RECT  2.225000 61.180000  2.425000 61.380000 ;
        RECT  2.225000 61.590000  2.425000 61.790000 ;
        RECT  2.225000 62.000000  2.425000 62.200000 ;
        RECT  2.225000 62.410000  2.425000 62.610000 ;
        RECT  2.635000 58.310000  2.835000 58.510000 ;
        RECT  2.635000 58.720000  2.835000 58.920000 ;
        RECT  2.635000 59.130000  2.835000 59.330000 ;
        RECT  2.635000 59.540000  2.835000 59.740000 ;
        RECT  2.635000 59.950000  2.835000 60.150000 ;
        RECT  2.635000 60.360000  2.835000 60.560000 ;
        RECT  2.635000 60.770000  2.835000 60.970000 ;
        RECT  2.635000 61.180000  2.835000 61.380000 ;
        RECT  2.635000 61.590000  2.835000 61.790000 ;
        RECT  2.635000 62.000000  2.835000 62.200000 ;
        RECT  2.635000 62.410000  2.835000 62.610000 ;
        RECT  3.045000 58.310000  3.245000 58.510000 ;
        RECT  3.045000 58.720000  3.245000 58.920000 ;
        RECT  3.045000 59.130000  3.245000 59.330000 ;
        RECT  3.045000 59.540000  3.245000 59.740000 ;
        RECT  3.045000 59.950000  3.245000 60.150000 ;
        RECT  3.045000 60.360000  3.245000 60.560000 ;
        RECT  3.045000 60.770000  3.245000 60.970000 ;
        RECT  3.045000 61.180000  3.245000 61.380000 ;
        RECT  3.045000 61.590000  3.245000 61.790000 ;
        RECT  3.045000 62.000000  3.245000 62.200000 ;
        RECT  3.045000 62.410000  3.245000 62.610000 ;
        RECT  3.450000 58.310000  3.650000 58.510000 ;
        RECT  3.450000 58.720000  3.650000 58.920000 ;
        RECT  3.450000 59.130000  3.650000 59.330000 ;
        RECT  3.450000 59.540000  3.650000 59.740000 ;
        RECT  3.450000 59.950000  3.650000 60.150000 ;
        RECT  3.450000 60.360000  3.650000 60.560000 ;
        RECT  3.450000 60.770000  3.650000 60.970000 ;
        RECT  3.450000 61.180000  3.650000 61.380000 ;
        RECT  3.450000 61.590000  3.650000 61.790000 ;
        RECT  3.450000 62.000000  3.650000 62.200000 ;
        RECT  3.450000 62.410000  3.650000 62.610000 ;
        RECT  3.855000 58.310000  4.055000 58.510000 ;
        RECT  3.855000 58.720000  4.055000 58.920000 ;
        RECT  3.855000 59.130000  4.055000 59.330000 ;
        RECT  3.855000 59.540000  4.055000 59.740000 ;
        RECT  3.855000 59.950000  4.055000 60.150000 ;
        RECT  3.855000 60.360000  4.055000 60.560000 ;
        RECT  3.855000 60.770000  4.055000 60.970000 ;
        RECT  3.855000 61.180000  4.055000 61.380000 ;
        RECT  3.855000 61.590000  4.055000 61.790000 ;
        RECT  3.855000 62.000000  4.055000 62.200000 ;
        RECT  3.855000 62.410000  4.055000 62.610000 ;
        RECT  4.260000 58.310000  4.460000 58.510000 ;
        RECT  4.260000 58.720000  4.460000 58.920000 ;
        RECT  4.260000 59.130000  4.460000 59.330000 ;
        RECT  4.260000 59.540000  4.460000 59.740000 ;
        RECT  4.260000 59.950000  4.460000 60.150000 ;
        RECT  4.260000 60.360000  4.460000 60.560000 ;
        RECT  4.260000 60.770000  4.460000 60.970000 ;
        RECT  4.260000 61.180000  4.460000 61.380000 ;
        RECT  4.260000 61.590000  4.460000 61.790000 ;
        RECT  4.260000 62.000000  4.460000 62.200000 ;
        RECT  4.260000 62.410000  4.460000 62.610000 ;
        RECT  4.665000 58.310000  4.865000 58.510000 ;
        RECT  4.665000 58.720000  4.865000 58.920000 ;
        RECT  4.665000 59.130000  4.865000 59.330000 ;
        RECT  4.665000 59.540000  4.865000 59.740000 ;
        RECT  4.665000 59.950000  4.865000 60.150000 ;
        RECT  4.665000 60.360000  4.865000 60.560000 ;
        RECT  4.665000 60.770000  4.865000 60.970000 ;
        RECT  4.665000 61.180000  4.865000 61.380000 ;
        RECT  4.665000 61.590000  4.865000 61.790000 ;
        RECT  4.665000 62.000000  4.865000 62.200000 ;
        RECT  4.665000 62.410000  4.865000 62.610000 ;
        RECT  5.070000 58.310000  5.270000 58.510000 ;
        RECT  5.070000 58.720000  5.270000 58.920000 ;
        RECT  5.070000 59.130000  5.270000 59.330000 ;
        RECT  5.070000 59.540000  5.270000 59.740000 ;
        RECT  5.070000 59.950000  5.270000 60.150000 ;
        RECT  5.070000 60.360000  5.270000 60.560000 ;
        RECT  5.070000 60.770000  5.270000 60.970000 ;
        RECT  5.070000 61.180000  5.270000 61.380000 ;
        RECT  5.070000 61.590000  5.270000 61.790000 ;
        RECT  5.070000 62.000000  5.270000 62.200000 ;
        RECT  5.070000 62.410000  5.270000 62.610000 ;
        RECT  5.475000 58.310000  5.675000 58.510000 ;
        RECT  5.475000 58.720000  5.675000 58.920000 ;
        RECT  5.475000 59.130000  5.675000 59.330000 ;
        RECT  5.475000 59.540000  5.675000 59.740000 ;
        RECT  5.475000 59.950000  5.675000 60.150000 ;
        RECT  5.475000 60.360000  5.675000 60.560000 ;
        RECT  5.475000 60.770000  5.675000 60.970000 ;
        RECT  5.475000 61.180000  5.675000 61.380000 ;
        RECT  5.475000 61.590000  5.675000 61.790000 ;
        RECT  5.475000 62.000000  5.675000 62.200000 ;
        RECT  5.475000 62.410000  5.675000 62.610000 ;
        RECT  5.880000 58.310000  6.080000 58.510000 ;
        RECT  5.880000 58.720000  6.080000 58.920000 ;
        RECT  5.880000 59.130000  6.080000 59.330000 ;
        RECT  5.880000 59.540000  6.080000 59.740000 ;
        RECT  5.880000 59.950000  6.080000 60.150000 ;
        RECT  5.880000 60.360000  6.080000 60.560000 ;
        RECT  5.880000 60.770000  6.080000 60.970000 ;
        RECT  5.880000 61.180000  6.080000 61.380000 ;
        RECT  5.880000 61.590000  6.080000 61.790000 ;
        RECT  5.880000 62.000000  6.080000 62.200000 ;
        RECT  5.880000 62.410000  6.080000 62.610000 ;
        RECT  6.285000 58.310000  6.485000 58.510000 ;
        RECT  6.285000 58.720000  6.485000 58.920000 ;
        RECT  6.285000 59.130000  6.485000 59.330000 ;
        RECT  6.285000 59.540000  6.485000 59.740000 ;
        RECT  6.285000 59.950000  6.485000 60.150000 ;
        RECT  6.285000 60.360000  6.485000 60.560000 ;
        RECT  6.285000 60.770000  6.485000 60.970000 ;
        RECT  6.285000 61.180000  6.485000 61.380000 ;
        RECT  6.285000 61.590000  6.485000 61.790000 ;
        RECT  6.285000 62.000000  6.485000 62.200000 ;
        RECT  6.285000 62.410000  6.485000 62.610000 ;
        RECT  6.690000 58.310000  6.890000 58.510000 ;
        RECT  6.690000 58.720000  6.890000 58.920000 ;
        RECT  6.690000 59.130000  6.890000 59.330000 ;
        RECT  6.690000 59.540000  6.890000 59.740000 ;
        RECT  6.690000 59.950000  6.890000 60.150000 ;
        RECT  6.690000 60.360000  6.890000 60.560000 ;
        RECT  6.690000 60.770000  6.890000 60.970000 ;
        RECT  6.690000 61.180000  6.890000 61.380000 ;
        RECT  6.690000 61.590000  6.890000 61.790000 ;
        RECT  6.690000 62.000000  6.890000 62.200000 ;
        RECT  6.690000 62.410000  6.890000 62.610000 ;
        RECT  7.095000 58.310000  7.295000 58.510000 ;
        RECT  7.095000 58.720000  7.295000 58.920000 ;
        RECT  7.095000 59.130000  7.295000 59.330000 ;
        RECT  7.095000 59.540000  7.295000 59.740000 ;
        RECT  7.095000 59.950000  7.295000 60.150000 ;
        RECT  7.095000 60.360000  7.295000 60.560000 ;
        RECT  7.095000 60.770000  7.295000 60.970000 ;
        RECT  7.095000 61.180000  7.295000 61.380000 ;
        RECT  7.095000 61.590000  7.295000 61.790000 ;
        RECT  7.095000 62.000000  7.295000 62.200000 ;
        RECT  7.095000 62.410000  7.295000 62.610000 ;
        RECT  7.500000 58.310000  7.700000 58.510000 ;
        RECT  7.500000 58.720000  7.700000 58.920000 ;
        RECT  7.500000 59.130000  7.700000 59.330000 ;
        RECT  7.500000 59.540000  7.700000 59.740000 ;
        RECT  7.500000 59.950000  7.700000 60.150000 ;
        RECT  7.500000 60.360000  7.700000 60.560000 ;
        RECT  7.500000 60.770000  7.700000 60.970000 ;
        RECT  7.500000 61.180000  7.700000 61.380000 ;
        RECT  7.500000 61.590000  7.700000 61.790000 ;
        RECT  7.500000 62.000000  7.700000 62.200000 ;
        RECT  7.500000 62.410000  7.700000 62.610000 ;
        RECT  7.905000 58.310000  8.105000 58.510000 ;
        RECT  7.905000 58.720000  8.105000 58.920000 ;
        RECT  7.905000 59.130000  8.105000 59.330000 ;
        RECT  7.905000 59.540000  8.105000 59.740000 ;
        RECT  7.905000 59.950000  8.105000 60.150000 ;
        RECT  7.905000 60.360000  8.105000 60.560000 ;
        RECT  7.905000 60.770000  8.105000 60.970000 ;
        RECT  7.905000 61.180000  8.105000 61.380000 ;
        RECT  7.905000 61.590000  8.105000 61.790000 ;
        RECT  7.905000 62.000000  8.105000 62.200000 ;
        RECT  7.905000 62.410000  8.105000 62.610000 ;
        RECT  8.310000 58.310000  8.510000 58.510000 ;
        RECT  8.310000 58.720000  8.510000 58.920000 ;
        RECT  8.310000 59.130000  8.510000 59.330000 ;
        RECT  8.310000 59.540000  8.510000 59.740000 ;
        RECT  8.310000 59.950000  8.510000 60.150000 ;
        RECT  8.310000 60.360000  8.510000 60.560000 ;
        RECT  8.310000 60.770000  8.510000 60.970000 ;
        RECT  8.310000 61.180000  8.510000 61.380000 ;
        RECT  8.310000 61.590000  8.510000 61.790000 ;
        RECT  8.310000 62.000000  8.510000 62.200000 ;
        RECT  8.310000 62.410000  8.510000 62.610000 ;
        RECT  8.715000 58.310000  8.915000 58.510000 ;
        RECT  8.715000 58.720000  8.915000 58.920000 ;
        RECT  8.715000 59.130000  8.915000 59.330000 ;
        RECT  8.715000 59.540000  8.915000 59.740000 ;
        RECT  8.715000 59.950000  8.915000 60.150000 ;
        RECT  8.715000 60.360000  8.915000 60.560000 ;
        RECT  8.715000 60.770000  8.915000 60.970000 ;
        RECT  8.715000 61.180000  8.915000 61.380000 ;
        RECT  8.715000 61.590000  8.915000 61.790000 ;
        RECT  8.715000 62.000000  8.915000 62.200000 ;
        RECT  8.715000 62.410000  8.915000 62.610000 ;
        RECT  9.120000 58.310000  9.320000 58.510000 ;
        RECT  9.120000 58.720000  9.320000 58.920000 ;
        RECT  9.120000 59.130000  9.320000 59.330000 ;
        RECT  9.120000 59.540000  9.320000 59.740000 ;
        RECT  9.120000 59.950000  9.320000 60.150000 ;
        RECT  9.120000 60.360000  9.320000 60.560000 ;
        RECT  9.120000 60.770000  9.320000 60.970000 ;
        RECT  9.120000 61.180000  9.320000 61.380000 ;
        RECT  9.120000 61.590000  9.320000 61.790000 ;
        RECT  9.120000 62.000000  9.320000 62.200000 ;
        RECT  9.120000 62.410000  9.320000 62.610000 ;
        RECT  9.525000 58.310000  9.725000 58.510000 ;
        RECT  9.525000 58.720000  9.725000 58.920000 ;
        RECT  9.525000 59.130000  9.725000 59.330000 ;
        RECT  9.525000 59.540000  9.725000 59.740000 ;
        RECT  9.525000 59.950000  9.725000 60.150000 ;
        RECT  9.525000 60.360000  9.725000 60.560000 ;
        RECT  9.525000 60.770000  9.725000 60.970000 ;
        RECT  9.525000 61.180000  9.725000 61.380000 ;
        RECT  9.525000 61.590000  9.725000 61.790000 ;
        RECT  9.525000 62.000000  9.725000 62.200000 ;
        RECT  9.525000 62.410000  9.725000 62.610000 ;
        RECT  9.930000 58.310000 10.130000 58.510000 ;
        RECT  9.930000 58.720000 10.130000 58.920000 ;
        RECT  9.930000 59.130000 10.130000 59.330000 ;
        RECT  9.930000 59.540000 10.130000 59.740000 ;
        RECT  9.930000 59.950000 10.130000 60.150000 ;
        RECT  9.930000 60.360000 10.130000 60.560000 ;
        RECT  9.930000 60.770000 10.130000 60.970000 ;
        RECT  9.930000 61.180000 10.130000 61.380000 ;
        RECT  9.930000 61.590000 10.130000 61.790000 ;
        RECT  9.930000 62.000000 10.130000 62.200000 ;
        RECT  9.930000 62.410000 10.130000 62.610000 ;
        RECT 10.335000 58.310000 10.535000 58.510000 ;
        RECT 10.335000 58.720000 10.535000 58.920000 ;
        RECT 10.335000 59.130000 10.535000 59.330000 ;
        RECT 10.335000 59.540000 10.535000 59.740000 ;
        RECT 10.335000 59.950000 10.535000 60.150000 ;
        RECT 10.335000 60.360000 10.535000 60.560000 ;
        RECT 10.335000 60.770000 10.535000 60.970000 ;
        RECT 10.335000 61.180000 10.535000 61.380000 ;
        RECT 10.335000 61.590000 10.535000 61.790000 ;
        RECT 10.335000 62.000000 10.535000 62.200000 ;
        RECT 10.335000 62.410000 10.535000 62.610000 ;
        RECT 10.740000 58.310000 10.940000 58.510000 ;
        RECT 10.740000 58.720000 10.940000 58.920000 ;
        RECT 10.740000 59.130000 10.940000 59.330000 ;
        RECT 10.740000 59.540000 10.940000 59.740000 ;
        RECT 10.740000 59.950000 10.940000 60.150000 ;
        RECT 10.740000 60.360000 10.940000 60.560000 ;
        RECT 10.740000 60.770000 10.940000 60.970000 ;
        RECT 10.740000 61.180000 10.940000 61.380000 ;
        RECT 10.740000 61.590000 10.940000 61.790000 ;
        RECT 10.740000 62.000000 10.940000 62.200000 ;
        RECT 10.740000 62.410000 10.940000 62.610000 ;
        RECT 11.145000 58.310000 11.345000 58.510000 ;
        RECT 11.145000 58.720000 11.345000 58.920000 ;
        RECT 11.145000 59.130000 11.345000 59.330000 ;
        RECT 11.145000 59.540000 11.345000 59.740000 ;
        RECT 11.145000 59.950000 11.345000 60.150000 ;
        RECT 11.145000 60.360000 11.345000 60.560000 ;
        RECT 11.145000 60.770000 11.345000 60.970000 ;
        RECT 11.145000 61.180000 11.345000 61.380000 ;
        RECT 11.145000 61.590000 11.345000 61.790000 ;
        RECT 11.145000 62.000000 11.345000 62.200000 ;
        RECT 11.145000 62.410000 11.345000 62.610000 ;
        RECT 11.550000 58.310000 11.750000 58.510000 ;
        RECT 11.550000 58.720000 11.750000 58.920000 ;
        RECT 11.550000 59.130000 11.750000 59.330000 ;
        RECT 11.550000 59.540000 11.750000 59.740000 ;
        RECT 11.550000 59.950000 11.750000 60.150000 ;
        RECT 11.550000 60.360000 11.750000 60.560000 ;
        RECT 11.550000 60.770000 11.750000 60.970000 ;
        RECT 11.550000 61.180000 11.750000 61.380000 ;
        RECT 11.550000 61.590000 11.750000 61.790000 ;
        RECT 11.550000 62.000000 11.750000 62.200000 ;
        RECT 11.550000 62.410000 11.750000 62.610000 ;
        RECT 11.955000 58.310000 12.155000 58.510000 ;
        RECT 11.955000 58.720000 12.155000 58.920000 ;
        RECT 11.955000 59.130000 12.155000 59.330000 ;
        RECT 11.955000 59.540000 12.155000 59.740000 ;
        RECT 11.955000 59.950000 12.155000 60.150000 ;
        RECT 11.955000 60.360000 12.155000 60.560000 ;
        RECT 11.955000 60.770000 12.155000 60.970000 ;
        RECT 11.955000 61.180000 12.155000 61.380000 ;
        RECT 11.955000 61.590000 12.155000 61.790000 ;
        RECT 11.955000 62.000000 12.155000 62.200000 ;
        RECT 11.955000 62.410000 12.155000 62.610000 ;
        RECT 12.360000 58.310000 12.560000 58.510000 ;
        RECT 12.360000 58.720000 12.560000 58.920000 ;
        RECT 12.360000 59.130000 12.560000 59.330000 ;
        RECT 12.360000 59.540000 12.560000 59.740000 ;
        RECT 12.360000 59.950000 12.560000 60.150000 ;
        RECT 12.360000 60.360000 12.560000 60.560000 ;
        RECT 12.360000 60.770000 12.560000 60.970000 ;
        RECT 12.360000 61.180000 12.560000 61.380000 ;
        RECT 12.360000 61.590000 12.560000 61.790000 ;
        RECT 12.360000 62.000000 12.560000 62.200000 ;
        RECT 12.360000 62.410000 12.560000 62.610000 ;
        RECT 12.765000 58.310000 12.965000 58.510000 ;
        RECT 12.765000 58.720000 12.965000 58.920000 ;
        RECT 12.765000 59.130000 12.965000 59.330000 ;
        RECT 12.765000 59.540000 12.965000 59.740000 ;
        RECT 12.765000 59.950000 12.965000 60.150000 ;
        RECT 12.765000 60.360000 12.965000 60.560000 ;
        RECT 12.765000 60.770000 12.965000 60.970000 ;
        RECT 12.765000 61.180000 12.965000 61.380000 ;
        RECT 12.765000 61.590000 12.965000 61.790000 ;
        RECT 12.765000 62.000000 12.965000 62.200000 ;
        RECT 12.765000 62.410000 12.965000 62.610000 ;
        RECT 13.170000 58.310000 13.370000 58.510000 ;
        RECT 13.170000 58.720000 13.370000 58.920000 ;
        RECT 13.170000 59.130000 13.370000 59.330000 ;
        RECT 13.170000 59.540000 13.370000 59.740000 ;
        RECT 13.170000 59.950000 13.370000 60.150000 ;
        RECT 13.170000 60.360000 13.370000 60.560000 ;
        RECT 13.170000 60.770000 13.370000 60.970000 ;
        RECT 13.170000 61.180000 13.370000 61.380000 ;
        RECT 13.170000 61.590000 13.370000 61.790000 ;
        RECT 13.170000 62.000000 13.370000 62.200000 ;
        RECT 13.170000 62.410000 13.370000 62.610000 ;
        RECT 13.575000 58.310000 13.775000 58.510000 ;
        RECT 13.575000 58.720000 13.775000 58.920000 ;
        RECT 13.575000 59.130000 13.775000 59.330000 ;
        RECT 13.575000 59.540000 13.775000 59.740000 ;
        RECT 13.575000 59.950000 13.775000 60.150000 ;
        RECT 13.575000 60.360000 13.775000 60.560000 ;
        RECT 13.575000 60.770000 13.775000 60.970000 ;
        RECT 13.575000 61.180000 13.775000 61.380000 ;
        RECT 13.575000 61.590000 13.775000 61.790000 ;
        RECT 13.575000 62.000000 13.775000 62.200000 ;
        RECT 13.575000 62.410000 13.775000 62.610000 ;
        RECT 13.980000 58.310000 14.180000 58.510000 ;
        RECT 13.980000 58.720000 14.180000 58.920000 ;
        RECT 13.980000 59.130000 14.180000 59.330000 ;
        RECT 13.980000 59.540000 14.180000 59.740000 ;
        RECT 13.980000 59.950000 14.180000 60.150000 ;
        RECT 13.980000 60.360000 14.180000 60.560000 ;
        RECT 13.980000 60.770000 14.180000 60.970000 ;
        RECT 13.980000 61.180000 14.180000 61.380000 ;
        RECT 13.980000 61.590000 14.180000 61.790000 ;
        RECT 13.980000 62.000000 14.180000 62.200000 ;
        RECT 13.980000 62.410000 14.180000 62.610000 ;
        RECT 14.385000 58.310000 14.585000 58.510000 ;
        RECT 14.385000 58.720000 14.585000 58.920000 ;
        RECT 14.385000 59.130000 14.585000 59.330000 ;
        RECT 14.385000 59.540000 14.585000 59.740000 ;
        RECT 14.385000 59.950000 14.585000 60.150000 ;
        RECT 14.385000 60.360000 14.585000 60.560000 ;
        RECT 14.385000 60.770000 14.585000 60.970000 ;
        RECT 14.385000 61.180000 14.585000 61.380000 ;
        RECT 14.385000 61.590000 14.585000 61.790000 ;
        RECT 14.385000 62.000000 14.585000 62.200000 ;
        RECT 14.385000 62.410000 14.585000 62.610000 ;
        RECT 14.790000 58.310000 14.990000 58.510000 ;
        RECT 14.790000 58.720000 14.990000 58.920000 ;
        RECT 14.790000 59.130000 14.990000 59.330000 ;
        RECT 14.790000 59.540000 14.990000 59.740000 ;
        RECT 14.790000 59.950000 14.990000 60.150000 ;
        RECT 14.790000 60.360000 14.990000 60.560000 ;
        RECT 14.790000 60.770000 14.990000 60.970000 ;
        RECT 14.790000 61.180000 14.990000 61.380000 ;
        RECT 14.790000 61.590000 14.990000 61.790000 ;
        RECT 14.790000 62.000000 14.990000 62.200000 ;
        RECT 14.790000 62.410000 14.990000 62.610000 ;
        RECT 15.195000 58.310000 15.395000 58.510000 ;
        RECT 15.195000 58.720000 15.395000 58.920000 ;
        RECT 15.195000 59.130000 15.395000 59.330000 ;
        RECT 15.195000 59.540000 15.395000 59.740000 ;
        RECT 15.195000 59.950000 15.395000 60.150000 ;
        RECT 15.195000 60.360000 15.395000 60.560000 ;
        RECT 15.195000 60.770000 15.395000 60.970000 ;
        RECT 15.195000 61.180000 15.395000 61.380000 ;
        RECT 15.195000 61.590000 15.395000 61.790000 ;
        RECT 15.195000 62.000000 15.395000 62.200000 ;
        RECT 15.195000 62.410000 15.395000 62.610000 ;
        RECT 15.600000 58.310000 15.800000 58.510000 ;
        RECT 15.600000 58.720000 15.800000 58.920000 ;
        RECT 15.600000 59.130000 15.800000 59.330000 ;
        RECT 15.600000 59.540000 15.800000 59.740000 ;
        RECT 15.600000 59.950000 15.800000 60.150000 ;
        RECT 15.600000 60.360000 15.800000 60.560000 ;
        RECT 15.600000 60.770000 15.800000 60.970000 ;
        RECT 15.600000 61.180000 15.800000 61.380000 ;
        RECT 15.600000 61.590000 15.800000 61.790000 ;
        RECT 15.600000 62.000000 15.800000 62.200000 ;
        RECT 15.600000 62.410000 15.800000 62.610000 ;
        RECT 16.005000 58.310000 16.205000 58.510000 ;
        RECT 16.005000 58.720000 16.205000 58.920000 ;
        RECT 16.005000 59.130000 16.205000 59.330000 ;
        RECT 16.005000 59.540000 16.205000 59.740000 ;
        RECT 16.005000 59.950000 16.205000 60.150000 ;
        RECT 16.005000 60.360000 16.205000 60.560000 ;
        RECT 16.005000 60.770000 16.205000 60.970000 ;
        RECT 16.005000 61.180000 16.205000 61.380000 ;
        RECT 16.005000 61.590000 16.205000 61.790000 ;
        RECT 16.005000 62.000000 16.205000 62.200000 ;
        RECT 16.005000 62.410000 16.205000 62.610000 ;
        RECT 16.410000 58.310000 16.610000 58.510000 ;
        RECT 16.410000 58.720000 16.610000 58.920000 ;
        RECT 16.410000 59.130000 16.610000 59.330000 ;
        RECT 16.410000 59.540000 16.610000 59.740000 ;
        RECT 16.410000 59.950000 16.610000 60.150000 ;
        RECT 16.410000 60.360000 16.610000 60.560000 ;
        RECT 16.410000 60.770000 16.610000 60.970000 ;
        RECT 16.410000 61.180000 16.610000 61.380000 ;
        RECT 16.410000 61.590000 16.610000 61.790000 ;
        RECT 16.410000 62.000000 16.610000 62.200000 ;
        RECT 16.410000 62.410000 16.610000 62.610000 ;
        RECT 16.815000 58.310000 17.015000 58.510000 ;
        RECT 16.815000 58.720000 17.015000 58.920000 ;
        RECT 16.815000 59.130000 17.015000 59.330000 ;
        RECT 16.815000 59.540000 17.015000 59.740000 ;
        RECT 16.815000 59.950000 17.015000 60.150000 ;
        RECT 16.815000 60.360000 17.015000 60.560000 ;
        RECT 16.815000 60.770000 17.015000 60.970000 ;
        RECT 16.815000 61.180000 17.015000 61.380000 ;
        RECT 16.815000 61.590000 17.015000 61.790000 ;
        RECT 16.815000 62.000000 17.015000 62.200000 ;
        RECT 16.815000 62.410000 17.015000 62.610000 ;
        RECT 17.220000 58.310000 17.420000 58.510000 ;
        RECT 17.220000 58.720000 17.420000 58.920000 ;
        RECT 17.220000 59.130000 17.420000 59.330000 ;
        RECT 17.220000 59.540000 17.420000 59.740000 ;
        RECT 17.220000 59.950000 17.420000 60.150000 ;
        RECT 17.220000 60.360000 17.420000 60.560000 ;
        RECT 17.220000 60.770000 17.420000 60.970000 ;
        RECT 17.220000 61.180000 17.420000 61.380000 ;
        RECT 17.220000 61.590000 17.420000 61.790000 ;
        RECT 17.220000 62.000000 17.420000 62.200000 ;
        RECT 17.220000 62.410000 17.420000 62.610000 ;
        RECT 17.625000 58.310000 17.825000 58.510000 ;
        RECT 17.625000 58.720000 17.825000 58.920000 ;
        RECT 17.625000 59.130000 17.825000 59.330000 ;
        RECT 17.625000 59.540000 17.825000 59.740000 ;
        RECT 17.625000 59.950000 17.825000 60.150000 ;
        RECT 17.625000 60.360000 17.825000 60.560000 ;
        RECT 17.625000 60.770000 17.825000 60.970000 ;
        RECT 17.625000 61.180000 17.825000 61.380000 ;
        RECT 17.625000 61.590000 17.825000 61.790000 ;
        RECT 17.625000 62.000000 17.825000 62.200000 ;
        RECT 17.625000 62.410000 17.825000 62.610000 ;
        RECT 18.030000 58.310000 18.230000 58.510000 ;
        RECT 18.030000 58.720000 18.230000 58.920000 ;
        RECT 18.030000 59.130000 18.230000 59.330000 ;
        RECT 18.030000 59.540000 18.230000 59.740000 ;
        RECT 18.030000 59.950000 18.230000 60.150000 ;
        RECT 18.030000 60.360000 18.230000 60.560000 ;
        RECT 18.030000 60.770000 18.230000 60.970000 ;
        RECT 18.030000 61.180000 18.230000 61.380000 ;
        RECT 18.030000 61.590000 18.230000 61.790000 ;
        RECT 18.030000 62.000000 18.230000 62.200000 ;
        RECT 18.030000 62.410000 18.230000 62.610000 ;
        RECT 18.435000 58.310000 18.635000 58.510000 ;
        RECT 18.435000 58.720000 18.635000 58.920000 ;
        RECT 18.435000 59.130000 18.635000 59.330000 ;
        RECT 18.435000 59.540000 18.635000 59.740000 ;
        RECT 18.435000 59.950000 18.635000 60.150000 ;
        RECT 18.435000 60.360000 18.635000 60.560000 ;
        RECT 18.435000 60.770000 18.635000 60.970000 ;
        RECT 18.435000 61.180000 18.635000 61.380000 ;
        RECT 18.435000 61.590000 18.635000 61.790000 ;
        RECT 18.435000 62.000000 18.635000 62.200000 ;
        RECT 18.435000 62.410000 18.635000 62.610000 ;
        RECT 18.840000 58.310000 19.040000 58.510000 ;
        RECT 18.840000 58.720000 19.040000 58.920000 ;
        RECT 18.840000 59.130000 19.040000 59.330000 ;
        RECT 18.840000 59.540000 19.040000 59.740000 ;
        RECT 18.840000 59.950000 19.040000 60.150000 ;
        RECT 18.840000 60.360000 19.040000 60.560000 ;
        RECT 18.840000 60.770000 19.040000 60.970000 ;
        RECT 18.840000 61.180000 19.040000 61.380000 ;
        RECT 18.840000 61.590000 19.040000 61.790000 ;
        RECT 18.840000 62.000000 19.040000 62.200000 ;
        RECT 18.840000 62.410000 19.040000 62.610000 ;
        RECT 19.245000 58.310000 19.445000 58.510000 ;
        RECT 19.245000 58.720000 19.445000 58.920000 ;
        RECT 19.245000 59.130000 19.445000 59.330000 ;
        RECT 19.245000 59.540000 19.445000 59.740000 ;
        RECT 19.245000 59.950000 19.445000 60.150000 ;
        RECT 19.245000 60.360000 19.445000 60.560000 ;
        RECT 19.245000 60.770000 19.445000 60.970000 ;
        RECT 19.245000 61.180000 19.445000 61.380000 ;
        RECT 19.245000 61.590000 19.445000 61.790000 ;
        RECT 19.245000 62.000000 19.445000 62.200000 ;
        RECT 19.245000 62.410000 19.445000 62.610000 ;
        RECT 19.650000 58.310000 19.850000 58.510000 ;
        RECT 19.650000 58.720000 19.850000 58.920000 ;
        RECT 19.650000 59.130000 19.850000 59.330000 ;
        RECT 19.650000 59.540000 19.850000 59.740000 ;
        RECT 19.650000 59.950000 19.850000 60.150000 ;
        RECT 19.650000 60.360000 19.850000 60.560000 ;
        RECT 19.650000 60.770000 19.850000 60.970000 ;
        RECT 19.650000 61.180000 19.850000 61.380000 ;
        RECT 19.650000 61.590000 19.850000 61.790000 ;
        RECT 19.650000 62.000000 19.850000 62.200000 ;
        RECT 19.650000 62.410000 19.850000 62.610000 ;
        RECT 20.055000 58.310000 20.255000 58.510000 ;
        RECT 20.055000 58.720000 20.255000 58.920000 ;
        RECT 20.055000 59.130000 20.255000 59.330000 ;
        RECT 20.055000 59.540000 20.255000 59.740000 ;
        RECT 20.055000 59.950000 20.255000 60.150000 ;
        RECT 20.055000 60.360000 20.255000 60.560000 ;
        RECT 20.055000 60.770000 20.255000 60.970000 ;
        RECT 20.055000 61.180000 20.255000 61.380000 ;
        RECT 20.055000 61.590000 20.255000 61.790000 ;
        RECT 20.055000 62.000000 20.255000 62.200000 ;
        RECT 20.055000 62.410000 20.255000 62.610000 ;
        RECT 20.460000 58.310000 20.660000 58.510000 ;
        RECT 20.460000 58.720000 20.660000 58.920000 ;
        RECT 20.460000 59.130000 20.660000 59.330000 ;
        RECT 20.460000 59.540000 20.660000 59.740000 ;
        RECT 20.460000 59.950000 20.660000 60.150000 ;
        RECT 20.460000 60.360000 20.660000 60.560000 ;
        RECT 20.460000 60.770000 20.660000 60.970000 ;
        RECT 20.460000 61.180000 20.660000 61.380000 ;
        RECT 20.460000 61.590000 20.660000 61.790000 ;
        RECT 20.460000 62.000000 20.660000 62.200000 ;
        RECT 20.460000 62.410000 20.660000 62.610000 ;
        RECT 20.865000 58.310000 21.065000 58.510000 ;
        RECT 20.865000 58.720000 21.065000 58.920000 ;
        RECT 20.865000 59.130000 21.065000 59.330000 ;
        RECT 20.865000 59.540000 21.065000 59.740000 ;
        RECT 20.865000 59.950000 21.065000 60.150000 ;
        RECT 20.865000 60.360000 21.065000 60.560000 ;
        RECT 20.865000 60.770000 21.065000 60.970000 ;
        RECT 20.865000 61.180000 21.065000 61.380000 ;
        RECT 20.865000 61.590000 21.065000 61.790000 ;
        RECT 20.865000 62.000000 21.065000 62.200000 ;
        RECT 20.865000 62.410000 21.065000 62.610000 ;
        RECT 21.270000 58.310000 21.470000 58.510000 ;
        RECT 21.270000 58.720000 21.470000 58.920000 ;
        RECT 21.270000 59.130000 21.470000 59.330000 ;
        RECT 21.270000 59.540000 21.470000 59.740000 ;
        RECT 21.270000 59.950000 21.470000 60.150000 ;
        RECT 21.270000 60.360000 21.470000 60.560000 ;
        RECT 21.270000 60.770000 21.470000 60.970000 ;
        RECT 21.270000 61.180000 21.470000 61.380000 ;
        RECT 21.270000 61.590000 21.470000 61.790000 ;
        RECT 21.270000 62.000000 21.470000 62.200000 ;
        RECT 21.270000 62.410000 21.470000 62.610000 ;
        RECT 21.675000 58.310000 21.875000 58.510000 ;
        RECT 21.675000 58.720000 21.875000 58.920000 ;
        RECT 21.675000 59.130000 21.875000 59.330000 ;
        RECT 21.675000 59.540000 21.875000 59.740000 ;
        RECT 21.675000 59.950000 21.875000 60.150000 ;
        RECT 21.675000 60.360000 21.875000 60.560000 ;
        RECT 21.675000 60.770000 21.875000 60.970000 ;
        RECT 21.675000 61.180000 21.875000 61.380000 ;
        RECT 21.675000 61.590000 21.875000 61.790000 ;
        RECT 21.675000 62.000000 21.875000 62.200000 ;
        RECT 21.675000 62.410000 21.875000 62.610000 ;
        RECT 22.080000 58.310000 22.280000 58.510000 ;
        RECT 22.080000 58.720000 22.280000 58.920000 ;
        RECT 22.080000 59.130000 22.280000 59.330000 ;
        RECT 22.080000 59.540000 22.280000 59.740000 ;
        RECT 22.080000 59.950000 22.280000 60.150000 ;
        RECT 22.080000 60.360000 22.280000 60.560000 ;
        RECT 22.080000 60.770000 22.280000 60.970000 ;
        RECT 22.080000 61.180000 22.280000 61.380000 ;
        RECT 22.080000 61.590000 22.280000 61.790000 ;
        RECT 22.080000 62.000000 22.280000 62.200000 ;
        RECT 22.080000 62.410000 22.280000 62.610000 ;
        RECT 22.485000 58.310000 22.685000 58.510000 ;
        RECT 22.485000 58.720000 22.685000 58.920000 ;
        RECT 22.485000 59.130000 22.685000 59.330000 ;
        RECT 22.485000 59.540000 22.685000 59.740000 ;
        RECT 22.485000 59.950000 22.685000 60.150000 ;
        RECT 22.485000 60.360000 22.685000 60.560000 ;
        RECT 22.485000 60.770000 22.685000 60.970000 ;
        RECT 22.485000 61.180000 22.685000 61.380000 ;
        RECT 22.485000 61.590000 22.685000 61.790000 ;
        RECT 22.485000 62.000000 22.685000 62.200000 ;
        RECT 22.485000 62.410000 22.685000 62.610000 ;
        RECT 22.890000 58.310000 23.090000 58.510000 ;
        RECT 22.890000 58.720000 23.090000 58.920000 ;
        RECT 22.890000 59.130000 23.090000 59.330000 ;
        RECT 22.890000 59.540000 23.090000 59.740000 ;
        RECT 22.890000 59.950000 23.090000 60.150000 ;
        RECT 22.890000 60.360000 23.090000 60.560000 ;
        RECT 22.890000 60.770000 23.090000 60.970000 ;
        RECT 22.890000 61.180000 23.090000 61.380000 ;
        RECT 22.890000 61.590000 23.090000 61.790000 ;
        RECT 22.890000 62.000000 23.090000 62.200000 ;
        RECT 22.890000 62.410000 23.090000 62.610000 ;
        RECT 23.295000 58.310000 23.495000 58.510000 ;
        RECT 23.295000 58.720000 23.495000 58.920000 ;
        RECT 23.295000 59.130000 23.495000 59.330000 ;
        RECT 23.295000 59.540000 23.495000 59.740000 ;
        RECT 23.295000 59.950000 23.495000 60.150000 ;
        RECT 23.295000 60.360000 23.495000 60.560000 ;
        RECT 23.295000 60.770000 23.495000 60.970000 ;
        RECT 23.295000 61.180000 23.495000 61.380000 ;
        RECT 23.295000 61.590000 23.495000 61.790000 ;
        RECT 23.295000 62.000000 23.495000 62.200000 ;
        RECT 23.295000 62.410000 23.495000 62.610000 ;
        RECT 23.700000 58.310000 23.900000 58.510000 ;
        RECT 23.700000 58.720000 23.900000 58.920000 ;
        RECT 23.700000 59.130000 23.900000 59.330000 ;
        RECT 23.700000 59.540000 23.900000 59.740000 ;
        RECT 23.700000 59.950000 23.900000 60.150000 ;
        RECT 23.700000 60.360000 23.900000 60.560000 ;
        RECT 23.700000 60.770000 23.900000 60.970000 ;
        RECT 23.700000 61.180000 23.900000 61.380000 ;
        RECT 23.700000 61.590000 23.900000 61.790000 ;
        RECT 23.700000 62.000000 23.900000 62.200000 ;
        RECT 23.700000 62.410000 23.900000 62.610000 ;
        RECT 24.105000 58.310000 24.305000 58.510000 ;
        RECT 24.105000 58.720000 24.305000 58.920000 ;
        RECT 24.105000 59.130000 24.305000 59.330000 ;
        RECT 24.105000 59.540000 24.305000 59.740000 ;
        RECT 24.105000 59.950000 24.305000 60.150000 ;
        RECT 24.105000 60.360000 24.305000 60.560000 ;
        RECT 24.105000 60.770000 24.305000 60.970000 ;
        RECT 24.105000 61.180000 24.305000 61.380000 ;
        RECT 24.105000 61.590000 24.305000 61.790000 ;
        RECT 24.105000 62.000000 24.305000 62.200000 ;
        RECT 24.105000 62.410000 24.305000 62.610000 ;
        RECT 50.480000 58.310000 50.680000 58.510000 ;
        RECT 50.480000 58.720000 50.680000 58.920000 ;
        RECT 50.480000 59.130000 50.680000 59.330000 ;
        RECT 50.480000 59.540000 50.680000 59.740000 ;
        RECT 50.480000 59.950000 50.680000 60.150000 ;
        RECT 50.480000 60.360000 50.680000 60.560000 ;
        RECT 50.480000 60.770000 50.680000 60.970000 ;
        RECT 50.480000 61.180000 50.680000 61.380000 ;
        RECT 50.480000 61.590000 50.680000 61.790000 ;
        RECT 50.480000 62.000000 50.680000 62.200000 ;
        RECT 50.480000 62.410000 50.680000 62.610000 ;
        RECT 50.890000 58.310000 51.090000 58.510000 ;
        RECT 50.890000 58.720000 51.090000 58.920000 ;
        RECT 50.890000 59.130000 51.090000 59.330000 ;
        RECT 50.890000 59.540000 51.090000 59.740000 ;
        RECT 50.890000 59.950000 51.090000 60.150000 ;
        RECT 50.890000 60.360000 51.090000 60.560000 ;
        RECT 50.890000 60.770000 51.090000 60.970000 ;
        RECT 50.890000 61.180000 51.090000 61.380000 ;
        RECT 50.890000 61.590000 51.090000 61.790000 ;
        RECT 50.890000 62.000000 51.090000 62.200000 ;
        RECT 50.890000 62.410000 51.090000 62.610000 ;
        RECT 51.300000 58.310000 51.500000 58.510000 ;
        RECT 51.300000 58.720000 51.500000 58.920000 ;
        RECT 51.300000 59.130000 51.500000 59.330000 ;
        RECT 51.300000 59.540000 51.500000 59.740000 ;
        RECT 51.300000 59.950000 51.500000 60.150000 ;
        RECT 51.300000 60.360000 51.500000 60.560000 ;
        RECT 51.300000 60.770000 51.500000 60.970000 ;
        RECT 51.300000 61.180000 51.500000 61.380000 ;
        RECT 51.300000 61.590000 51.500000 61.790000 ;
        RECT 51.300000 62.000000 51.500000 62.200000 ;
        RECT 51.300000 62.410000 51.500000 62.610000 ;
        RECT 51.710000 58.310000 51.910000 58.510000 ;
        RECT 51.710000 58.720000 51.910000 58.920000 ;
        RECT 51.710000 59.130000 51.910000 59.330000 ;
        RECT 51.710000 59.540000 51.910000 59.740000 ;
        RECT 51.710000 59.950000 51.910000 60.150000 ;
        RECT 51.710000 60.360000 51.910000 60.560000 ;
        RECT 51.710000 60.770000 51.910000 60.970000 ;
        RECT 51.710000 61.180000 51.910000 61.380000 ;
        RECT 51.710000 61.590000 51.910000 61.790000 ;
        RECT 51.710000 62.000000 51.910000 62.200000 ;
        RECT 51.710000 62.410000 51.910000 62.610000 ;
        RECT 52.120000 58.310000 52.320000 58.510000 ;
        RECT 52.120000 58.720000 52.320000 58.920000 ;
        RECT 52.120000 59.130000 52.320000 59.330000 ;
        RECT 52.120000 59.540000 52.320000 59.740000 ;
        RECT 52.120000 59.950000 52.320000 60.150000 ;
        RECT 52.120000 60.360000 52.320000 60.560000 ;
        RECT 52.120000 60.770000 52.320000 60.970000 ;
        RECT 52.120000 61.180000 52.320000 61.380000 ;
        RECT 52.120000 61.590000 52.320000 61.790000 ;
        RECT 52.120000 62.000000 52.320000 62.200000 ;
        RECT 52.120000 62.410000 52.320000 62.610000 ;
        RECT 52.530000 58.310000 52.730000 58.510000 ;
        RECT 52.530000 58.720000 52.730000 58.920000 ;
        RECT 52.530000 59.130000 52.730000 59.330000 ;
        RECT 52.530000 59.540000 52.730000 59.740000 ;
        RECT 52.530000 59.950000 52.730000 60.150000 ;
        RECT 52.530000 60.360000 52.730000 60.560000 ;
        RECT 52.530000 60.770000 52.730000 60.970000 ;
        RECT 52.530000 61.180000 52.730000 61.380000 ;
        RECT 52.530000 61.590000 52.730000 61.790000 ;
        RECT 52.530000 62.000000 52.730000 62.200000 ;
        RECT 52.530000 62.410000 52.730000 62.610000 ;
        RECT 52.940000 58.310000 53.140000 58.510000 ;
        RECT 52.940000 58.720000 53.140000 58.920000 ;
        RECT 52.940000 59.130000 53.140000 59.330000 ;
        RECT 52.940000 59.540000 53.140000 59.740000 ;
        RECT 52.940000 59.950000 53.140000 60.150000 ;
        RECT 52.940000 60.360000 53.140000 60.560000 ;
        RECT 52.940000 60.770000 53.140000 60.970000 ;
        RECT 52.940000 61.180000 53.140000 61.380000 ;
        RECT 52.940000 61.590000 53.140000 61.790000 ;
        RECT 52.940000 62.000000 53.140000 62.200000 ;
        RECT 52.940000 62.410000 53.140000 62.610000 ;
        RECT 53.345000 58.310000 53.545000 58.510000 ;
        RECT 53.345000 58.720000 53.545000 58.920000 ;
        RECT 53.345000 59.130000 53.545000 59.330000 ;
        RECT 53.345000 59.540000 53.545000 59.740000 ;
        RECT 53.345000 59.950000 53.545000 60.150000 ;
        RECT 53.345000 60.360000 53.545000 60.560000 ;
        RECT 53.345000 60.770000 53.545000 60.970000 ;
        RECT 53.345000 61.180000 53.545000 61.380000 ;
        RECT 53.345000 61.590000 53.545000 61.790000 ;
        RECT 53.345000 62.000000 53.545000 62.200000 ;
        RECT 53.345000 62.410000 53.545000 62.610000 ;
        RECT 53.750000 58.310000 53.950000 58.510000 ;
        RECT 53.750000 58.720000 53.950000 58.920000 ;
        RECT 53.750000 59.130000 53.950000 59.330000 ;
        RECT 53.750000 59.540000 53.950000 59.740000 ;
        RECT 53.750000 59.950000 53.950000 60.150000 ;
        RECT 53.750000 60.360000 53.950000 60.560000 ;
        RECT 53.750000 60.770000 53.950000 60.970000 ;
        RECT 53.750000 61.180000 53.950000 61.380000 ;
        RECT 53.750000 61.590000 53.950000 61.790000 ;
        RECT 53.750000 62.000000 53.950000 62.200000 ;
        RECT 53.750000 62.410000 53.950000 62.610000 ;
        RECT 54.155000 58.310000 54.355000 58.510000 ;
        RECT 54.155000 58.720000 54.355000 58.920000 ;
        RECT 54.155000 59.130000 54.355000 59.330000 ;
        RECT 54.155000 59.540000 54.355000 59.740000 ;
        RECT 54.155000 59.950000 54.355000 60.150000 ;
        RECT 54.155000 60.360000 54.355000 60.560000 ;
        RECT 54.155000 60.770000 54.355000 60.970000 ;
        RECT 54.155000 61.180000 54.355000 61.380000 ;
        RECT 54.155000 61.590000 54.355000 61.790000 ;
        RECT 54.155000 62.000000 54.355000 62.200000 ;
        RECT 54.155000 62.410000 54.355000 62.610000 ;
        RECT 54.560000 58.310000 54.760000 58.510000 ;
        RECT 54.560000 58.720000 54.760000 58.920000 ;
        RECT 54.560000 59.130000 54.760000 59.330000 ;
        RECT 54.560000 59.540000 54.760000 59.740000 ;
        RECT 54.560000 59.950000 54.760000 60.150000 ;
        RECT 54.560000 60.360000 54.760000 60.560000 ;
        RECT 54.560000 60.770000 54.760000 60.970000 ;
        RECT 54.560000 61.180000 54.760000 61.380000 ;
        RECT 54.560000 61.590000 54.760000 61.790000 ;
        RECT 54.560000 62.000000 54.760000 62.200000 ;
        RECT 54.560000 62.410000 54.760000 62.610000 ;
        RECT 54.965000 58.310000 55.165000 58.510000 ;
        RECT 54.965000 58.720000 55.165000 58.920000 ;
        RECT 54.965000 59.130000 55.165000 59.330000 ;
        RECT 54.965000 59.540000 55.165000 59.740000 ;
        RECT 54.965000 59.950000 55.165000 60.150000 ;
        RECT 54.965000 60.360000 55.165000 60.560000 ;
        RECT 54.965000 60.770000 55.165000 60.970000 ;
        RECT 54.965000 61.180000 55.165000 61.380000 ;
        RECT 54.965000 61.590000 55.165000 61.790000 ;
        RECT 54.965000 62.000000 55.165000 62.200000 ;
        RECT 54.965000 62.410000 55.165000 62.610000 ;
        RECT 55.370000 58.310000 55.570000 58.510000 ;
        RECT 55.370000 58.720000 55.570000 58.920000 ;
        RECT 55.370000 59.130000 55.570000 59.330000 ;
        RECT 55.370000 59.540000 55.570000 59.740000 ;
        RECT 55.370000 59.950000 55.570000 60.150000 ;
        RECT 55.370000 60.360000 55.570000 60.560000 ;
        RECT 55.370000 60.770000 55.570000 60.970000 ;
        RECT 55.370000 61.180000 55.570000 61.380000 ;
        RECT 55.370000 61.590000 55.570000 61.790000 ;
        RECT 55.370000 62.000000 55.570000 62.200000 ;
        RECT 55.370000 62.410000 55.570000 62.610000 ;
        RECT 55.775000 58.310000 55.975000 58.510000 ;
        RECT 55.775000 58.720000 55.975000 58.920000 ;
        RECT 55.775000 59.130000 55.975000 59.330000 ;
        RECT 55.775000 59.540000 55.975000 59.740000 ;
        RECT 55.775000 59.950000 55.975000 60.150000 ;
        RECT 55.775000 60.360000 55.975000 60.560000 ;
        RECT 55.775000 60.770000 55.975000 60.970000 ;
        RECT 55.775000 61.180000 55.975000 61.380000 ;
        RECT 55.775000 61.590000 55.975000 61.790000 ;
        RECT 55.775000 62.000000 55.975000 62.200000 ;
        RECT 55.775000 62.410000 55.975000 62.610000 ;
        RECT 56.180000 58.310000 56.380000 58.510000 ;
        RECT 56.180000 58.720000 56.380000 58.920000 ;
        RECT 56.180000 59.130000 56.380000 59.330000 ;
        RECT 56.180000 59.540000 56.380000 59.740000 ;
        RECT 56.180000 59.950000 56.380000 60.150000 ;
        RECT 56.180000 60.360000 56.380000 60.560000 ;
        RECT 56.180000 60.770000 56.380000 60.970000 ;
        RECT 56.180000 61.180000 56.380000 61.380000 ;
        RECT 56.180000 61.590000 56.380000 61.790000 ;
        RECT 56.180000 62.000000 56.380000 62.200000 ;
        RECT 56.180000 62.410000 56.380000 62.610000 ;
        RECT 56.585000 58.310000 56.785000 58.510000 ;
        RECT 56.585000 58.720000 56.785000 58.920000 ;
        RECT 56.585000 59.130000 56.785000 59.330000 ;
        RECT 56.585000 59.540000 56.785000 59.740000 ;
        RECT 56.585000 59.950000 56.785000 60.150000 ;
        RECT 56.585000 60.360000 56.785000 60.560000 ;
        RECT 56.585000 60.770000 56.785000 60.970000 ;
        RECT 56.585000 61.180000 56.785000 61.380000 ;
        RECT 56.585000 61.590000 56.785000 61.790000 ;
        RECT 56.585000 62.000000 56.785000 62.200000 ;
        RECT 56.585000 62.410000 56.785000 62.610000 ;
        RECT 56.990000 58.310000 57.190000 58.510000 ;
        RECT 56.990000 58.720000 57.190000 58.920000 ;
        RECT 56.990000 59.130000 57.190000 59.330000 ;
        RECT 56.990000 59.540000 57.190000 59.740000 ;
        RECT 56.990000 59.950000 57.190000 60.150000 ;
        RECT 56.990000 60.360000 57.190000 60.560000 ;
        RECT 56.990000 60.770000 57.190000 60.970000 ;
        RECT 56.990000 61.180000 57.190000 61.380000 ;
        RECT 56.990000 61.590000 57.190000 61.790000 ;
        RECT 56.990000 62.000000 57.190000 62.200000 ;
        RECT 56.990000 62.410000 57.190000 62.610000 ;
        RECT 57.395000 58.310000 57.595000 58.510000 ;
        RECT 57.395000 58.720000 57.595000 58.920000 ;
        RECT 57.395000 59.130000 57.595000 59.330000 ;
        RECT 57.395000 59.540000 57.595000 59.740000 ;
        RECT 57.395000 59.950000 57.595000 60.150000 ;
        RECT 57.395000 60.360000 57.595000 60.560000 ;
        RECT 57.395000 60.770000 57.595000 60.970000 ;
        RECT 57.395000 61.180000 57.595000 61.380000 ;
        RECT 57.395000 61.590000 57.595000 61.790000 ;
        RECT 57.395000 62.000000 57.595000 62.200000 ;
        RECT 57.395000 62.410000 57.595000 62.610000 ;
        RECT 57.800000 58.310000 58.000000 58.510000 ;
        RECT 57.800000 58.720000 58.000000 58.920000 ;
        RECT 57.800000 59.130000 58.000000 59.330000 ;
        RECT 57.800000 59.540000 58.000000 59.740000 ;
        RECT 57.800000 59.950000 58.000000 60.150000 ;
        RECT 57.800000 60.360000 58.000000 60.560000 ;
        RECT 57.800000 60.770000 58.000000 60.970000 ;
        RECT 57.800000 61.180000 58.000000 61.380000 ;
        RECT 57.800000 61.590000 58.000000 61.790000 ;
        RECT 57.800000 62.000000 58.000000 62.200000 ;
        RECT 57.800000 62.410000 58.000000 62.610000 ;
        RECT 58.205000 58.310000 58.405000 58.510000 ;
        RECT 58.205000 58.720000 58.405000 58.920000 ;
        RECT 58.205000 59.130000 58.405000 59.330000 ;
        RECT 58.205000 59.540000 58.405000 59.740000 ;
        RECT 58.205000 59.950000 58.405000 60.150000 ;
        RECT 58.205000 60.360000 58.405000 60.560000 ;
        RECT 58.205000 60.770000 58.405000 60.970000 ;
        RECT 58.205000 61.180000 58.405000 61.380000 ;
        RECT 58.205000 61.590000 58.405000 61.790000 ;
        RECT 58.205000 62.000000 58.405000 62.200000 ;
        RECT 58.205000 62.410000 58.405000 62.610000 ;
        RECT 58.610000 58.310000 58.810000 58.510000 ;
        RECT 58.610000 58.720000 58.810000 58.920000 ;
        RECT 58.610000 59.130000 58.810000 59.330000 ;
        RECT 58.610000 59.540000 58.810000 59.740000 ;
        RECT 58.610000 59.950000 58.810000 60.150000 ;
        RECT 58.610000 60.360000 58.810000 60.560000 ;
        RECT 58.610000 60.770000 58.810000 60.970000 ;
        RECT 58.610000 61.180000 58.810000 61.380000 ;
        RECT 58.610000 61.590000 58.810000 61.790000 ;
        RECT 58.610000 62.000000 58.810000 62.200000 ;
        RECT 58.610000 62.410000 58.810000 62.610000 ;
        RECT 59.015000 58.310000 59.215000 58.510000 ;
        RECT 59.015000 58.720000 59.215000 58.920000 ;
        RECT 59.015000 59.130000 59.215000 59.330000 ;
        RECT 59.015000 59.540000 59.215000 59.740000 ;
        RECT 59.015000 59.950000 59.215000 60.150000 ;
        RECT 59.015000 60.360000 59.215000 60.560000 ;
        RECT 59.015000 60.770000 59.215000 60.970000 ;
        RECT 59.015000 61.180000 59.215000 61.380000 ;
        RECT 59.015000 61.590000 59.215000 61.790000 ;
        RECT 59.015000 62.000000 59.215000 62.200000 ;
        RECT 59.015000 62.410000 59.215000 62.610000 ;
        RECT 59.420000 58.310000 59.620000 58.510000 ;
        RECT 59.420000 58.720000 59.620000 58.920000 ;
        RECT 59.420000 59.130000 59.620000 59.330000 ;
        RECT 59.420000 59.540000 59.620000 59.740000 ;
        RECT 59.420000 59.950000 59.620000 60.150000 ;
        RECT 59.420000 60.360000 59.620000 60.560000 ;
        RECT 59.420000 60.770000 59.620000 60.970000 ;
        RECT 59.420000 61.180000 59.620000 61.380000 ;
        RECT 59.420000 61.590000 59.620000 61.790000 ;
        RECT 59.420000 62.000000 59.620000 62.200000 ;
        RECT 59.420000 62.410000 59.620000 62.610000 ;
        RECT 59.825000 58.310000 60.025000 58.510000 ;
        RECT 59.825000 58.720000 60.025000 58.920000 ;
        RECT 59.825000 59.130000 60.025000 59.330000 ;
        RECT 59.825000 59.540000 60.025000 59.740000 ;
        RECT 59.825000 59.950000 60.025000 60.150000 ;
        RECT 59.825000 60.360000 60.025000 60.560000 ;
        RECT 59.825000 60.770000 60.025000 60.970000 ;
        RECT 59.825000 61.180000 60.025000 61.380000 ;
        RECT 59.825000 61.590000 60.025000 61.790000 ;
        RECT 59.825000 62.000000 60.025000 62.200000 ;
        RECT 59.825000 62.410000 60.025000 62.610000 ;
        RECT 60.230000 58.310000 60.430000 58.510000 ;
        RECT 60.230000 58.720000 60.430000 58.920000 ;
        RECT 60.230000 59.130000 60.430000 59.330000 ;
        RECT 60.230000 59.540000 60.430000 59.740000 ;
        RECT 60.230000 59.950000 60.430000 60.150000 ;
        RECT 60.230000 60.360000 60.430000 60.560000 ;
        RECT 60.230000 60.770000 60.430000 60.970000 ;
        RECT 60.230000 61.180000 60.430000 61.380000 ;
        RECT 60.230000 61.590000 60.430000 61.790000 ;
        RECT 60.230000 62.000000 60.430000 62.200000 ;
        RECT 60.230000 62.410000 60.430000 62.610000 ;
        RECT 60.635000 58.310000 60.835000 58.510000 ;
        RECT 60.635000 58.720000 60.835000 58.920000 ;
        RECT 60.635000 59.130000 60.835000 59.330000 ;
        RECT 60.635000 59.540000 60.835000 59.740000 ;
        RECT 60.635000 59.950000 60.835000 60.150000 ;
        RECT 60.635000 60.360000 60.835000 60.560000 ;
        RECT 60.635000 60.770000 60.835000 60.970000 ;
        RECT 60.635000 61.180000 60.835000 61.380000 ;
        RECT 60.635000 61.590000 60.835000 61.790000 ;
        RECT 60.635000 62.000000 60.835000 62.200000 ;
        RECT 60.635000 62.410000 60.835000 62.610000 ;
        RECT 61.040000 58.310000 61.240000 58.510000 ;
        RECT 61.040000 58.720000 61.240000 58.920000 ;
        RECT 61.040000 59.130000 61.240000 59.330000 ;
        RECT 61.040000 59.540000 61.240000 59.740000 ;
        RECT 61.040000 59.950000 61.240000 60.150000 ;
        RECT 61.040000 60.360000 61.240000 60.560000 ;
        RECT 61.040000 60.770000 61.240000 60.970000 ;
        RECT 61.040000 61.180000 61.240000 61.380000 ;
        RECT 61.040000 61.590000 61.240000 61.790000 ;
        RECT 61.040000 62.000000 61.240000 62.200000 ;
        RECT 61.040000 62.410000 61.240000 62.610000 ;
        RECT 61.445000 58.310000 61.645000 58.510000 ;
        RECT 61.445000 58.720000 61.645000 58.920000 ;
        RECT 61.445000 59.130000 61.645000 59.330000 ;
        RECT 61.445000 59.540000 61.645000 59.740000 ;
        RECT 61.445000 59.950000 61.645000 60.150000 ;
        RECT 61.445000 60.360000 61.645000 60.560000 ;
        RECT 61.445000 60.770000 61.645000 60.970000 ;
        RECT 61.445000 61.180000 61.645000 61.380000 ;
        RECT 61.445000 61.590000 61.645000 61.790000 ;
        RECT 61.445000 62.000000 61.645000 62.200000 ;
        RECT 61.445000 62.410000 61.645000 62.610000 ;
        RECT 61.850000 58.310000 62.050000 58.510000 ;
        RECT 61.850000 58.720000 62.050000 58.920000 ;
        RECT 61.850000 59.130000 62.050000 59.330000 ;
        RECT 61.850000 59.540000 62.050000 59.740000 ;
        RECT 61.850000 59.950000 62.050000 60.150000 ;
        RECT 61.850000 60.360000 62.050000 60.560000 ;
        RECT 61.850000 60.770000 62.050000 60.970000 ;
        RECT 61.850000 61.180000 62.050000 61.380000 ;
        RECT 61.850000 61.590000 62.050000 61.790000 ;
        RECT 61.850000 62.000000 62.050000 62.200000 ;
        RECT 61.850000 62.410000 62.050000 62.610000 ;
        RECT 62.255000 58.310000 62.455000 58.510000 ;
        RECT 62.255000 58.720000 62.455000 58.920000 ;
        RECT 62.255000 59.130000 62.455000 59.330000 ;
        RECT 62.255000 59.540000 62.455000 59.740000 ;
        RECT 62.255000 59.950000 62.455000 60.150000 ;
        RECT 62.255000 60.360000 62.455000 60.560000 ;
        RECT 62.255000 60.770000 62.455000 60.970000 ;
        RECT 62.255000 61.180000 62.455000 61.380000 ;
        RECT 62.255000 61.590000 62.455000 61.790000 ;
        RECT 62.255000 62.000000 62.455000 62.200000 ;
        RECT 62.255000 62.410000 62.455000 62.610000 ;
        RECT 62.660000 58.310000 62.860000 58.510000 ;
        RECT 62.660000 58.720000 62.860000 58.920000 ;
        RECT 62.660000 59.130000 62.860000 59.330000 ;
        RECT 62.660000 59.540000 62.860000 59.740000 ;
        RECT 62.660000 59.950000 62.860000 60.150000 ;
        RECT 62.660000 60.360000 62.860000 60.560000 ;
        RECT 62.660000 60.770000 62.860000 60.970000 ;
        RECT 62.660000 61.180000 62.860000 61.380000 ;
        RECT 62.660000 61.590000 62.860000 61.790000 ;
        RECT 62.660000 62.000000 62.860000 62.200000 ;
        RECT 62.660000 62.410000 62.860000 62.610000 ;
        RECT 63.065000 58.310000 63.265000 58.510000 ;
        RECT 63.065000 58.720000 63.265000 58.920000 ;
        RECT 63.065000 59.130000 63.265000 59.330000 ;
        RECT 63.065000 59.540000 63.265000 59.740000 ;
        RECT 63.065000 59.950000 63.265000 60.150000 ;
        RECT 63.065000 60.360000 63.265000 60.560000 ;
        RECT 63.065000 60.770000 63.265000 60.970000 ;
        RECT 63.065000 61.180000 63.265000 61.380000 ;
        RECT 63.065000 61.590000 63.265000 61.790000 ;
        RECT 63.065000 62.000000 63.265000 62.200000 ;
        RECT 63.065000 62.410000 63.265000 62.610000 ;
        RECT 63.470000 58.310000 63.670000 58.510000 ;
        RECT 63.470000 58.720000 63.670000 58.920000 ;
        RECT 63.470000 59.130000 63.670000 59.330000 ;
        RECT 63.470000 59.540000 63.670000 59.740000 ;
        RECT 63.470000 59.950000 63.670000 60.150000 ;
        RECT 63.470000 60.360000 63.670000 60.560000 ;
        RECT 63.470000 60.770000 63.670000 60.970000 ;
        RECT 63.470000 61.180000 63.670000 61.380000 ;
        RECT 63.470000 61.590000 63.670000 61.790000 ;
        RECT 63.470000 62.000000 63.670000 62.200000 ;
        RECT 63.470000 62.410000 63.670000 62.610000 ;
        RECT 63.875000 58.310000 64.075000 58.510000 ;
        RECT 63.875000 58.720000 64.075000 58.920000 ;
        RECT 63.875000 59.130000 64.075000 59.330000 ;
        RECT 63.875000 59.540000 64.075000 59.740000 ;
        RECT 63.875000 59.950000 64.075000 60.150000 ;
        RECT 63.875000 60.360000 64.075000 60.560000 ;
        RECT 63.875000 60.770000 64.075000 60.970000 ;
        RECT 63.875000 61.180000 64.075000 61.380000 ;
        RECT 63.875000 61.590000 64.075000 61.790000 ;
        RECT 63.875000 62.000000 64.075000 62.200000 ;
        RECT 63.875000 62.410000 64.075000 62.610000 ;
        RECT 64.280000 58.310000 64.480000 58.510000 ;
        RECT 64.280000 58.720000 64.480000 58.920000 ;
        RECT 64.280000 59.130000 64.480000 59.330000 ;
        RECT 64.280000 59.540000 64.480000 59.740000 ;
        RECT 64.280000 59.950000 64.480000 60.150000 ;
        RECT 64.280000 60.360000 64.480000 60.560000 ;
        RECT 64.280000 60.770000 64.480000 60.970000 ;
        RECT 64.280000 61.180000 64.480000 61.380000 ;
        RECT 64.280000 61.590000 64.480000 61.790000 ;
        RECT 64.280000 62.000000 64.480000 62.200000 ;
        RECT 64.280000 62.410000 64.480000 62.610000 ;
        RECT 64.685000 58.310000 64.885000 58.510000 ;
        RECT 64.685000 58.720000 64.885000 58.920000 ;
        RECT 64.685000 59.130000 64.885000 59.330000 ;
        RECT 64.685000 59.540000 64.885000 59.740000 ;
        RECT 64.685000 59.950000 64.885000 60.150000 ;
        RECT 64.685000 60.360000 64.885000 60.560000 ;
        RECT 64.685000 60.770000 64.885000 60.970000 ;
        RECT 64.685000 61.180000 64.885000 61.380000 ;
        RECT 64.685000 61.590000 64.885000 61.790000 ;
        RECT 64.685000 62.000000 64.885000 62.200000 ;
        RECT 64.685000 62.410000 64.885000 62.610000 ;
        RECT 65.090000 58.310000 65.290000 58.510000 ;
        RECT 65.090000 58.720000 65.290000 58.920000 ;
        RECT 65.090000 59.130000 65.290000 59.330000 ;
        RECT 65.090000 59.540000 65.290000 59.740000 ;
        RECT 65.090000 59.950000 65.290000 60.150000 ;
        RECT 65.090000 60.360000 65.290000 60.560000 ;
        RECT 65.090000 60.770000 65.290000 60.970000 ;
        RECT 65.090000 61.180000 65.290000 61.380000 ;
        RECT 65.090000 61.590000 65.290000 61.790000 ;
        RECT 65.090000 62.000000 65.290000 62.200000 ;
        RECT 65.090000 62.410000 65.290000 62.610000 ;
        RECT 65.495000 58.310000 65.695000 58.510000 ;
        RECT 65.495000 58.720000 65.695000 58.920000 ;
        RECT 65.495000 59.130000 65.695000 59.330000 ;
        RECT 65.495000 59.540000 65.695000 59.740000 ;
        RECT 65.495000 59.950000 65.695000 60.150000 ;
        RECT 65.495000 60.360000 65.695000 60.560000 ;
        RECT 65.495000 60.770000 65.695000 60.970000 ;
        RECT 65.495000 61.180000 65.695000 61.380000 ;
        RECT 65.495000 61.590000 65.695000 61.790000 ;
        RECT 65.495000 62.000000 65.695000 62.200000 ;
        RECT 65.495000 62.410000 65.695000 62.610000 ;
        RECT 65.900000 58.310000 66.100000 58.510000 ;
        RECT 65.900000 58.720000 66.100000 58.920000 ;
        RECT 65.900000 59.130000 66.100000 59.330000 ;
        RECT 65.900000 59.540000 66.100000 59.740000 ;
        RECT 65.900000 59.950000 66.100000 60.150000 ;
        RECT 65.900000 60.360000 66.100000 60.560000 ;
        RECT 65.900000 60.770000 66.100000 60.970000 ;
        RECT 65.900000 61.180000 66.100000 61.380000 ;
        RECT 65.900000 61.590000 66.100000 61.790000 ;
        RECT 65.900000 62.000000 66.100000 62.200000 ;
        RECT 65.900000 62.410000 66.100000 62.610000 ;
        RECT 66.305000 58.310000 66.505000 58.510000 ;
        RECT 66.305000 58.720000 66.505000 58.920000 ;
        RECT 66.305000 59.130000 66.505000 59.330000 ;
        RECT 66.305000 59.540000 66.505000 59.740000 ;
        RECT 66.305000 59.950000 66.505000 60.150000 ;
        RECT 66.305000 60.360000 66.505000 60.560000 ;
        RECT 66.305000 60.770000 66.505000 60.970000 ;
        RECT 66.305000 61.180000 66.505000 61.380000 ;
        RECT 66.305000 61.590000 66.505000 61.790000 ;
        RECT 66.305000 62.000000 66.505000 62.200000 ;
        RECT 66.305000 62.410000 66.505000 62.610000 ;
        RECT 66.710000 58.310000 66.910000 58.510000 ;
        RECT 66.710000 58.720000 66.910000 58.920000 ;
        RECT 66.710000 59.130000 66.910000 59.330000 ;
        RECT 66.710000 59.540000 66.910000 59.740000 ;
        RECT 66.710000 59.950000 66.910000 60.150000 ;
        RECT 66.710000 60.360000 66.910000 60.560000 ;
        RECT 66.710000 60.770000 66.910000 60.970000 ;
        RECT 66.710000 61.180000 66.910000 61.380000 ;
        RECT 66.710000 61.590000 66.910000 61.790000 ;
        RECT 66.710000 62.000000 66.910000 62.200000 ;
        RECT 66.710000 62.410000 66.910000 62.610000 ;
        RECT 67.115000 58.310000 67.315000 58.510000 ;
        RECT 67.115000 58.720000 67.315000 58.920000 ;
        RECT 67.115000 59.130000 67.315000 59.330000 ;
        RECT 67.115000 59.540000 67.315000 59.740000 ;
        RECT 67.115000 59.950000 67.315000 60.150000 ;
        RECT 67.115000 60.360000 67.315000 60.560000 ;
        RECT 67.115000 60.770000 67.315000 60.970000 ;
        RECT 67.115000 61.180000 67.315000 61.380000 ;
        RECT 67.115000 61.590000 67.315000 61.790000 ;
        RECT 67.115000 62.000000 67.315000 62.200000 ;
        RECT 67.115000 62.410000 67.315000 62.610000 ;
        RECT 67.520000 58.310000 67.720000 58.510000 ;
        RECT 67.520000 58.720000 67.720000 58.920000 ;
        RECT 67.520000 59.130000 67.720000 59.330000 ;
        RECT 67.520000 59.540000 67.720000 59.740000 ;
        RECT 67.520000 59.950000 67.720000 60.150000 ;
        RECT 67.520000 60.360000 67.720000 60.560000 ;
        RECT 67.520000 60.770000 67.720000 60.970000 ;
        RECT 67.520000 61.180000 67.720000 61.380000 ;
        RECT 67.520000 61.590000 67.720000 61.790000 ;
        RECT 67.520000 62.000000 67.720000 62.200000 ;
        RECT 67.520000 62.410000 67.720000 62.610000 ;
        RECT 67.925000 58.310000 68.125000 58.510000 ;
        RECT 67.925000 58.720000 68.125000 58.920000 ;
        RECT 67.925000 59.130000 68.125000 59.330000 ;
        RECT 67.925000 59.540000 68.125000 59.740000 ;
        RECT 67.925000 59.950000 68.125000 60.150000 ;
        RECT 67.925000 60.360000 68.125000 60.560000 ;
        RECT 67.925000 60.770000 68.125000 60.970000 ;
        RECT 67.925000 61.180000 68.125000 61.380000 ;
        RECT 67.925000 61.590000 68.125000 61.790000 ;
        RECT 67.925000 62.000000 68.125000 62.200000 ;
        RECT 67.925000 62.410000 68.125000 62.610000 ;
        RECT 68.330000 58.310000 68.530000 58.510000 ;
        RECT 68.330000 58.720000 68.530000 58.920000 ;
        RECT 68.330000 59.130000 68.530000 59.330000 ;
        RECT 68.330000 59.540000 68.530000 59.740000 ;
        RECT 68.330000 59.950000 68.530000 60.150000 ;
        RECT 68.330000 60.360000 68.530000 60.560000 ;
        RECT 68.330000 60.770000 68.530000 60.970000 ;
        RECT 68.330000 61.180000 68.530000 61.380000 ;
        RECT 68.330000 61.590000 68.530000 61.790000 ;
        RECT 68.330000 62.000000 68.530000 62.200000 ;
        RECT 68.330000 62.410000 68.530000 62.610000 ;
        RECT 68.735000 58.310000 68.935000 58.510000 ;
        RECT 68.735000 58.720000 68.935000 58.920000 ;
        RECT 68.735000 59.130000 68.935000 59.330000 ;
        RECT 68.735000 59.540000 68.935000 59.740000 ;
        RECT 68.735000 59.950000 68.935000 60.150000 ;
        RECT 68.735000 60.360000 68.935000 60.560000 ;
        RECT 68.735000 60.770000 68.935000 60.970000 ;
        RECT 68.735000 61.180000 68.935000 61.380000 ;
        RECT 68.735000 61.590000 68.935000 61.790000 ;
        RECT 68.735000 62.000000 68.935000 62.200000 ;
        RECT 68.735000 62.410000 68.935000 62.610000 ;
        RECT 69.140000 58.310000 69.340000 58.510000 ;
        RECT 69.140000 58.720000 69.340000 58.920000 ;
        RECT 69.140000 59.130000 69.340000 59.330000 ;
        RECT 69.140000 59.540000 69.340000 59.740000 ;
        RECT 69.140000 59.950000 69.340000 60.150000 ;
        RECT 69.140000 60.360000 69.340000 60.560000 ;
        RECT 69.140000 60.770000 69.340000 60.970000 ;
        RECT 69.140000 61.180000 69.340000 61.380000 ;
        RECT 69.140000 61.590000 69.340000 61.790000 ;
        RECT 69.140000 62.000000 69.340000 62.200000 ;
        RECT 69.140000 62.410000 69.340000 62.610000 ;
        RECT 69.545000 58.310000 69.745000 58.510000 ;
        RECT 69.545000 58.720000 69.745000 58.920000 ;
        RECT 69.545000 59.130000 69.745000 59.330000 ;
        RECT 69.545000 59.540000 69.745000 59.740000 ;
        RECT 69.545000 59.950000 69.745000 60.150000 ;
        RECT 69.545000 60.360000 69.745000 60.560000 ;
        RECT 69.545000 60.770000 69.745000 60.970000 ;
        RECT 69.545000 61.180000 69.745000 61.380000 ;
        RECT 69.545000 61.590000 69.745000 61.790000 ;
        RECT 69.545000 62.000000 69.745000 62.200000 ;
        RECT 69.545000 62.410000 69.745000 62.610000 ;
        RECT 69.950000 58.310000 70.150000 58.510000 ;
        RECT 69.950000 58.720000 70.150000 58.920000 ;
        RECT 69.950000 59.130000 70.150000 59.330000 ;
        RECT 69.950000 59.540000 70.150000 59.740000 ;
        RECT 69.950000 59.950000 70.150000 60.150000 ;
        RECT 69.950000 60.360000 70.150000 60.560000 ;
        RECT 69.950000 60.770000 70.150000 60.970000 ;
        RECT 69.950000 61.180000 70.150000 61.380000 ;
        RECT 69.950000 61.590000 70.150000 61.790000 ;
        RECT 69.950000 62.000000 70.150000 62.200000 ;
        RECT 69.950000 62.410000 70.150000 62.610000 ;
        RECT 70.355000 58.310000 70.555000 58.510000 ;
        RECT 70.355000 58.720000 70.555000 58.920000 ;
        RECT 70.355000 59.130000 70.555000 59.330000 ;
        RECT 70.355000 59.540000 70.555000 59.740000 ;
        RECT 70.355000 59.950000 70.555000 60.150000 ;
        RECT 70.355000 60.360000 70.555000 60.560000 ;
        RECT 70.355000 60.770000 70.555000 60.970000 ;
        RECT 70.355000 61.180000 70.555000 61.380000 ;
        RECT 70.355000 61.590000 70.555000 61.790000 ;
        RECT 70.355000 62.000000 70.555000 62.200000 ;
        RECT 70.355000 62.410000 70.555000 62.610000 ;
        RECT 70.760000 58.310000 70.960000 58.510000 ;
        RECT 70.760000 58.720000 70.960000 58.920000 ;
        RECT 70.760000 59.130000 70.960000 59.330000 ;
        RECT 70.760000 59.540000 70.960000 59.740000 ;
        RECT 70.760000 59.950000 70.960000 60.150000 ;
        RECT 70.760000 60.360000 70.960000 60.560000 ;
        RECT 70.760000 60.770000 70.960000 60.970000 ;
        RECT 70.760000 61.180000 70.960000 61.380000 ;
        RECT 70.760000 61.590000 70.960000 61.790000 ;
        RECT 70.760000 62.000000 70.960000 62.200000 ;
        RECT 70.760000 62.410000 70.960000 62.610000 ;
        RECT 71.165000 58.310000 71.365000 58.510000 ;
        RECT 71.165000 58.720000 71.365000 58.920000 ;
        RECT 71.165000 59.130000 71.365000 59.330000 ;
        RECT 71.165000 59.540000 71.365000 59.740000 ;
        RECT 71.165000 59.950000 71.365000 60.150000 ;
        RECT 71.165000 60.360000 71.365000 60.560000 ;
        RECT 71.165000 60.770000 71.365000 60.970000 ;
        RECT 71.165000 61.180000 71.365000 61.380000 ;
        RECT 71.165000 61.590000 71.365000 61.790000 ;
        RECT 71.165000 62.000000 71.365000 62.200000 ;
        RECT 71.165000 62.410000 71.365000 62.610000 ;
        RECT 71.570000 58.310000 71.770000 58.510000 ;
        RECT 71.570000 58.720000 71.770000 58.920000 ;
        RECT 71.570000 59.130000 71.770000 59.330000 ;
        RECT 71.570000 59.540000 71.770000 59.740000 ;
        RECT 71.570000 59.950000 71.770000 60.150000 ;
        RECT 71.570000 60.360000 71.770000 60.560000 ;
        RECT 71.570000 60.770000 71.770000 60.970000 ;
        RECT 71.570000 61.180000 71.770000 61.380000 ;
        RECT 71.570000 61.590000 71.770000 61.790000 ;
        RECT 71.570000 62.000000 71.770000 62.200000 ;
        RECT 71.570000 62.410000 71.770000 62.610000 ;
        RECT 71.975000 58.310000 72.175000 58.510000 ;
        RECT 71.975000 58.720000 72.175000 58.920000 ;
        RECT 71.975000 59.130000 72.175000 59.330000 ;
        RECT 71.975000 59.540000 72.175000 59.740000 ;
        RECT 71.975000 59.950000 72.175000 60.150000 ;
        RECT 71.975000 60.360000 72.175000 60.560000 ;
        RECT 71.975000 60.770000 72.175000 60.970000 ;
        RECT 71.975000 61.180000 72.175000 61.380000 ;
        RECT 71.975000 61.590000 72.175000 61.790000 ;
        RECT 71.975000 62.000000 72.175000 62.200000 ;
        RECT 71.975000 62.410000 72.175000 62.610000 ;
        RECT 72.380000 58.310000 72.580000 58.510000 ;
        RECT 72.380000 58.720000 72.580000 58.920000 ;
        RECT 72.380000 59.130000 72.580000 59.330000 ;
        RECT 72.380000 59.540000 72.580000 59.740000 ;
        RECT 72.380000 59.950000 72.580000 60.150000 ;
        RECT 72.380000 60.360000 72.580000 60.560000 ;
        RECT 72.380000 60.770000 72.580000 60.970000 ;
        RECT 72.380000 61.180000 72.580000 61.380000 ;
        RECT 72.380000 61.590000 72.580000 61.790000 ;
        RECT 72.380000 62.000000 72.580000 62.200000 ;
        RECT 72.380000 62.410000 72.580000 62.610000 ;
        RECT 72.785000 58.310000 72.985000 58.510000 ;
        RECT 72.785000 58.720000 72.985000 58.920000 ;
        RECT 72.785000 59.130000 72.985000 59.330000 ;
        RECT 72.785000 59.540000 72.985000 59.740000 ;
        RECT 72.785000 59.950000 72.985000 60.150000 ;
        RECT 72.785000 60.360000 72.985000 60.560000 ;
        RECT 72.785000 60.770000 72.985000 60.970000 ;
        RECT 72.785000 61.180000 72.985000 61.380000 ;
        RECT 72.785000 61.590000 72.985000 61.790000 ;
        RECT 72.785000 62.000000 72.985000 62.200000 ;
        RECT 72.785000 62.410000 72.985000 62.610000 ;
        RECT 73.190000 58.310000 73.390000 58.510000 ;
        RECT 73.190000 58.720000 73.390000 58.920000 ;
        RECT 73.190000 59.130000 73.390000 59.330000 ;
        RECT 73.190000 59.540000 73.390000 59.740000 ;
        RECT 73.190000 59.950000 73.390000 60.150000 ;
        RECT 73.190000 60.360000 73.390000 60.560000 ;
        RECT 73.190000 60.770000 73.390000 60.970000 ;
        RECT 73.190000 61.180000 73.390000 61.380000 ;
        RECT 73.190000 61.590000 73.390000 61.790000 ;
        RECT 73.190000 62.000000 73.390000 62.200000 ;
        RECT 73.190000 62.410000 73.390000 62.610000 ;
        RECT 73.595000 58.310000 73.795000 58.510000 ;
        RECT 73.595000 58.720000 73.795000 58.920000 ;
        RECT 73.595000 59.130000 73.795000 59.330000 ;
        RECT 73.595000 59.540000 73.795000 59.740000 ;
        RECT 73.595000 59.950000 73.795000 60.150000 ;
        RECT 73.595000 60.360000 73.795000 60.560000 ;
        RECT 73.595000 60.770000 73.795000 60.970000 ;
        RECT 73.595000 61.180000 73.795000 61.380000 ;
        RECT 73.595000 61.590000 73.795000 61.790000 ;
        RECT 73.595000 62.000000 73.795000 62.200000 ;
        RECT 73.595000 62.410000 73.795000 62.610000 ;
        RECT 74.000000 58.310000 74.200000 58.510000 ;
        RECT 74.000000 58.720000 74.200000 58.920000 ;
        RECT 74.000000 59.130000 74.200000 59.330000 ;
        RECT 74.000000 59.540000 74.200000 59.740000 ;
        RECT 74.000000 59.950000 74.200000 60.150000 ;
        RECT 74.000000 60.360000 74.200000 60.560000 ;
        RECT 74.000000 60.770000 74.200000 60.970000 ;
        RECT 74.000000 61.180000 74.200000 61.380000 ;
        RECT 74.000000 61.590000 74.200000 61.790000 ;
        RECT 74.000000 62.000000 74.200000 62.200000 ;
        RECT 74.000000 62.410000 74.200000 62.610000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730000 31.885000 75.000000 35.335000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 31.985000 1.270000 35.235000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met1 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 75.000000 200.000000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000 75.000000  25.440000 ;
      RECT  0.000000  30.880000 75.000000  57.840000 ;
      RECT  0.000000  63.080000 75.000000 172.755000 ;
      RECT 13.900000  63.080000 61.100000 195.174000 ;
      RECT 13.900000  63.080000 75.000000 172.920000 ;
      RECT 13.900000 172.755000 75.000000 172.920000 ;
      RECT 13.900000 172.920000 61.100000 195.144000 ;
      RECT 13.900000 195.144000 61.084000 195.160000 ;
      RECT 13.900000 195.144000 61.084000 195.160000 ;
      RECT 13.900000 195.160000 61.069000 195.175000 ;
      RECT 13.900000 195.160000 61.069000 195.175000 ;
      RECT 14.051000 195.174000 60.919000 195.325000 ;
      RECT 14.051000 195.174000 60.919000 195.325000 ;
      RECT 14.201000 195.325000 60.769000 195.475000 ;
      RECT 14.201000 195.325000 60.769000 195.475000 ;
      RECT 14.351000 195.475000 60.619000 195.625000 ;
      RECT 14.351000 195.475000 60.619000 195.625000 ;
      RECT 14.501000 195.625000 60.469000 195.775000 ;
      RECT 14.501000 195.625000 60.469000 195.775000 ;
      RECT 14.651000 195.775000 60.319000 195.925000 ;
      RECT 14.651000 195.775000 60.319000 195.925000 ;
      RECT 14.801000 195.925000 60.169000 196.075000 ;
      RECT 14.801000 195.925000 60.169000 196.075000 ;
      RECT 14.951000 196.075000 60.019000 196.225000 ;
      RECT 14.951000 196.075000 60.019000 196.225000 ;
      RECT 15.101000 196.225000 59.869000 196.375000 ;
      RECT 15.101000 196.225000 59.869000 196.375000 ;
      RECT 15.251000 196.375000 59.719000 196.525000 ;
      RECT 15.251000 196.375000 59.719000 196.525000 ;
      RECT 15.401000 196.525000 59.569000 196.675000 ;
      RECT 15.401000 196.525000 59.569000 196.675000 ;
      RECT 15.501000 196.675000 59.469000 196.775000 ;
      RECT 15.501000 196.675000 59.469000 196.775000 ;
      RECT 24.795000   0.000000 49.990000  63.080000 ;
      RECT 24.795000   0.000000 49.990000 172.920000 ;
      RECT 24.795000  25.440000 49.990000  30.880000 ;
      RECT 24.795000  57.840000 49.990000  63.080000 ;
      RECT 74.690000  25.440000 75.000000  30.880000 ;
      RECT 74.690000  57.840000 75.000000  63.080000 ;
      RECT 74.690000 172.920000 75.000000 200.000000 ;
    LAYER met4 ;
      RECT  0.000000   0.000000  1.670000   1.635000 ;
      RECT  0.000000   7.885000  1.670000   8.485000 ;
      RECT  0.000000  13.935000  1.365000  14.535000 ;
      RECT  0.000000  18.785000  1.365000  19.385000 ;
      RECT  0.000000  24.835000  1.670000  25.435000 ;
      RECT  0.000000  30.885000  1.670000  31.485000 ;
      RECT  0.000000  35.735000  1.670000  36.335000 ;
      RECT  0.000000  40.585000  1.670000  41.185000 ;
      RECT  0.000000  46.635000  1.670000  47.335000 ;
      RECT  0.000000  57.135000  1.670000  57.835000 ;
      RECT  0.000000  63.085000  1.670000  63.685000 ;
      RECT  0.000000  68.935000  1.670000  69.635000 ;
      RECT  0.000000  95.400000 75.000000 175.385000 ;
      RECT  1.365000  13.935000 73.635000  19.385000 ;
      RECT  1.365000  13.935000 73.635000  19.385000 ;
      RECT  1.670000   0.000000 73.330000  13.935000 ;
      RECT  1.670000   0.000000 73.330000  25.435000 ;
      RECT  1.670000   0.000000 73.330000  25.435000 ;
      RECT  1.670000   0.000000 73.330000  25.435000 ;
      RECT  1.670000  19.385000 73.330000  25.435000 ;
      RECT  1.670000  30.885000 73.330000  57.835000 ;
      RECT  1.670000  30.885000 73.330000  57.835000 ;
      RECT  1.670000  30.885000 73.330000  57.835000 ;
      RECT  1.670000  30.885000 73.330000  57.835000 ;
      RECT  1.670000  30.885000 73.330000  57.835000 ;
      RECT  1.670000  63.085000 73.330000  95.400000 ;
      RECT  1.670000  63.085000 73.330000 175.530000 ;
      RECT  1.670000  63.085000 73.330000 175.530000 ;
      RECT  1.670000  63.085000 73.330000 175.530000 ;
      RECT  1.670000 175.385000 73.330000 175.530000 ;
      RECT 13.875000  63.085000 61.105000 195.830000 ;
      RECT 13.875000 175.530000 61.105000 195.830000 ;
      RECT 14.655000  63.085000 60.280000 196.770000 ;
      RECT 14.655000 195.830000 60.280000 196.770000 ;
      RECT 24.770000   0.000000 50.015000  63.085000 ;
      RECT 24.770000   0.000000 50.015000 196.770000 ;
      RECT 24.770000  25.435000 50.015000  30.885000 ;
      RECT 24.770000  57.835000 50.015000  63.085000 ;
      RECT 73.330000   0.000000 75.000000   1.635000 ;
      RECT 73.330000   7.885000 75.000000   8.485000 ;
      RECT 73.330000  24.835000 75.000000  25.435000 ;
      RECT 73.330000  30.885000 75.000000  31.485000 ;
      RECT 73.330000  35.735000 75.000000  36.335000 ;
      RECT 73.330000  40.585000 75.000000  41.185000 ;
      RECT 73.330000  46.635000 75.000000  47.335000 ;
      RECT 73.330000  57.135000 75.000000  57.835000 ;
      RECT 73.330000  63.085000 75.000000  63.685000 ;
      RECT 73.330000  68.935000 75.000000  69.635000 ;
      RECT 73.635000  13.935000 75.000000  14.535000 ;
      RECT 73.635000  18.785000 75.000000  19.385000 ;
    LAYER met5 ;
      RECT 0.000000   0.000000 75.000000   1.335000 ;
      RECT 0.000000  95.785000 75.000000 174.985000 ;
      RECT 1.765000  14.235000 73.235000  19.085000 ;
      RECT 2.070000   1.335000 72.930000  14.235000 ;
      RECT 2.070000  19.085000 72.930000  95.785000 ;
      RECT 2.070000 174.985000 72.930000 200.000000 ;
  END
END sky130_fd_io__overlay_vssio_hvc
END LIBRARY
