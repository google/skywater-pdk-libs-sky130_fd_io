# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__overlay_vdda_lvc
  CLASS BLOCK ;
  FOREIGN sky130_fd_io__overlay_vdda_lvc ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  75.00000 BY  198.0000 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 51.125000 75.000000 54.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 46.365000 75.000000 49.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 6.985000 75.000000 11.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 0.135000 75.000000 5.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.630000 12.960000 0.950000 13.280000 ;
      LAYER met4 ;
        RECT 0.630000 12.960000 0.950000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 13.400000 0.950000 13.720000 ;
      LAYER met4 ;
        RECT 0.630000 13.400000 0.950000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 13.840000 0.950000 14.160000 ;
      LAYER met4 ;
        RECT 0.630000 13.840000 0.950000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 14.280000 0.950000 14.600000 ;
      LAYER met4 ;
        RECT 0.630000 14.280000 0.950000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 14.720000 0.950000 15.040000 ;
      LAYER met4 ;
        RECT 0.630000 14.720000 0.950000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 15.160000 0.950000 15.480000 ;
      LAYER met4 ;
        RECT 0.630000 15.160000 0.950000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 15.600000 0.950000 15.920000 ;
      LAYER met4 ;
        RECT 0.630000 15.600000 0.950000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630000 16.040000 0.950000 16.360000 ;
      LAYER met4 ;
        RECT 0.630000 16.040000 0.950000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040000 12.960000 1.360000 13.280000 ;
      LAYER met4 ;
        RECT 1.040000 12.960000 1.360000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040000 13.400000 1.360000 13.720000 ;
      LAYER met4 ;
        RECT 1.040000 13.400000 1.360000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040000 13.840000 1.360000 14.160000 ;
      LAYER met4 ;
        RECT 1.040000 13.840000 1.360000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040000 14.280000 1.360000 14.600000 ;
      LAYER met4 ;
        RECT 1.040000 14.280000 1.360000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040000 14.720000 1.360000 15.040000 ;
      LAYER met4 ;
        RECT 1.040000 14.720000 1.360000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040000 15.160000 1.360000 15.480000 ;
      LAYER met4 ;
        RECT 1.040000 15.160000 1.360000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040000 15.600000 1.360000 15.920000 ;
      LAYER met4 ;
        RECT 1.040000 15.600000 1.360000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040000 16.040000 1.360000 16.360000 ;
      LAYER met4 ;
        RECT 1.040000 16.040000 1.360000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450000 12.960000 1.770000 13.280000 ;
      LAYER met4 ;
        RECT 1.450000 12.960000 1.770000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450000 13.400000 1.770000 13.720000 ;
      LAYER met4 ;
        RECT 1.450000 13.400000 1.770000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450000 13.840000 1.770000 14.160000 ;
      LAYER met4 ;
        RECT 1.450000 13.840000 1.770000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450000 14.280000 1.770000 14.600000 ;
      LAYER met4 ;
        RECT 1.450000 14.280000 1.770000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450000 14.720000 1.770000 15.040000 ;
      LAYER met4 ;
        RECT 1.450000 14.720000 1.770000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450000 15.160000 1.770000 15.480000 ;
      LAYER met4 ;
        RECT 1.450000 15.160000 1.770000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450000 15.600000 1.770000 15.920000 ;
      LAYER met4 ;
        RECT 1.450000 15.600000 1.770000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450000 16.040000 1.770000 16.360000 ;
      LAYER met4 ;
        RECT 1.450000 16.040000 1.770000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860000 12.960000 2.180000 13.280000 ;
      LAYER met4 ;
        RECT 1.860000 12.960000 2.180000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860000 13.400000 2.180000 13.720000 ;
      LAYER met4 ;
        RECT 1.860000 13.400000 2.180000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860000 13.840000 2.180000 14.160000 ;
      LAYER met4 ;
        RECT 1.860000 13.840000 2.180000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860000 14.280000 2.180000 14.600000 ;
      LAYER met4 ;
        RECT 1.860000 14.280000 2.180000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860000 14.720000 2.180000 15.040000 ;
      LAYER met4 ;
        RECT 1.860000 14.720000 2.180000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860000 15.160000 2.180000 15.480000 ;
      LAYER met4 ;
        RECT 1.860000 15.160000 2.180000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860000 15.600000 2.180000 15.920000 ;
      LAYER met4 ;
        RECT 1.860000 15.600000 2.180000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860000 16.040000 2.180000 16.360000 ;
      LAYER met4 ;
        RECT 1.860000 16.040000 2.180000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380000 12.960000 10.700000 13.280000 ;
      LAYER met4 ;
        RECT 10.380000 12.960000 10.700000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380000 13.400000 10.700000 13.720000 ;
      LAYER met4 ;
        RECT 10.380000 13.400000 10.700000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380000 13.840000 10.700000 14.160000 ;
      LAYER met4 ;
        RECT 10.380000 13.840000 10.700000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380000 14.280000 10.700000 14.600000 ;
      LAYER met4 ;
        RECT 10.380000 14.280000 10.700000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380000 14.720000 10.700000 15.040000 ;
      LAYER met4 ;
        RECT 10.380000 14.720000 10.700000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380000 15.160000 10.700000 15.480000 ;
      LAYER met4 ;
        RECT 10.380000 15.160000 10.700000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380000 15.600000 10.700000 15.920000 ;
      LAYER met4 ;
        RECT 10.380000 15.600000 10.700000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380000 16.040000 10.700000 16.360000 ;
      LAYER met4 ;
        RECT 10.380000 16.040000 10.700000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 12.960000 11.105000 13.280000 ;
      LAYER met4 ;
        RECT 10.785000 12.960000 11.105000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 13.400000 11.105000 13.720000 ;
      LAYER met4 ;
        RECT 10.785000 13.400000 11.105000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 13.840000 11.105000 14.160000 ;
      LAYER met4 ;
        RECT 10.785000 13.840000 11.105000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 14.280000 11.105000 14.600000 ;
      LAYER met4 ;
        RECT 10.785000 14.280000 11.105000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 14.720000 11.105000 15.040000 ;
      LAYER met4 ;
        RECT 10.785000 14.720000 11.105000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 15.160000 11.105000 15.480000 ;
      LAYER met4 ;
        RECT 10.785000 15.160000 11.105000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 15.600000 11.105000 15.920000 ;
      LAYER met4 ;
        RECT 10.785000 15.600000 11.105000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785000 16.040000 11.105000 16.360000 ;
      LAYER met4 ;
        RECT 10.785000 16.040000 11.105000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190000 12.960000 11.510000 13.280000 ;
      LAYER met4 ;
        RECT 11.190000 12.960000 11.510000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190000 13.400000 11.510000 13.720000 ;
      LAYER met4 ;
        RECT 11.190000 13.400000 11.510000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190000 13.840000 11.510000 14.160000 ;
      LAYER met4 ;
        RECT 11.190000 13.840000 11.510000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190000 14.280000 11.510000 14.600000 ;
      LAYER met4 ;
        RECT 11.190000 14.280000 11.510000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190000 14.720000 11.510000 15.040000 ;
      LAYER met4 ;
        RECT 11.190000 14.720000 11.510000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190000 15.160000 11.510000 15.480000 ;
      LAYER met4 ;
        RECT 11.190000 15.160000 11.510000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190000 15.600000 11.510000 15.920000 ;
      LAYER met4 ;
        RECT 11.190000 15.600000 11.510000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190000 16.040000 11.510000 16.360000 ;
      LAYER met4 ;
        RECT 11.190000 16.040000 11.510000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595000 12.960000 11.915000 13.280000 ;
      LAYER met4 ;
        RECT 11.595000 12.960000 11.915000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595000 13.400000 11.915000 13.720000 ;
      LAYER met4 ;
        RECT 11.595000 13.400000 11.915000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595000 13.840000 11.915000 14.160000 ;
      LAYER met4 ;
        RECT 11.595000 13.840000 11.915000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595000 14.280000 11.915000 14.600000 ;
      LAYER met4 ;
        RECT 11.595000 14.280000 11.915000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595000 14.720000 11.915000 15.040000 ;
      LAYER met4 ;
        RECT 11.595000 14.720000 11.915000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595000 15.160000 11.915000 15.480000 ;
      LAYER met4 ;
        RECT 11.595000 15.160000 11.915000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595000 15.600000 11.915000 15.920000 ;
      LAYER met4 ;
        RECT 11.595000 15.600000 11.915000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595000 16.040000 11.915000 16.360000 ;
      LAYER met4 ;
        RECT 11.595000 16.040000 11.915000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000000 12.960000 12.320000 13.280000 ;
      LAYER met4 ;
        RECT 12.000000 12.960000 12.320000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000000 13.400000 12.320000 13.720000 ;
      LAYER met4 ;
        RECT 12.000000 13.400000 12.320000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000000 13.840000 12.320000 14.160000 ;
      LAYER met4 ;
        RECT 12.000000 13.840000 12.320000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000000 14.280000 12.320000 14.600000 ;
      LAYER met4 ;
        RECT 12.000000 14.280000 12.320000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000000 14.720000 12.320000 15.040000 ;
      LAYER met4 ;
        RECT 12.000000 14.720000 12.320000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000000 15.160000 12.320000 15.480000 ;
      LAYER met4 ;
        RECT 12.000000 15.160000 12.320000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000000 15.600000 12.320000 15.920000 ;
      LAYER met4 ;
        RECT 12.000000 15.600000 12.320000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000000 16.040000 12.320000 16.360000 ;
      LAYER met4 ;
        RECT 12.000000 16.040000 12.320000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405000 12.960000 12.725000 13.280000 ;
      LAYER met4 ;
        RECT 12.405000 12.960000 12.725000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405000 13.400000 12.725000 13.720000 ;
      LAYER met4 ;
        RECT 12.405000 13.400000 12.725000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405000 13.840000 12.725000 14.160000 ;
      LAYER met4 ;
        RECT 12.405000 13.840000 12.725000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405000 14.280000 12.725000 14.600000 ;
      LAYER met4 ;
        RECT 12.405000 14.280000 12.725000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405000 14.720000 12.725000 15.040000 ;
      LAYER met4 ;
        RECT 12.405000 14.720000 12.725000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405000 15.160000 12.725000 15.480000 ;
      LAYER met4 ;
        RECT 12.405000 15.160000 12.725000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405000 15.600000 12.725000 15.920000 ;
      LAYER met4 ;
        RECT 12.405000 15.600000 12.725000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405000 16.040000 12.725000 16.360000 ;
      LAYER met4 ;
        RECT 12.405000 16.040000 12.725000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810000 12.960000 13.130000 13.280000 ;
      LAYER met4 ;
        RECT 12.810000 12.960000 13.130000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810000 13.400000 13.130000 13.720000 ;
      LAYER met4 ;
        RECT 12.810000 13.400000 13.130000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810000 13.840000 13.130000 14.160000 ;
      LAYER met4 ;
        RECT 12.810000 13.840000 13.130000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810000 14.280000 13.130000 14.600000 ;
      LAYER met4 ;
        RECT 12.810000 14.280000 13.130000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810000 14.720000 13.130000 15.040000 ;
      LAYER met4 ;
        RECT 12.810000 14.720000 13.130000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810000 15.160000 13.130000 15.480000 ;
      LAYER met4 ;
        RECT 12.810000 15.160000 13.130000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810000 15.600000 13.130000 15.920000 ;
      LAYER met4 ;
        RECT 12.810000 15.600000 13.130000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810000 16.040000 13.130000 16.360000 ;
      LAYER met4 ;
        RECT 12.810000 16.040000 13.130000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215000 12.960000 13.535000 13.280000 ;
      LAYER met4 ;
        RECT 13.215000 12.960000 13.535000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215000 13.400000 13.535000 13.720000 ;
      LAYER met4 ;
        RECT 13.215000 13.400000 13.535000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215000 13.840000 13.535000 14.160000 ;
      LAYER met4 ;
        RECT 13.215000 13.840000 13.535000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215000 14.280000 13.535000 14.600000 ;
      LAYER met4 ;
        RECT 13.215000 14.280000 13.535000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215000 14.720000 13.535000 15.040000 ;
      LAYER met4 ;
        RECT 13.215000 14.720000 13.535000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215000 15.160000 13.535000 15.480000 ;
      LAYER met4 ;
        RECT 13.215000 15.160000 13.535000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215000 15.600000 13.535000 15.920000 ;
      LAYER met4 ;
        RECT 13.215000 15.600000 13.535000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215000 16.040000 13.535000 16.360000 ;
      LAYER met4 ;
        RECT 13.215000 16.040000 13.535000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620000 12.960000 13.940000 13.280000 ;
      LAYER met4 ;
        RECT 13.620000 12.960000 13.940000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620000 13.400000 13.940000 13.720000 ;
      LAYER met4 ;
        RECT 13.620000 13.400000 13.940000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620000 13.840000 13.940000 14.160000 ;
      LAYER met4 ;
        RECT 13.620000 13.840000 13.940000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620000 14.280000 13.940000 14.600000 ;
      LAYER met4 ;
        RECT 13.620000 14.280000 13.940000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620000 14.720000 13.940000 15.040000 ;
      LAYER met4 ;
        RECT 13.620000 14.720000 13.940000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620000 15.160000 13.940000 15.480000 ;
      LAYER met4 ;
        RECT 13.620000 15.160000 13.940000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620000 15.600000 13.940000 15.920000 ;
      LAYER met4 ;
        RECT 13.620000 15.600000 13.940000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620000 16.040000 13.940000 16.360000 ;
      LAYER met4 ;
        RECT 13.620000 16.040000 13.940000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025000 12.960000 14.345000 13.280000 ;
      LAYER met4 ;
        RECT 14.025000 12.960000 14.345000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025000 13.400000 14.345000 13.720000 ;
      LAYER met4 ;
        RECT 14.025000 13.400000 14.345000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025000 13.840000 14.345000 14.160000 ;
      LAYER met4 ;
        RECT 14.025000 13.840000 14.345000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025000 14.280000 14.345000 14.600000 ;
      LAYER met4 ;
        RECT 14.025000 14.280000 14.345000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025000 14.720000 14.345000 15.040000 ;
      LAYER met4 ;
        RECT 14.025000 14.720000 14.345000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025000 15.160000 14.345000 15.480000 ;
      LAYER met4 ;
        RECT 14.025000 15.160000 14.345000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025000 15.600000 14.345000 15.920000 ;
      LAYER met4 ;
        RECT 14.025000 15.600000 14.345000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025000 16.040000 14.345000 16.360000 ;
      LAYER met4 ;
        RECT 14.025000 16.040000 14.345000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430000 12.960000 14.750000 13.280000 ;
      LAYER met4 ;
        RECT 14.430000 12.960000 14.750000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430000 13.400000 14.750000 13.720000 ;
      LAYER met4 ;
        RECT 14.430000 13.400000 14.750000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430000 13.840000 14.750000 14.160000 ;
      LAYER met4 ;
        RECT 14.430000 13.840000 14.750000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430000 14.280000 14.750000 14.600000 ;
      LAYER met4 ;
        RECT 14.430000 14.280000 14.750000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430000 14.720000 14.750000 15.040000 ;
      LAYER met4 ;
        RECT 14.430000 14.720000 14.750000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430000 15.160000 14.750000 15.480000 ;
      LAYER met4 ;
        RECT 14.430000 15.160000 14.750000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430000 15.600000 14.750000 15.920000 ;
      LAYER met4 ;
        RECT 14.430000 15.600000 14.750000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430000 16.040000 14.750000 16.360000 ;
      LAYER met4 ;
        RECT 14.430000 16.040000 14.750000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835000 12.960000 15.155000 13.280000 ;
      LAYER met4 ;
        RECT 14.835000 12.960000 15.155000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835000 13.400000 15.155000 13.720000 ;
      LAYER met4 ;
        RECT 14.835000 13.400000 15.155000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835000 13.840000 15.155000 14.160000 ;
      LAYER met4 ;
        RECT 14.835000 13.840000 15.155000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835000 14.280000 15.155000 14.600000 ;
      LAYER met4 ;
        RECT 14.835000 14.280000 15.155000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835000 14.720000 15.155000 15.040000 ;
      LAYER met4 ;
        RECT 14.835000 14.720000 15.155000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835000 15.160000 15.155000 15.480000 ;
      LAYER met4 ;
        RECT 14.835000 15.160000 15.155000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835000 15.600000 15.155000 15.920000 ;
      LAYER met4 ;
        RECT 14.835000 15.600000 15.155000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835000 16.040000 15.155000 16.360000 ;
      LAYER met4 ;
        RECT 14.835000 16.040000 15.155000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240000 12.960000 15.560000 13.280000 ;
      LAYER met4 ;
        RECT 15.240000 12.960000 15.560000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240000 13.400000 15.560000 13.720000 ;
      LAYER met4 ;
        RECT 15.240000 13.400000 15.560000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240000 13.840000 15.560000 14.160000 ;
      LAYER met4 ;
        RECT 15.240000 13.840000 15.560000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240000 14.280000 15.560000 14.600000 ;
      LAYER met4 ;
        RECT 15.240000 14.280000 15.560000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240000 14.720000 15.560000 15.040000 ;
      LAYER met4 ;
        RECT 15.240000 14.720000 15.560000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240000 15.160000 15.560000 15.480000 ;
      LAYER met4 ;
        RECT 15.240000 15.160000 15.560000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240000 15.600000 15.560000 15.920000 ;
      LAYER met4 ;
        RECT 15.240000 15.600000 15.560000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240000 16.040000 15.560000 16.360000 ;
      LAYER met4 ;
        RECT 15.240000 16.040000 15.560000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645000 12.960000 15.965000 13.280000 ;
      LAYER met4 ;
        RECT 15.645000 12.960000 15.965000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645000 13.400000 15.965000 13.720000 ;
      LAYER met4 ;
        RECT 15.645000 13.400000 15.965000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645000 13.840000 15.965000 14.160000 ;
      LAYER met4 ;
        RECT 15.645000 13.840000 15.965000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645000 14.280000 15.965000 14.600000 ;
      LAYER met4 ;
        RECT 15.645000 14.280000 15.965000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645000 14.720000 15.965000 15.040000 ;
      LAYER met4 ;
        RECT 15.645000 14.720000 15.965000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645000 15.160000 15.965000 15.480000 ;
      LAYER met4 ;
        RECT 15.645000 15.160000 15.965000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645000 15.600000 15.965000 15.920000 ;
      LAYER met4 ;
        RECT 15.645000 15.600000 15.965000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645000 16.040000 15.965000 16.360000 ;
      LAYER met4 ;
        RECT 15.645000 16.040000 15.965000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050000 12.960000 16.370000 13.280000 ;
      LAYER met4 ;
        RECT 16.050000 12.960000 16.370000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050000 13.400000 16.370000 13.720000 ;
      LAYER met4 ;
        RECT 16.050000 13.400000 16.370000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050000 13.840000 16.370000 14.160000 ;
      LAYER met4 ;
        RECT 16.050000 13.840000 16.370000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050000 14.280000 16.370000 14.600000 ;
      LAYER met4 ;
        RECT 16.050000 14.280000 16.370000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050000 14.720000 16.370000 15.040000 ;
      LAYER met4 ;
        RECT 16.050000 14.720000 16.370000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050000 15.160000 16.370000 15.480000 ;
      LAYER met4 ;
        RECT 16.050000 15.160000 16.370000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050000 15.600000 16.370000 15.920000 ;
      LAYER met4 ;
        RECT 16.050000 15.600000 16.370000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050000 16.040000 16.370000 16.360000 ;
      LAYER met4 ;
        RECT 16.050000 16.040000 16.370000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 12.960000 16.775000 13.280000 ;
      LAYER met4 ;
        RECT 16.455000 12.960000 16.775000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 13.400000 16.775000 13.720000 ;
      LAYER met4 ;
        RECT 16.455000 13.400000 16.775000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 13.840000 16.775000 14.160000 ;
      LAYER met4 ;
        RECT 16.455000 13.840000 16.775000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 14.280000 16.775000 14.600000 ;
      LAYER met4 ;
        RECT 16.455000 14.280000 16.775000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 14.720000 16.775000 15.040000 ;
      LAYER met4 ;
        RECT 16.455000 14.720000 16.775000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 15.160000 16.775000 15.480000 ;
      LAYER met4 ;
        RECT 16.455000 15.160000 16.775000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 15.600000 16.775000 15.920000 ;
      LAYER met4 ;
        RECT 16.455000 15.600000 16.775000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455000 16.040000 16.775000 16.360000 ;
      LAYER met4 ;
        RECT 16.455000 16.040000 16.775000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860000 12.960000 17.180000 13.280000 ;
      LAYER met4 ;
        RECT 16.860000 12.960000 17.180000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860000 13.400000 17.180000 13.720000 ;
      LAYER met4 ;
        RECT 16.860000 13.400000 17.180000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860000 13.840000 17.180000 14.160000 ;
      LAYER met4 ;
        RECT 16.860000 13.840000 17.180000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860000 14.280000 17.180000 14.600000 ;
      LAYER met4 ;
        RECT 16.860000 14.280000 17.180000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860000 14.720000 17.180000 15.040000 ;
      LAYER met4 ;
        RECT 16.860000 14.720000 17.180000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860000 15.160000 17.180000 15.480000 ;
      LAYER met4 ;
        RECT 16.860000 15.160000 17.180000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860000 15.600000 17.180000 15.920000 ;
      LAYER met4 ;
        RECT 16.860000 15.600000 17.180000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860000 16.040000 17.180000 16.360000 ;
      LAYER met4 ;
        RECT 16.860000 16.040000 17.180000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265000 12.960000 17.585000 13.280000 ;
      LAYER met4 ;
        RECT 17.265000 12.960000 17.585000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265000 13.400000 17.585000 13.720000 ;
      LAYER met4 ;
        RECT 17.265000 13.400000 17.585000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265000 13.840000 17.585000 14.160000 ;
      LAYER met4 ;
        RECT 17.265000 13.840000 17.585000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265000 14.280000 17.585000 14.600000 ;
      LAYER met4 ;
        RECT 17.265000 14.280000 17.585000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265000 14.720000 17.585000 15.040000 ;
      LAYER met4 ;
        RECT 17.265000 14.720000 17.585000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265000 15.160000 17.585000 15.480000 ;
      LAYER met4 ;
        RECT 17.265000 15.160000 17.585000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265000 15.600000 17.585000 15.920000 ;
      LAYER met4 ;
        RECT 17.265000 15.600000 17.585000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265000 16.040000 17.585000 16.360000 ;
      LAYER met4 ;
        RECT 17.265000 16.040000 17.585000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670000 12.960000 17.990000 13.280000 ;
      LAYER met4 ;
        RECT 17.670000 12.960000 17.990000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670000 13.400000 17.990000 13.720000 ;
      LAYER met4 ;
        RECT 17.670000 13.400000 17.990000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670000 13.840000 17.990000 14.160000 ;
      LAYER met4 ;
        RECT 17.670000 13.840000 17.990000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670000 14.280000 17.990000 14.600000 ;
      LAYER met4 ;
        RECT 17.670000 14.280000 17.990000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670000 14.720000 17.990000 15.040000 ;
      LAYER met4 ;
        RECT 17.670000 14.720000 17.990000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670000 15.160000 17.990000 15.480000 ;
      LAYER met4 ;
        RECT 17.670000 15.160000 17.990000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670000 15.600000 17.990000 15.920000 ;
      LAYER met4 ;
        RECT 17.670000 15.600000 17.990000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670000 16.040000 17.990000 16.360000 ;
      LAYER met4 ;
        RECT 17.670000 16.040000 17.990000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075000 12.960000 18.395000 13.280000 ;
      LAYER met4 ;
        RECT 18.075000 12.960000 18.395000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075000 13.400000 18.395000 13.720000 ;
      LAYER met4 ;
        RECT 18.075000 13.400000 18.395000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075000 13.840000 18.395000 14.160000 ;
      LAYER met4 ;
        RECT 18.075000 13.840000 18.395000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075000 14.280000 18.395000 14.600000 ;
      LAYER met4 ;
        RECT 18.075000 14.280000 18.395000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075000 14.720000 18.395000 15.040000 ;
      LAYER met4 ;
        RECT 18.075000 14.720000 18.395000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075000 15.160000 18.395000 15.480000 ;
      LAYER met4 ;
        RECT 18.075000 15.160000 18.395000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075000 15.600000 18.395000 15.920000 ;
      LAYER met4 ;
        RECT 18.075000 15.600000 18.395000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075000 16.040000 18.395000 16.360000 ;
      LAYER met4 ;
        RECT 18.075000 16.040000 18.395000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480000 12.960000 18.800000 13.280000 ;
      LAYER met4 ;
        RECT 18.480000 12.960000 18.800000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480000 13.400000 18.800000 13.720000 ;
      LAYER met4 ;
        RECT 18.480000 13.400000 18.800000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480000 13.840000 18.800000 14.160000 ;
      LAYER met4 ;
        RECT 18.480000 13.840000 18.800000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480000 14.280000 18.800000 14.600000 ;
      LAYER met4 ;
        RECT 18.480000 14.280000 18.800000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480000 14.720000 18.800000 15.040000 ;
      LAYER met4 ;
        RECT 18.480000 14.720000 18.800000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480000 15.160000 18.800000 15.480000 ;
      LAYER met4 ;
        RECT 18.480000 15.160000 18.800000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480000 15.600000 18.800000 15.920000 ;
      LAYER met4 ;
        RECT 18.480000 15.600000 18.800000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480000 16.040000 18.800000 16.360000 ;
      LAYER met4 ;
        RECT 18.480000 16.040000 18.800000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885000 12.960000 19.205000 13.280000 ;
      LAYER met4 ;
        RECT 18.885000 12.960000 19.205000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885000 13.400000 19.205000 13.720000 ;
      LAYER met4 ;
        RECT 18.885000 13.400000 19.205000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885000 13.840000 19.205000 14.160000 ;
      LAYER met4 ;
        RECT 18.885000 13.840000 19.205000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885000 14.280000 19.205000 14.600000 ;
      LAYER met4 ;
        RECT 18.885000 14.280000 19.205000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885000 14.720000 19.205000 15.040000 ;
      LAYER met4 ;
        RECT 18.885000 14.720000 19.205000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885000 15.160000 19.205000 15.480000 ;
      LAYER met4 ;
        RECT 18.885000 15.160000 19.205000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885000 15.600000 19.205000 15.920000 ;
      LAYER met4 ;
        RECT 18.885000 15.600000 19.205000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885000 16.040000 19.205000 16.360000 ;
      LAYER met4 ;
        RECT 18.885000 16.040000 19.205000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290000 12.960000 19.610000 13.280000 ;
      LAYER met4 ;
        RECT 19.290000 12.960000 19.610000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290000 13.400000 19.610000 13.720000 ;
      LAYER met4 ;
        RECT 19.290000 13.400000 19.610000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290000 13.840000 19.610000 14.160000 ;
      LAYER met4 ;
        RECT 19.290000 13.840000 19.610000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290000 14.280000 19.610000 14.600000 ;
      LAYER met4 ;
        RECT 19.290000 14.280000 19.610000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290000 14.720000 19.610000 15.040000 ;
      LAYER met4 ;
        RECT 19.290000 14.720000 19.610000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290000 15.160000 19.610000 15.480000 ;
      LAYER met4 ;
        RECT 19.290000 15.160000 19.610000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290000 15.600000 19.610000 15.920000 ;
      LAYER met4 ;
        RECT 19.290000 15.600000 19.610000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290000 16.040000 19.610000 16.360000 ;
      LAYER met4 ;
        RECT 19.290000 16.040000 19.610000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695000 12.960000 20.015000 13.280000 ;
      LAYER met4 ;
        RECT 19.695000 12.960000 20.015000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695000 13.400000 20.015000 13.720000 ;
      LAYER met4 ;
        RECT 19.695000 13.400000 20.015000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695000 13.840000 20.015000 14.160000 ;
      LAYER met4 ;
        RECT 19.695000 13.840000 20.015000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695000 14.280000 20.015000 14.600000 ;
      LAYER met4 ;
        RECT 19.695000 14.280000 20.015000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695000 14.720000 20.015000 15.040000 ;
      LAYER met4 ;
        RECT 19.695000 14.720000 20.015000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695000 15.160000 20.015000 15.480000 ;
      LAYER met4 ;
        RECT 19.695000 15.160000 20.015000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695000 15.600000 20.015000 15.920000 ;
      LAYER met4 ;
        RECT 19.695000 15.600000 20.015000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695000 16.040000 20.015000 16.360000 ;
      LAYER met4 ;
        RECT 19.695000 16.040000 20.015000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270000 12.960000 2.590000 13.280000 ;
      LAYER met4 ;
        RECT 2.270000 12.960000 2.590000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270000 13.400000 2.590000 13.720000 ;
      LAYER met4 ;
        RECT 2.270000 13.400000 2.590000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270000 13.840000 2.590000 14.160000 ;
      LAYER met4 ;
        RECT 2.270000 13.840000 2.590000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270000 14.280000 2.590000 14.600000 ;
      LAYER met4 ;
        RECT 2.270000 14.280000 2.590000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270000 14.720000 2.590000 15.040000 ;
      LAYER met4 ;
        RECT 2.270000 14.720000 2.590000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270000 15.160000 2.590000 15.480000 ;
      LAYER met4 ;
        RECT 2.270000 15.160000 2.590000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270000 15.600000 2.590000 15.920000 ;
      LAYER met4 ;
        RECT 2.270000 15.600000 2.590000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270000 16.040000 2.590000 16.360000 ;
      LAYER met4 ;
        RECT 2.270000 16.040000 2.590000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680000 12.960000 3.000000 13.280000 ;
      LAYER met4 ;
        RECT 2.680000 12.960000 3.000000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680000 13.400000 3.000000 13.720000 ;
      LAYER met4 ;
        RECT 2.680000 13.400000 3.000000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680000 13.840000 3.000000 14.160000 ;
      LAYER met4 ;
        RECT 2.680000 13.840000 3.000000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680000 14.280000 3.000000 14.600000 ;
      LAYER met4 ;
        RECT 2.680000 14.280000 3.000000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680000 14.720000 3.000000 15.040000 ;
      LAYER met4 ;
        RECT 2.680000 14.720000 3.000000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680000 15.160000 3.000000 15.480000 ;
      LAYER met4 ;
        RECT 2.680000 15.160000 3.000000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680000 15.600000 3.000000 15.920000 ;
      LAYER met4 ;
        RECT 2.680000 15.600000 3.000000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680000 16.040000 3.000000 16.360000 ;
      LAYER met4 ;
        RECT 2.680000 16.040000 3.000000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100000 12.960000 20.420000 13.280000 ;
      LAYER met4 ;
        RECT 20.100000 12.960000 20.420000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100000 13.400000 20.420000 13.720000 ;
      LAYER met4 ;
        RECT 20.100000 13.400000 20.420000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100000 13.840000 20.420000 14.160000 ;
      LAYER met4 ;
        RECT 20.100000 13.840000 20.420000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100000 14.280000 20.420000 14.600000 ;
      LAYER met4 ;
        RECT 20.100000 14.280000 20.420000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100000 14.720000 20.420000 15.040000 ;
      LAYER met4 ;
        RECT 20.100000 14.720000 20.420000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100000 15.160000 20.420000 15.480000 ;
      LAYER met4 ;
        RECT 20.100000 15.160000 20.420000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100000 15.600000 20.420000 15.920000 ;
      LAYER met4 ;
        RECT 20.100000 15.600000 20.420000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100000 16.040000 20.420000 16.360000 ;
      LAYER met4 ;
        RECT 20.100000 16.040000 20.420000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505000 12.960000 20.825000 13.280000 ;
      LAYER met4 ;
        RECT 20.505000 12.960000 20.825000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505000 13.400000 20.825000 13.720000 ;
      LAYER met4 ;
        RECT 20.505000 13.400000 20.825000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505000 13.840000 20.825000 14.160000 ;
      LAYER met4 ;
        RECT 20.505000 13.840000 20.825000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505000 14.280000 20.825000 14.600000 ;
      LAYER met4 ;
        RECT 20.505000 14.280000 20.825000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505000 14.720000 20.825000 15.040000 ;
      LAYER met4 ;
        RECT 20.505000 14.720000 20.825000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505000 15.160000 20.825000 15.480000 ;
      LAYER met4 ;
        RECT 20.505000 15.160000 20.825000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505000 15.600000 20.825000 15.920000 ;
      LAYER met4 ;
        RECT 20.505000 15.600000 20.825000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505000 16.040000 20.825000 16.360000 ;
      LAYER met4 ;
        RECT 20.505000 16.040000 20.825000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910000 12.960000 21.230000 13.280000 ;
      LAYER met4 ;
        RECT 20.910000 12.960000 21.230000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910000 13.400000 21.230000 13.720000 ;
      LAYER met4 ;
        RECT 20.910000 13.400000 21.230000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910000 13.840000 21.230000 14.160000 ;
      LAYER met4 ;
        RECT 20.910000 13.840000 21.230000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910000 14.280000 21.230000 14.600000 ;
      LAYER met4 ;
        RECT 20.910000 14.280000 21.230000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910000 14.720000 21.230000 15.040000 ;
      LAYER met4 ;
        RECT 20.910000 14.720000 21.230000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910000 15.160000 21.230000 15.480000 ;
      LAYER met4 ;
        RECT 20.910000 15.160000 21.230000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910000 15.600000 21.230000 15.920000 ;
      LAYER met4 ;
        RECT 20.910000 15.600000 21.230000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910000 16.040000 21.230000 16.360000 ;
      LAYER met4 ;
        RECT 20.910000 16.040000 21.230000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315000 12.960000 21.635000 13.280000 ;
      LAYER met4 ;
        RECT 21.315000 12.960000 21.635000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315000 13.400000 21.635000 13.720000 ;
      LAYER met4 ;
        RECT 21.315000 13.400000 21.635000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315000 13.840000 21.635000 14.160000 ;
      LAYER met4 ;
        RECT 21.315000 13.840000 21.635000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315000 14.280000 21.635000 14.600000 ;
      LAYER met4 ;
        RECT 21.315000 14.280000 21.635000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315000 14.720000 21.635000 15.040000 ;
      LAYER met4 ;
        RECT 21.315000 14.720000 21.635000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315000 15.160000 21.635000 15.480000 ;
      LAYER met4 ;
        RECT 21.315000 15.160000 21.635000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315000 15.600000 21.635000 15.920000 ;
      LAYER met4 ;
        RECT 21.315000 15.600000 21.635000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315000 16.040000 21.635000 16.360000 ;
      LAYER met4 ;
        RECT 21.315000 16.040000 21.635000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720000 12.960000 22.040000 13.280000 ;
      LAYER met4 ;
        RECT 21.720000 12.960000 22.040000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720000 13.400000 22.040000 13.720000 ;
      LAYER met4 ;
        RECT 21.720000 13.400000 22.040000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720000 13.840000 22.040000 14.160000 ;
      LAYER met4 ;
        RECT 21.720000 13.840000 22.040000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720000 14.280000 22.040000 14.600000 ;
      LAYER met4 ;
        RECT 21.720000 14.280000 22.040000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720000 14.720000 22.040000 15.040000 ;
      LAYER met4 ;
        RECT 21.720000 14.720000 22.040000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720000 15.160000 22.040000 15.480000 ;
      LAYER met4 ;
        RECT 21.720000 15.160000 22.040000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720000 15.600000 22.040000 15.920000 ;
      LAYER met4 ;
        RECT 21.720000 15.600000 22.040000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720000 16.040000 22.040000 16.360000 ;
      LAYER met4 ;
        RECT 21.720000 16.040000 22.040000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125000 12.960000 22.445000 13.280000 ;
      LAYER met4 ;
        RECT 22.125000 12.960000 22.445000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125000 13.400000 22.445000 13.720000 ;
      LAYER met4 ;
        RECT 22.125000 13.400000 22.445000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125000 13.840000 22.445000 14.160000 ;
      LAYER met4 ;
        RECT 22.125000 13.840000 22.445000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125000 14.280000 22.445000 14.600000 ;
      LAYER met4 ;
        RECT 22.125000 14.280000 22.445000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125000 14.720000 22.445000 15.040000 ;
      LAYER met4 ;
        RECT 22.125000 14.720000 22.445000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125000 15.160000 22.445000 15.480000 ;
      LAYER met4 ;
        RECT 22.125000 15.160000 22.445000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125000 15.600000 22.445000 15.920000 ;
      LAYER met4 ;
        RECT 22.125000 15.600000 22.445000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125000 16.040000 22.445000 16.360000 ;
      LAYER met4 ;
        RECT 22.125000 16.040000 22.445000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530000 12.960000 22.850000 13.280000 ;
      LAYER met4 ;
        RECT 22.530000 12.960000 22.850000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530000 13.400000 22.850000 13.720000 ;
      LAYER met4 ;
        RECT 22.530000 13.400000 22.850000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530000 13.840000 22.850000 14.160000 ;
      LAYER met4 ;
        RECT 22.530000 13.840000 22.850000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530000 14.280000 22.850000 14.600000 ;
      LAYER met4 ;
        RECT 22.530000 14.280000 22.850000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530000 14.720000 22.850000 15.040000 ;
      LAYER met4 ;
        RECT 22.530000 14.720000 22.850000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530000 15.160000 22.850000 15.480000 ;
      LAYER met4 ;
        RECT 22.530000 15.160000 22.850000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530000 15.600000 22.850000 15.920000 ;
      LAYER met4 ;
        RECT 22.530000 15.600000 22.850000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530000 16.040000 22.850000 16.360000 ;
      LAYER met4 ;
        RECT 22.530000 16.040000 22.850000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935000 12.960000 23.255000 13.280000 ;
      LAYER met4 ;
        RECT 22.935000 12.960000 23.255000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935000 13.400000 23.255000 13.720000 ;
      LAYER met4 ;
        RECT 22.935000 13.400000 23.255000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935000 13.840000 23.255000 14.160000 ;
      LAYER met4 ;
        RECT 22.935000 13.840000 23.255000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935000 14.280000 23.255000 14.600000 ;
      LAYER met4 ;
        RECT 22.935000 14.280000 23.255000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935000 14.720000 23.255000 15.040000 ;
      LAYER met4 ;
        RECT 22.935000 14.720000 23.255000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935000 15.160000 23.255000 15.480000 ;
      LAYER met4 ;
        RECT 22.935000 15.160000 23.255000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935000 15.600000 23.255000 15.920000 ;
      LAYER met4 ;
        RECT 22.935000 15.600000 23.255000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935000 16.040000 23.255000 16.360000 ;
      LAYER met4 ;
        RECT 22.935000 16.040000 23.255000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340000 12.960000 23.660000 13.280000 ;
      LAYER met4 ;
        RECT 23.340000 12.960000 23.660000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340000 13.400000 23.660000 13.720000 ;
      LAYER met4 ;
        RECT 23.340000 13.400000 23.660000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340000 13.840000 23.660000 14.160000 ;
      LAYER met4 ;
        RECT 23.340000 13.840000 23.660000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340000 14.280000 23.660000 14.600000 ;
      LAYER met4 ;
        RECT 23.340000 14.280000 23.660000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340000 14.720000 23.660000 15.040000 ;
      LAYER met4 ;
        RECT 23.340000 14.720000 23.660000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340000 15.160000 23.660000 15.480000 ;
      LAYER met4 ;
        RECT 23.340000 15.160000 23.660000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340000 15.600000 23.660000 15.920000 ;
      LAYER met4 ;
        RECT 23.340000 15.600000 23.660000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340000 16.040000 23.660000 16.360000 ;
      LAYER met4 ;
        RECT 23.340000 16.040000 23.660000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 12.960000 24.065000 13.280000 ;
      LAYER met4 ;
        RECT 23.745000 12.960000 24.065000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 13.400000 24.065000 13.720000 ;
      LAYER met4 ;
        RECT 23.745000 13.400000 24.065000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 13.840000 24.065000 14.160000 ;
      LAYER met4 ;
        RECT 23.745000 13.840000 24.065000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 14.280000 24.065000 14.600000 ;
      LAYER met4 ;
        RECT 23.745000 14.280000 24.065000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 14.720000 24.065000 15.040000 ;
      LAYER met4 ;
        RECT 23.745000 14.720000 24.065000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 15.160000 24.065000 15.480000 ;
      LAYER met4 ;
        RECT 23.745000 15.160000 24.065000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 15.600000 24.065000 15.920000 ;
      LAYER met4 ;
        RECT 23.745000 15.600000 24.065000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745000 16.040000 24.065000 16.360000 ;
      LAYER met4 ;
        RECT 23.745000 16.040000 24.065000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 12.960000 24.470000 13.280000 ;
      LAYER met4 ;
        RECT 24.150000 12.960000 24.470000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 13.400000 24.470000 13.720000 ;
      LAYER met4 ;
        RECT 24.150000 13.400000 24.470000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 13.840000 24.470000 14.160000 ;
      LAYER met4 ;
        RECT 24.150000 13.840000 24.470000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 14.280000 24.470000 14.600000 ;
      LAYER met4 ;
        RECT 24.150000 14.280000 24.470000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 14.720000 24.470000 15.040000 ;
      LAYER met4 ;
        RECT 24.150000 14.720000 24.470000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 15.160000 24.470000 15.480000 ;
      LAYER met4 ;
        RECT 24.150000 15.160000 24.470000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 15.600000 24.470000 15.920000 ;
      LAYER met4 ;
        RECT 24.150000 15.600000 24.470000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150000 16.040000 24.470000 16.360000 ;
      LAYER met4 ;
        RECT 24.150000 16.040000 24.470000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090000 12.960000 3.410000 13.280000 ;
      LAYER met4 ;
        RECT 3.090000 12.960000 3.410000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090000 13.400000 3.410000 13.720000 ;
      LAYER met4 ;
        RECT 3.090000 13.400000 3.410000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090000 13.840000 3.410000 14.160000 ;
      LAYER met4 ;
        RECT 3.090000 13.840000 3.410000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090000 14.280000 3.410000 14.600000 ;
      LAYER met4 ;
        RECT 3.090000 14.280000 3.410000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090000 14.720000 3.410000 15.040000 ;
      LAYER met4 ;
        RECT 3.090000 14.720000 3.410000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090000 15.160000 3.410000 15.480000 ;
      LAYER met4 ;
        RECT 3.090000 15.160000 3.410000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090000 15.600000 3.410000 15.920000 ;
      LAYER met4 ;
        RECT 3.090000 15.600000 3.410000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090000 16.040000 3.410000 16.360000 ;
      LAYER met4 ;
        RECT 3.090000 16.040000 3.410000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495000 12.960000 3.815000 13.280000 ;
      LAYER met4 ;
        RECT 3.495000 12.960000 3.815000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495000 13.400000 3.815000 13.720000 ;
      LAYER met4 ;
        RECT 3.495000 13.400000 3.815000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495000 13.840000 3.815000 14.160000 ;
      LAYER met4 ;
        RECT 3.495000 13.840000 3.815000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495000 14.280000 3.815000 14.600000 ;
      LAYER met4 ;
        RECT 3.495000 14.280000 3.815000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495000 14.720000 3.815000 15.040000 ;
      LAYER met4 ;
        RECT 3.495000 14.720000 3.815000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495000 15.160000 3.815000 15.480000 ;
      LAYER met4 ;
        RECT 3.495000 15.160000 3.815000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495000 15.600000 3.815000 15.920000 ;
      LAYER met4 ;
        RECT 3.495000 15.600000 3.815000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495000 16.040000 3.815000 16.360000 ;
      LAYER met4 ;
        RECT 3.495000 16.040000 3.815000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900000 12.960000 4.220000 13.280000 ;
      LAYER met4 ;
        RECT 3.900000 12.960000 4.220000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900000 13.400000 4.220000 13.720000 ;
      LAYER met4 ;
        RECT 3.900000 13.400000 4.220000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900000 13.840000 4.220000 14.160000 ;
      LAYER met4 ;
        RECT 3.900000 13.840000 4.220000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900000 14.280000 4.220000 14.600000 ;
      LAYER met4 ;
        RECT 3.900000 14.280000 4.220000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900000 14.720000 4.220000 15.040000 ;
      LAYER met4 ;
        RECT 3.900000 14.720000 4.220000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900000 15.160000 4.220000 15.480000 ;
      LAYER met4 ;
        RECT 3.900000 15.160000 4.220000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900000 15.600000 4.220000 15.920000 ;
      LAYER met4 ;
        RECT 3.900000 15.600000 4.220000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900000 16.040000 4.220000 16.360000 ;
      LAYER met4 ;
        RECT 3.900000 16.040000 4.220000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305000 12.960000 4.625000 13.280000 ;
      LAYER met4 ;
        RECT 4.305000 12.960000 4.625000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305000 13.400000 4.625000 13.720000 ;
      LAYER met4 ;
        RECT 4.305000 13.400000 4.625000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305000 13.840000 4.625000 14.160000 ;
      LAYER met4 ;
        RECT 4.305000 13.840000 4.625000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305000 14.280000 4.625000 14.600000 ;
      LAYER met4 ;
        RECT 4.305000 14.280000 4.625000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305000 14.720000 4.625000 15.040000 ;
      LAYER met4 ;
        RECT 4.305000 14.720000 4.625000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305000 15.160000 4.625000 15.480000 ;
      LAYER met4 ;
        RECT 4.305000 15.160000 4.625000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305000 15.600000 4.625000 15.920000 ;
      LAYER met4 ;
        RECT 4.305000 15.600000 4.625000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305000 16.040000 4.625000 16.360000 ;
      LAYER met4 ;
        RECT 4.305000 16.040000 4.625000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710000 12.960000 5.030000 13.280000 ;
      LAYER met4 ;
        RECT 4.710000 12.960000 5.030000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710000 13.400000 5.030000 13.720000 ;
      LAYER met4 ;
        RECT 4.710000 13.400000 5.030000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710000 13.840000 5.030000 14.160000 ;
      LAYER met4 ;
        RECT 4.710000 13.840000 5.030000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710000 14.280000 5.030000 14.600000 ;
      LAYER met4 ;
        RECT 4.710000 14.280000 5.030000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710000 14.720000 5.030000 15.040000 ;
      LAYER met4 ;
        RECT 4.710000 14.720000 5.030000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710000 15.160000 5.030000 15.480000 ;
      LAYER met4 ;
        RECT 4.710000 15.160000 5.030000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710000 15.600000 5.030000 15.920000 ;
      LAYER met4 ;
        RECT 4.710000 15.600000 5.030000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710000 16.040000 5.030000 16.360000 ;
      LAYER met4 ;
        RECT 4.710000 16.040000 5.030000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115000 12.960000 5.435000 13.280000 ;
      LAYER met4 ;
        RECT 5.115000 12.960000 5.435000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115000 13.400000 5.435000 13.720000 ;
      LAYER met4 ;
        RECT 5.115000 13.400000 5.435000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115000 13.840000 5.435000 14.160000 ;
      LAYER met4 ;
        RECT 5.115000 13.840000 5.435000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115000 14.280000 5.435000 14.600000 ;
      LAYER met4 ;
        RECT 5.115000 14.280000 5.435000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115000 14.720000 5.435000 15.040000 ;
      LAYER met4 ;
        RECT 5.115000 14.720000 5.435000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115000 15.160000 5.435000 15.480000 ;
      LAYER met4 ;
        RECT 5.115000 15.160000 5.435000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115000 15.600000 5.435000 15.920000 ;
      LAYER met4 ;
        RECT 5.115000 15.600000 5.435000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115000 16.040000 5.435000 16.360000 ;
      LAYER met4 ;
        RECT 5.115000 16.040000 5.435000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520000 12.960000 5.840000 13.280000 ;
      LAYER met4 ;
        RECT 5.520000 12.960000 5.840000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520000 13.400000 5.840000 13.720000 ;
      LAYER met4 ;
        RECT 5.520000 13.400000 5.840000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520000 13.840000 5.840000 14.160000 ;
      LAYER met4 ;
        RECT 5.520000 13.840000 5.840000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520000 14.280000 5.840000 14.600000 ;
      LAYER met4 ;
        RECT 5.520000 14.280000 5.840000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520000 14.720000 5.840000 15.040000 ;
      LAYER met4 ;
        RECT 5.520000 14.720000 5.840000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520000 15.160000 5.840000 15.480000 ;
      LAYER met4 ;
        RECT 5.520000 15.160000 5.840000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520000 15.600000 5.840000 15.920000 ;
      LAYER met4 ;
        RECT 5.520000 15.600000 5.840000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520000 16.040000 5.840000 16.360000 ;
      LAYER met4 ;
        RECT 5.520000 16.040000 5.840000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925000 12.960000 6.245000 13.280000 ;
      LAYER met4 ;
        RECT 5.925000 12.960000 6.245000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925000 13.400000 6.245000 13.720000 ;
      LAYER met4 ;
        RECT 5.925000 13.400000 6.245000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925000 13.840000 6.245000 14.160000 ;
      LAYER met4 ;
        RECT 5.925000 13.840000 6.245000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925000 14.280000 6.245000 14.600000 ;
      LAYER met4 ;
        RECT 5.925000 14.280000 6.245000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925000 14.720000 6.245000 15.040000 ;
      LAYER met4 ;
        RECT 5.925000 14.720000 6.245000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925000 15.160000 6.245000 15.480000 ;
      LAYER met4 ;
        RECT 5.925000 15.160000 6.245000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925000 15.600000 6.245000 15.920000 ;
      LAYER met4 ;
        RECT 5.925000 15.600000 6.245000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925000 16.040000 6.245000 16.360000 ;
      LAYER met4 ;
        RECT 5.925000 16.040000 6.245000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 12.960000 51.105000 13.280000 ;
      LAYER met4 ;
        RECT 50.785000 12.960000 51.105000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 13.400000 51.105000 13.720000 ;
      LAYER met4 ;
        RECT 50.785000 13.400000 51.105000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 13.840000 51.105000 14.160000 ;
      LAYER met4 ;
        RECT 50.785000 13.840000 51.105000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 14.280000 51.105000 14.600000 ;
      LAYER met4 ;
        RECT 50.785000 14.280000 51.105000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 14.720000 51.105000 15.040000 ;
      LAYER met4 ;
        RECT 50.785000 14.720000 51.105000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 15.160000 51.105000 15.480000 ;
      LAYER met4 ;
        RECT 50.785000 15.160000 51.105000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 15.600000 51.105000 15.920000 ;
      LAYER met4 ;
        RECT 50.785000 15.600000 51.105000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.785000 16.040000 51.105000 16.360000 ;
      LAYER met4 ;
        RECT 50.785000 16.040000 51.105000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 12.960000 51.515000 13.280000 ;
      LAYER met4 ;
        RECT 51.195000 12.960000 51.515000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 13.400000 51.515000 13.720000 ;
      LAYER met4 ;
        RECT 51.195000 13.400000 51.515000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 13.840000 51.515000 14.160000 ;
      LAYER met4 ;
        RECT 51.195000 13.840000 51.515000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 14.280000 51.515000 14.600000 ;
      LAYER met4 ;
        RECT 51.195000 14.280000 51.515000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 14.720000 51.515000 15.040000 ;
      LAYER met4 ;
        RECT 51.195000 14.720000 51.515000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 15.160000 51.515000 15.480000 ;
      LAYER met4 ;
        RECT 51.195000 15.160000 51.515000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 15.600000 51.515000 15.920000 ;
      LAYER met4 ;
        RECT 51.195000 15.600000 51.515000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.195000 16.040000 51.515000 16.360000 ;
      LAYER met4 ;
        RECT 51.195000 16.040000 51.515000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 12.960000 51.925000 13.280000 ;
      LAYER met4 ;
        RECT 51.605000 12.960000 51.925000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 13.400000 51.925000 13.720000 ;
      LAYER met4 ;
        RECT 51.605000 13.400000 51.925000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 13.840000 51.925000 14.160000 ;
      LAYER met4 ;
        RECT 51.605000 13.840000 51.925000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 14.280000 51.925000 14.600000 ;
      LAYER met4 ;
        RECT 51.605000 14.280000 51.925000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 14.720000 51.925000 15.040000 ;
      LAYER met4 ;
        RECT 51.605000 14.720000 51.925000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 15.160000 51.925000 15.480000 ;
      LAYER met4 ;
        RECT 51.605000 15.160000 51.925000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 15.600000 51.925000 15.920000 ;
      LAYER met4 ;
        RECT 51.605000 15.600000 51.925000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.605000 16.040000 51.925000 16.360000 ;
      LAYER met4 ;
        RECT 51.605000 16.040000 51.925000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 12.960000 52.335000 13.280000 ;
      LAYER met4 ;
        RECT 52.015000 12.960000 52.335000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 13.400000 52.335000 13.720000 ;
      LAYER met4 ;
        RECT 52.015000 13.400000 52.335000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 13.840000 52.335000 14.160000 ;
      LAYER met4 ;
        RECT 52.015000 13.840000 52.335000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 14.280000 52.335000 14.600000 ;
      LAYER met4 ;
        RECT 52.015000 14.280000 52.335000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 14.720000 52.335000 15.040000 ;
      LAYER met4 ;
        RECT 52.015000 14.720000 52.335000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 15.160000 52.335000 15.480000 ;
      LAYER met4 ;
        RECT 52.015000 15.160000 52.335000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 15.600000 52.335000 15.920000 ;
      LAYER met4 ;
        RECT 52.015000 15.600000 52.335000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.015000 16.040000 52.335000 16.360000 ;
      LAYER met4 ;
        RECT 52.015000 16.040000 52.335000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 12.960000 52.745000 13.280000 ;
      LAYER met4 ;
        RECT 52.425000 12.960000 52.745000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 13.400000 52.745000 13.720000 ;
      LAYER met4 ;
        RECT 52.425000 13.400000 52.745000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 13.840000 52.745000 14.160000 ;
      LAYER met4 ;
        RECT 52.425000 13.840000 52.745000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 14.280000 52.745000 14.600000 ;
      LAYER met4 ;
        RECT 52.425000 14.280000 52.745000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 14.720000 52.745000 15.040000 ;
      LAYER met4 ;
        RECT 52.425000 14.720000 52.745000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 15.160000 52.745000 15.480000 ;
      LAYER met4 ;
        RECT 52.425000 15.160000 52.745000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 15.600000 52.745000 15.920000 ;
      LAYER met4 ;
        RECT 52.425000 15.600000 52.745000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.425000 16.040000 52.745000 16.360000 ;
      LAYER met4 ;
        RECT 52.425000 16.040000 52.745000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 12.960000 53.155000 13.280000 ;
      LAYER met4 ;
        RECT 52.835000 12.960000 53.155000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 13.400000 53.155000 13.720000 ;
      LAYER met4 ;
        RECT 52.835000 13.400000 53.155000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 13.840000 53.155000 14.160000 ;
      LAYER met4 ;
        RECT 52.835000 13.840000 53.155000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 14.280000 53.155000 14.600000 ;
      LAYER met4 ;
        RECT 52.835000 14.280000 53.155000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 14.720000 53.155000 15.040000 ;
      LAYER met4 ;
        RECT 52.835000 14.720000 53.155000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 15.160000 53.155000 15.480000 ;
      LAYER met4 ;
        RECT 52.835000 15.160000 53.155000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 15.600000 53.155000 15.920000 ;
      LAYER met4 ;
        RECT 52.835000 15.600000 53.155000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.835000 16.040000 53.155000 16.360000 ;
      LAYER met4 ;
        RECT 52.835000 16.040000 53.155000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 12.960000 53.565000 13.280000 ;
      LAYER met4 ;
        RECT 53.245000 12.960000 53.565000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 13.400000 53.565000 13.720000 ;
      LAYER met4 ;
        RECT 53.245000 13.400000 53.565000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 13.840000 53.565000 14.160000 ;
      LAYER met4 ;
        RECT 53.245000 13.840000 53.565000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 14.280000 53.565000 14.600000 ;
      LAYER met4 ;
        RECT 53.245000 14.280000 53.565000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 14.720000 53.565000 15.040000 ;
      LAYER met4 ;
        RECT 53.245000 14.720000 53.565000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 15.160000 53.565000 15.480000 ;
      LAYER met4 ;
        RECT 53.245000 15.160000 53.565000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 15.600000 53.565000 15.920000 ;
      LAYER met4 ;
        RECT 53.245000 15.600000 53.565000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.245000 16.040000 53.565000 16.360000 ;
      LAYER met4 ;
        RECT 53.245000 16.040000 53.565000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 12.960000 53.970000 13.280000 ;
      LAYER met4 ;
        RECT 53.650000 12.960000 53.970000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 13.400000 53.970000 13.720000 ;
      LAYER met4 ;
        RECT 53.650000 13.400000 53.970000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 13.840000 53.970000 14.160000 ;
      LAYER met4 ;
        RECT 53.650000 13.840000 53.970000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 14.280000 53.970000 14.600000 ;
      LAYER met4 ;
        RECT 53.650000 14.280000 53.970000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 14.720000 53.970000 15.040000 ;
      LAYER met4 ;
        RECT 53.650000 14.720000 53.970000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 15.160000 53.970000 15.480000 ;
      LAYER met4 ;
        RECT 53.650000 15.160000 53.970000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 15.600000 53.970000 15.920000 ;
      LAYER met4 ;
        RECT 53.650000 15.600000 53.970000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.650000 16.040000 53.970000 16.360000 ;
      LAYER met4 ;
        RECT 53.650000 16.040000 53.970000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 12.960000 54.375000 13.280000 ;
      LAYER met4 ;
        RECT 54.055000 12.960000 54.375000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 13.400000 54.375000 13.720000 ;
      LAYER met4 ;
        RECT 54.055000 13.400000 54.375000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 13.840000 54.375000 14.160000 ;
      LAYER met4 ;
        RECT 54.055000 13.840000 54.375000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 14.280000 54.375000 14.600000 ;
      LAYER met4 ;
        RECT 54.055000 14.280000 54.375000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 14.720000 54.375000 15.040000 ;
      LAYER met4 ;
        RECT 54.055000 14.720000 54.375000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 15.160000 54.375000 15.480000 ;
      LAYER met4 ;
        RECT 54.055000 15.160000 54.375000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 15.600000 54.375000 15.920000 ;
      LAYER met4 ;
        RECT 54.055000 15.600000 54.375000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.055000 16.040000 54.375000 16.360000 ;
      LAYER met4 ;
        RECT 54.055000 16.040000 54.375000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 12.960000 54.780000 13.280000 ;
      LAYER met4 ;
        RECT 54.460000 12.960000 54.780000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 13.400000 54.780000 13.720000 ;
      LAYER met4 ;
        RECT 54.460000 13.400000 54.780000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 13.840000 54.780000 14.160000 ;
      LAYER met4 ;
        RECT 54.460000 13.840000 54.780000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 14.280000 54.780000 14.600000 ;
      LAYER met4 ;
        RECT 54.460000 14.280000 54.780000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 14.720000 54.780000 15.040000 ;
      LAYER met4 ;
        RECT 54.460000 14.720000 54.780000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 15.160000 54.780000 15.480000 ;
      LAYER met4 ;
        RECT 54.460000 15.160000 54.780000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 15.600000 54.780000 15.920000 ;
      LAYER met4 ;
        RECT 54.460000 15.600000 54.780000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.460000 16.040000 54.780000 16.360000 ;
      LAYER met4 ;
        RECT 54.460000 16.040000 54.780000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 12.960000 55.185000 13.280000 ;
      LAYER met4 ;
        RECT 54.865000 12.960000 55.185000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 13.400000 55.185000 13.720000 ;
      LAYER met4 ;
        RECT 54.865000 13.400000 55.185000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 13.840000 55.185000 14.160000 ;
      LAYER met4 ;
        RECT 54.865000 13.840000 55.185000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 14.280000 55.185000 14.600000 ;
      LAYER met4 ;
        RECT 54.865000 14.280000 55.185000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 14.720000 55.185000 15.040000 ;
      LAYER met4 ;
        RECT 54.865000 14.720000 55.185000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 15.160000 55.185000 15.480000 ;
      LAYER met4 ;
        RECT 54.865000 15.160000 55.185000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 15.600000 55.185000 15.920000 ;
      LAYER met4 ;
        RECT 54.865000 15.600000 55.185000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.865000 16.040000 55.185000 16.360000 ;
      LAYER met4 ;
        RECT 54.865000 16.040000 55.185000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 12.960000 55.590000 13.280000 ;
      LAYER met4 ;
        RECT 55.270000 12.960000 55.590000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 13.400000 55.590000 13.720000 ;
      LAYER met4 ;
        RECT 55.270000 13.400000 55.590000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 13.840000 55.590000 14.160000 ;
      LAYER met4 ;
        RECT 55.270000 13.840000 55.590000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 14.280000 55.590000 14.600000 ;
      LAYER met4 ;
        RECT 55.270000 14.280000 55.590000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 14.720000 55.590000 15.040000 ;
      LAYER met4 ;
        RECT 55.270000 14.720000 55.590000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 15.160000 55.590000 15.480000 ;
      LAYER met4 ;
        RECT 55.270000 15.160000 55.590000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 15.600000 55.590000 15.920000 ;
      LAYER met4 ;
        RECT 55.270000 15.600000 55.590000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.270000 16.040000 55.590000 16.360000 ;
      LAYER met4 ;
        RECT 55.270000 16.040000 55.590000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 12.960000 55.995000 13.280000 ;
      LAYER met4 ;
        RECT 55.675000 12.960000 55.995000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 13.400000 55.995000 13.720000 ;
      LAYER met4 ;
        RECT 55.675000 13.400000 55.995000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 13.840000 55.995000 14.160000 ;
      LAYER met4 ;
        RECT 55.675000 13.840000 55.995000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 14.280000 55.995000 14.600000 ;
      LAYER met4 ;
        RECT 55.675000 14.280000 55.995000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 14.720000 55.995000 15.040000 ;
      LAYER met4 ;
        RECT 55.675000 14.720000 55.995000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 15.160000 55.995000 15.480000 ;
      LAYER met4 ;
        RECT 55.675000 15.160000 55.995000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 15.600000 55.995000 15.920000 ;
      LAYER met4 ;
        RECT 55.675000 15.600000 55.995000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.675000 16.040000 55.995000 16.360000 ;
      LAYER met4 ;
        RECT 55.675000 16.040000 55.995000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 12.960000 56.400000 13.280000 ;
      LAYER met4 ;
        RECT 56.080000 12.960000 56.400000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 13.400000 56.400000 13.720000 ;
      LAYER met4 ;
        RECT 56.080000 13.400000 56.400000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 13.840000 56.400000 14.160000 ;
      LAYER met4 ;
        RECT 56.080000 13.840000 56.400000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 14.280000 56.400000 14.600000 ;
      LAYER met4 ;
        RECT 56.080000 14.280000 56.400000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 14.720000 56.400000 15.040000 ;
      LAYER met4 ;
        RECT 56.080000 14.720000 56.400000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 15.160000 56.400000 15.480000 ;
      LAYER met4 ;
        RECT 56.080000 15.160000 56.400000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 15.600000 56.400000 15.920000 ;
      LAYER met4 ;
        RECT 56.080000 15.600000 56.400000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.080000 16.040000 56.400000 16.360000 ;
      LAYER met4 ;
        RECT 56.080000 16.040000 56.400000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 12.960000 56.805000 13.280000 ;
      LAYER met4 ;
        RECT 56.485000 12.960000 56.805000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 13.400000 56.805000 13.720000 ;
      LAYER met4 ;
        RECT 56.485000 13.400000 56.805000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 13.840000 56.805000 14.160000 ;
      LAYER met4 ;
        RECT 56.485000 13.840000 56.805000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 14.280000 56.805000 14.600000 ;
      LAYER met4 ;
        RECT 56.485000 14.280000 56.805000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 14.720000 56.805000 15.040000 ;
      LAYER met4 ;
        RECT 56.485000 14.720000 56.805000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 15.160000 56.805000 15.480000 ;
      LAYER met4 ;
        RECT 56.485000 15.160000 56.805000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 15.600000 56.805000 15.920000 ;
      LAYER met4 ;
        RECT 56.485000 15.600000 56.805000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.485000 16.040000 56.805000 16.360000 ;
      LAYER met4 ;
        RECT 56.485000 16.040000 56.805000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 12.960000 57.210000 13.280000 ;
      LAYER met4 ;
        RECT 56.890000 12.960000 57.210000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 13.400000 57.210000 13.720000 ;
      LAYER met4 ;
        RECT 56.890000 13.400000 57.210000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 13.840000 57.210000 14.160000 ;
      LAYER met4 ;
        RECT 56.890000 13.840000 57.210000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 14.280000 57.210000 14.600000 ;
      LAYER met4 ;
        RECT 56.890000 14.280000 57.210000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 14.720000 57.210000 15.040000 ;
      LAYER met4 ;
        RECT 56.890000 14.720000 57.210000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 15.160000 57.210000 15.480000 ;
      LAYER met4 ;
        RECT 56.890000 15.160000 57.210000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 15.600000 57.210000 15.920000 ;
      LAYER met4 ;
        RECT 56.890000 15.600000 57.210000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.890000 16.040000 57.210000 16.360000 ;
      LAYER met4 ;
        RECT 56.890000 16.040000 57.210000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 12.960000 57.615000 13.280000 ;
      LAYER met4 ;
        RECT 57.295000 12.960000 57.615000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 13.400000 57.615000 13.720000 ;
      LAYER met4 ;
        RECT 57.295000 13.400000 57.615000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 13.840000 57.615000 14.160000 ;
      LAYER met4 ;
        RECT 57.295000 13.840000 57.615000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 14.280000 57.615000 14.600000 ;
      LAYER met4 ;
        RECT 57.295000 14.280000 57.615000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 14.720000 57.615000 15.040000 ;
      LAYER met4 ;
        RECT 57.295000 14.720000 57.615000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 15.160000 57.615000 15.480000 ;
      LAYER met4 ;
        RECT 57.295000 15.160000 57.615000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 15.600000 57.615000 15.920000 ;
      LAYER met4 ;
        RECT 57.295000 15.600000 57.615000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.295000 16.040000 57.615000 16.360000 ;
      LAYER met4 ;
        RECT 57.295000 16.040000 57.615000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 12.960000 58.020000 13.280000 ;
      LAYER met4 ;
        RECT 57.700000 12.960000 58.020000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 13.400000 58.020000 13.720000 ;
      LAYER met4 ;
        RECT 57.700000 13.400000 58.020000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 13.840000 58.020000 14.160000 ;
      LAYER met4 ;
        RECT 57.700000 13.840000 58.020000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 14.280000 58.020000 14.600000 ;
      LAYER met4 ;
        RECT 57.700000 14.280000 58.020000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 14.720000 58.020000 15.040000 ;
      LAYER met4 ;
        RECT 57.700000 14.720000 58.020000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 15.160000 58.020000 15.480000 ;
      LAYER met4 ;
        RECT 57.700000 15.160000 58.020000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 15.600000 58.020000 15.920000 ;
      LAYER met4 ;
        RECT 57.700000 15.600000 58.020000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.700000 16.040000 58.020000 16.360000 ;
      LAYER met4 ;
        RECT 57.700000 16.040000 58.020000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 12.960000 58.425000 13.280000 ;
      LAYER met4 ;
        RECT 58.105000 12.960000 58.425000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 13.400000 58.425000 13.720000 ;
      LAYER met4 ;
        RECT 58.105000 13.400000 58.425000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 13.840000 58.425000 14.160000 ;
      LAYER met4 ;
        RECT 58.105000 13.840000 58.425000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 14.280000 58.425000 14.600000 ;
      LAYER met4 ;
        RECT 58.105000 14.280000 58.425000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 14.720000 58.425000 15.040000 ;
      LAYER met4 ;
        RECT 58.105000 14.720000 58.425000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 15.160000 58.425000 15.480000 ;
      LAYER met4 ;
        RECT 58.105000 15.160000 58.425000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 15.600000 58.425000 15.920000 ;
      LAYER met4 ;
        RECT 58.105000 15.600000 58.425000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.105000 16.040000 58.425000 16.360000 ;
      LAYER met4 ;
        RECT 58.105000 16.040000 58.425000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 12.960000 58.830000 13.280000 ;
      LAYER met4 ;
        RECT 58.510000 12.960000 58.830000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 13.400000 58.830000 13.720000 ;
      LAYER met4 ;
        RECT 58.510000 13.400000 58.830000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 13.840000 58.830000 14.160000 ;
      LAYER met4 ;
        RECT 58.510000 13.840000 58.830000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 14.280000 58.830000 14.600000 ;
      LAYER met4 ;
        RECT 58.510000 14.280000 58.830000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 14.720000 58.830000 15.040000 ;
      LAYER met4 ;
        RECT 58.510000 14.720000 58.830000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 15.160000 58.830000 15.480000 ;
      LAYER met4 ;
        RECT 58.510000 15.160000 58.830000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 15.600000 58.830000 15.920000 ;
      LAYER met4 ;
        RECT 58.510000 15.600000 58.830000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.510000 16.040000 58.830000 16.360000 ;
      LAYER met4 ;
        RECT 58.510000 16.040000 58.830000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 12.960000 59.235000 13.280000 ;
      LAYER met4 ;
        RECT 58.915000 12.960000 59.235000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 13.400000 59.235000 13.720000 ;
      LAYER met4 ;
        RECT 58.915000 13.400000 59.235000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 13.840000 59.235000 14.160000 ;
      LAYER met4 ;
        RECT 58.915000 13.840000 59.235000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 14.280000 59.235000 14.600000 ;
      LAYER met4 ;
        RECT 58.915000 14.280000 59.235000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 14.720000 59.235000 15.040000 ;
      LAYER met4 ;
        RECT 58.915000 14.720000 59.235000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 15.160000 59.235000 15.480000 ;
      LAYER met4 ;
        RECT 58.915000 15.160000 59.235000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 15.600000 59.235000 15.920000 ;
      LAYER met4 ;
        RECT 58.915000 15.600000 59.235000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.915000 16.040000 59.235000 16.360000 ;
      LAYER met4 ;
        RECT 58.915000 16.040000 59.235000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 12.960000 59.640000 13.280000 ;
      LAYER met4 ;
        RECT 59.320000 12.960000 59.640000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 13.400000 59.640000 13.720000 ;
      LAYER met4 ;
        RECT 59.320000 13.400000 59.640000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 13.840000 59.640000 14.160000 ;
      LAYER met4 ;
        RECT 59.320000 13.840000 59.640000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 14.280000 59.640000 14.600000 ;
      LAYER met4 ;
        RECT 59.320000 14.280000 59.640000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 14.720000 59.640000 15.040000 ;
      LAYER met4 ;
        RECT 59.320000 14.720000 59.640000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 15.160000 59.640000 15.480000 ;
      LAYER met4 ;
        RECT 59.320000 15.160000 59.640000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 15.600000 59.640000 15.920000 ;
      LAYER met4 ;
        RECT 59.320000 15.600000 59.640000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.320000 16.040000 59.640000 16.360000 ;
      LAYER met4 ;
        RECT 59.320000 16.040000 59.640000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 12.960000 60.045000 13.280000 ;
      LAYER met4 ;
        RECT 59.725000 12.960000 60.045000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 13.400000 60.045000 13.720000 ;
      LAYER met4 ;
        RECT 59.725000 13.400000 60.045000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 13.840000 60.045000 14.160000 ;
      LAYER met4 ;
        RECT 59.725000 13.840000 60.045000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 14.280000 60.045000 14.600000 ;
      LAYER met4 ;
        RECT 59.725000 14.280000 60.045000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 14.720000 60.045000 15.040000 ;
      LAYER met4 ;
        RECT 59.725000 14.720000 60.045000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 15.160000 60.045000 15.480000 ;
      LAYER met4 ;
        RECT 59.725000 15.160000 60.045000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 15.600000 60.045000 15.920000 ;
      LAYER met4 ;
        RECT 59.725000 15.600000 60.045000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.725000 16.040000 60.045000 16.360000 ;
      LAYER met4 ;
        RECT 59.725000 16.040000 60.045000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330000 12.960000 6.650000 13.280000 ;
      LAYER met4 ;
        RECT 6.330000 12.960000 6.650000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330000 13.400000 6.650000 13.720000 ;
      LAYER met4 ;
        RECT 6.330000 13.400000 6.650000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330000 13.840000 6.650000 14.160000 ;
      LAYER met4 ;
        RECT 6.330000 13.840000 6.650000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330000 14.280000 6.650000 14.600000 ;
      LAYER met4 ;
        RECT 6.330000 14.280000 6.650000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330000 14.720000 6.650000 15.040000 ;
      LAYER met4 ;
        RECT 6.330000 14.720000 6.650000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330000 15.160000 6.650000 15.480000 ;
      LAYER met4 ;
        RECT 6.330000 15.160000 6.650000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330000 15.600000 6.650000 15.920000 ;
      LAYER met4 ;
        RECT 6.330000 15.600000 6.650000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330000 16.040000 6.650000 16.360000 ;
      LAYER met4 ;
        RECT 6.330000 16.040000 6.650000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735000 12.960000 7.055000 13.280000 ;
      LAYER met4 ;
        RECT 6.735000 12.960000 7.055000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735000 13.400000 7.055000 13.720000 ;
      LAYER met4 ;
        RECT 6.735000 13.400000 7.055000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735000 13.840000 7.055000 14.160000 ;
      LAYER met4 ;
        RECT 6.735000 13.840000 7.055000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735000 14.280000 7.055000 14.600000 ;
      LAYER met4 ;
        RECT 6.735000 14.280000 7.055000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735000 14.720000 7.055000 15.040000 ;
      LAYER met4 ;
        RECT 6.735000 14.720000 7.055000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735000 15.160000 7.055000 15.480000 ;
      LAYER met4 ;
        RECT 6.735000 15.160000 7.055000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735000 15.600000 7.055000 15.920000 ;
      LAYER met4 ;
        RECT 6.735000 15.600000 7.055000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735000 16.040000 7.055000 16.360000 ;
      LAYER met4 ;
        RECT 6.735000 16.040000 7.055000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 12.960000 60.450000 13.280000 ;
      LAYER met4 ;
        RECT 60.130000 12.960000 60.450000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 13.400000 60.450000 13.720000 ;
      LAYER met4 ;
        RECT 60.130000 13.400000 60.450000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 13.840000 60.450000 14.160000 ;
      LAYER met4 ;
        RECT 60.130000 13.840000 60.450000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 14.280000 60.450000 14.600000 ;
      LAYER met4 ;
        RECT 60.130000 14.280000 60.450000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 14.720000 60.450000 15.040000 ;
      LAYER met4 ;
        RECT 60.130000 14.720000 60.450000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 15.160000 60.450000 15.480000 ;
      LAYER met4 ;
        RECT 60.130000 15.160000 60.450000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 15.600000 60.450000 15.920000 ;
      LAYER met4 ;
        RECT 60.130000 15.600000 60.450000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.130000 16.040000 60.450000 16.360000 ;
      LAYER met4 ;
        RECT 60.130000 16.040000 60.450000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 12.960000 60.855000 13.280000 ;
      LAYER met4 ;
        RECT 60.535000 12.960000 60.855000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 13.400000 60.855000 13.720000 ;
      LAYER met4 ;
        RECT 60.535000 13.400000 60.855000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 13.840000 60.855000 14.160000 ;
      LAYER met4 ;
        RECT 60.535000 13.840000 60.855000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 14.280000 60.855000 14.600000 ;
      LAYER met4 ;
        RECT 60.535000 14.280000 60.855000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 14.720000 60.855000 15.040000 ;
      LAYER met4 ;
        RECT 60.535000 14.720000 60.855000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 15.160000 60.855000 15.480000 ;
      LAYER met4 ;
        RECT 60.535000 15.160000 60.855000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 15.600000 60.855000 15.920000 ;
      LAYER met4 ;
        RECT 60.535000 15.600000 60.855000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.535000 16.040000 60.855000 16.360000 ;
      LAYER met4 ;
        RECT 60.535000 16.040000 60.855000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 12.960000 61.260000 13.280000 ;
      LAYER met4 ;
        RECT 60.940000 12.960000 61.260000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 13.400000 61.260000 13.720000 ;
      LAYER met4 ;
        RECT 60.940000 13.400000 61.260000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 13.840000 61.260000 14.160000 ;
      LAYER met4 ;
        RECT 60.940000 13.840000 61.260000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 14.280000 61.260000 14.600000 ;
      LAYER met4 ;
        RECT 60.940000 14.280000 61.260000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 14.720000 61.260000 15.040000 ;
      LAYER met4 ;
        RECT 60.940000 14.720000 61.260000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 15.160000 61.260000 15.480000 ;
      LAYER met4 ;
        RECT 60.940000 15.160000 61.260000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 15.600000 61.260000 15.920000 ;
      LAYER met4 ;
        RECT 60.940000 15.600000 61.260000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.940000 16.040000 61.260000 16.360000 ;
      LAYER met4 ;
        RECT 60.940000 16.040000 61.260000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 12.960000 61.665000 13.280000 ;
      LAYER met4 ;
        RECT 61.345000 12.960000 61.665000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 13.400000 61.665000 13.720000 ;
      LAYER met4 ;
        RECT 61.345000 13.400000 61.665000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 13.840000 61.665000 14.160000 ;
      LAYER met4 ;
        RECT 61.345000 13.840000 61.665000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 14.280000 61.665000 14.600000 ;
      LAYER met4 ;
        RECT 61.345000 14.280000 61.665000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 14.720000 61.665000 15.040000 ;
      LAYER met4 ;
        RECT 61.345000 14.720000 61.665000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 15.160000 61.665000 15.480000 ;
      LAYER met4 ;
        RECT 61.345000 15.160000 61.665000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 15.600000 61.665000 15.920000 ;
      LAYER met4 ;
        RECT 61.345000 15.600000 61.665000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.345000 16.040000 61.665000 16.360000 ;
      LAYER met4 ;
        RECT 61.345000 16.040000 61.665000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 12.960000 62.070000 13.280000 ;
      LAYER met4 ;
        RECT 61.750000 12.960000 62.070000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 13.400000 62.070000 13.720000 ;
      LAYER met4 ;
        RECT 61.750000 13.400000 62.070000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 13.840000 62.070000 14.160000 ;
      LAYER met4 ;
        RECT 61.750000 13.840000 62.070000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 14.280000 62.070000 14.600000 ;
      LAYER met4 ;
        RECT 61.750000 14.280000 62.070000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 14.720000 62.070000 15.040000 ;
      LAYER met4 ;
        RECT 61.750000 14.720000 62.070000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 15.160000 62.070000 15.480000 ;
      LAYER met4 ;
        RECT 61.750000 15.160000 62.070000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 15.600000 62.070000 15.920000 ;
      LAYER met4 ;
        RECT 61.750000 15.600000 62.070000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.750000 16.040000 62.070000 16.360000 ;
      LAYER met4 ;
        RECT 61.750000 16.040000 62.070000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 12.960000 62.475000 13.280000 ;
      LAYER met4 ;
        RECT 62.155000 12.960000 62.475000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 13.400000 62.475000 13.720000 ;
      LAYER met4 ;
        RECT 62.155000 13.400000 62.475000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 13.840000 62.475000 14.160000 ;
      LAYER met4 ;
        RECT 62.155000 13.840000 62.475000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 14.280000 62.475000 14.600000 ;
      LAYER met4 ;
        RECT 62.155000 14.280000 62.475000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 14.720000 62.475000 15.040000 ;
      LAYER met4 ;
        RECT 62.155000 14.720000 62.475000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 15.160000 62.475000 15.480000 ;
      LAYER met4 ;
        RECT 62.155000 15.160000 62.475000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 15.600000 62.475000 15.920000 ;
      LAYER met4 ;
        RECT 62.155000 15.600000 62.475000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.155000 16.040000 62.475000 16.360000 ;
      LAYER met4 ;
        RECT 62.155000 16.040000 62.475000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 12.960000 62.880000 13.280000 ;
      LAYER met4 ;
        RECT 62.560000 12.960000 62.880000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 13.400000 62.880000 13.720000 ;
      LAYER met4 ;
        RECT 62.560000 13.400000 62.880000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 13.840000 62.880000 14.160000 ;
      LAYER met4 ;
        RECT 62.560000 13.840000 62.880000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 14.280000 62.880000 14.600000 ;
      LAYER met4 ;
        RECT 62.560000 14.280000 62.880000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 14.720000 62.880000 15.040000 ;
      LAYER met4 ;
        RECT 62.560000 14.720000 62.880000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 15.160000 62.880000 15.480000 ;
      LAYER met4 ;
        RECT 62.560000 15.160000 62.880000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 15.600000 62.880000 15.920000 ;
      LAYER met4 ;
        RECT 62.560000 15.600000 62.880000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.560000 16.040000 62.880000 16.360000 ;
      LAYER met4 ;
        RECT 62.560000 16.040000 62.880000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 12.960000 63.285000 13.280000 ;
      LAYER met4 ;
        RECT 62.965000 12.960000 63.285000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 13.400000 63.285000 13.720000 ;
      LAYER met4 ;
        RECT 62.965000 13.400000 63.285000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 13.840000 63.285000 14.160000 ;
      LAYER met4 ;
        RECT 62.965000 13.840000 63.285000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 14.280000 63.285000 14.600000 ;
      LAYER met4 ;
        RECT 62.965000 14.280000 63.285000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 14.720000 63.285000 15.040000 ;
      LAYER met4 ;
        RECT 62.965000 14.720000 63.285000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 15.160000 63.285000 15.480000 ;
      LAYER met4 ;
        RECT 62.965000 15.160000 63.285000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 15.600000 63.285000 15.920000 ;
      LAYER met4 ;
        RECT 62.965000 15.600000 63.285000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.965000 16.040000 63.285000 16.360000 ;
      LAYER met4 ;
        RECT 62.965000 16.040000 63.285000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 12.960000 63.690000 13.280000 ;
      LAYER met4 ;
        RECT 63.370000 12.960000 63.690000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 13.400000 63.690000 13.720000 ;
      LAYER met4 ;
        RECT 63.370000 13.400000 63.690000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 13.840000 63.690000 14.160000 ;
      LAYER met4 ;
        RECT 63.370000 13.840000 63.690000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 14.280000 63.690000 14.600000 ;
      LAYER met4 ;
        RECT 63.370000 14.280000 63.690000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 14.720000 63.690000 15.040000 ;
      LAYER met4 ;
        RECT 63.370000 14.720000 63.690000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 15.160000 63.690000 15.480000 ;
      LAYER met4 ;
        RECT 63.370000 15.160000 63.690000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 15.600000 63.690000 15.920000 ;
      LAYER met4 ;
        RECT 63.370000 15.600000 63.690000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370000 16.040000 63.690000 16.360000 ;
      LAYER met4 ;
        RECT 63.370000 16.040000 63.690000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 12.960000 64.095000 13.280000 ;
      LAYER met4 ;
        RECT 63.775000 12.960000 64.095000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 13.400000 64.095000 13.720000 ;
      LAYER met4 ;
        RECT 63.775000 13.400000 64.095000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 13.840000 64.095000 14.160000 ;
      LAYER met4 ;
        RECT 63.775000 13.840000 64.095000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 14.280000 64.095000 14.600000 ;
      LAYER met4 ;
        RECT 63.775000 14.280000 64.095000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 14.720000 64.095000 15.040000 ;
      LAYER met4 ;
        RECT 63.775000 14.720000 64.095000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 15.160000 64.095000 15.480000 ;
      LAYER met4 ;
        RECT 63.775000 15.160000 64.095000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 15.600000 64.095000 15.920000 ;
      LAYER met4 ;
        RECT 63.775000 15.600000 64.095000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.775000 16.040000 64.095000 16.360000 ;
      LAYER met4 ;
        RECT 63.775000 16.040000 64.095000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 12.960000 64.500000 13.280000 ;
      LAYER met4 ;
        RECT 64.180000 12.960000 64.500000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 13.400000 64.500000 13.720000 ;
      LAYER met4 ;
        RECT 64.180000 13.400000 64.500000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 13.840000 64.500000 14.160000 ;
      LAYER met4 ;
        RECT 64.180000 13.840000 64.500000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 14.280000 64.500000 14.600000 ;
      LAYER met4 ;
        RECT 64.180000 14.280000 64.500000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 14.720000 64.500000 15.040000 ;
      LAYER met4 ;
        RECT 64.180000 14.720000 64.500000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 15.160000 64.500000 15.480000 ;
      LAYER met4 ;
        RECT 64.180000 15.160000 64.500000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 15.600000 64.500000 15.920000 ;
      LAYER met4 ;
        RECT 64.180000 15.600000 64.500000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.180000 16.040000 64.500000 16.360000 ;
      LAYER met4 ;
        RECT 64.180000 16.040000 64.500000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 12.960000 64.905000 13.280000 ;
      LAYER met4 ;
        RECT 64.585000 12.960000 64.905000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 13.400000 64.905000 13.720000 ;
      LAYER met4 ;
        RECT 64.585000 13.400000 64.905000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 13.840000 64.905000 14.160000 ;
      LAYER met4 ;
        RECT 64.585000 13.840000 64.905000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 14.280000 64.905000 14.600000 ;
      LAYER met4 ;
        RECT 64.585000 14.280000 64.905000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 14.720000 64.905000 15.040000 ;
      LAYER met4 ;
        RECT 64.585000 14.720000 64.905000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 15.160000 64.905000 15.480000 ;
      LAYER met4 ;
        RECT 64.585000 15.160000 64.905000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 15.600000 64.905000 15.920000 ;
      LAYER met4 ;
        RECT 64.585000 15.600000 64.905000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.585000 16.040000 64.905000 16.360000 ;
      LAYER met4 ;
        RECT 64.585000 16.040000 64.905000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 12.960000 65.310000 13.280000 ;
      LAYER met4 ;
        RECT 64.990000 12.960000 65.310000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 13.400000 65.310000 13.720000 ;
      LAYER met4 ;
        RECT 64.990000 13.400000 65.310000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 13.840000 65.310000 14.160000 ;
      LAYER met4 ;
        RECT 64.990000 13.840000 65.310000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 14.280000 65.310000 14.600000 ;
      LAYER met4 ;
        RECT 64.990000 14.280000 65.310000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 14.720000 65.310000 15.040000 ;
      LAYER met4 ;
        RECT 64.990000 14.720000 65.310000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 15.160000 65.310000 15.480000 ;
      LAYER met4 ;
        RECT 64.990000 15.160000 65.310000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 15.600000 65.310000 15.920000 ;
      LAYER met4 ;
        RECT 64.990000 15.600000 65.310000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.990000 16.040000 65.310000 16.360000 ;
      LAYER met4 ;
        RECT 64.990000 16.040000 65.310000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 12.960000 65.715000 13.280000 ;
      LAYER met4 ;
        RECT 65.395000 12.960000 65.715000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 13.400000 65.715000 13.720000 ;
      LAYER met4 ;
        RECT 65.395000 13.400000 65.715000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 13.840000 65.715000 14.160000 ;
      LAYER met4 ;
        RECT 65.395000 13.840000 65.715000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 14.280000 65.715000 14.600000 ;
      LAYER met4 ;
        RECT 65.395000 14.280000 65.715000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 14.720000 65.715000 15.040000 ;
      LAYER met4 ;
        RECT 65.395000 14.720000 65.715000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 15.160000 65.715000 15.480000 ;
      LAYER met4 ;
        RECT 65.395000 15.160000 65.715000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 15.600000 65.715000 15.920000 ;
      LAYER met4 ;
        RECT 65.395000 15.600000 65.715000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.395000 16.040000 65.715000 16.360000 ;
      LAYER met4 ;
        RECT 65.395000 16.040000 65.715000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 12.960000 66.120000 13.280000 ;
      LAYER met4 ;
        RECT 65.800000 12.960000 66.120000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 13.400000 66.120000 13.720000 ;
      LAYER met4 ;
        RECT 65.800000 13.400000 66.120000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 13.840000 66.120000 14.160000 ;
      LAYER met4 ;
        RECT 65.800000 13.840000 66.120000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 14.280000 66.120000 14.600000 ;
      LAYER met4 ;
        RECT 65.800000 14.280000 66.120000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 14.720000 66.120000 15.040000 ;
      LAYER met4 ;
        RECT 65.800000 14.720000 66.120000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 15.160000 66.120000 15.480000 ;
      LAYER met4 ;
        RECT 65.800000 15.160000 66.120000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 15.600000 66.120000 15.920000 ;
      LAYER met4 ;
        RECT 65.800000 15.600000 66.120000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.800000 16.040000 66.120000 16.360000 ;
      LAYER met4 ;
        RECT 65.800000 16.040000 66.120000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 12.960000 66.525000 13.280000 ;
      LAYER met4 ;
        RECT 66.205000 12.960000 66.525000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 13.400000 66.525000 13.720000 ;
      LAYER met4 ;
        RECT 66.205000 13.400000 66.525000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 13.840000 66.525000 14.160000 ;
      LAYER met4 ;
        RECT 66.205000 13.840000 66.525000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 14.280000 66.525000 14.600000 ;
      LAYER met4 ;
        RECT 66.205000 14.280000 66.525000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 14.720000 66.525000 15.040000 ;
      LAYER met4 ;
        RECT 66.205000 14.720000 66.525000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 15.160000 66.525000 15.480000 ;
      LAYER met4 ;
        RECT 66.205000 15.160000 66.525000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 15.600000 66.525000 15.920000 ;
      LAYER met4 ;
        RECT 66.205000 15.600000 66.525000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.205000 16.040000 66.525000 16.360000 ;
      LAYER met4 ;
        RECT 66.205000 16.040000 66.525000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 12.960000 66.930000 13.280000 ;
      LAYER met4 ;
        RECT 66.610000 12.960000 66.930000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 13.400000 66.930000 13.720000 ;
      LAYER met4 ;
        RECT 66.610000 13.400000 66.930000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 13.840000 66.930000 14.160000 ;
      LAYER met4 ;
        RECT 66.610000 13.840000 66.930000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 14.280000 66.930000 14.600000 ;
      LAYER met4 ;
        RECT 66.610000 14.280000 66.930000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 14.720000 66.930000 15.040000 ;
      LAYER met4 ;
        RECT 66.610000 14.720000 66.930000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 15.160000 66.930000 15.480000 ;
      LAYER met4 ;
        RECT 66.610000 15.160000 66.930000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 15.600000 66.930000 15.920000 ;
      LAYER met4 ;
        RECT 66.610000 15.600000 66.930000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610000 16.040000 66.930000 16.360000 ;
      LAYER met4 ;
        RECT 66.610000 16.040000 66.930000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 12.960000 67.335000 13.280000 ;
      LAYER met4 ;
        RECT 67.015000 12.960000 67.335000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 13.400000 67.335000 13.720000 ;
      LAYER met4 ;
        RECT 67.015000 13.400000 67.335000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 13.840000 67.335000 14.160000 ;
      LAYER met4 ;
        RECT 67.015000 13.840000 67.335000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 14.280000 67.335000 14.600000 ;
      LAYER met4 ;
        RECT 67.015000 14.280000 67.335000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 14.720000 67.335000 15.040000 ;
      LAYER met4 ;
        RECT 67.015000 14.720000 67.335000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 15.160000 67.335000 15.480000 ;
      LAYER met4 ;
        RECT 67.015000 15.160000 67.335000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 15.600000 67.335000 15.920000 ;
      LAYER met4 ;
        RECT 67.015000 15.600000 67.335000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.015000 16.040000 67.335000 16.360000 ;
      LAYER met4 ;
        RECT 67.015000 16.040000 67.335000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 12.960000 67.740000 13.280000 ;
      LAYER met4 ;
        RECT 67.420000 12.960000 67.740000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 13.400000 67.740000 13.720000 ;
      LAYER met4 ;
        RECT 67.420000 13.400000 67.740000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 13.840000 67.740000 14.160000 ;
      LAYER met4 ;
        RECT 67.420000 13.840000 67.740000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 14.280000 67.740000 14.600000 ;
      LAYER met4 ;
        RECT 67.420000 14.280000 67.740000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 14.720000 67.740000 15.040000 ;
      LAYER met4 ;
        RECT 67.420000 14.720000 67.740000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 15.160000 67.740000 15.480000 ;
      LAYER met4 ;
        RECT 67.420000 15.160000 67.740000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 15.600000 67.740000 15.920000 ;
      LAYER met4 ;
        RECT 67.420000 15.600000 67.740000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.420000 16.040000 67.740000 16.360000 ;
      LAYER met4 ;
        RECT 67.420000 16.040000 67.740000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 12.960000 68.145000 13.280000 ;
      LAYER met4 ;
        RECT 67.825000 12.960000 68.145000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 13.400000 68.145000 13.720000 ;
      LAYER met4 ;
        RECT 67.825000 13.400000 68.145000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 13.840000 68.145000 14.160000 ;
      LAYER met4 ;
        RECT 67.825000 13.840000 68.145000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 14.280000 68.145000 14.600000 ;
      LAYER met4 ;
        RECT 67.825000 14.280000 68.145000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 14.720000 68.145000 15.040000 ;
      LAYER met4 ;
        RECT 67.825000 14.720000 68.145000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 15.160000 68.145000 15.480000 ;
      LAYER met4 ;
        RECT 67.825000 15.160000 68.145000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 15.600000 68.145000 15.920000 ;
      LAYER met4 ;
        RECT 67.825000 15.600000 68.145000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.825000 16.040000 68.145000 16.360000 ;
      LAYER met4 ;
        RECT 67.825000 16.040000 68.145000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 12.960000 68.550000 13.280000 ;
      LAYER met4 ;
        RECT 68.230000 12.960000 68.550000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 13.400000 68.550000 13.720000 ;
      LAYER met4 ;
        RECT 68.230000 13.400000 68.550000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 13.840000 68.550000 14.160000 ;
      LAYER met4 ;
        RECT 68.230000 13.840000 68.550000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 14.280000 68.550000 14.600000 ;
      LAYER met4 ;
        RECT 68.230000 14.280000 68.550000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 14.720000 68.550000 15.040000 ;
      LAYER met4 ;
        RECT 68.230000 14.720000 68.550000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 15.160000 68.550000 15.480000 ;
      LAYER met4 ;
        RECT 68.230000 15.160000 68.550000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 15.600000 68.550000 15.920000 ;
      LAYER met4 ;
        RECT 68.230000 15.600000 68.550000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.230000 16.040000 68.550000 16.360000 ;
      LAYER met4 ;
        RECT 68.230000 16.040000 68.550000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 12.960000 68.955000 13.280000 ;
      LAYER met4 ;
        RECT 68.635000 12.960000 68.955000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 13.400000 68.955000 13.720000 ;
      LAYER met4 ;
        RECT 68.635000 13.400000 68.955000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 13.840000 68.955000 14.160000 ;
      LAYER met4 ;
        RECT 68.635000 13.840000 68.955000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 14.280000 68.955000 14.600000 ;
      LAYER met4 ;
        RECT 68.635000 14.280000 68.955000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 14.720000 68.955000 15.040000 ;
      LAYER met4 ;
        RECT 68.635000 14.720000 68.955000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 15.160000 68.955000 15.480000 ;
      LAYER met4 ;
        RECT 68.635000 15.160000 68.955000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 15.600000 68.955000 15.920000 ;
      LAYER met4 ;
        RECT 68.635000 15.600000 68.955000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.635000 16.040000 68.955000 16.360000 ;
      LAYER met4 ;
        RECT 68.635000 16.040000 68.955000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 12.960000 69.360000 13.280000 ;
      LAYER met4 ;
        RECT 69.040000 12.960000 69.360000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 13.400000 69.360000 13.720000 ;
      LAYER met4 ;
        RECT 69.040000 13.400000 69.360000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 13.840000 69.360000 14.160000 ;
      LAYER met4 ;
        RECT 69.040000 13.840000 69.360000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 14.280000 69.360000 14.600000 ;
      LAYER met4 ;
        RECT 69.040000 14.280000 69.360000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 14.720000 69.360000 15.040000 ;
      LAYER met4 ;
        RECT 69.040000 14.720000 69.360000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 15.160000 69.360000 15.480000 ;
      LAYER met4 ;
        RECT 69.040000 15.160000 69.360000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 15.600000 69.360000 15.920000 ;
      LAYER met4 ;
        RECT 69.040000 15.600000 69.360000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.040000 16.040000 69.360000 16.360000 ;
      LAYER met4 ;
        RECT 69.040000 16.040000 69.360000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 12.960000 69.765000 13.280000 ;
      LAYER met4 ;
        RECT 69.445000 12.960000 69.765000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 13.400000 69.765000 13.720000 ;
      LAYER met4 ;
        RECT 69.445000 13.400000 69.765000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 13.840000 69.765000 14.160000 ;
      LAYER met4 ;
        RECT 69.445000 13.840000 69.765000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 14.280000 69.765000 14.600000 ;
      LAYER met4 ;
        RECT 69.445000 14.280000 69.765000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 14.720000 69.765000 15.040000 ;
      LAYER met4 ;
        RECT 69.445000 14.720000 69.765000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 15.160000 69.765000 15.480000 ;
      LAYER met4 ;
        RECT 69.445000 15.160000 69.765000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 15.600000 69.765000 15.920000 ;
      LAYER met4 ;
        RECT 69.445000 15.600000 69.765000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.445000 16.040000 69.765000 16.360000 ;
      LAYER met4 ;
        RECT 69.445000 16.040000 69.765000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 12.960000 70.170000 13.280000 ;
      LAYER met4 ;
        RECT 69.850000 12.960000 70.170000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 13.400000 70.170000 13.720000 ;
      LAYER met4 ;
        RECT 69.850000 13.400000 70.170000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 13.840000 70.170000 14.160000 ;
      LAYER met4 ;
        RECT 69.850000 13.840000 70.170000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 14.280000 70.170000 14.600000 ;
      LAYER met4 ;
        RECT 69.850000 14.280000 70.170000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 14.720000 70.170000 15.040000 ;
      LAYER met4 ;
        RECT 69.850000 14.720000 70.170000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 15.160000 70.170000 15.480000 ;
      LAYER met4 ;
        RECT 69.850000 15.160000 70.170000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 15.600000 70.170000 15.920000 ;
      LAYER met4 ;
        RECT 69.850000 15.600000 70.170000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.850000 16.040000 70.170000 16.360000 ;
      LAYER met4 ;
        RECT 69.850000 16.040000 70.170000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140000 12.960000 7.460000 13.280000 ;
      LAYER met4 ;
        RECT 7.140000 12.960000 7.460000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140000 13.400000 7.460000 13.720000 ;
      LAYER met4 ;
        RECT 7.140000 13.400000 7.460000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140000 13.840000 7.460000 14.160000 ;
      LAYER met4 ;
        RECT 7.140000 13.840000 7.460000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140000 14.280000 7.460000 14.600000 ;
      LAYER met4 ;
        RECT 7.140000 14.280000 7.460000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140000 14.720000 7.460000 15.040000 ;
      LAYER met4 ;
        RECT 7.140000 14.720000 7.460000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140000 15.160000 7.460000 15.480000 ;
      LAYER met4 ;
        RECT 7.140000 15.160000 7.460000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140000 15.600000 7.460000 15.920000 ;
      LAYER met4 ;
        RECT 7.140000 15.600000 7.460000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140000 16.040000 7.460000 16.360000 ;
      LAYER met4 ;
        RECT 7.140000 16.040000 7.460000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545000 12.960000 7.865000 13.280000 ;
      LAYER met4 ;
        RECT 7.545000 12.960000 7.865000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545000 13.400000 7.865000 13.720000 ;
      LAYER met4 ;
        RECT 7.545000 13.400000 7.865000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545000 13.840000 7.865000 14.160000 ;
      LAYER met4 ;
        RECT 7.545000 13.840000 7.865000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545000 14.280000 7.865000 14.600000 ;
      LAYER met4 ;
        RECT 7.545000 14.280000 7.865000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545000 14.720000 7.865000 15.040000 ;
      LAYER met4 ;
        RECT 7.545000 14.720000 7.865000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545000 15.160000 7.865000 15.480000 ;
      LAYER met4 ;
        RECT 7.545000 15.160000 7.865000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545000 15.600000 7.865000 15.920000 ;
      LAYER met4 ;
        RECT 7.545000 15.600000 7.865000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545000 16.040000 7.865000 16.360000 ;
      LAYER met4 ;
        RECT 7.545000 16.040000 7.865000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950000 12.960000 8.270000 13.280000 ;
      LAYER met4 ;
        RECT 7.950000 12.960000 8.270000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950000 13.400000 8.270000 13.720000 ;
      LAYER met4 ;
        RECT 7.950000 13.400000 8.270000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950000 13.840000 8.270000 14.160000 ;
      LAYER met4 ;
        RECT 7.950000 13.840000 8.270000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950000 14.280000 8.270000 14.600000 ;
      LAYER met4 ;
        RECT 7.950000 14.280000 8.270000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950000 14.720000 8.270000 15.040000 ;
      LAYER met4 ;
        RECT 7.950000 14.720000 8.270000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950000 15.160000 8.270000 15.480000 ;
      LAYER met4 ;
        RECT 7.950000 15.160000 8.270000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950000 15.600000 8.270000 15.920000 ;
      LAYER met4 ;
        RECT 7.950000 15.600000 8.270000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950000 16.040000 8.270000 16.360000 ;
      LAYER met4 ;
        RECT 7.950000 16.040000 8.270000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 12.960000 70.575000 13.280000 ;
      LAYER met4 ;
        RECT 70.255000 12.960000 70.575000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 13.400000 70.575000 13.720000 ;
      LAYER met4 ;
        RECT 70.255000 13.400000 70.575000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 13.840000 70.575000 14.160000 ;
      LAYER met4 ;
        RECT 70.255000 13.840000 70.575000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 14.280000 70.575000 14.600000 ;
      LAYER met4 ;
        RECT 70.255000 14.280000 70.575000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 14.720000 70.575000 15.040000 ;
      LAYER met4 ;
        RECT 70.255000 14.720000 70.575000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 15.160000 70.575000 15.480000 ;
      LAYER met4 ;
        RECT 70.255000 15.160000 70.575000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 15.600000 70.575000 15.920000 ;
      LAYER met4 ;
        RECT 70.255000 15.600000 70.575000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.255000 16.040000 70.575000 16.360000 ;
      LAYER met4 ;
        RECT 70.255000 16.040000 70.575000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 12.960000 70.980000 13.280000 ;
      LAYER met4 ;
        RECT 70.660000 12.960000 70.980000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 13.400000 70.980000 13.720000 ;
      LAYER met4 ;
        RECT 70.660000 13.400000 70.980000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 13.840000 70.980000 14.160000 ;
      LAYER met4 ;
        RECT 70.660000 13.840000 70.980000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 14.280000 70.980000 14.600000 ;
      LAYER met4 ;
        RECT 70.660000 14.280000 70.980000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 14.720000 70.980000 15.040000 ;
      LAYER met4 ;
        RECT 70.660000 14.720000 70.980000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 15.160000 70.980000 15.480000 ;
      LAYER met4 ;
        RECT 70.660000 15.160000 70.980000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 15.600000 70.980000 15.920000 ;
      LAYER met4 ;
        RECT 70.660000 15.600000 70.980000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.660000 16.040000 70.980000 16.360000 ;
      LAYER met4 ;
        RECT 70.660000 16.040000 70.980000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 12.960000 71.385000 13.280000 ;
      LAYER met4 ;
        RECT 71.065000 12.960000 71.385000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 13.400000 71.385000 13.720000 ;
      LAYER met4 ;
        RECT 71.065000 13.400000 71.385000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 13.840000 71.385000 14.160000 ;
      LAYER met4 ;
        RECT 71.065000 13.840000 71.385000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 14.280000 71.385000 14.600000 ;
      LAYER met4 ;
        RECT 71.065000 14.280000 71.385000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 14.720000 71.385000 15.040000 ;
      LAYER met4 ;
        RECT 71.065000 14.720000 71.385000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 15.160000 71.385000 15.480000 ;
      LAYER met4 ;
        RECT 71.065000 15.160000 71.385000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 15.600000 71.385000 15.920000 ;
      LAYER met4 ;
        RECT 71.065000 15.600000 71.385000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.065000 16.040000 71.385000 16.360000 ;
      LAYER met4 ;
        RECT 71.065000 16.040000 71.385000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 12.960000 71.790000 13.280000 ;
      LAYER met4 ;
        RECT 71.470000 12.960000 71.790000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 13.400000 71.790000 13.720000 ;
      LAYER met4 ;
        RECT 71.470000 13.400000 71.790000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 13.840000 71.790000 14.160000 ;
      LAYER met4 ;
        RECT 71.470000 13.840000 71.790000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 14.280000 71.790000 14.600000 ;
      LAYER met4 ;
        RECT 71.470000 14.280000 71.790000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 14.720000 71.790000 15.040000 ;
      LAYER met4 ;
        RECT 71.470000 14.720000 71.790000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 15.160000 71.790000 15.480000 ;
      LAYER met4 ;
        RECT 71.470000 15.160000 71.790000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 15.600000 71.790000 15.920000 ;
      LAYER met4 ;
        RECT 71.470000 15.600000 71.790000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.470000 16.040000 71.790000 16.360000 ;
      LAYER met4 ;
        RECT 71.470000 16.040000 71.790000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 12.960000 72.195000 13.280000 ;
      LAYER met4 ;
        RECT 71.875000 12.960000 72.195000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 13.400000 72.195000 13.720000 ;
      LAYER met4 ;
        RECT 71.875000 13.400000 72.195000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 13.840000 72.195000 14.160000 ;
      LAYER met4 ;
        RECT 71.875000 13.840000 72.195000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 14.280000 72.195000 14.600000 ;
      LAYER met4 ;
        RECT 71.875000 14.280000 72.195000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 14.720000 72.195000 15.040000 ;
      LAYER met4 ;
        RECT 71.875000 14.720000 72.195000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 15.160000 72.195000 15.480000 ;
      LAYER met4 ;
        RECT 71.875000 15.160000 72.195000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 15.600000 72.195000 15.920000 ;
      LAYER met4 ;
        RECT 71.875000 15.600000 72.195000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.875000 16.040000 72.195000 16.360000 ;
      LAYER met4 ;
        RECT 71.875000 16.040000 72.195000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 12.960000 72.600000 13.280000 ;
      LAYER met4 ;
        RECT 72.280000 12.960000 72.600000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 13.400000 72.600000 13.720000 ;
      LAYER met4 ;
        RECT 72.280000 13.400000 72.600000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 13.840000 72.600000 14.160000 ;
      LAYER met4 ;
        RECT 72.280000 13.840000 72.600000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 14.280000 72.600000 14.600000 ;
      LAYER met4 ;
        RECT 72.280000 14.280000 72.600000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 14.720000 72.600000 15.040000 ;
      LAYER met4 ;
        RECT 72.280000 14.720000 72.600000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 15.160000 72.600000 15.480000 ;
      LAYER met4 ;
        RECT 72.280000 15.160000 72.600000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 15.600000 72.600000 15.920000 ;
      LAYER met4 ;
        RECT 72.280000 15.600000 72.600000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.280000 16.040000 72.600000 16.360000 ;
      LAYER met4 ;
        RECT 72.280000 16.040000 72.600000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 12.960000 73.005000 13.280000 ;
      LAYER met4 ;
        RECT 72.685000 12.960000 73.005000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 13.400000 73.005000 13.720000 ;
      LAYER met4 ;
        RECT 72.685000 13.400000 73.005000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 13.840000 73.005000 14.160000 ;
      LAYER met4 ;
        RECT 72.685000 13.840000 73.005000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 14.280000 73.005000 14.600000 ;
      LAYER met4 ;
        RECT 72.685000 14.280000 73.005000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 14.720000 73.005000 15.040000 ;
      LAYER met4 ;
        RECT 72.685000 14.720000 73.005000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 15.160000 73.005000 15.480000 ;
      LAYER met4 ;
        RECT 72.685000 15.160000 73.005000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 15.600000 73.005000 15.920000 ;
      LAYER met4 ;
        RECT 72.685000 15.600000 73.005000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.685000 16.040000 73.005000 16.360000 ;
      LAYER met4 ;
        RECT 72.685000 16.040000 73.005000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 12.960000 73.410000 13.280000 ;
      LAYER met4 ;
        RECT 73.090000 12.960000 73.410000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 13.400000 73.410000 13.720000 ;
      LAYER met4 ;
        RECT 73.090000 13.400000 73.410000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 13.840000 73.410000 14.160000 ;
      LAYER met4 ;
        RECT 73.090000 13.840000 73.410000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 14.280000 73.410000 14.600000 ;
      LAYER met4 ;
        RECT 73.090000 14.280000 73.410000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 14.720000 73.410000 15.040000 ;
      LAYER met4 ;
        RECT 73.090000 14.720000 73.410000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 15.160000 73.410000 15.480000 ;
      LAYER met4 ;
        RECT 73.090000 15.160000 73.410000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 15.600000 73.410000 15.920000 ;
      LAYER met4 ;
        RECT 73.090000 15.600000 73.410000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090000 16.040000 73.410000 16.360000 ;
      LAYER met4 ;
        RECT 73.090000 16.040000 73.410000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 12.960000 73.815000 13.280000 ;
      LAYER met4 ;
        RECT 73.495000 12.960000 73.815000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 13.400000 73.815000 13.720000 ;
      LAYER met4 ;
        RECT 73.495000 13.400000 73.815000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 13.840000 73.815000 14.160000 ;
      LAYER met4 ;
        RECT 73.495000 13.840000 73.815000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 14.280000 73.815000 14.600000 ;
      LAYER met4 ;
        RECT 73.495000 14.280000 73.815000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 14.720000 73.815000 15.040000 ;
      LAYER met4 ;
        RECT 73.495000 14.720000 73.815000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 15.160000 73.815000 15.480000 ;
      LAYER met4 ;
        RECT 73.495000 15.160000 73.815000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 15.600000 73.815000 15.920000 ;
      LAYER met4 ;
        RECT 73.495000 15.600000 73.815000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.495000 16.040000 73.815000 16.360000 ;
      LAYER met4 ;
        RECT 73.495000 16.040000 73.815000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 12.960000 74.220000 13.280000 ;
      LAYER met4 ;
        RECT 73.900000 12.960000 74.220000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 13.400000 74.220000 13.720000 ;
      LAYER met4 ;
        RECT 73.900000 13.400000 74.220000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 13.840000 74.220000 14.160000 ;
      LAYER met4 ;
        RECT 73.900000 13.840000 74.220000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 14.280000 74.220000 14.600000 ;
      LAYER met4 ;
        RECT 73.900000 14.280000 74.220000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 14.720000 74.220000 15.040000 ;
      LAYER met4 ;
        RECT 73.900000 14.720000 74.220000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 15.160000 74.220000 15.480000 ;
      LAYER met4 ;
        RECT 73.900000 15.160000 74.220000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 15.600000 74.220000 15.920000 ;
      LAYER met4 ;
        RECT 73.900000 15.600000 74.220000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.900000 16.040000 74.220000 16.360000 ;
      LAYER met4 ;
        RECT 73.900000 16.040000 74.220000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 12.960000 74.625000 13.280000 ;
      LAYER met4 ;
        RECT 74.305000 12.960000 74.625000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 13.400000 74.625000 13.720000 ;
      LAYER met4 ;
        RECT 74.305000 13.400000 74.625000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 13.840000 74.625000 14.160000 ;
      LAYER met4 ;
        RECT 74.305000 13.840000 74.625000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 14.280000 74.625000 14.600000 ;
      LAYER met4 ;
        RECT 74.305000 14.280000 74.625000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 14.720000 74.625000 15.040000 ;
      LAYER met4 ;
        RECT 74.305000 14.720000 74.625000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 15.160000 74.625000 15.480000 ;
      LAYER met4 ;
        RECT 74.305000 15.160000 74.625000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 15.600000 74.625000 15.920000 ;
      LAYER met4 ;
        RECT 74.305000 15.600000 74.625000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.305000 16.040000 74.625000 16.360000 ;
      LAYER met4 ;
        RECT 74.305000 16.040000 74.625000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355000 12.960000 8.675000 13.280000 ;
      LAYER met4 ;
        RECT 8.355000 12.960000 8.675000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355000 13.400000 8.675000 13.720000 ;
      LAYER met4 ;
        RECT 8.355000 13.400000 8.675000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355000 13.840000 8.675000 14.160000 ;
      LAYER met4 ;
        RECT 8.355000 13.840000 8.675000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355000 14.280000 8.675000 14.600000 ;
      LAYER met4 ;
        RECT 8.355000 14.280000 8.675000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355000 14.720000 8.675000 15.040000 ;
      LAYER met4 ;
        RECT 8.355000 14.720000 8.675000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355000 15.160000 8.675000 15.480000 ;
      LAYER met4 ;
        RECT 8.355000 15.160000 8.675000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355000 15.600000 8.675000 15.920000 ;
      LAYER met4 ;
        RECT 8.355000 15.600000 8.675000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355000 16.040000 8.675000 16.360000 ;
      LAYER met4 ;
        RECT 8.355000 16.040000 8.675000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760000 12.960000 9.080000 13.280000 ;
      LAYER met4 ;
        RECT 8.760000 12.960000 9.080000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760000 13.400000 9.080000 13.720000 ;
      LAYER met4 ;
        RECT 8.760000 13.400000 9.080000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760000 13.840000 9.080000 14.160000 ;
      LAYER met4 ;
        RECT 8.760000 13.840000 9.080000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760000 14.280000 9.080000 14.600000 ;
      LAYER met4 ;
        RECT 8.760000 14.280000 9.080000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760000 14.720000 9.080000 15.040000 ;
      LAYER met4 ;
        RECT 8.760000 14.720000 9.080000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760000 15.160000 9.080000 15.480000 ;
      LAYER met4 ;
        RECT 8.760000 15.160000 9.080000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760000 15.600000 9.080000 15.920000 ;
      LAYER met4 ;
        RECT 8.760000 15.600000 9.080000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760000 16.040000 9.080000 16.360000 ;
      LAYER met4 ;
        RECT 8.760000 16.040000 9.080000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165000 12.960000 9.485000 13.280000 ;
      LAYER met4 ;
        RECT 9.165000 12.960000 9.485000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165000 13.400000 9.485000 13.720000 ;
      LAYER met4 ;
        RECT 9.165000 13.400000 9.485000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165000 13.840000 9.485000 14.160000 ;
      LAYER met4 ;
        RECT 9.165000 13.840000 9.485000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165000 14.280000 9.485000 14.600000 ;
      LAYER met4 ;
        RECT 9.165000 14.280000 9.485000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165000 14.720000 9.485000 15.040000 ;
      LAYER met4 ;
        RECT 9.165000 14.720000 9.485000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165000 15.160000 9.485000 15.480000 ;
      LAYER met4 ;
        RECT 9.165000 15.160000 9.485000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165000 15.600000 9.485000 15.920000 ;
      LAYER met4 ;
        RECT 9.165000 15.600000 9.485000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165000 16.040000 9.485000 16.360000 ;
      LAYER met4 ;
        RECT 9.165000 16.040000 9.485000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570000 12.960000 9.890000 13.280000 ;
      LAYER met4 ;
        RECT 9.570000 12.960000 9.890000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570000 13.400000 9.890000 13.720000 ;
      LAYER met4 ;
        RECT 9.570000 13.400000 9.890000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570000 13.840000 9.890000 14.160000 ;
      LAYER met4 ;
        RECT 9.570000 13.840000 9.890000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570000 14.280000 9.890000 14.600000 ;
      LAYER met4 ;
        RECT 9.570000 14.280000 9.890000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570000 14.720000 9.890000 15.040000 ;
      LAYER met4 ;
        RECT 9.570000 14.720000 9.890000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570000 15.160000 9.890000 15.480000 ;
      LAYER met4 ;
        RECT 9.570000 15.160000 9.890000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570000 15.600000 9.890000 15.920000 ;
      LAYER met4 ;
        RECT 9.570000 15.600000 9.890000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570000 16.040000 9.890000 16.360000 ;
      LAYER met4 ;
        RECT 9.570000 16.040000 9.890000 16.360000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975000 12.960000 10.295000 13.280000 ;
      LAYER met4 ;
        RECT 9.975000 12.960000 10.295000 13.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975000 13.400000 10.295000 13.720000 ;
      LAYER met4 ;
        RECT 9.975000 13.400000 10.295000 13.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975000 13.840000 10.295000 14.160000 ;
      LAYER met4 ;
        RECT 9.975000 13.840000 10.295000 14.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975000 14.280000 10.295000 14.600000 ;
      LAYER met4 ;
        RECT 9.975000 14.280000 10.295000 14.600000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975000 14.720000 10.295000 15.040000 ;
      LAYER met4 ;
        RECT 9.975000 14.720000 10.295000 15.040000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975000 15.160000 10.295000 15.480000 ;
      LAYER met4 ;
        RECT 9.975000 15.160000 10.295000 15.480000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975000 15.600000 10.295000 15.920000 ;
      LAYER met4 ;
        RECT 9.975000 15.600000 10.295000 15.920000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975000 16.040000 10.295000 16.360000 ;
      LAYER met4 ;
        RECT 9.975000 16.040000 10.295000 16.360000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 68.035000 75.000000 92.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 62.185000 75.000000 66.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 45.735000 75.000000 54.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 39.685000 75.000000 44.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 23.935000 75.000000 28.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 56.335000 75.000000 60.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 29.985000 75.000000 33.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met3 ;
      RECT 0.600000 12.940000 74.655000 16.380000 ;
    LAYER met4 ;
      RECT 0.000000  0.035000 75.000000  45.965000 ;
      RECT 0.000000 49.745000 75.000000  50.725000 ;
      RECT 0.000000 54.505000 75.000000 198.000000 ;
    LAYER met5 ;
      RECT 0.000000  0.135000 72.130000  13.035000 ;
      RECT 0.000000 13.035000 75.000000  22.335000 ;
      RECT 0.000000 22.335000 72.130000  34.835000 ;
      RECT 0.000000 34.835000 75.000000  38.085000 ;
      RECT 0.000000 38.085000 72.130000  94.585000 ;
      RECT 0.000000 94.585000 75.000000 198.000000 ;
  END
END sky130_fd_io__overlay_vdda_lvc
END LIBRARY
