# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__overlay_vccd_hvc
  CLASS BLOCK ;
  FOREIGN sky130_fd_io__overlay_vccd_hvc ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  75.00000 BY  200.0000 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.525000 10.190000 0.845000 10.510000 ;
      LAYER met4 ;
        RECT 0.525000 10.190000 0.845000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 10.620000 0.845000 10.940000 ;
      LAYER met4 ;
        RECT 0.525000 10.620000 0.845000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 11.050000 0.845000 11.370000 ;
      LAYER met4 ;
        RECT 0.525000 11.050000 0.845000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 11.480000 0.845000 11.800000 ;
      LAYER met4 ;
        RECT 0.525000 11.480000 0.845000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 11.910000 0.845000 12.230000 ;
      LAYER met4 ;
        RECT 0.525000 11.910000 0.845000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 12.340000 0.845000 12.660000 ;
      LAYER met4 ;
        RECT 0.525000 12.340000 0.845000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 12.770000 0.845000 13.090000 ;
      LAYER met4 ;
        RECT 0.525000 12.770000 0.845000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 13.200000 0.845000 13.520000 ;
      LAYER met4 ;
        RECT 0.525000 13.200000 0.845000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 8.900000 0.845000 9.220000 ;
      LAYER met4 ;
        RECT 0.525000 8.900000 0.845000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 9.330000 0.845000 9.650000 ;
      LAYER met4 ;
        RECT 0.525000 9.330000 0.845000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 9.760000 0.845000 10.080000 ;
      LAYER met4 ;
        RECT 0.525000 9.760000 0.845000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 10.190000 1.255000 10.510000 ;
      LAYER met4 ;
        RECT 0.935000 10.190000 1.255000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 10.620000 1.255000 10.940000 ;
      LAYER met4 ;
        RECT 0.935000 10.620000 1.255000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 11.050000 1.255000 11.370000 ;
      LAYER met4 ;
        RECT 0.935000 11.050000 1.255000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 11.480000 1.255000 11.800000 ;
      LAYER met4 ;
        RECT 0.935000 11.480000 1.255000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 11.910000 1.255000 12.230000 ;
      LAYER met4 ;
        RECT 0.935000 11.910000 1.255000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 12.340000 1.255000 12.660000 ;
      LAYER met4 ;
        RECT 0.935000 12.340000 1.255000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 12.770000 1.255000 13.090000 ;
      LAYER met4 ;
        RECT 0.935000 12.770000 1.255000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 13.200000 1.255000 13.520000 ;
      LAYER met4 ;
        RECT 0.935000 13.200000 1.255000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 8.900000 1.255000 9.220000 ;
      LAYER met4 ;
        RECT 0.935000 8.900000 1.255000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 9.330000 1.255000 9.650000 ;
      LAYER met4 ;
        RECT 0.935000 9.330000 1.255000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 9.760000 1.255000 10.080000 ;
      LAYER met4 ;
        RECT 0.935000 9.760000 1.255000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 10.190000 1.665000 10.510000 ;
      LAYER met4 ;
        RECT 1.345000 10.190000 1.665000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 10.620000 1.665000 10.940000 ;
      LAYER met4 ;
        RECT 1.345000 10.620000 1.665000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 11.050000 1.665000 11.370000 ;
      LAYER met4 ;
        RECT 1.345000 11.050000 1.665000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 11.480000 1.665000 11.800000 ;
      LAYER met4 ;
        RECT 1.345000 11.480000 1.665000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 11.910000 1.665000 12.230000 ;
      LAYER met4 ;
        RECT 1.345000 11.910000 1.665000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 12.340000 1.665000 12.660000 ;
      LAYER met4 ;
        RECT 1.345000 12.340000 1.665000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 12.770000 1.665000 13.090000 ;
      LAYER met4 ;
        RECT 1.345000 12.770000 1.665000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 13.200000 1.665000 13.520000 ;
      LAYER met4 ;
        RECT 1.345000 13.200000 1.665000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 8.900000 1.665000 9.220000 ;
      LAYER met4 ;
        RECT 1.345000 8.900000 1.665000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 9.330000 1.665000 9.650000 ;
      LAYER met4 ;
        RECT 1.345000 9.330000 1.665000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 9.760000 1.665000 10.080000 ;
      LAYER met4 ;
        RECT 1.345000 9.760000 1.665000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 10.190000 2.075000 10.510000 ;
      LAYER met4 ;
        RECT 1.755000 10.190000 2.075000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 10.620000 2.075000 10.940000 ;
      LAYER met4 ;
        RECT 1.755000 10.620000 2.075000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 11.050000 2.075000 11.370000 ;
      LAYER met4 ;
        RECT 1.755000 11.050000 2.075000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 11.480000 2.075000 11.800000 ;
      LAYER met4 ;
        RECT 1.755000 11.480000 2.075000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 11.910000 2.075000 12.230000 ;
      LAYER met4 ;
        RECT 1.755000 11.910000 2.075000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 12.340000 2.075000 12.660000 ;
      LAYER met4 ;
        RECT 1.755000 12.340000 2.075000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 12.770000 2.075000 13.090000 ;
      LAYER met4 ;
        RECT 1.755000 12.770000 2.075000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 13.200000 2.075000 13.520000 ;
      LAYER met4 ;
        RECT 1.755000 13.200000 2.075000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 8.900000 2.075000 9.220000 ;
      LAYER met4 ;
        RECT 1.755000 8.900000 2.075000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 9.330000 2.075000 9.650000 ;
      LAYER met4 ;
        RECT 1.755000 9.330000 2.075000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 9.760000 2.075000 10.080000 ;
      LAYER met4 ;
        RECT 1.755000 9.760000 2.075000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 10.190000 10.595000 10.510000 ;
      LAYER met4 ;
        RECT 10.275000 10.190000 10.595000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 10.620000 10.595000 10.940000 ;
      LAYER met4 ;
        RECT 10.275000 10.620000 10.595000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 11.050000 10.595000 11.370000 ;
      LAYER met4 ;
        RECT 10.275000 11.050000 10.595000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 11.480000 10.595000 11.800000 ;
      LAYER met4 ;
        RECT 10.275000 11.480000 10.595000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 11.910000 10.595000 12.230000 ;
      LAYER met4 ;
        RECT 10.275000 11.910000 10.595000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 12.340000 10.595000 12.660000 ;
      LAYER met4 ;
        RECT 10.275000 12.340000 10.595000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 12.770000 10.595000 13.090000 ;
      LAYER met4 ;
        RECT 10.275000 12.770000 10.595000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 13.200000 10.595000 13.520000 ;
      LAYER met4 ;
        RECT 10.275000 13.200000 10.595000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 8.900000 10.595000 9.220000 ;
      LAYER met4 ;
        RECT 10.275000 8.900000 10.595000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 9.330000 10.595000 9.650000 ;
      LAYER met4 ;
        RECT 10.275000 9.330000 10.595000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 9.760000 10.595000 10.080000 ;
      LAYER met4 ;
        RECT 10.275000 9.760000 10.595000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 10.190000 11.000000 10.510000 ;
      LAYER met4 ;
        RECT 10.680000 10.190000 11.000000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 10.620000 11.000000 10.940000 ;
      LAYER met4 ;
        RECT 10.680000 10.620000 11.000000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 11.050000 11.000000 11.370000 ;
      LAYER met4 ;
        RECT 10.680000 11.050000 11.000000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 11.480000 11.000000 11.800000 ;
      LAYER met4 ;
        RECT 10.680000 11.480000 11.000000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 11.910000 11.000000 12.230000 ;
      LAYER met4 ;
        RECT 10.680000 11.910000 11.000000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 12.340000 11.000000 12.660000 ;
      LAYER met4 ;
        RECT 10.680000 12.340000 11.000000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 12.770000 11.000000 13.090000 ;
      LAYER met4 ;
        RECT 10.680000 12.770000 11.000000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 13.200000 11.000000 13.520000 ;
      LAYER met4 ;
        RECT 10.680000 13.200000 11.000000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 8.900000 11.000000 9.220000 ;
      LAYER met4 ;
        RECT 10.680000 8.900000 11.000000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 9.330000 11.000000 9.650000 ;
      LAYER met4 ;
        RECT 10.680000 9.330000 11.000000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 9.760000 11.000000 10.080000 ;
      LAYER met4 ;
        RECT 10.680000 9.760000 11.000000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 10.190000 11.405000 10.510000 ;
      LAYER met4 ;
        RECT 11.085000 10.190000 11.405000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 10.620000 11.405000 10.940000 ;
      LAYER met4 ;
        RECT 11.085000 10.620000 11.405000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 11.050000 11.405000 11.370000 ;
      LAYER met4 ;
        RECT 11.085000 11.050000 11.405000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 11.480000 11.405000 11.800000 ;
      LAYER met4 ;
        RECT 11.085000 11.480000 11.405000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 11.910000 11.405000 12.230000 ;
      LAYER met4 ;
        RECT 11.085000 11.910000 11.405000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 12.340000 11.405000 12.660000 ;
      LAYER met4 ;
        RECT 11.085000 12.340000 11.405000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 12.770000 11.405000 13.090000 ;
      LAYER met4 ;
        RECT 11.085000 12.770000 11.405000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 13.200000 11.405000 13.520000 ;
      LAYER met4 ;
        RECT 11.085000 13.200000 11.405000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 8.900000 11.405000 9.220000 ;
      LAYER met4 ;
        RECT 11.085000 8.900000 11.405000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 9.330000 11.405000 9.650000 ;
      LAYER met4 ;
        RECT 11.085000 9.330000 11.405000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 9.760000 11.405000 10.080000 ;
      LAYER met4 ;
        RECT 11.085000 9.760000 11.405000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 10.190000 11.810000 10.510000 ;
      LAYER met4 ;
        RECT 11.490000 10.190000 11.810000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 10.620000 11.810000 10.940000 ;
      LAYER met4 ;
        RECT 11.490000 10.620000 11.810000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 11.050000 11.810000 11.370000 ;
      LAYER met4 ;
        RECT 11.490000 11.050000 11.810000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 11.480000 11.810000 11.800000 ;
      LAYER met4 ;
        RECT 11.490000 11.480000 11.810000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 11.910000 11.810000 12.230000 ;
      LAYER met4 ;
        RECT 11.490000 11.910000 11.810000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 12.340000 11.810000 12.660000 ;
      LAYER met4 ;
        RECT 11.490000 12.340000 11.810000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 12.770000 11.810000 13.090000 ;
      LAYER met4 ;
        RECT 11.490000 12.770000 11.810000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 13.200000 11.810000 13.520000 ;
      LAYER met4 ;
        RECT 11.490000 13.200000 11.810000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 8.900000 11.810000 9.220000 ;
      LAYER met4 ;
        RECT 11.490000 8.900000 11.810000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 9.330000 11.810000 9.650000 ;
      LAYER met4 ;
        RECT 11.490000 9.330000 11.810000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 9.760000 11.810000 10.080000 ;
      LAYER met4 ;
        RECT 11.490000 9.760000 11.810000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 10.190000 12.215000 10.510000 ;
      LAYER met4 ;
        RECT 11.895000 10.190000 12.215000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 10.620000 12.215000 10.940000 ;
      LAYER met4 ;
        RECT 11.895000 10.620000 12.215000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 11.050000 12.215000 11.370000 ;
      LAYER met4 ;
        RECT 11.895000 11.050000 12.215000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 11.480000 12.215000 11.800000 ;
      LAYER met4 ;
        RECT 11.895000 11.480000 12.215000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 11.910000 12.215000 12.230000 ;
      LAYER met4 ;
        RECT 11.895000 11.910000 12.215000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 12.340000 12.215000 12.660000 ;
      LAYER met4 ;
        RECT 11.895000 12.340000 12.215000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 12.770000 12.215000 13.090000 ;
      LAYER met4 ;
        RECT 11.895000 12.770000 12.215000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 13.200000 12.215000 13.520000 ;
      LAYER met4 ;
        RECT 11.895000 13.200000 12.215000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 8.900000 12.215000 9.220000 ;
      LAYER met4 ;
        RECT 11.895000 8.900000 12.215000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 9.330000 12.215000 9.650000 ;
      LAYER met4 ;
        RECT 11.895000 9.330000 12.215000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 9.760000 12.215000 10.080000 ;
      LAYER met4 ;
        RECT 11.895000 9.760000 12.215000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 10.190000 12.620000 10.510000 ;
      LAYER met4 ;
        RECT 12.300000 10.190000 12.620000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 10.620000 12.620000 10.940000 ;
      LAYER met4 ;
        RECT 12.300000 10.620000 12.620000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 11.050000 12.620000 11.370000 ;
      LAYER met4 ;
        RECT 12.300000 11.050000 12.620000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 11.480000 12.620000 11.800000 ;
      LAYER met4 ;
        RECT 12.300000 11.480000 12.620000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 11.910000 12.620000 12.230000 ;
      LAYER met4 ;
        RECT 12.300000 11.910000 12.620000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 12.340000 12.620000 12.660000 ;
      LAYER met4 ;
        RECT 12.300000 12.340000 12.620000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 12.770000 12.620000 13.090000 ;
      LAYER met4 ;
        RECT 12.300000 12.770000 12.620000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 13.200000 12.620000 13.520000 ;
      LAYER met4 ;
        RECT 12.300000 13.200000 12.620000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 8.900000 12.620000 9.220000 ;
      LAYER met4 ;
        RECT 12.300000 8.900000 12.620000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 9.330000 12.620000 9.650000 ;
      LAYER met4 ;
        RECT 12.300000 9.330000 12.620000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 9.760000 12.620000 10.080000 ;
      LAYER met4 ;
        RECT 12.300000 9.760000 12.620000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 10.190000 13.025000 10.510000 ;
      LAYER met4 ;
        RECT 12.705000 10.190000 13.025000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 10.620000 13.025000 10.940000 ;
      LAYER met4 ;
        RECT 12.705000 10.620000 13.025000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 11.050000 13.025000 11.370000 ;
      LAYER met4 ;
        RECT 12.705000 11.050000 13.025000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 11.480000 13.025000 11.800000 ;
      LAYER met4 ;
        RECT 12.705000 11.480000 13.025000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 11.910000 13.025000 12.230000 ;
      LAYER met4 ;
        RECT 12.705000 11.910000 13.025000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 12.340000 13.025000 12.660000 ;
      LAYER met4 ;
        RECT 12.705000 12.340000 13.025000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 12.770000 13.025000 13.090000 ;
      LAYER met4 ;
        RECT 12.705000 12.770000 13.025000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 13.200000 13.025000 13.520000 ;
      LAYER met4 ;
        RECT 12.705000 13.200000 13.025000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 8.900000 13.025000 9.220000 ;
      LAYER met4 ;
        RECT 12.705000 8.900000 13.025000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 9.330000 13.025000 9.650000 ;
      LAYER met4 ;
        RECT 12.705000 9.330000 13.025000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 9.760000 13.025000 10.080000 ;
      LAYER met4 ;
        RECT 12.705000 9.760000 13.025000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 10.190000 13.430000 10.510000 ;
      LAYER met4 ;
        RECT 13.110000 10.190000 13.430000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 10.620000 13.430000 10.940000 ;
      LAYER met4 ;
        RECT 13.110000 10.620000 13.430000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 11.050000 13.430000 11.370000 ;
      LAYER met4 ;
        RECT 13.110000 11.050000 13.430000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 11.480000 13.430000 11.800000 ;
      LAYER met4 ;
        RECT 13.110000 11.480000 13.430000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 11.910000 13.430000 12.230000 ;
      LAYER met4 ;
        RECT 13.110000 11.910000 13.430000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 12.340000 13.430000 12.660000 ;
      LAYER met4 ;
        RECT 13.110000 12.340000 13.430000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 12.770000 13.430000 13.090000 ;
      LAYER met4 ;
        RECT 13.110000 12.770000 13.430000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 13.200000 13.430000 13.520000 ;
      LAYER met4 ;
        RECT 13.110000 13.200000 13.430000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 8.900000 13.430000 9.220000 ;
      LAYER met4 ;
        RECT 13.110000 8.900000 13.430000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 9.330000 13.430000 9.650000 ;
      LAYER met4 ;
        RECT 13.110000 9.330000 13.430000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 9.760000 13.430000 10.080000 ;
      LAYER met4 ;
        RECT 13.110000 9.760000 13.430000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 10.190000 13.835000 10.510000 ;
      LAYER met4 ;
        RECT 13.515000 10.190000 13.835000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 10.620000 13.835000 10.940000 ;
      LAYER met4 ;
        RECT 13.515000 10.620000 13.835000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 11.050000 13.835000 11.370000 ;
      LAYER met4 ;
        RECT 13.515000 11.050000 13.835000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 11.480000 13.835000 11.800000 ;
      LAYER met4 ;
        RECT 13.515000 11.480000 13.835000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 11.910000 13.835000 12.230000 ;
      LAYER met4 ;
        RECT 13.515000 11.910000 13.835000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 12.340000 13.835000 12.660000 ;
      LAYER met4 ;
        RECT 13.515000 12.340000 13.835000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 12.770000 13.835000 13.090000 ;
      LAYER met4 ;
        RECT 13.515000 12.770000 13.835000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 13.200000 13.835000 13.520000 ;
      LAYER met4 ;
        RECT 13.515000 13.200000 13.835000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 8.900000 13.835000 9.220000 ;
      LAYER met4 ;
        RECT 13.515000 8.900000 13.835000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 9.330000 13.835000 9.650000 ;
      LAYER met4 ;
        RECT 13.515000 9.330000 13.835000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 9.760000 13.835000 10.080000 ;
      LAYER met4 ;
        RECT 13.515000 9.760000 13.835000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 10.190000 14.240000 10.510000 ;
      LAYER met4 ;
        RECT 13.920000 10.190000 14.240000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 10.620000 14.240000 10.940000 ;
      LAYER met4 ;
        RECT 13.920000 10.620000 14.240000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 11.050000 14.240000 11.370000 ;
      LAYER met4 ;
        RECT 13.920000 11.050000 14.240000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 11.480000 14.240000 11.800000 ;
      LAYER met4 ;
        RECT 13.920000 11.480000 14.240000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 11.910000 14.240000 12.230000 ;
      LAYER met4 ;
        RECT 13.920000 11.910000 14.240000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 12.340000 14.240000 12.660000 ;
      LAYER met4 ;
        RECT 13.920000 12.340000 14.240000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 12.770000 14.240000 13.090000 ;
      LAYER met4 ;
        RECT 13.920000 12.770000 14.240000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 13.200000 14.240000 13.520000 ;
      LAYER met4 ;
        RECT 13.920000 13.200000 14.240000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 8.900000 14.240000 9.220000 ;
      LAYER met4 ;
        RECT 13.920000 8.900000 14.240000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 9.330000 14.240000 9.650000 ;
      LAYER met4 ;
        RECT 13.920000 9.330000 14.240000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 9.760000 14.240000 10.080000 ;
      LAYER met4 ;
        RECT 13.920000 9.760000 14.240000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 10.190000 14.645000 10.510000 ;
      LAYER met4 ;
        RECT 14.325000 10.190000 14.645000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 10.620000 14.645000 10.940000 ;
      LAYER met4 ;
        RECT 14.325000 10.620000 14.645000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 11.050000 14.645000 11.370000 ;
      LAYER met4 ;
        RECT 14.325000 11.050000 14.645000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 11.480000 14.645000 11.800000 ;
      LAYER met4 ;
        RECT 14.325000 11.480000 14.645000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 11.910000 14.645000 12.230000 ;
      LAYER met4 ;
        RECT 14.325000 11.910000 14.645000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 12.340000 14.645000 12.660000 ;
      LAYER met4 ;
        RECT 14.325000 12.340000 14.645000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 12.770000 14.645000 13.090000 ;
      LAYER met4 ;
        RECT 14.325000 12.770000 14.645000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 13.200000 14.645000 13.520000 ;
      LAYER met4 ;
        RECT 14.325000 13.200000 14.645000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 8.900000 14.645000 9.220000 ;
      LAYER met4 ;
        RECT 14.325000 8.900000 14.645000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 9.330000 14.645000 9.650000 ;
      LAYER met4 ;
        RECT 14.325000 9.330000 14.645000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 9.760000 14.645000 10.080000 ;
      LAYER met4 ;
        RECT 14.325000 9.760000 14.645000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 10.190000 15.050000 10.510000 ;
      LAYER met4 ;
        RECT 14.730000 10.190000 15.050000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 10.620000 15.050000 10.940000 ;
      LAYER met4 ;
        RECT 14.730000 10.620000 15.050000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 11.050000 15.050000 11.370000 ;
      LAYER met4 ;
        RECT 14.730000 11.050000 15.050000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 11.480000 15.050000 11.800000 ;
      LAYER met4 ;
        RECT 14.730000 11.480000 15.050000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 11.910000 15.050000 12.230000 ;
      LAYER met4 ;
        RECT 14.730000 11.910000 15.050000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 12.340000 15.050000 12.660000 ;
      LAYER met4 ;
        RECT 14.730000 12.340000 15.050000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 12.770000 15.050000 13.090000 ;
      LAYER met4 ;
        RECT 14.730000 12.770000 15.050000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 13.200000 15.050000 13.520000 ;
      LAYER met4 ;
        RECT 14.730000 13.200000 15.050000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 8.900000 15.050000 9.220000 ;
      LAYER met4 ;
        RECT 14.730000 8.900000 15.050000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 9.330000 15.050000 9.650000 ;
      LAYER met4 ;
        RECT 14.730000 9.330000 15.050000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 9.760000 15.050000 10.080000 ;
      LAYER met4 ;
        RECT 14.730000 9.760000 15.050000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 10.190000 15.455000 10.510000 ;
      LAYER met4 ;
        RECT 15.135000 10.190000 15.455000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 10.620000 15.455000 10.940000 ;
      LAYER met4 ;
        RECT 15.135000 10.620000 15.455000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 11.050000 15.455000 11.370000 ;
      LAYER met4 ;
        RECT 15.135000 11.050000 15.455000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 11.480000 15.455000 11.800000 ;
      LAYER met4 ;
        RECT 15.135000 11.480000 15.455000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 11.910000 15.455000 12.230000 ;
      LAYER met4 ;
        RECT 15.135000 11.910000 15.455000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 12.340000 15.455000 12.660000 ;
      LAYER met4 ;
        RECT 15.135000 12.340000 15.455000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 12.770000 15.455000 13.090000 ;
      LAYER met4 ;
        RECT 15.135000 12.770000 15.455000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 13.200000 15.455000 13.520000 ;
      LAYER met4 ;
        RECT 15.135000 13.200000 15.455000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 8.900000 15.455000 9.220000 ;
      LAYER met4 ;
        RECT 15.135000 8.900000 15.455000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 9.330000 15.455000 9.650000 ;
      LAYER met4 ;
        RECT 15.135000 9.330000 15.455000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 9.760000 15.455000 10.080000 ;
      LAYER met4 ;
        RECT 15.135000 9.760000 15.455000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 10.190000 15.860000 10.510000 ;
      LAYER met4 ;
        RECT 15.540000 10.190000 15.860000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 10.620000 15.860000 10.940000 ;
      LAYER met4 ;
        RECT 15.540000 10.620000 15.860000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 11.050000 15.860000 11.370000 ;
      LAYER met4 ;
        RECT 15.540000 11.050000 15.860000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 11.480000 15.860000 11.800000 ;
      LAYER met4 ;
        RECT 15.540000 11.480000 15.860000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 11.910000 15.860000 12.230000 ;
      LAYER met4 ;
        RECT 15.540000 11.910000 15.860000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 12.340000 15.860000 12.660000 ;
      LAYER met4 ;
        RECT 15.540000 12.340000 15.860000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 12.770000 15.860000 13.090000 ;
      LAYER met4 ;
        RECT 15.540000 12.770000 15.860000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 13.200000 15.860000 13.520000 ;
      LAYER met4 ;
        RECT 15.540000 13.200000 15.860000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 8.900000 15.860000 9.220000 ;
      LAYER met4 ;
        RECT 15.540000 8.900000 15.860000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 9.330000 15.860000 9.650000 ;
      LAYER met4 ;
        RECT 15.540000 9.330000 15.860000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 9.760000 15.860000 10.080000 ;
      LAYER met4 ;
        RECT 15.540000 9.760000 15.860000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 10.190000 16.265000 10.510000 ;
      LAYER met4 ;
        RECT 15.945000 10.190000 16.265000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 10.620000 16.265000 10.940000 ;
      LAYER met4 ;
        RECT 15.945000 10.620000 16.265000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 11.050000 16.265000 11.370000 ;
      LAYER met4 ;
        RECT 15.945000 11.050000 16.265000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 11.480000 16.265000 11.800000 ;
      LAYER met4 ;
        RECT 15.945000 11.480000 16.265000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 11.910000 16.265000 12.230000 ;
      LAYER met4 ;
        RECT 15.945000 11.910000 16.265000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 12.340000 16.265000 12.660000 ;
      LAYER met4 ;
        RECT 15.945000 12.340000 16.265000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 12.770000 16.265000 13.090000 ;
      LAYER met4 ;
        RECT 15.945000 12.770000 16.265000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 13.200000 16.265000 13.520000 ;
      LAYER met4 ;
        RECT 15.945000 13.200000 16.265000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 8.900000 16.265000 9.220000 ;
      LAYER met4 ;
        RECT 15.945000 8.900000 16.265000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 9.330000 16.265000 9.650000 ;
      LAYER met4 ;
        RECT 15.945000 9.330000 16.265000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 9.760000 16.265000 10.080000 ;
      LAYER met4 ;
        RECT 15.945000 9.760000 16.265000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 10.190000 16.670000 10.510000 ;
      LAYER met4 ;
        RECT 16.350000 10.190000 16.670000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 10.620000 16.670000 10.940000 ;
      LAYER met4 ;
        RECT 16.350000 10.620000 16.670000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 11.050000 16.670000 11.370000 ;
      LAYER met4 ;
        RECT 16.350000 11.050000 16.670000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 11.480000 16.670000 11.800000 ;
      LAYER met4 ;
        RECT 16.350000 11.480000 16.670000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 11.910000 16.670000 12.230000 ;
      LAYER met4 ;
        RECT 16.350000 11.910000 16.670000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 12.340000 16.670000 12.660000 ;
      LAYER met4 ;
        RECT 16.350000 12.340000 16.670000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 12.770000 16.670000 13.090000 ;
      LAYER met4 ;
        RECT 16.350000 12.770000 16.670000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 13.200000 16.670000 13.520000 ;
      LAYER met4 ;
        RECT 16.350000 13.200000 16.670000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 8.900000 16.670000 9.220000 ;
      LAYER met4 ;
        RECT 16.350000 8.900000 16.670000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 9.330000 16.670000 9.650000 ;
      LAYER met4 ;
        RECT 16.350000 9.330000 16.670000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 9.760000 16.670000 10.080000 ;
      LAYER met4 ;
        RECT 16.350000 9.760000 16.670000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 10.190000 17.075000 10.510000 ;
      LAYER met4 ;
        RECT 16.755000 10.190000 17.075000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 10.620000 17.075000 10.940000 ;
      LAYER met4 ;
        RECT 16.755000 10.620000 17.075000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 11.050000 17.075000 11.370000 ;
      LAYER met4 ;
        RECT 16.755000 11.050000 17.075000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 11.480000 17.075000 11.800000 ;
      LAYER met4 ;
        RECT 16.755000 11.480000 17.075000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 11.910000 17.075000 12.230000 ;
      LAYER met4 ;
        RECT 16.755000 11.910000 17.075000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 12.340000 17.075000 12.660000 ;
      LAYER met4 ;
        RECT 16.755000 12.340000 17.075000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 12.770000 17.075000 13.090000 ;
      LAYER met4 ;
        RECT 16.755000 12.770000 17.075000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 13.200000 17.075000 13.520000 ;
      LAYER met4 ;
        RECT 16.755000 13.200000 17.075000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 8.900000 17.075000 9.220000 ;
      LAYER met4 ;
        RECT 16.755000 8.900000 17.075000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 9.330000 17.075000 9.650000 ;
      LAYER met4 ;
        RECT 16.755000 9.330000 17.075000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 9.760000 17.075000 10.080000 ;
      LAYER met4 ;
        RECT 16.755000 9.760000 17.075000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 10.190000 17.480000 10.510000 ;
      LAYER met4 ;
        RECT 17.160000 10.190000 17.480000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 10.620000 17.480000 10.940000 ;
      LAYER met4 ;
        RECT 17.160000 10.620000 17.480000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 11.050000 17.480000 11.370000 ;
      LAYER met4 ;
        RECT 17.160000 11.050000 17.480000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 11.480000 17.480000 11.800000 ;
      LAYER met4 ;
        RECT 17.160000 11.480000 17.480000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 11.910000 17.480000 12.230000 ;
      LAYER met4 ;
        RECT 17.160000 11.910000 17.480000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 12.340000 17.480000 12.660000 ;
      LAYER met4 ;
        RECT 17.160000 12.340000 17.480000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 12.770000 17.480000 13.090000 ;
      LAYER met4 ;
        RECT 17.160000 12.770000 17.480000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 13.200000 17.480000 13.520000 ;
      LAYER met4 ;
        RECT 17.160000 13.200000 17.480000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 8.900000 17.480000 9.220000 ;
      LAYER met4 ;
        RECT 17.160000 8.900000 17.480000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 9.330000 17.480000 9.650000 ;
      LAYER met4 ;
        RECT 17.160000 9.330000 17.480000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 9.760000 17.480000 10.080000 ;
      LAYER met4 ;
        RECT 17.160000 9.760000 17.480000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 10.190000 17.885000 10.510000 ;
      LAYER met4 ;
        RECT 17.565000 10.190000 17.885000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 10.620000 17.885000 10.940000 ;
      LAYER met4 ;
        RECT 17.565000 10.620000 17.885000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 11.050000 17.885000 11.370000 ;
      LAYER met4 ;
        RECT 17.565000 11.050000 17.885000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 11.480000 17.885000 11.800000 ;
      LAYER met4 ;
        RECT 17.565000 11.480000 17.885000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 11.910000 17.885000 12.230000 ;
      LAYER met4 ;
        RECT 17.565000 11.910000 17.885000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 12.340000 17.885000 12.660000 ;
      LAYER met4 ;
        RECT 17.565000 12.340000 17.885000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 12.770000 17.885000 13.090000 ;
      LAYER met4 ;
        RECT 17.565000 12.770000 17.885000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 13.200000 17.885000 13.520000 ;
      LAYER met4 ;
        RECT 17.565000 13.200000 17.885000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 8.900000 17.885000 9.220000 ;
      LAYER met4 ;
        RECT 17.565000 8.900000 17.885000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 9.330000 17.885000 9.650000 ;
      LAYER met4 ;
        RECT 17.565000 9.330000 17.885000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 9.760000 17.885000 10.080000 ;
      LAYER met4 ;
        RECT 17.565000 9.760000 17.885000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 10.190000 18.290000 10.510000 ;
      LAYER met4 ;
        RECT 17.970000 10.190000 18.290000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 10.620000 18.290000 10.940000 ;
      LAYER met4 ;
        RECT 17.970000 10.620000 18.290000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 11.050000 18.290000 11.370000 ;
      LAYER met4 ;
        RECT 17.970000 11.050000 18.290000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 11.480000 18.290000 11.800000 ;
      LAYER met4 ;
        RECT 17.970000 11.480000 18.290000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 11.910000 18.290000 12.230000 ;
      LAYER met4 ;
        RECT 17.970000 11.910000 18.290000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 12.340000 18.290000 12.660000 ;
      LAYER met4 ;
        RECT 17.970000 12.340000 18.290000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 12.770000 18.290000 13.090000 ;
      LAYER met4 ;
        RECT 17.970000 12.770000 18.290000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 13.200000 18.290000 13.520000 ;
      LAYER met4 ;
        RECT 17.970000 13.200000 18.290000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 8.900000 18.290000 9.220000 ;
      LAYER met4 ;
        RECT 17.970000 8.900000 18.290000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 9.330000 18.290000 9.650000 ;
      LAYER met4 ;
        RECT 17.970000 9.330000 18.290000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 9.760000 18.290000 10.080000 ;
      LAYER met4 ;
        RECT 17.970000 9.760000 18.290000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 10.190000 18.695000 10.510000 ;
      LAYER met4 ;
        RECT 18.375000 10.190000 18.695000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 10.620000 18.695000 10.940000 ;
      LAYER met4 ;
        RECT 18.375000 10.620000 18.695000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 11.050000 18.695000 11.370000 ;
      LAYER met4 ;
        RECT 18.375000 11.050000 18.695000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 11.480000 18.695000 11.800000 ;
      LAYER met4 ;
        RECT 18.375000 11.480000 18.695000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 11.910000 18.695000 12.230000 ;
      LAYER met4 ;
        RECT 18.375000 11.910000 18.695000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 12.340000 18.695000 12.660000 ;
      LAYER met4 ;
        RECT 18.375000 12.340000 18.695000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 12.770000 18.695000 13.090000 ;
      LAYER met4 ;
        RECT 18.375000 12.770000 18.695000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 13.200000 18.695000 13.520000 ;
      LAYER met4 ;
        RECT 18.375000 13.200000 18.695000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 8.900000 18.695000 9.220000 ;
      LAYER met4 ;
        RECT 18.375000 8.900000 18.695000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 9.330000 18.695000 9.650000 ;
      LAYER met4 ;
        RECT 18.375000 9.330000 18.695000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 9.760000 18.695000 10.080000 ;
      LAYER met4 ;
        RECT 18.375000 9.760000 18.695000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 10.190000 19.100000 10.510000 ;
      LAYER met4 ;
        RECT 18.780000 10.190000 19.100000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 10.620000 19.100000 10.940000 ;
      LAYER met4 ;
        RECT 18.780000 10.620000 19.100000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 11.050000 19.100000 11.370000 ;
      LAYER met4 ;
        RECT 18.780000 11.050000 19.100000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 11.480000 19.100000 11.800000 ;
      LAYER met4 ;
        RECT 18.780000 11.480000 19.100000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 11.910000 19.100000 12.230000 ;
      LAYER met4 ;
        RECT 18.780000 11.910000 19.100000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 12.340000 19.100000 12.660000 ;
      LAYER met4 ;
        RECT 18.780000 12.340000 19.100000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 12.770000 19.100000 13.090000 ;
      LAYER met4 ;
        RECT 18.780000 12.770000 19.100000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 13.200000 19.100000 13.520000 ;
      LAYER met4 ;
        RECT 18.780000 13.200000 19.100000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 8.900000 19.100000 9.220000 ;
      LAYER met4 ;
        RECT 18.780000 8.900000 19.100000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 9.330000 19.100000 9.650000 ;
      LAYER met4 ;
        RECT 18.780000 9.330000 19.100000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 9.760000 19.100000 10.080000 ;
      LAYER met4 ;
        RECT 18.780000 9.760000 19.100000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 10.190000 19.505000 10.510000 ;
      LAYER met4 ;
        RECT 19.185000 10.190000 19.505000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 10.620000 19.505000 10.940000 ;
      LAYER met4 ;
        RECT 19.185000 10.620000 19.505000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 11.050000 19.505000 11.370000 ;
      LAYER met4 ;
        RECT 19.185000 11.050000 19.505000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 11.480000 19.505000 11.800000 ;
      LAYER met4 ;
        RECT 19.185000 11.480000 19.505000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 11.910000 19.505000 12.230000 ;
      LAYER met4 ;
        RECT 19.185000 11.910000 19.505000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 12.340000 19.505000 12.660000 ;
      LAYER met4 ;
        RECT 19.185000 12.340000 19.505000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 12.770000 19.505000 13.090000 ;
      LAYER met4 ;
        RECT 19.185000 12.770000 19.505000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 13.200000 19.505000 13.520000 ;
      LAYER met4 ;
        RECT 19.185000 13.200000 19.505000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 8.900000 19.505000 9.220000 ;
      LAYER met4 ;
        RECT 19.185000 8.900000 19.505000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 9.330000 19.505000 9.650000 ;
      LAYER met4 ;
        RECT 19.185000 9.330000 19.505000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 9.760000 19.505000 10.080000 ;
      LAYER met4 ;
        RECT 19.185000 9.760000 19.505000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 10.190000 19.910000 10.510000 ;
      LAYER met4 ;
        RECT 19.590000 10.190000 19.910000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 10.620000 19.910000 10.940000 ;
      LAYER met4 ;
        RECT 19.590000 10.620000 19.910000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 11.050000 19.910000 11.370000 ;
      LAYER met4 ;
        RECT 19.590000 11.050000 19.910000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 11.480000 19.910000 11.800000 ;
      LAYER met4 ;
        RECT 19.590000 11.480000 19.910000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 11.910000 19.910000 12.230000 ;
      LAYER met4 ;
        RECT 19.590000 11.910000 19.910000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 12.340000 19.910000 12.660000 ;
      LAYER met4 ;
        RECT 19.590000 12.340000 19.910000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 12.770000 19.910000 13.090000 ;
      LAYER met4 ;
        RECT 19.590000 12.770000 19.910000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 13.200000 19.910000 13.520000 ;
      LAYER met4 ;
        RECT 19.590000 13.200000 19.910000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 8.900000 19.910000 9.220000 ;
      LAYER met4 ;
        RECT 19.590000 8.900000 19.910000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 9.330000 19.910000 9.650000 ;
      LAYER met4 ;
        RECT 19.590000 9.330000 19.910000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 9.760000 19.910000 10.080000 ;
      LAYER met4 ;
        RECT 19.590000 9.760000 19.910000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 10.190000 20.315000 10.510000 ;
      LAYER met4 ;
        RECT 19.995000 10.190000 20.315000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 10.620000 20.315000 10.940000 ;
      LAYER met4 ;
        RECT 19.995000 10.620000 20.315000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 11.050000 20.315000 11.370000 ;
      LAYER met4 ;
        RECT 19.995000 11.050000 20.315000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 11.480000 20.315000 11.800000 ;
      LAYER met4 ;
        RECT 19.995000 11.480000 20.315000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 11.910000 20.315000 12.230000 ;
      LAYER met4 ;
        RECT 19.995000 11.910000 20.315000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 12.340000 20.315000 12.660000 ;
      LAYER met4 ;
        RECT 19.995000 12.340000 20.315000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 12.770000 20.315000 13.090000 ;
      LAYER met4 ;
        RECT 19.995000 12.770000 20.315000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 13.200000 20.315000 13.520000 ;
      LAYER met4 ;
        RECT 19.995000 13.200000 20.315000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 8.900000 20.315000 9.220000 ;
      LAYER met4 ;
        RECT 19.995000 8.900000 20.315000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 9.330000 20.315000 9.650000 ;
      LAYER met4 ;
        RECT 19.995000 9.330000 20.315000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 9.760000 20.315000 10.080000 ;
      LAYER met4 ;
        RECT 19.995000 9.760000 20.315000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 10.190000 2.485000 10.510000 ;
      LAYER met4 ;
        RECT 2.165000 10.190000 2.485000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 10.620000 2.485000 10.940000 ;
      LAYER met4 ;
        RECT 2.165000 10.620000 2.485000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 11.050000 2.485000 11.370000 ;
      LAYER met4 ;
        RECT 2.165000 11.050000 2.485000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 11.480000 2.485000 11.800000 ;
      LAYER met4 ;
        RECT 2.165000 11.480000 2.485000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 11.910000 2.485000 12.230000 ;
      LAYER met4 ;
        RECT 2.165000 11.910000 2.485000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 12.340000 2.485000 12.660000 ;
      LAYER met4 ;
        RECT 2.165000 12.340000 2.485000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 12.770000 2.485000 13.090000 ;
      LAYER met4 ;
        RECT 2.165000 12.770000 2.485000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 13.200000 2.485000 13.520000 ;
      LAYER met4 ;
        RECT 2.165000 13.200000 2.485000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 8.900000 2.485000 9.220000 ;
      LAYER met4 ;
        RECT 2.165000 8.900000 2.485000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 9.330000 2.485000 9.650000 ;
      LAYER met4 ;
        RECT 2.165000 9.330000 2.485000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 9.760000 2.485000 10.080000 ;
      LAYER met4 ;
        RECT 2.165000 9.760000 2.485000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 10.190000 2.895000 10.510000 ;
      LAYER met4 ;
        RECT 2.575000 10.190000 2.895000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 10.620000 2.895000 10.940000 ;
      LAYER met4 ;
        RECT 2.575000 10.620000 2.895000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 11.050000 2.895000 11.370000 ;
      LAYER met4 ;
        RECT 2.575000 11.050000 2.895000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 11.480000 2.895000 11.800000 ;
      LAYER met4 ;
        RECT 2.575000 11.480000 2.895000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 11.910000 2.895000 12.230000 ;
      LAYER met4 ;
        RECT 2.575000 11.910000 2.895000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 12.340000 2.895000 12.660000 ;
      LAYER met4 ;
        RECT 2.575000 12.340000 2.895000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 12.770000 2.895000 13.090000 ;
      LAYER met4 ;
        RECT 2.575000 12.770000 2.895000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 13.200000 2.895000 13.520000 ;
      LAYER met4 ;
        RECT 2.575000 13.200000 2.895000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 8.900000 2.895000 9.220000 ;
      LAYER met4 ;
        RECT 2.575000 8.900000 2.895000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 9.330000 2.895000 9.650000 ;
      LAYER met4 ;
        RECT 2.575000 9.330000 2.895000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 9.760000 2.895000 10.080000 ;
      LAYER met4 ;
        RECT 2.575000 9.760000 2.895000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 10.190000 3.305000 10.510000 ;
      LAYER met4 ;
        RECT 2.985000 10.190000 3.305000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 10.620000 3.305000 10.940000 ;
      LAYER met4 ;
        RECT 2.985000 10.620000 3.305000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 11.050000 3.305000 11.370000 ;
      LAYER met4 ;
        RECT 2.985000 11.050000 3.305000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 11.480000 3.305000 11.800000 ;
      LAYER met4 ;
        RECT 2.985000 11.480000 3.305000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 11.910000 3.305000 12.230000 ;
      LAYER met4 ;
        RECT 2.985000 11.910000 3.305000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 12.340000 3.305000 12.660000 ;
      LAYER met4 ;
        RECT 2.985000 12.340000 3.305000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 12.770000 3.305000 13.090000 ;
      LAYER met4 ;
        RECT 2.985000 12.770000 3.305000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 13.200000 3.305000 13.520000 ;
      LAYER met4 ;
        RECT 2.985000 13.200000 3.305000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 8.900000 3.305000 9.220000 ;
      LAYER met4 ;
        RECT 2.985000 8.900000 3.305000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 9.330000 3.305000 9.650000 ;
      LAYER met4 ;
        RECT 2.985000 9.330000 3.305000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 9.760000 3.305000 10.080000 ;
      LAYER met4 ;
        RECT 2.985000 9.760000 3.305000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 10.190000 20.720000 10.510000 ;
      LAYER met4 ;
        RECT 20.400000 10.190000 20.720000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 10.620000 20.720000 10.940000 ;
      LAYER met4 ;
        RECT 20.400000 10.620000 20.720000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 11.050000 20.720000 11.370000 ;
      LAYER met4 ;
        RECT 20.400000 11.050000 20.720000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 11.480000 20.720000 11.800000 ;
      LAYER met4 ;
        RECT 20.400000 11.480000 20.720000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 11.910000 20.720000 12.230000 ;
      LAYER met4 ;
        RECT 20.400000 11.910000 20.720000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 12.340000 20.720000 12.660000 ;
      LAYER met4 ;
        RECT 20.400000 12.340000 20.720000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 12.770000 20.720000 13.090000 ;
      LAYER met4 ;
        RECT 20.400000 12.770000 20.720000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 13.200000 20.720000 13.520000 ;
      LAYER met4 ;
        RECT 20.400000 13.200000 20.720000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 8.900000 20.720000 9.220000 ;
      LAYER met4 ;
        RECT 20.400000 8.900000 20.720000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 9.330000 20.720000 9.650000 ;
      LAYER met4 ;
        RECT 20.400000 9.330000 20.720000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 9.760000 20.720000 10.080000 ;
      LAYER met4 ;
        RECT 20.400000 9.760000 20.720000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 10.190000 21.125000 10.510000 ;
      LAYER met4 ;
        RECT 20.805000 10.190000 21.125000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 10.620000 21.125000 10.940000 ;
      LAYER met4 ;
        RECT 20.805000 10.620000 21.125000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 11.050000 21.125000 11.370000 ;
      LAYER met4 ;
        RECT 20.805000 11.050000 21.125000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 11.480000 21.125000 11.800000 ;
      LAYER met4 ;
        RECT 20.805000 11.480000 21.125000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 11.910000 21.125000 12.230000 ;
      LAYER met4 ;
        RECT 20.805000 11.910000 21.125000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 12.340000 21.125000 12.660000 ;
      LAYER met4 ;
        RECT 20.805000 12.340000 21.125000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 12.770000 21.125000 13.090000 ;
      LAYER met4 ;
        RECT 20.805000 12.770000 21.125000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 13.200000 21.125000 13.520000 ;
      LAYER met4 ;
        RECT 20.805000 13.200000 21.125000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 8.900000 21.125000 9.220000 ;
      LAYER met4 ;
        RECT 20.805000 8.900000 21.125000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 9.330000 21.125000 9.650000 ;
      LAYER met4 ;
        RECT 20.805000 9.330000 21.125000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 9.760000 21.125000 10.080000 ;
      LAYER met4 ;
        RECT 20.805000 9.760000 21.125000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 10.190000 21.530000 10.510000 ;
      LAYER met4 ;
        RECT 21.210000 10.190000 21.530000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 10.620000 21.530000 10.940000 ;
      LAYER met4 ;
        RECT 21.210000 10.620000 21.530000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 11.050000 21.530000 11.370000 ;
      LAYER met4 ;
        RECT 21.210000 11.050000 21.530000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 11.480000 21.530000 11.800000 ;
      LAYER met4 ;
        RECT 21.210000 11.480000 21.530000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 11.910000 21.530000 12.230000 ;
      LAYER met4 ;
        RECT 21.210000 11.910000 21.530000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 12.340000 21.530000 12.660000 ;
      LAYER met4 ;
        RECT 21.210000 12.340000 21.530000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 12.770000 21.530000 13.090000 ;
      LAYER met4 ;
        RECT 21.210000 12.770000 21.530000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 13.200000 21.530000 13.520000 ;
      LAYER met4 ;
        RECT 21.210000 13.200000 21.530000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 8.900000 21.530000 9.220000 ;
      LAYER met4 ;
        RECT 21.210000 8.900000 21.530000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 9.330000 21.530000 9.650000 ;
      LAYER met4 ;
        RECT 21.210000 9.330000 21.530000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 9.760000 21.530000 10.080000 ;
      LAYER met4 ;
        RECT 21.210000 9.760000 21.530000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 10.190000 21.935000 10.510000 ;
      LAYER met4 ;
        RECT 21.615000 10.190000 21.935000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 10.620000 21.935000 10.940000 ;
      LAYER met4 ;
        RECT 21.615000 10.620000 21.935000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 11.050000 21.935000 11.370000 ;
      LAYER met4 ;
        RECT 21.615000 11.050000 21.935000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 11.480000 21.935000 11.800000 ;
      LAYER met4 ;
        RECT 21.615000 11.480000 21.935000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 11.910000 21.935000 12.230000 ;
      LAYER met4 ;
        RECT 21.615000 11.910000 21.935000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 12.340000 21.935000 12.660000 ;
      LAYER met4 ;
        RECT 21.615000 12.340000 21.935000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 12.770000 21.935000 13.090000 ;
      LAYER met4 ;
        RECT 21.615000 12.770000 21.935000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 13.200000 21.935000 13.520000 ;
      LAYER met4 ;
        RECT 21.615000 13.200000 21.935000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 8.900000 21.935000 9.220000 ;
      LAYER met4 ;
        RECT 21.615000 8.900000 21.935000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 9.330000 21.935000 9.650000 ;
      LAYER met4 ;
        RECT 21.615000 9.330000 21.935000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 9.760000 21.935000 10.080000 ;
      LAYER met4 ;
        RECT 21.615000 9.760000 21.935000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 10.190000 22.340000 10.510000 ;
      LAYER met4 ;
        RECT 22.020000 10.190000 22.340000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 10.620000 22.340000 10.940000 ;
      LAYER met4 ;
        RECT 22.020000 10.620000 22.340000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 11.050000 22.340000 11.370000 ;
      LAYER met4 ;
        RECT 22.020000 11.050000 22.340000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 11.480000 22.340000 11.800000 ;
      LAYER met4 ;
        RECT 22.020000 11.480000 22.340000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 11.910000 22.340000 12.230000 ;
      LAYER met4 ;
        RECT 22.020000 11.910000 22.340000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 12.340000 22.340000 12.660000 ;
      LAYER met4 ;
        RECT 22.020000 12.340000 22.340000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 12.770000 22.340000 13.090000 ;
      LAYER met4 ;
        RECT 22.020000 12.770000 22.340000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 13.200000 22.340000 13.520000 ;
      LAYER met4 ;
        RECT 22.020000 13.200000 22.340000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 8.900000 22.340000 9.220000 ;
      LAYER met4 ;
        RECT 22.020000 8.900000 22.340000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 9.330000 22.340000 9.650000 ;
      LAYER met4 ;
        RECT 22.020000 9.330000 22.340000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 9.760000 22.340000 10.080000 ;
      LAYER met4 ;
        RECT 22.020000 9.760000 22.340000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 10.190000 22.745000 10.510000 ;
      LAYER met4 ;
        RECT 22.425000 10.190000 22.745000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 10.620000 22.745000 10.940000 ;
      LAYER met4 ;
        RECT 22.425000 10.620000 22.745000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 11.050000 22.745000 11.370000 ;
      LAYER met4 ;
        RECT 22.425000 11.050000 22.745000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 11.480000 22.745000 11.800000 ;
      LAYER met4 ;
        RECT 22.425000 11.480000 22.745000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 11.910000 22.745000 12.230000 ;
      LAYER met4 ;
        RECT 22.425000 11.910000 22.745000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 12.340000 22.745000 12.660000 ;
      LAYER met4 ;
        RECT 22.425000 12.340000 22.745000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 12.770000 22.745000 13.090000 ;
      LAYER met4 ;
        RECT 22.425000 12.770000 22.745000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 13.200000 22.745000 13.520000 ;
      LAYER met4 ;
        RECT 22.425000 13.200000 22.745000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 8.900000 22.745000 9.220000 ;
      LAYER met4 ;
        RECT 22.425000 8.900000 22.745000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 9.330000 22.745000 9.650000 ;
      LAYER met4 ;
        RECT 22.425000 9.330000 22.745000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 9.760000 22.745000 10.080000 ;
      LAYER met4 ;
        RECT 22.425000 9.760000 22.745000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 10.190000 23.150000 10.510000 ;
      LAYER met4 ;
        RECT 22.830000 10.190000 23.150000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 10.620000 23.150000 10.940000 ;
      LAYER met4 ;
        RECT 22.830000 10.620000 23.150000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 11.050000 23.150000 11.370000 ;
      LAYER met4 ;
        RECT 22.830000 11.050000 23.150000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 11.480000 23.150000 11.800000 ;
      LAYER met4 ;
        RECT 22.830000 11.480000 23.150000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 11.910000 23.150000 12.230000 ;
      LAYER met4 ;
        RECT 22.830000 11.910000 23.150000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 12.340000 23.150000 12.660000 ;
      LAYER met4 ;
        RECT 22.830000 12.340000 23.150000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 12.770000 23.150000 13.090000 ;
      LAYER met4 ;
        RECT 22.830000 12.770000 23.150000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 13.200000 23.150000 13.520000 ;
      LAYER met4 ;
        RECT 22.830000 13.200000 23.150000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 8.900000 23.150000 9.220000 ;
      LAYER met4 ;
        RECT 22.830000 8.900000 23.150000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 9.330000 23.150000 9.650000 ;
      LAYER met4 ;
        RECT 22.830000 9.330000 23.150000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 9.760000 23.150000 10.080000 ;
      LAYER met4 ;
        RECT 22.830000 9.760000 23.150000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 10.190000 23.555000 10.510000 ;
      LAYER met4 ;
        RECT 23.235000 10.190000 23.555000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 10.620000 23.555000 10.940000 ;
      LAYER met4 ;
        RECT 23.235000 10.620000 23.555000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 11.050000 23.555000 11.370000 ;
      LAYER met4 ;
        RECT 23.235000 11.050000 23.555000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 11.480000 23.555000 11.800000 ;
      LAYER met4 ;
        RECT 23.235000 11.480000 23.555000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 11.910000 23.555000 12.230000 ;
      LAYER met4 ;
        RECT 23.235000 11.910000 23.555000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 12.340000 23.555000 12.660000 ;
      LAYER met4 ;
        RECT 23.235000 12.340000 23.555000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 12.770000 23.555000 13.090000 ;
      LAYER met4 ;
        RECT 23.235000 12.770000 23.555000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 13.200000 23.555000 13.520000 ;
      LAYER met4 ;
        RECT 23.235000 13.200000 23.555000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 8.900000 23.555000 9.220000 ;
      LAYER met4 ;
        RECT 23.235000 8.900000 23.555000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 9.330000 23.555000 9.650000 ;
      LAYER met4 ;
        RECT 23.235000 9.330000 23.555000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 9.760000 23.555000 10.080000 ;
      LAYER met4 ;
        RECT 23.235000 9.760000 23.555000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 10.190000 23.960000 10.510000 ;
      LAYER met4 ;
        RECT 23.640000 10.190000 23.960000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 10.620000 23.960000 10.940000 ;
      LAYER met4 ;
        RECT 23.640000 10.620000 23.960000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 11.050000 23.960000 11.370000 ;
      LAYER met4 ;
        RECT 23.640000 11.050000 23.960000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 11.480000 23.960000 11.800000 ;
      LAYER met4 ;
        RECT 23.640000 11.480000 23.960000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 11.910000 23.960000 12.230000 ;
      LAYER met4 ;
        RECT 23.640000 11.910000 23.960000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 12.340000 23.960000 12.660000 ;
      LAYER met4 ;
        RECT 23.640000 12.340000 23.960000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 12.770000 23.960000 13.090000 ;
      LAYER met4 ;
        RECT 23.640000 12.770000 23.960000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 13.200000 23.960000 13.520000 ;
      LAYER met4 ;
        RECT 23.640000 13.200000 23.960000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 8.900000 23.960000 9.220000 ;
      LAYER met4 ;
        RECT 23.640000 8.900000 23.960000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 9.330000 23.960000 9.650000 ;
      LAYER met4 ;
        RECT 23.640000 9.330000 23.960000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 9.760000 23.960000 10.080000 ;
      LAYER met4 ;
        RECT 23.640000 9.760000 23.960000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 10.190000 24.365000 10.510000 ;
      LAYER met4 ;
        RECT 24.045000 10.190000 24.365000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 10.620000 24.365000 10.940000 ;
      LAYER met4 ;
        RECT 24.045000 10.620000 24.365000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 11.050000 24.365000 11.370000 ;
      LAYER met4 ;
        RECT 24.045000 11.050000 24.365000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 11.480000 24.365000 11.800000 ;
      LAYER met4 ;
        RECT 24.045000 11.480000 24.365000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 11.910000 24.365000 12.230000 ;
      LAYER met4 ;
        RECT 24.045000 11.910000 24.365000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 12.340000 24.365000 12.660000 ;
      LAYER met4 ;
        RECT 24.045000 12.340000 24.365000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 12.770000 24.365000 13.090000 ;
      LAYER met4 ;
        RECT 24.045000 12.770000 24.365000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 13.200000 24.365000 13.520000 ;
      LAYER met4 ;
        RECT 24.045000 13.200000 24.365000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 8.900000 24.365000 9.220000 ;
      LAYER met4 ;
        RECT 24.045000 8.900000 24.365000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 9.330000 24.365000 9.650000 ;
      LAYER met4 ;
        RECT 24.045000 9.330000 24.365000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 9.760000 24.365000 10.080000 ;
      LAYER met4 ;
        RECT 24.045000 9.760000 24.365000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 10.190000 3.710000 10.510000 ;
      LAYER met4 ;
        RECT 3.390000 10.190000 3.710000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 10.620000 3.710000 10.940000 ;
      LAYER met4 ;
        RECT 3.390000 10.620000 3.710000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 11.050000 3.710000 11.370000 ;
      LAYER met4 ;
        RECT 3.390000 11.050000 3.710000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 11.480000 3.710000 11.800000 ;
      LAYER met4 ;
        RECT 3.390000 11.480000 3.710000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 11.910000 3.710000 12.230000 ;
      LAYER met4 ;
        RECT 3.390000 11.910000 3.710000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 12.340000 3.710000 12.660000 ;
      LAYER met4 ;
        RECT 3.390000 12.340000 3.710000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 12.770000 3.710000 13.090000 ;
      LAYER met4 ;
        RECT 3.390000 12.770000 3.710000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 13.200000 3.710000 13.520000 ;
      LAYER met4 ;
        RECT 3.390000 13.200000 3.710000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 8.900000 3.710000 9.220000 ;
      LAYER met4 ;
        RECT 3.390000 8.900000 3.710000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 9.330000 3.710000 9.650000 ;
      LAYER met4 ;
        RECT 3.390000 9.330000 3.710000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 9.760000 3.710000 10.080000 ;
      LAYER met4 ;
        RECT 3.390000 9.760000 3.710000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 10.190000 4.115000 10.510000 ;
      LAYER met4 ;
        RECT 3.795000 10.190000 4.115000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 10.620000 4.115000 10.940000 ;
      LAYER met4 ;
        RECT 3.795000 10.620000 4.115000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 11.050000 4.115000 11.370000 ;
      LAYER met4 ;
        RECT 3.795000 11.050000 4.115000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 11.480000 4.115000 11.800000 ;
      LAYER met4 ;
        RECT 3.795000 11.480000 4.115000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 11.910000 4.115000 12.230000 ;
      LAYER met4 ;
        RECT 3.795000 11.910000 4.115000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 12.340000 4.115000 12.660000 ;
      LAYER met4 ;
        RECT 3.795000 12.340000 4.115000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 12.770000 4.115000 13.090000 ;
      LAYER met4 ;
        RECT 3.795000 12.770000 4.115000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 13.200000 4.115000 13.520000 ;
      LAYER met4 ;
        RECT 3.795000 13.200000 4.115000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 8.900000 4.115000 9.220000 ;
      LAYER met4 ;
        RECT 3.795000 8.900000 4.115000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 9.330000 4.115000 9.650000 ;
      LAYER met4 ;
        RECT 3.795000 9.330000 4.115000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 9.760000 4.115000 10.080000 ;
      LAYER met4 ;
        RECT 3.795000 9.760000 4.115000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 10.190000 4.520000 10.510000 ;
      LAYER met4 ;
        RECT 4.200000 10.190000 4.520000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 10.620000 4.520000 10.940000 ;
      LAYER met4 ;
        RECT 4.200000 10.620000 4.520000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 11.050000 4.520000 11.370000 ;
      LAYER met4 ;
        RECT 4.200000 11.050000 4.520000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 11.480000 4.520000 11.800000 ;
      LAYER met4 ;
        RECT 4.200000 11.480000 4.520000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 11.910000 4.520000 12.230000 ;
      LAYER met4 ;
        RECT 4.200000 11.910000 4.520000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 12.340000 4.520000 12.660000 ;
      LAYER met4 ;
        RECT 4.200000 12.340000 4.520000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 12.770000 4.520000 13.090000 ;
      LAYER met4 ;
        RECT 4.200000 12.770000 4.520000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 13.200000 4.520000 13.520000 ;
      LAYER met4 ;
        RECT 4.200000 13.200000 4.520000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 8.900000 4.520000 9.220000 ;
      LAYER met4 ;
        RECT 4.200000 8.900000 4.520000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 9.330000 4.520000 9.650000 ;
      LAYER met4 ;
        RECT 4.200000 9.330000 4.520000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 9.760000 4.520000 10.080000 ;
      LAYER met4 ;
        RECT 4.200000 9.760000 4.520000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 10.190000 4.925000 10.510000 ;
      LAYER met4 ;
        RECT 4.605000 10.190000 4.925000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 10.620000 4.925000 10.940000 ;
      LAYER met4 ;
        RECT 4.605000 10.620000 4.925000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 11.050000 4.925000 11.370000 ;
      LAYER met4 ;
        RECT 4.605000 11.050000 4.925000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 11.480000 4.925000 11.800000 ;
      LAYER met4 ;
        RECT 4.605000 11.480000 4.925000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 11.910000 4.925000 12.230000 ;
      LAYER met4 ;
        RECT 4.605000 11.910000 4.925000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 12.340000 4.925000 12.660000 ;
      LAYER met4 ;
        RECT 4.605000 12.340000 4.925000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 12.770000 4.925000 13.090000 ;
      LAYER met4 ;
        RECT 4.605000 12.770000 4.925000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 13.200000 4.925000 13.520000 ;
      LAYER met4 ;
        RECT 4.605000 13.200000 4.925000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 8.900000 4.925000 9.220000 ;
      LAYER met4 ;
        RECT 4.605000 8.900000 4.925000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 9.330000 4.925000 9.650000 ;
      LAYER met4 ;
        RECT 4.605000 9.330000 4.925000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 9.760000 4.925000 10.080000 ;
      LAYER met4 ;
        RECT 4.605000 9.760000 4.925000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 10.190000 5.330000 10.510000 ;
      LAYER met4 ;
        RECT 5.010000 10.190000 5.330000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 10.620000 5.330000 10.940000 ;
      LAYER met4 ;
        RECT 5.010000 10.620000 5.330000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 11.050000 5.330000 11.370000 ;
      LAYER met4 ;
        RECT 5.010000 11.050000 5.330000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 11.480000 5.330000 11.800000 ;
      LAYER met4 ;
        RECT 5.010000 11.480000 5.330000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 11.910000 5.330000 12.230000 ;
      LAYER met4 ;
        RECT 5.010000 11.910000 5.330000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 12.340000 5.330000 12.660000 ;
      LAYER met4 ;
        RECT 5.010000 12.340000 5.330000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 12.770000 5.330000 13.090000 ;
      LAYER met4 ;
        RECT 5.010000 12.770000 5.330000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 13.200000 5.330000 13.520000 ;
      LAYER met4 ;
        RECT 5.010000 13.200000 5.330000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 8.900000 5.330000 9.220000 ;
      LAYER met4 ;
        RECT 5.010000 8.900000 5.330000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 9.330000 5.330000 9.650000 ;
      LAYER met4 ;
        RECT 5.010000 9.330000 5.330000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 9.760000 5.330000 10.080000 ;
      LAYER met4 ;
        RECT 5.010000 9.760000 5.330000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 10.190000 5.735000 10.510000 ;
      LAYER met4 ;
        RECT 5.415000 10.190000 5.735000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 10.620000 5.735000 10.940000 ;
      LAYER met4 ;
        RECT 5.415000 10.620000 5.735000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 11.050000 5.735000 11.370000 ;
      LAYER met4 ;
        RECT 5.415000 11.050000 5.735000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 11.480000 5.735000 11.800000 ;
      LAYER met4 ;
        RECT 5.415000 11.480000 5.735000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 11.910000 5.735000 12.230000 ;
      LAYER met4 ;
        RECT 5.415000 11.910000 5.735000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 12.340000 5.735000 12.660000 ;
      LAYER met4 ;
        RECT 5.415000 12.340000 5.735000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 12.770000 5.735000 13.090000 ;
      LAYER met4 ;
        RECT 5.415000 12.770000 5.735000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 13.200000 5.735000 13.520000 ;
      LAYER met4 ;
        RECT 5.415000 13.200000 5.735000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 8.900000 5.735000 9.220000 ;
      LAYER met4 ;
        RECT 5.415000 8.900000 5.735000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 9.330000 5.735000 9.650000 ;
      LAYER met4 ;
        RECT 5.415000 9.330000 5.735000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 9.760000 5.735000 10.080000 ;
      LAYER met4 ;
        RECT 5.415000 9.760000 5.735000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 10.190000 6.140000 10.510000 ;
      LAYER met4 ;
        RECT 5.820000 10.190000 6.140000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 10.620000 6.140000 10.940000 ;
      LAYER met4 ;
        RECT 5.820000 10.620000 6.140000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 11.050000 6.140000 11.370000 ;
      LAYER met4 ;
        RECT 5.820000 11.050000 6.140000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 11.480000 6.140000 11.800000 ;
      LAYER met4 ;
        RECT 5.820000 11.480000 6.140000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 11.910000 6.140000 12.230000 ;
      LAYER met4 ;
        RECT 5.820000 11.910000 6.140000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 12.340000 6.140000 12.660000 ;
      LAYER met4 ;
        RECT 5.820000 12.340000 6.140000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 12.770000 6.140000 13.090000 ;
      LAYER met4 ;
        RECT 5.820000 12.770000 6.140000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 13.200000 6.140000 13.520000 ;
      LAYER met4 ;
        RECT 5.820000 13.200000 6.140000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 8.900000 6.140000 9.220000 ;
      LAYER met4 ;
        RECT 5.820000 8.900000 6.140000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 9.330000 6.140000 9.650000 ;
      LAYER met4 ;
        RECT 5.820000 9.330000 6.140000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 9.760000 6.140000 10.080000 ;
      LAYER met4 ;
        RECT 5.820000 9.760000 6.140000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 10.190000 50.740000 10.510000 ;
      LAYER met4 ;
        RECT 50.420000 10.190000 50.740000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 10.620000 50.740000 10.940000 ;
      LAYER met4 ;
        RECT 50.420000 10.620000 50.740000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 11.050000 50.740000 11.370000 ;
      LAYER met4 ;
        RECT 50.420000 11.050000 50.740000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 11.480000 50.740000 11.800000 ;
      LAYER met4 ;
        RECT 50.420000 11.480000 50.740000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 11.910000 50.740000 12.230000 ;
      LAYER met4 ;
        RECT 50.420000 11.910000 50.740000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 12.340000 50.740000 12.660000 ;
      LAYER met4 ;
        RECT 50.420000 12.340000 50.740000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 12.770000 50.740000 13.090000 ;
      LAYER met4 ;
        RECT 50.420000 12.770000 50.740000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 13.200000 50.740000 13.520000 ;
      LAYER met4 ;
        RECT 50.420000 13.200000 50.740000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 8.900000 50.740000 9.220000 ;
      LAYER met4 ;
        RECT 50.420000 8.900000 50.740000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 9.330000 50.740000 9.650000 ;
      LAYER met4 ;
        RECT 50.420000 9.330000 50.740000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 9.760000 50.740000 10.080000 ;
      LAYER met4 ;
        RECT 50.420000 9.760000 50.740000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 10.190000 51.150000 10.510000 ;
      LAYER met4 ;
        RECT 50.830000 10.190000 51.150000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 10.620000 51.150000 10.940000 ;
      LAYER met4 ;
        RECT 50.830000 10.620000 51.150000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 11.050000 51.150000 11.370000 ;
      LAYER met4 ;
        RECT 50.830000 11.050000 51.150000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 11.480000 51.150000 11.800000 ;
      LAYER met4 ;
        RECT 50.830000 11.480000 51.150000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 11.910000 51.150000 12.230000 ;
      LAYER met4 ;
        RECT 50.830000 11.910000 51.150000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 12.340000 51.150000 12.660000 ;
      LAYER met4 ;
        RECT 50.830000 12.340000 51.150000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 12.770000 51.150000 13.090000 ;
      LAYER met4 ;
        RECT 50.830000 12.770000 51.150000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 13.200000 51.150000 13.520000 ;
      LAYER met4 ;
        RECT 50.830000 13.200000 51.150000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 8.900000 51.150000 9.220000 ;
      LAYER met4 ;
        RECT 50.830000 8.900000 51.150000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 9.330000 51.150000 9.650000 ;
      LAYER met4 ;
        RECT 50.830000 9.330000 51.150000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 9.760000 51.150000 10.080000 ;
      LAYER met4 ;
        RECT 50.830000 9.760000 51.150000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 10.190000 51.560000 10.510000 ;
      LAYER met4 ;
        RECT 51.240000 10.190000 51.560000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 10.620000 51.560000 10.940000 ;
      LAYER met4 ;
        RECT 51.240000 10.620000 51.560000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 11.050000 51.560000 11.370000 ;
      LAYER met4 ;
        RECT 51.240000 11.050000 51.560000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 11.480000 51.560000 11.800000 ;
      LAYER met4 ;
        RECT 51.240000 11.480000 51.560000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 11.910000 51.560000 12.230000 ;
      LAYER met4 ;
        RECT 51.240000 11.910000 51.560000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 12.340000 51.560000 12.660000 ;
      LAYER met4 ;
        RECT 51.240000 12.340000 51.560000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 12.770000 51.560000 13.090000 ;
      LAYER met4 ;
        RECT 51.240000 12.770000 51.560000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 13.200000 51.560000 13.520000 ;
      LAYER met4 ;
        RECT 51.240000 13.200000 51.560000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 8.900000 51.560000 9.220000 ;
      LAYER met4 ;
        RECT 51.240000 8.900000 51.560000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 9.330000 51.560000 9.650000 ;
      LAYER met4 ;
        RECT 51.240000 9.330000 51.560000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 9.760000 51.560000 10.080000 ;
      LAYER met4 ;
        RECT 51.240000 9.760000 51.560000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 10.190000 51.970000 10.510000 ;
      LAYER met4 ;
        RECT 51.650000 10.190000 51.970000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 10.620000 51.970000 10.940000 ;
      LAYER met4 ;
        RECT 51.650000 10.620000 51.970000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 11.050000 51.970000 11.370000 ;
      LAYER met4 ;
        RECT 51.650000 11.050000 51.970000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 11.480000 51.970000 11.800000 ;
      LAYER met4 ;
        RECT 51.650000 11.480000 51.970000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 11.910000 51.970000 12.230000 ;
      LAYER met4 ;
        RECT 51.650000 11.910000 51.970000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 12.340000 51.970000 12.660000 ;
      LAYER met4 ;
        RECT 51.650000 12.340000 51.970000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 12.770000 51.970000 13.090000 ;
      LAYER met4 ;
        RECT 51.650000 12.770000 51.970000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 13.200000 51.970000 13.520000 ;
      LAYER met4 ;
        RECT 51.650000 13.200000 51.970000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 8.900000 51.970000 9.220000 ;
      LAYER met4 ;
        RECT 51.650000 8.900000 51.970000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 9.330000 51.970000 9.650000 ;
      LAYER met4 ;
        RECT 51.650000 9.330000 51.970000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 9.760000 51.970000 10.080000 ;
      LAYER met4 ;
        RECT 51.650000 9.760000 51.970000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 10.190000 52.380000 10.510000 ;
      LAYER met4 ;
        RECT 52.060000 10.190000 52.380000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 10.620000 52.380000 10.940000 ;
      LAYER met4 ;
        RECT 52.060000 10.620000 52.380000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 11.050000 52.380000 11.370000 ;
      LAYER met4 ;
        RECT 52.060000 11.050000 52.380000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 11.480000 52.380000 11.800000 ;
      LAYER met4 ;
        RECT 52.060000 11.480000 52.380000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 11.910000 52.380000 12.230000 ;
      LAYER met4 ;
        RECT 52.060000 11.910000 52.380000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 12.340000 52.380000 12.660000 ;
      LAYER met4 ;
        RECT 52.060000 12.340000 52.380000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 12.770000 52.380000 13.090000 ;
      LAYER met4 ;
        RECT 52.060000 12.770000 52.380000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 13.200000 52.380000 13.520000 ;
      LAYER met4 ;
        RECT 52.060000 13.200000 52.380000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 8.900000 52.380000 9.220000 ;
      LAYER met4 ;
        RECT 52.060000 8.900000 52.380000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 9.330000 52.380000 9.650000 ;
      LAYER met4 ;
        RECT 52.060000 9.330000 52.380000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 9.760000 52.380000 10.080000 ;
      LAYER met4 ;
        RECT 52.060000 9.760000 52.380000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 10.190000 52.790000 10.510000 ;
      LAYER met4 ;
        RECT 52.470000 10.190000 52.790000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 10.620000 52.790000 10.940000 ;
      LAYER met4 ;
        RECT 52.470000 10.620000 52.790000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 11.050000 52.790000 11.370000 ;
      LAYER met4 ;
        RECT 52.470000 11.050000 52.790000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 11.480000 52.790000 11.800000 ;
      LAYER met4 ;
        RECT 52.470000 11.480000 52.790000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 11.910000 52.790000 12.230000 ;
      LAYER met4 ;
        RECT 52.470000 11.910000 52.790000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 12.340000 52.790000 12.660000 ;
      LAYER met4 ;
        RECT 52.470000 12.340000 52.790000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 12.770000 52.790000 13.090000 ;
      LAYER met4 ;
        RECT 52.470000 12.770000 52.790000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 13.200000 52.790000 13.520000 ;
      LAYER met4 ;
        RECT 52.470000 13.200000 52.790000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 8.900000 52.790000 9.220000 ;
      LAYER met4 ;
        RECT 52.470000 8.900000 52.790000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 9.330000 52.790000 9.650000 ;
      LAYER met4 ;
        RECT 52.470000 9.330000 52.790000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 9.760000 52.790000 10.080000 ;
      LAYER met4 ;
        RECT 52.470000 9.760000 52.790000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 10.190000 53.200000 10.510000 ;
      LAYER met4 ;
        RECT 52.880000 10.190000 53.200000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 10.620000 53.200000 10.940000 ;
      LAYER met4 ;
        RECT 52.880000 10.620000 53.200000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 11.050000 53.200000 11.370000 ;
      LAYER met4 ;
        RECT 52.880000 11.050000 53.200000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 11.480000 53.200000 11.800000 ;
      LAYER met4 ;
        RECT 52.880000 11.480000 53.200000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 11.910000 53.200000 12.230000 ;
      LAYER met4 ;
        RECT 52.880000 11.910000 53.200000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 12.340000 53.200000 12.660000 ;
      LAYER met4 ;
        RECT 52.880000 12.340000 53.200000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 12.770000 53.200000 13.090000 ;
      LAYER met4 ;
        RECT 52.880000 12.770000 53.200000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 13.200000 53.200000 13.520000 ;
      LAYER met4 ;
        RECT 52.880000 13.200000 53.200000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 8.900000 53.200000 9.220000 ;
      LAYER met4 ;
        RECT 52.880000 8.900000 53.200000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 9.330000 53.200000 9.650000 ;
      LAYER met4 ;
        RECT 52.880000 9.330000 53.200000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 9.760000 53.200000 10.080000 ;
      LAYER met4 ;
        RECT 52.880000 9.760000 53.200000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 10.190000 53.605000 10.510000 ;
      LAYER met4 ;
        RECT 53.285000 10.190000 53.605000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 10.620000 53.605000 10.940000 ;
      LAYER met4 ;
        RECT 53.285000 10.620000 53.605000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 11.050000 53.605000 11.370000 ;
      LAYER met4 ;
        RECT 53.285000 11.050000 53.605000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 11.480000 53.605000 11.800000 ;
      LAYER met4 ;
        RECT 53.285000 11.480000 53.605000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 11.910000 53.605000 12.230000 ;
      LAYER met4 ;
        RECT 53.285000 11.910000 53.605000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 12.340000 53.605000 12.660000 ;
      LAYER met4 ;
        RECT 53.285000 12.340000 53.605000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 12.770000 53.605000 13.090000 ;
      LAYER met4 ;
        RECT 53.285000 12.770000 53.605000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 13.200000 53.605000 13.520000 ;
      LAYER met4 ;
        RECT 53.285000 13.200000 53.605000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 8.900000 53.605000 9.220000 ;
      LAYER met4 ;
        RECT 53.285000 8.900000 53.605000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 9.330000 53.605000 9.650000 ;
      LAYER met4 ;
        RECT 53.285000 9.330000 53.605000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 9.760000 53.605000 10.080000 ;
      LAYER met4 ;
        RECT 53.285000 9.760000 53.605000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 10.190000 54.010000 10.510000 ;
      LAYER met4 ;
        RECT 53.690000 10.190000 54.010000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 10.620000 54.010000 10.940000 ;
      LAYER met4 ;
        RECT 53.690000 10.620000 54.010000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 11.050000 54.010000 11.370000 ;
      LAYER met4 ;
        RECT 53.690000 11.050000 54.010000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 11.480000 54.010000 11.800000 ;
      LAYER met4 ;
        RECT 53.690000 11.480000 54.010000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 11.910000 54.010000 12.230000 ;
      LAYER met4 ;
        RECT 53.690000 11.910000 54.010000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 12.340000 54.010000 12.660000 ;
      LAYER met4 ;
        RECT 53.690000 12.340000 54.010000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 12.770000 54.010000 13.090000 ;
      LAYER met4 ;
        RECT 53.690000 12.770000 54.010000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 13.200000 54.010000 13.520000 ;
      LAYER met4 ;
        RECT 53.690000 13.200000 54.010000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 8.900000 54.010000 9.220000 ;
      LAYER met4 ;
        RECT 53.690000 8.900000 54.010000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 9.330000 54.010000 9.650000 ;
      LAYER met4 ;
        RECT 53.690000 9.330000 54.010000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 9.760000 54.010000 10.080000 ;
      LAYER met4 ;
        RECT 53.690000 9.760000 54.010000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 10.190000 54.415000 10.510000 ;
      LAYER met4 ;
        RECT 54.095000 10.190000 54.415000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 10.620000 54.415000 10.940000 ;
      LAYER met4 ;
        RECT 54.095000 10.620000 54.415000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 11.050000 54.415000 11.370000 ;
      LAYER met4 ;
        RECT 54.095000 11.050000 54.415000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 11.480000 54.415000 11.800000 ;
      LAYER met4 ;
        RECT 54.095000 11.480000 54.415000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 11.910000 54.415000 12.230000 ;
      LAYER met4 ;
        RECT 54.095000 11.910000 54.415000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 12.340000 54.415000 12.660000 ;
      LAYER met4 ;
        RECT 54.095000 12.340000 54.415000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 12.770000 54.415000 13.090000 ;
      LAYER met4 ;
        RECT 54.095000 12.770000 54.415000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 13.200000 54.415000 13.520000 ;
      LAYER met4 ;
        RECT 54.095000 13.200000 54.415000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 8.900000 54.415000 9.220000 ;
      LAYER met4 ;
        RECT 54.095000 8.900000 54.415000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 9.330000 54.415000 9.650000 ;
      LAYER met4 ;
        RECT 54.095000 9.330000 54.415000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 9.760000 54.415000 10.080000 ;
      LAYER met4 ;
        RECT 54.095000 9.760000 54.415000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 10.190000 54.820000 10.510000 ;
      LAYER met4 ;
        RECT 54.500000 10.190000 54.820000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 10.620000 54.820000 10.940000 ;
      LAYER met4 ;
        RECT 54.500000 10.620000 54.820000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 11.050000 54.820000 11.370000 ;
      LAYER met4 ;
        RECT 54.500000 11.050000 54.820000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 11.480000 54.820000 11.800000 ;
      LAYER met4 ;
        RECT 54.500000 11.480000 54.820000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 11.910000 54.820000 12.230000 ;
      LAYER met4 ;
        RECT 54.500000 11.910000 54.820000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 12.340000 54.820000 12.660000 ;
      LAYER met4 ;
        RECT 54.500000 12.340000 54.820000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 12.770000 54.820000 13.090000 ;
      LAYER met4 ;
        RECT 54.500000 12.770000 54.820000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 13.200000 54.820000 13.520000 ;
      LAYER met4 ;
        RECT 54.500000 13.200000 54.820000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 8.900000 54.820000 9.220000 ;
      LAYER met4 ;
        RECT 54.500000 8.900000 54.820000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 9.330000 54.820000 9.650000 ;
      LAYER met4 ;
        RECT 54.500000 9.330000 54.820000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 9.760000 54.820000 10.080000 ;
      LAYER met4 ;
        RECT 54.500000 9.760000 54.820000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 10.190000 55.225000 10.510000 ;
      LAYER met4 ;
        RECT 54.905000 10.190000 55.225000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 10.620000 55.225000 10.940000 ;
      LAYER met4 ;
        RECT 54.905000 10.620000 55.225000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 11.050000 55.225000 11.370000 ;
      LAYER met4 ;
        RECT 54.905000 11.050000 55.225000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 11.480000 55.225000 11.800000 ;
      LAYER met4 ;
        RECT 54.905000 11.480000 55.225000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 11.910000 55.225000 12.230000 ;
      LAYER met4 ;
        RECT 54.905000 11.910000 55.225000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 12.340000 55.225000 12.660000 ;
      LAYER met4 ;
        RECT 54.905000 12.340000 55.225000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 12.770000 55.225000 13.090000 ;
      LAYER met4 ;
        RECT 54.905000 12.770000 55.225000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 13.200000 55.225000 13.520000 ;
      LAYER met4 ;
        RECT 54.905000 13.200000 55.225000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 8.900000 55.225000 9.220000 ;
      LAYER met4 ;
        RECT 54.905000 8.900000 55.225000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 9.330000 55.225000 9.650000 ;
      LAYER met4 ;
        RECT 54.905000 9.330000 55.225000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 9.760000 55.225000 10.080000 ;
      LAYER met4 ;
        RECT 54.905000 9.760000 55.225000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 10.190000 55.630000 10.510000 ;
      LAYER met4 ;
        RECT 55.310000 10.190000 55.630000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 10.620000 55.630000 10.940000 ;
      LAYER met4 ;
        RECT 55.310000 10.620000 55.630000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 11.050000 55.630000 11.370000 ;
      LAYER met4 ;
        RECT 55.310000 11.050000 55.630000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 11.480000 55.630000 11.800000 ;
      LAYER met4 ;
        RECT 55.310000 11.480000 55.630000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 11.910000 55.630000 12.230000 ;
      LAYER met4 ;
        RECT 55.310000 11.910000 55.630000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 12.340000 55.630000 12.660000 ;
      LAYER met4 ;
        RECT 55.310000 12.340000 55.630000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 12.770000 55.630000 13.090000 ;
      LAYER met4 ;
        RECT 55.310000 12.770000 55.630000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 13.200000 55.630000 13.520000 ;
      LAYER met4 ;
        RECT 55.310000 13.200000 55.630000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 8.900000 55.630000 9.220000 ;
      LAYER met4 ;
        RECT 55.310000 8.900000 55.630000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 9.330000 55.630000 9.650000 ;
      LAYER met4 ;
        RECT 55.310000 9.330000 55.630000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 9.760000 55.630000 10.080000 ;
      LAYER met4 ;
        RECT 55.310000 9.760000 55.630000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 10.190000 56.035000 10.510000 ;
      LAYER met4 ;
        RECT 55.715000 10.190000 56.035000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 10.620000 56.035000 10.940000 ;
      LAYER met4 ;
        RECT 55.715000 10.620000 56.035000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 11.050000 56.035000 11.370000 ;
      LAYER met4 ;
        RECT 55.715000 11.050000 56.035000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 11.480000 56.035000 11.800000 ;
      LAYER met4 ;
        RECT 55.715000 11.480000 56.035000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 11.910000 56.035000 12.230000 ;
      LAYER met4 ;
        RECT 55.715000 11.910000 56.035000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 12.340000 56.035000 12.660000 ;
      LAYER met4 ;
        RECT 55.715000 12.340000 56.035000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 12.770000 56.035000 13.090000 ;
      LAYER met4 ;
        RECT 55.715000 12.770000 56.035000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 13.200000 56.035000 13.520000 ;
      LAYER met4 ;
        RECT 55.715000 13.200000 56.035000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 8.900000 56.035000 9.220000 ;
      LAYER met4 ;
        RECT 55.715000 8.900000 56.035000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 9.330000 56.035000 9.650000 ;
      LAYER met4 ;
        RECT 55.715000 9.330000 56.035000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 9.760000 56.035000 10.080000 ;
      LAYER met4 ;
        RECT 55.715000 9.760000 56.035000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 10.190000 56.440000 10.510000 ;
      LAYER met4 ;
        RECT 56.120000 10.190000 56.440000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 10.620000 56.440000 10.940000 ;
      LAYER met4 ;
        RECT 56.120000 10.620000 56.440000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 11.050000 56.440000 11.370000 ;
      LAYER met4 ;
        RECT 56.120000 11.050000 56.440000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 11.480000 56.440000 11.800000 ;
      LAYER met4 ;
        RECT 56.120000 11.480000 56.440000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 11.910000 56.440000 12.230000 ;
      LAYER met4 ;
        RECT 56.120000 11.910000 56.440000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 12.340000 56.440000 12.660000 ;
      LAYER met4 ;
        RECT 56.120000 12.340000 56.440000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 12.770000 56.440000 13.090000 ;
      LAYER met4 ;
        RECT 56.120000 12.770000 56.440000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 13.200000 56.440000 13.520000 ;
      LAYER met4 ;
        RECT 56.120000 13.200000 56.440000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 8.900000 56.440000 9.220000 ;
      LAYER met4 ;
        RECT 56.120000 8.900000 56.440000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 9.330000 56.440000 9.650000 ;
      LAYER met4 ;
        RECT 56.120000 9.330000 56.440000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 9.760000 56.440000 10.080000 ;
      LAYER met4 ;
        RECT 56.120000 9.760000 56.440000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 10.190000 56.845000 10.510000 ;
      LAYER met4 ;
        RECT 56.525000 10.190000 56.845000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 10.620000 56.845000 10.940000 ;
      LAYER met4 ;
        RECT 56.525000 10.620000 56.845000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 11.050000 56.845000 11.370000 ;
      LAYER met4 ;
        RECT 56.525000 11.050000 56.845000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 11.480000 56.845000 11.800000 ;
      LAYER met4 ;
        RECT 56.525000 11.480000 56.845000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 11.910000 56.845000 12.230000 ;
      LAYER met4 ;
        RECT 56.525000 11.910000 56.845000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 12.340000 56.845000 12.660000 ;
      LAYER met4 ;
        RECT 56.525000 12.340000 56.845000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 12.770000 56.845000 13.090000 ;
      LAYER met4 ;
        RECT 56.525000 12.770000 56.845000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 13.200000 56.845000 13.520000 ;
      LAYER met4 ;
        RECT 56.525000 13.200000 56.845000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 8.900000 56.845000 9.220000 ;
      LAYER met4 ;
        RECT 56.525000 8.900000 56.845000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 9.330000 56.845000 9.650000 ;
      LAYER met4 ;
        RECT 56.525000 9.330000 56.845000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 9.760000 56.845000 10.080000 ;
      LAYER met4 ;
        RECT 56.525000 9.760000 56.845000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 10.190000 57.250000 10.510000 ;
      LAYER met4 ;
        RECT 56.930000 10.190000 57.250000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 10.620000 57.250000 10.940000 ;
      LAYER met4 ;
        RECT 56.930000 10.620000 57.250000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 11.050000 57.250000 11.370000 ;
      LAYER met4 ;
        RECT 56.930000 11.050000 57.250000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 11.480000 57.250000 11.800000 ;
      LAYER met4 ;
        RECT 56.930000 11.480000 57.250000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 11.910000 57.250000 12.230000 ;
      LAYER met4 ;
        RECT 56.930000 11.910000 57.250000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 12.340000 57.250000 12.660000 ;
      LAYER met4 ;
        RECT 56.930000 12.340000 57.250000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 12.770000 57.250000 13.090000 ;
      LAYER met4 ;
        RECT 56.930000 12.770000 57.250000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 13.200000 57.250000 13.520000 ;
      LAYER met4 ;
        RECT 56.930000 13.200000 57.250000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 8.900000 57.250000 9.220000 ;
      LAYER met4 ;
        RECT 56.930000 8.900000 57.250000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 9.330000 57.250000 9.650000 ;
      LAYER met4 ;
        RECT 56.930000 9.330000 57.250000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 9.760000 57.250000 10.080000 ;
      LAYER met4 ;
        RECT 56.930000 9.760000 57.250000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 10.190000 57.655000 10.510000 ;
      LAYER met4 ;
        RECT 57.335000 10.190000 57.655000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 10.620000 57.655000 10.940000 ;
      LAYER met4 ;
        RECT 57.335000 10.620000 57.655000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 11.050000 57.655000 11.370000 ;
      LAYER met4 ;
        RECT 57.335000 11.050000 57.655000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 11.480000 57.655000 11.800000 ;
      LAYER met4 ;
        RECT 57.335000 11.480000 57.655000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 11.910000 57.655000 12.230000 ;
      LAYER met4 ;
        RECT 57.335000 11.910000 57.655000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 12.340000 57.655000 12.660000 ;
      LAYER met4 ;
        RECT 57.335000 12.340000 57.655000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 12.770000 57.655000 13.090000 ;
      LAYER met4 ;
        RECT 57.335000 12.770000 57.655000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 13.200000 57.655000 13.520000 ;
      LAYER met4 ;
        RECT 57.335000 13.200000 57.655000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 8.900000 57.655000 9.220000 ;
      LAYER met4 ;
        RECT 57.335000 8.900000 57.655000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 9.330000 57.655000 9.650000 ;
      LAYER met4 ;
        RECT 57.335000 9.330000 57.655000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 9.760000 57.655000 10.080000 ;
      LAYER met4 ;
        RECT 57.335000 9.760000 57.655000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 10.190000 58.060000 10.510000 ;
      LAYER met4 ;
        RECT 57.740000 10.190000 58.060000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 10.620000 58.060000 10.940000 ;
      LAYER met4 ;
        RECT 57.740000 10.620000 58.060000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 11.050000 58.060000 11.370000 ;
      LAYER met4 ;
        RECT 57.740000 11.050000 58.060000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 11.480000 58.060000 11.800000 ;
      LAYER met4 ;
        RECT 57.740000 11.480000 58.060000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 11.910000 58.060000 12.230000 ;
      LAYER met4 ;
        RECT 57.740000 11.910000 58.060000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 12.340000 58.060000 12.660000 ;
      LAYER met4 ;
        RECT 57.740000 12.340000 58.060000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 12.770000 58.060000 13.090000 ;
      LAYER met4 ;
        RECT 57.740000 12.770000 58.060000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 13.200000 58.060000 13.520000 ;
      LAYER met4 ;
        RECT 57.740000 13.200000 58.060000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 8.900000 58.060000 9.220000 ;
      LAYER met4 ;
        RECT 57.740000 8.900000 58.060000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 9.330000 58.060000 9.650000 ;
      LAYER met4 ;
        RECT 57.740000 9.330000 58.060000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 9.760000 58.060000 10.080000 ;
      LAYER met4 ;
        RECT 57.740000 9.760000 58.060000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 10.190000 58.465000 10.510000 ;
      LAYER met4 ;
        RECT 58.145000 10.190000 58.465000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 10.620000 58.465000 10.940000 ;
      LAYER met4 ;
        RECT 58.145000 10.620000 58.465000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 11.050000 58.465000 11.370000 ;
      LAYER met4 ;
        RECT 58.145000 11.050000 58.465000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 11.480000 58.465000 11.800000 ;
      LAYER met4 ;
        RECT 58.145000 11.480000 58.465000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 11.910000 58.465000 12.230000 ;
      LAYER met4 ;
        RECT 58.145000 11.910000 58.465000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 12.340000 58.465000 12.660000 ;
      LAYER met4 ;
        RECT 58.145000 12.340000 58.465000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 12.770000 58.465000 13.090000 ;
      LAYER met4 ;
        RECT 58.145000 12.770000 58.465000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 13.200000 58.465000 13.520000 ;
      LAYER met4 ;
        RECT 58.145000 13.200000 58.465000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 8.900000 58.465000 9.220000 ;
      LAYER met4 ;
        RECT 58.145000 8.900000 58.465000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 9.330000 58.465000 9.650000 ;
      LAYER met4 ;
        RECT 58.145000 9.330000 58.465000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 9.760000 58.465000 10.080000 ;
      LAYER met4 ;
        RECT 58.145000 9.760000 58.465000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 10.190000 58.870000 10.510000 ;
      LAYER met4 ;
        RECT 58.550000 10.190000 58.870000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 10.620000 58.870000 10.940000 ;
      LAYER met4 ;
        RECT 58.550000 10.620000 58.870000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 11.050000 58.870000 11.370000 ;
      LAYER met4 ;
        RECT 58.550000 11.050000 58.870000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 11.480000 58.870000 11.800000 ;
      LAYER met4 ;
        RECT 58.550000 11.480000 58.870000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 11.910000 58.870000 12.230000 ;
      LAYER met4 ;
        RECT 58.550000 11.910000 58.870000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 12.340000 58.870000 12.660000 ;
      LAYER met4 ;
        RECT 58.550000 12.340000 58.870000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 12.770000 58.870000 13.090000 ;
      LAYER met4 ;
        RECT 58.550000 12.770000 58.870000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 13.200000 58.870000 13.520000 ;
      LAYER met4 ;
        RECT 58.550000 13.200000 58.870000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 8.900000 58.870000 9.220000 ;
      LAYER met4 ;
        RECT 58.550000 8.900000 58.870000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 9.330000 58.870000 9.650000 ;
      LAYER met4 ;
        RECT 58.550000 9.330000 58.870000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 9.760000 58.870000 10.080000 ;
      LAYER met4 ;
        RECT 58.550000 9.760000 58.870000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 10.190000 59.275000 10.510000 ;
      LAYER met4 ;
        RECT 58.955000 10.190000 59.275000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 10.620000 59.275000 10.940000 ;
      LAYER met4 ;
        RECT 58.955000 10.620000 59.275000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 11.050000 59.275000 11.370000 ;
      LAYER met4 ;
        RECT 58.955000 11.050000 59.275000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 11.480000 59.275000 11.800000 ;
      LAYER met4 ;
        RECT 58.955000 11.480000 59.275000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 11.910000 59.275000 12.230000 ;
      LAYER met4 ;
        RECT 58.955000 11.910000 59.275000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 12.340000 59.275000 12.660000 ;
      LAYER met4 ;
        RECT 58.955000 12.340000 59.275000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 12.770000 59.275000 13.090000 ;
      LAYER met4 ;
        RECT 58.955000 12.770000 59.275000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 13.200000 59.275000 13.520000 ;
      LAYER met4 ;
        RECT 58.955000 13.200000 59.275000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 8.900000 59.275000 9.220000 ;
      LAYER met4 ;
        RECT 58.955000 8.900000 59.275000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 9.330000 59.275000 9.650000 ;
      LAYER met4 ;
        RECT 58.955000 9.330000 59.275000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 9.760000 59.275000 10.080000 ;
      LAYER met4 ;
        RECT 58.955000 9.760000 59.275000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 10.190000 59.680000 10.510000 ;
      LAYER met4 ;
        RECT 59.360000 10.190000 59.680000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 10.620000 59.680000 10.940000 ;
      LAYER met4 ;
        RECT 59.360000 10.620000 59.680000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 11.050000 59.680000 11.370000 ;
      LAYER met4 ;
        RECT 59.360000 11.050000 59.680000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 11.480000 59.680000 11.800000 ;
      LAYER met4 ;
        RECT 59.360000 11.480000 59.680000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 11.910000 59.680000 12.230000 ;
      LAYER met4 ;
        RECT 59.360000 11.910000 59.680000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 12.340000 59.680000 12.660000 ;
      LAYER met4 ;
        RECT 59.360000 12.340000 59.680000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 12.770000 59.680000 13.090000 ;
      LAYER met4 ;
        RECT 59.360000 12.770000 59.680000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 13.200000 59.680000 13.520000 ;
      LAYER met4 ;
        RECT 59.360000 13.200000 59.680000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 8.900000 59.680000 9.220000 ;
      LAYER met4 ;
        RECT 59.360000 8.900000 59.680000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 9.330000 59.680000 9.650000 ;
      LAYER met4 ;
        RECT 59.360000 9.330000 59.680000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 9.760000 59.680000 10.080000 ;
      LAYER met4 ;
        RECT 59.360000 9.760000 59.680000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 10.190000 60.085000 10.510000 ;
      LAYER met4 ;
        RECT 59.765000 10.190000 60.085000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 10.620000 60.085000 10.940000 ;
      LAYER met4 ;
        RECT 59.765000 10.620000 60.085000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 11.050000 60.085000 11.370000 ;
      LAYER met4 ;
        RECT 59.765000 11.050000 60.085000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 11.480000 60.085000 11.800000 ;
      LAYER met4 ;
        RECT 59.765000 11.480000 60.085000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 11.910000 60.085000 12.230000 ;
      LAYER met4 ;
        RECT 59.765000 11.910000 60.085000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 12.340000 60.085000 12.660000 ;
      LAYER met4 ;
        RECT 59.765000 12.340000 60.085000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 12.770000 60.085000 13.090000 ;
      LAYER met4 ;
        RECT 59.765000 12.770000 60.085000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 13.200000 60.085000 13.520000 ;
      LAYER met4 ;
        RECT 59.765000 13.200000 60.085000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 8.900000 60.085000 9.220000 ;
      LAYER met4 ;
        RECT 59.765000 8.900000 60.085000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 9.330000 60.085000 9.650000 ;
      LAYER met4 ;
        RECT 59.765000 9.330000 60.085000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 9.760000 60.085000 10.080000 ;
      LAYER met4 ;
        RECT 59.765000 9.760000 60.085000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 10.190000 6.545000 10.510000 ;
      LAYER met4 ;
        RECT 6.225000 10.190000 6.545000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 10.620000 6.545000 10.940000 ;
      LAYER met4 ;
        RECT 6.225000 10.620000 6.545000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 11.050000 6.545000 11.370000 ;
      LAYER met4 ;
        RECT 6.225000 11.050000 6.545000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 11.480000 6.545000 11.800000 ;
      LAYER met4 ;
        RECT 6.225000 11.480000 6.545000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 11.910000 6.545000 12.230000 ;
      LAYER met4 ;
        RECT 6.225000 11.910000 6.545000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 12.340000 6.545000 12.660000 ;
      LAYER met4 ;
        RECT 6.225000 12.340000 6.545000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 12.770000 6.545000 13.090000 ;
      LAYER met4 ;
        RECT 6.225000 12.770000 6.545000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 13.200000 6.545000 13.520000 ;
      LAYER met4 ;
        RECT 6.225000 13.200000 6.545000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 8.900000 6.545000 9.220000 ;
      LAYER met4 ;
        RECT 6.225000 8.900000 6.545000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 9.330000 6.545000 9.650000 ;
      LAYER met4 ;
        RECT 6.225000 9.330000 6.545000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 9.760000 6.545000 10.080000 ;
      LAYER met4 ;
        RECT 6.225000 9.760000 6.545000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 10.190000 6.950000 10.510000 ;
      LAYER met4 ;
        RECT 6.630000 10.190000 6.950000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 10.620000 6.950000 10.940000 ;
      LAYER met4 ;
        RECT 6.630000 10.620000 6.950000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 11.050000 6.950000 11.370000 ;
      LAYER met4 ;
        RECT 6.630000 11.050000 6.950000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 11.480000 6.950000 11.800000 ;
      LAYER met4 ;
        RECT 6.630000 11.480000 6.950000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 11.910000 6.950000 12.230000 ;
      LAYER met4 ;
        RECT 6.630000 11.910000 6.950000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 12.340000 6.950000 12.660000 ;
      LAYER met4 ;
        RECT 6.630000 12.340000 6.950000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 12.770000 6.950000 13.090000 ;
      LAYER met4 ;
        RECT 6.630000 12.770000 6.950000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 13.200000 6.950000 13.520000 ;
      LAYER met4 ;
        RECT 6.630000 13.200000 6.950000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 8.900000 6.950000 9.220000 ;
      LAYER met4 ;
        RECT 6.630000 8.900000 6.950000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 9.330000 6.950000 9.650000 ;
      LAYER met4 ;
        RECT 6.630000 9.330000 6.950000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 9.760000 6.950000 10.080000 ;
      LAYER met4 ;
        RECT 6.630000 9.760000 6.950000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 10.190000 60.490000 10.510000 ;
      LAYER met4 ;
        RECT 60.170000 10.190000 60.490000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 10.620000 60.490000 10.940000 ;
      LAYER met4 ;
        RECT 60.170000 10.620000 60.490000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 11.050000 60.490000 11.370000 ;
      LAYER met4 ;
        RECT 60.170000 11.050000 60.490000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 11.480000 60.490000 11.800000 ;
      LAYER met4 ;
        RECT 60.170000 11.480000 60.490000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 11.910000 60.490000 12.230000 ;
      LAYER met4 ;
        RECT 60.170000 11.910000 60.490000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 12.340000 60.490000 12.660000 ;
      LAYER met4 ;
        RECT 60.170000 12.340000 60.490000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 12.770000 60.490000 13.090000 ;
      LAYER met4 ;
        RECT 60.170000 12.770000 60.490000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 13.200000 60.490000 13.520000 ;
      LAYER met4 ;
        RECT 60.170000 13.200000 60.490000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 8.900000 60.490000 9.220000 ;
      LAYER met4 ;
        RECT 60.170000 8.900000 60.490000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 9.330000 60.490000 9.650000 ;
      LAYER met4 ;
        RECT 60.170000 9.330000 60.490000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 9.760000 60.490000 10.080000 ;
      LAYER met4 ;
        RECT 60.170000 9.760000 60.490000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 10.190000 60.895000 10.510000 ;
      LAYER met4 ;
        RECT 60.575000 10.190000 60.895000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 10.620000 60.895000 10.940000 ;
      LAYER met4 ;
        RECT 60.575000 10.620000 60.895000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 11.050000 60.895000 11.370000 ;
      LAYER met4 ;
        RECT 60.575000 11.050000 60.895000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 11.480000 60.895000 11.800000 ;
      LAYER met4 ;
        RECT 60.575000 11.480000 60.895000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 11.910000 60.895000 12.230000 ;
      LAYER met4 ;
        RECT 60.575000 11.910000 60.895000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 12.340000 60.895000 12.660000 ;
      LAYER met4 ;
        RECT 60.575000 12.340000 60.895000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 12.770000 60.895000 13.090000 ;
      LAYER met4 ;
        RECT 60.575000 12.770000 60.895000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 13.200000 60.895000 13.520000 ;
      LAYER met4 ;
        RECT 60.575000 13.200000 60.895000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 8.900000 60.895000 9.220000 ;
      LAYER met4 ;
        RECT 60.575000 8.900000 60.895000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 9.330000 60.895000 9.650000 ;
      LAYER met4 ;
        RECT 60.575000 9.330000 60.895000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 9.760000 60.895000 10.080000 ;
      LAYER met4 ;
        RECT 60.575000 9.760000 60.895000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 10.190000 61.300000 10.510000 ;
      LAYER met4 ;
        RECT 60.980000 10.190000 61.300000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 10.620000 61.300000 10.940000 ;
      LAYER met4 ;
        RECT 60.980000 10.620000 61.300000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 11.050000 61.300000 11.370000 ;
      LAYER met4 ;
        RECT 60.980000 11.050000 61.300000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 11.480000 61.300000 11.800000 ;
      LAYER met4 ;
        RECT 60.980000 11.480000 61.300000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 11.910000 61.300000 12.230000 ;
      LAYER met4 ;
        RECT 60.980000 11.910000 61.300000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 12.340000 61.300000 12.660000 ;
      LAYER met4 ;
        RECT 60.980000 12.340000 61.300000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 12.770000 61.300000 13.090000 ;
      LAYER met4 ;
        RECT 60.980000 12.770000 61.300000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 13.200000 61.300000 13.520000 ;
      LAYER met4 ;
        RECT 60.980000 13.200000 61.300000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 8.900000 61.300000 9.220000 ;
      LAYER met4 ;
        RECT 60.980000 8.900000 61.300000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 9.330000 61.300000 9.650000 ;
      LAYER met4 ;
        RECT 60.980000 9.330000 61.300000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 9.760000 61.300000 10.080000 ;
      LAYER met4 ;
        RECT 60.980000 9.760000 61.300000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 10.190000 61.705000 10.510000 ;
      LAYER met4 ;
        RECT 61.385000 10.190000 61.705000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 10.620000 61.705000 10.940000 ;
      LAYER met4 ;
        RECT 61.385000 10.620000 61.705000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 11.050000 61.705000 11.370000 ;
      LAYER met4 ;
        RECT 61.385000 11.050000 61.705000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 11.480000 61.705000 11.800000 ;
      LAYER met4 ;
        RECT 61.385000 11.480000 61.705000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 11.910000 61.705000 12.230000 ;
      LAYER met4 ;
        RECT 61.385000 11.910000 61.705000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 12.340000 61.705000 12.660000 ;
      LAYER met4 ;
        RECT 61.385000 12.340000 61.705000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 12.770000 61.705000 13.090000 ;
      LAYER met4 ;
        RECT 61.385000 12.770000 61.705000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 13.200000 61.705000 13.520000 ;
      LAYER met4 ;
        RECT 61.385000 13.200000 61.705000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 8.900000 61.705000 9.220000 ;
      LAYER met4 ;
        RECT 61.385000 8.900000 61.705000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 9.330000 61.705000 9.650000 ;
      LAYER met4 ;
        RECT 61.385000 9.330000 61.705000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 9.760000 61.705000 10.080000 ;
      LAYER met4 ;
        RECT 61.385000 9.760000 61.705000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 10.190000 62.110000 10.510000 ;
      LAYER met4 ;
        RECT 61.790000 10.190000 62.110000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 10.620000 62.110000 10.940000 ;
      LAYER met4 ;
        RECT 61.790000 10.620000 62.110000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 11.050000 62.110000 11.370000 ;
      LAYER met4 ;
        RECT 61.790000 11.050000 62.110000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 11.480000 62.110000 11.800000 ;
      LAYER met4 ;
        RECT 61.790000 11.480000 62.110000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 11.910000 62.110000 12.230000 ;
      LAYER met4 ;
        RECT 61.790000 11.910000 62.110000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 12.340000 62.110000 12.660000 ;
      LAYER met4 ;
        RECT 61.790000 12.340000 62.110000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 12.770000 62.110000 13.090000 ;
      LAYER met4 ;
        RECT 61.790000 12.770000 62.110000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 13.200000 62.110000 13.520000 ;
      LAYER met4 ;
        RECT 61.790000 13.200000 62.110000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 8.900000 62.110000 9.220000 ;
      LAYER met4 ;
        RECT 61.790000 8.900000 62.110000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 9.330000 62.110000 9.650000 ;
      LAYER met4 ;
        RECT 61.790000 9.330000 62.110000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 9.760000 62.110000 10.080000 ;
      LAYER met4 ;
        RECT 61.790000 9.760000 62.110000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 10.190000 62.515000 10.510000 ;
      LAYER met4 ;
        RECT 62.195000 10.190000 62.515000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 10.620000 62.515000 10.940000 ;
      LAYER met4 ;
        RECT 62.195000 10.620000 62.515000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 11.050000 62.515000 11.370000 ;
      LAYER met4 ;
        RECT 62.195000 11.050000 62.515000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 11.480000 62.515000 11.800000 ;
      LAYER met4 ;
        RECT 62.195000 11.480000 62.515000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 11.910000 62.515000 12.230000 ;
      LAYER met4 ;
        RECT 62.195000 11.910000 62.515000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 12.340000 62.515000 12.660000 ;
      LAYER met4 ;
        RECT 62.195000 12.340000 62.515000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 12.770000 62.515000 13.090000 ;
      LAYER met4 ;
        RECT 62.195000 12.770000 62.515000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 13.200000 62.515000 13.520000 ;
      LAYER met4 ;
        RECT 62.195000 13.200000 62.515000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 8.900000 62.515000 9.220000 ;
      LAYER met4 ;
        RECT 62.195000 8.900000 62.515000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 9.330000 62.515000 9.650000 ;
      LAYER met4 ;
        RECT 62.195000 9.330000 62.515000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 9.760000 62.515000 10.080000 ;
      LAYER met4 ;
        RECT 62.195000 9.760000 62.515000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 10.190000 62.920000 10.510000 ;
      LAYER met4 ;
        RECT 62.600000 10.190000 62.920000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 10.620000 62.920000 10.940000 ;
      LAYER met4 ;
        RECT 62.600000 10.620000 62.920000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 11.050000 62.920000 11.370000 ;
      LAYER met4 ;
        RECT 62.600000 11.050000 62.920000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 11.480000 62.920000 11.800000 ;
      LAYER met4 ;
        RECT 62.600000 11.480000 62.920000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 11.910000 62.920000 12.230000 ;
      LAYER met4 ;
        RECT 62.600000 11.910000 62.920000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 12.340000 62.920000 12.660000 ;
      LAYER met4 ;
        RECT 62.600000 12.340000 62.920000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 12.770000 62.920000 13.090000 ;
      LAYER met4 ;
        RECT 62.600000 12.770000 62.920000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 13.200000 62.920000 13.520000 ;
      LAYER met4 ;
        RECT 62.600000 13.200000 62.920000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 8.900000 62.920000 9.220000 ;
      LAYER met4 ;
        RECT 62.600000 8.900000 62.920000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 9.330000 62.920000 9.650000 ;
      LAYER met4 ;
        RECT 62.600000 9.330000 62.920000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 9.760000 62.920000 10.080000 ;
      LAYER met4 ;
        RECT 62.600000 9.760000 62.920000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 10.190000 63.325000 10.510000 ;
      LAYER met4 ;
        RECT 63.005000 10.190000 63.325000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 10.620000 63.325000 10.940000 ;
      LAYER met4 ;
        RECT 63.005000 10.620000 63.325000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 11.050000 63.325000 11.370000 ;
      LAYER met4 ;
        RECT 63.005000 11.050000 63.325000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 11.480000 63.325000 11.800000 ;
      LAYER met4 ;
        RECT 63.005000 11.480000 63.325000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 11.910000 63.325000 12.230000 ;
      LAYER met4 ;
        RECT 63.005000 11.910000 63.325000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 12.340000 63.325000 12.660000 ;
      LAYER met4 ;
        RECT 63.005000 12.340000 63.325000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 12.770000 63.325000 13.090000 ;
      LAYER met4 ;
        RECT 63.005000 12.770000 63.325000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 13.200000 63.325000 13.520000 ;
      LAYER met4 ;
        RECT 63.005000 13.200000 63.325000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 8.900000 63.325000 9.220000 ;
      LAYER met4 ;
        RECT 63.005000 8.900000 63.325000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 9.330000 63.325000 9.650000 ;
      LAYER met4 ;
        RECT 63.005000 9.330000 63.325000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 9.760000 63.325000 10.080000 ;
      LAYER met4 ;
        RECT 63.005000 9.760000 63.325000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 10.190000 63.730000 10.510000 ;
      LAYER met4 ;
        RECT 63.410000 10.190000 63.730000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 10.620000 63.730000 10.940000 ;
      LAYER met4 ;
        RECT 63.410000 10.620000 63.730000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 11.050000 63.730000 11.370000 ;
      LAYER met4 ;
        RECT 63.410000 11.050000 63.730000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 11.480000 63.730000 11.800000 ;
      LAYER met4 ;
        RECT 63.410000 11.480000 63.730000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 11.910000 63.730000 12.230000 ;
      LAYER met4 ;
        RECT 63.410000 11.910000 63.730000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 12.340000 63.730000 12.660000 ;
      LAYER met4 ;
        RECT 63.410000 12.340000 63.730000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 12.770000 63.730000 13.090000 ;
      LAYER met4 ;
        RECT 63.410000 12.770000 63.730000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 13.200000 63.730000 13.520000 ;
      LAYER met4 ;
        RECT 63.410000 13.200000 63.730000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 8.900000 63.730000 9.220000 ;
      LAYER met4 ;
        RECT 63.410000 8.900000 63.730000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 9.330000 63.730000 9.650000 ;
      LAYER met4 ;
        RECT 63.410000 9.330000 63.730000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 9.760000 63.730000 10.080000 ;
      LAYER met4 ;
        RECT 63.410000 9.760000 63.730000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 10.190000 64.135000 10.510000 ;
      LAYER met4 ;
        RECT 63.815000 10.190000 64.135000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 10.620000 64.135000 10.940000 ;
      LAYER met4 ;
        RECT 63.815000 10.620000 64.135000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 11.050000 64.135000 11.370000 ;
      LAYER met4 ;
        RECT 63.815000 11.050000 64.135000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 11.480000 64.135000 11.800000 ;
      LAYER met4 ;
        RECT 63.815000 11.480000 64.135000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 11.910000 64.135000 12.230000 ;
      LAYER met4 ;
        RECT 63.815000 11.910000 64.135000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 12.340000 64.135000 12.660000 ;
      LAYER met4 ;
        RECT 63.815000 12.340000 64.135000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 12.770000 64.135000 13.090000 ;
      LAYER met4 ;
        RECT 63.815000 12.770000 64.135000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 13.200000 64.135000 13.520000 ;
      LAYER met4 ;
        RECT 63.815000 13.200000 64.135000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 8.900000 64.135000 9.220000 ;
      LAYER met4 ;
        RECT 63.815000 8.900000 64.135000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 9.330000 64.135000 9.650000 ;
      LAYER met4 ;
        RECT 63.815000 9.330000 64.135000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 9.760000 64.135000 10.080000 ;
      LAYER met4 ;
        RECT 63.815000 9.760000 64.135000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 10.190000 64.540000 10.510000 ;
      LAYER met4 ;
        RECT 64.220000 10.190000 64.540000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 10.620000 64.540000 10.940000 ;
      LAYER met4 ;
        RECT 64.220000 10.620000 64.540000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 11.050000 64.540000 11.370000 ;
      LAYER met4 ;
        RECT 64.220000 11.050000 64.540000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 11.480000 64.540000 11.800000 ;
      LAYER met4 ;
        RECT 64.220000 11.480000 64.540000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 11.910000 64.540000 12.230000 ;
      LAYER met4 ;
        RECT 64.220000 11.910000 64.540000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 12.340000 64.540000 12.660000 ;
      LAYER met4 ;
        RECT 64.220000 12.340000 64.540000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 12.770000 64.540000 13.090000 ;
      LAYER met4 ;
        RECT 64.220000 12.770000 64.540000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 13.200000 64.540000 13.520000 ;
      LAYER met4 ;
        RECT 64.220000 13.200000 64.540000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 8.900000 64.540000 9.220000 ;
      LAYER met4 ;
        RECT 64.220000 8.900000 64.540000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 9.330000 64.540000 9.650000 ;
      LAYER met4 ;
        RECT 64.220000 9.330000 64.540000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 9.760000 64.540000 10.080000 ;
      LAYER met4 ;
        RECT 64.220000 9.760000 64.540000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 10.190000 64.945000 10.510000 ;
      LAYER met4 ;
        RECT 64.625000 10.190000 64.945000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 10.620000 64.945000 10.940000 ;
      LAYER met4 ;
        RECT 64.625000 10.620000 64.945000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 11.050000 64.945000 11.370000 ;
      LAYER met4 ;
        RECT 64.625000 11.050000 64.945000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 11.480000 64.945000 11.800000 ;
      LAYER met4 ;
        RECT 64.625000 11.480000 64.945000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 11.910000 64.945000 12.230000 ;
      LAYER met4 ;
        RECT 64.625000 11.910000 64.945000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 12.340000 64.945000 12.660000 ;
      LAYER met4 ;
        RECT 64.625000 12.340000 64.945000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 12.770000 64.945000 13.090000 ;
      LAYER met4 ;
        RECT 64.625000 12.770000 64.945000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 13.200000 64.945000 13.520000 ;
      LAYER met4 ;
        RECT 64.625000 13.200000 64.945000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 8.900000 64.945000 9.220000 ;
      LAYER met4 ;
        RECT 64.625000 8.900000 64.945000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 9.330000 64.945000 9.650000 ;
      LAYER met4 ;
        RECT 64.625000 9.330000 64.945000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 9.760000 64.945000 10.080000 ;
      LAYER met4 ;
        RECT 64.625000 9.760000 64.945000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 10.190000 65.350000 10.510000 ;
      LAYER met4 ;
        RECT 65.030000 10.190000 65.350000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 10.620000 65.350000 10.940000 ;
      LAYER met4 ;
        RECT 65.030000 10.620000 65.350000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 11.050000 65.350000 11.370000 ;
      LAYER met4 ;
        RECT 65.030000 11.050000 65.350000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 11.480000 65.350000 11.800000 ;
      LAYER met4 ;
        RECT 65.030000 11.480000 65.350000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 11.910000 65.350000 12.230000 ;
      LAYER met4 ;
        RECT 65.030000 11.910000 65.350000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 12.340000 65.350000 12.660000 ;
      LAYER met4 ;
        RECT 65.030000 12.340000 65.350000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 12.770000 65.350000 13.090000 ;
      LAYER met4 ;
        RECT 65.030000 12.770000 65.350000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 13.200000 65.350000 13.520000 ;
      LAYER met4 ;
        RECT 65.030000 13.200000 65.350000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 8.900000 65.350000 9.220000 ;
      LAYER met4 ;
        RECT 65.030000 8.900000 65.350000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 9.330000 65.350000 9.650000 ;
      LAYER met4 ;
        RECT 65.030000 9.330000 65.350000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 9.760000 65.350000 10.080000 ;
      LAYER met4 ;
        RECT 65.030000 9.760000 65.350000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 10.190000 65.755000 10.510000 ;
      LAYER met4 ;
        RECT 65.435000 10.190000 65.755000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 10.620000 65.755000 10.940000 ;
      LAYER met4 ;
        RECT 65.435000 10.620000 65.755000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 11.050000 65.755000 11.370000 ;
      LAYER met4 ;
        RECT 65.435000 11.050000 65.755000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 11.480000 65.755000 11.800000 ;
      LAYER met4 ;
        RECT 65.435000 11.480000 65.755000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 11.910000 65.755000 12.230000 ;
      LAYER met4 ;
        RECT 65.435000 11.910000 65.755000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 12.340000 65.755000 12.660000 ;
      LAYER met4 ;
        RECT 65.435000 12.340000 65.755000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 12.770000 65.755000 13.090000 ;
      LAYER met4 ;
        RECT 65.435000 12.770000 65.755000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 13.200000 65.755000 13.520000 ;
      LAYER met4 ;
        RECT 65.435000 13.200000 65.755000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 8.900000 65.755000 9.220000 ;
      LAYER met4 ;
        RECT 65.435000 8.900000 65.755000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 9.330000 65.755000 9.650000 ;
      LAYER met4 ;
        RECT 65.435000 9.330000 65.755000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 9.760000 65.755000 10.080000 ;
      LAYER met4 ;
        RECT 65.435000 9.760000 65.755000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 10.190000 66.160000 10.510000 ;
      LAYER met4 ;
        RECT 65.840000 10.190000 66.160000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 10.620000 66.160000 10.940000 ;
      LAYER met4 ;
        RECT 65.840000 10.620000 66.160000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 11.050000 66.160000 11.370000 ;
      LAYER met4 ;
        RECT 65.840000 11.050000 66.160000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 11.480000 66.160000 11.800000 ;
      LAYER met4 ;
        RECT 65.840000 11.480000 66.160000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 11.910000 66.160000 12.230000 ;
      LAYER met4 ;
        RECT 65.840000 11.910000 66.160000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 12.340000 66.160000 12.660000 ;
      LAYER met4 ;
        RECT 65.840000 12.340000 66.160000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 12.770000 66.160000 13.090000 ;
      LAYER met4 ;
        RECT 65.840000 12.770000 66.160000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 13.200000 66.160000 13.520000 ;
      LAYER met4 ;
        RECT 65.840000 13.200000 66.160000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 8.900000 66.160000 9.220000 ;
      LAYER met4 ;
        RECT 65.840000 8.900000 66.160000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 9.330000 66.160000 9.650000 ;
      LAYER met4 ;
        RECT 65.840000 9.330000 66.160000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 9.760000 66.160000 10.080000 ;
      LAYER met4 ;
        RECT 65.840000 9.760000 66.160000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 10.190000 66.565000 10.510000 ;
      LAYER met4 ;
        RECT 66.245000 10.190000 66.565000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 10.620000 66.565000 10.940000 ;
      LAYER met4 ;
        RECT 66.245000 10.620000 66.565000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 11.050000 66.565000 11.370000 ;
      LAYER met4 ;
        RECT 66.245000 11.050000 66.565000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 11.480000 66.565000 11.800000 ;
      LAYER met4 ;
        RECT 66.245000 11.480000 66.565000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 11.910000 66.565000 12.230000 ;
      LAYER met4 ;
        RECT 66.245000 11.910000 66.565000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 12.340000 66.565000 12.660000 ;
      LAYER met4 ;
        RECT 66.245000 12.340000 66.565000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 12.770000 66.565000 13.090000 ;
      LAYER met4 ;
        RECT 66.245000 12.770000 66.565000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 13.200000 66.565000 13.520000 ;
      LAYER met4 ;
        RECT 66.245000 13.200000 66.565000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 8.900000 66.565000 9.220000 ;
      LAYER met4 ;
        RECT 66.245000 8.900000 66.565000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 9.330000 66.565000 9.650000 ;
      LAYER met4 ;
        RECT 66.245000 9.330000 66.565000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 9.760000 66.565000 10.080000 ;
      LAYER met4 ;
        RECT 66.245000 9.760000 66.565000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 10.190000 66.970000 10.510000 ;
      LAYER met4 ;
        RECT 66.650000 10.190000 66.970000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 10.620000 66.970000 10.940000 ;
      LAYER met4 ;
        RECT 66.650000 10.620000 66.970000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 11.050000 66.970000 11.370000 ;
      LAYER met4 ;
        RECT 66.650000 11.050000 66.970000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 11.480000 66.970000 11.800000 ;
      LAYER met4 ;
        RECT 66.650000 11.480000 66.970000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 11.910000 66.970000 12.230000 ;
      LAYER met4 ;
        RECT 66.650000 11.910000 66.970000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 12.340000 66.970000 12.660000 ;
      LAYER met4 ;
        RECT 66.650000 12.340000 66.970000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 12.770000 66.970000 13.090000 ;
      LAYER met4 ;
        RECT 66.650000 12.770000 66.970000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 13.200000 66.970000 13.520000 ;
      LAYER met4 ;
        RECT 66.650000 13.200000 66.970000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 8.900000 66.970000 9.220000 ;
      LAYER met4 ;
        RECT 66.650000 8.900000 66.970000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 9.330000 66.970000 9.650000 ;
      LAYER met4 ;
        RECT 66.650000 9.330000 66.970000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 9.760000 66.970000 10.080000 ;
      LAYER met4 ;
        RECT 66.650000 9.760000 66.970000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 10.190000 67.375000 10.510000 ;
      LAYER met4 ;
        RECT 67.055000 10.190000 67.375000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 10.620000 67.375000 10.940000 ;
      LAYER met4 ;
        RECT 67.055000 10.620000 67.375000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 11.050000 67.375000 11.370000 ;
      LAYER met4 ;
        RECT 67.055000 11.050000 67.375000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 11.480000 67.375000 11.800000 ;
      LAYER met4 ;
        RECT 67.055000 11.480000 67.375000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 11.910000 67.375000 12.230000 ;
      LAYER met4 ;
        RECT 67.055000 11.910000 67.375000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 12.340000 67.375000 12.660000 ;
      LAYER met4 ;
        RECT 67.055000 12.340000 67.375000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 12.770000 67.375000 13.090000 ;
      LAYER met4 ;
        RECT 67.055000 12.770000 67.375000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 13.200000 67.375000 13.520000 ;
      LAYER met4 ;
        RECT 67.055000 13.200000 67.375000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 8.900000 67.375000 9.220000 ;
      LAYER met4 ;
        RECT 67.055000 8.900000 67.375000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 9.330000 67.375000 9.650000 ;
      LAYER met4 ;
        RECT 67.055000 9.330000 67.375000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 9.760000 67.375000 10.080000 ;
      LAYER met4 ;
        RECT 67.055000 9.760000 67.375000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 10.190000 67.780000 10.510000 ;
      LAYER met4 ;
        RECT 67.460000 10.190000 67.780000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 10.620000 67.780000 10.940000 ;
      LAYER met4 ;
        RECT 67.460000 10.620000 67.780000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 11.050000 67.780000 11.370000 ;
      LAYER met4 ;
        RECT 67.460000 11.050000 67.780000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 11.480000 67.780000 11.800000 ;
      LAYER met4 ;
        RECT 67.460000 11.480000 67.780000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 11.910000 67.780000 12.230000 ;
      LAYER met4 ;
        RECT 67.460000 11.910000 67.780000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 12.340000 67.780000 12.660000 ;
      LAYER met4 ;
        RECT 67.460000 12.340000 67.780000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 12.770000 67.780000 13.090000 ;
      LAYER met4 ;
        RECT 67.460000 12.770000 67.780000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 13.200000 67.780000 13.520000 ;
      LAYER met4 ;
        RECT 67.460000 13.200000 67.780000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 8.900000 67.780000 9.220000 ;
      LAYER met4 ;
        RECT 67.460000 8.900000 67.780000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 9.330000 67.780000 9.650000 ;
      LAYER met4 ;
        RECT 67.460000 9.330000 67.780000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 9.760000 67.780000 10.080000 ;
      LAYER met4 ;
        RECT 67.460000 9.760000 67.780000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 10.190000 68.185000 10.510000 ;
      LAYER met4 ;
        RECT 67.865000 10.190000 68.185000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 10.620000 68.185000 10.940000 ;
      LAYER met4 ;
        RECT 67.865000 10.620000 68.185000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 11.050000 68.185000 11.370000 ;
      LAYER met4 ;
        RECT 67.865000 11.050000 68.185000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 11.480000 68.185000 11.800000 ;
      LAYER met4 ;
        RECT 67.865000 11.480000 68.185000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 11.910000 68.185000 12.230000 ;
      LAYER met4 ;
        RECT 67.865000 11.910000 68.185000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 12.340000 68.185000 12.660000 ;
      LAYER met4 ;
        RECT 67.865000 12.340000 68.185000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 12.770000 68.185000 13.090000 ;
      LAYER met4 ;
        RECT 67.865000 12.770000 68.185000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 13.200000 68.185000 13.520000 ;
      LAYER met4 ;
        RECT 67.865000 13.200000 68.185000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 8.900000 68.185000 9.220000 ;
      LAYER met4 ;
        RECT 67.865000 8.900000 68.185000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 9.330000 68.185000 9.650000 ;
      LAYER met4 ;
        RECT 67.865000 9.330000 68.185000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 9.760000 68.185000 10.080000 ;
      LAYER met4 ;
        RECT 67.865000 9.760000 68.185000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 10.190000 68.590000 10.510000 ;
      LAYER met4 ;
        RECT 68.270000 10.190000 68.590000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 10.620000 68.590000 10.940000 ;
      LAYER met4 ;
        RECT 68.270000 10.620000 68.590000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 11.050000 68.590000 11.370000 ;
      LAYER met4 ;
        RECT 68.270000 11.050000 68.590000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 11.480000 68.590000 11.800000 ;
      LAYER met4 ;
        RECT 68.270000 11.480000 68.590000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 11.910000 68.590000 12.230000 ;
      LAYER met4 ;
        RECT 68.270000 11.910000 68.590000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 12.340000 68.590000 12.660000 ;
      LAYER met4 ;
        RECT 68.270000 12.340000 68.590000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 12.770000 68.590000 13.090000 ;
      LAYER met4 ;
        RECT 68.270000 12.770000 68.590000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 13.200000 68.590000 13.520000 ;
      LAYER met4 ;
        RECT 68.270000 13.200000 68.590000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 8.900000 68.590000 9.220000 ;
      LAYER met4 ;
        RECT 68.270000 8.900000 68.590000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 9.330000 68.590000 9.650000 ;
      LAYER met4 ;
        RECT 68.270000 9.330000 68.590000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 9.760000 68.590000 10.080000 ;
      LAYER met4 ;
        RECT 68.270000 9.760000 68.590000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 10.190000 68.995000 10.510000 ;
      LAYER met4 ;
        RECT 68.675000 10.190000 68.995000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 10.620000 68.995000 10.940000 ;
      LAYER met4 ;
        RECT 68.675000 10.620000 68.995000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 11.050000 68.995000 11.370000 ;
      LAYER met4 ;
        RECT 68.675000 11.050000 68.995000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 11.480000 68.995000 11.800000 ;
      LAYER met4 ;
        RECT 68.675000 11.480000 68.995000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 11.910000 68.995000 12.230000 ;
      LAYER met4 ;
        RECT 68.675000 11.910000 68.995000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 12.340000 68.995000 12.660000 ;
      LAYER met4 ;
        RECT 68.675000 12.340000 68.995000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 12.770000 68.995000 13.090000 ;
      LAYER met4 ;
        RECT 68.675000 12.770000 68.995000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 13.200000 68.995000 13.520000 ;
      LAYER met4 ;
        RECT 68.675000 13.200000 68.995000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 8.900000 68.995000 9.220000 ;
      LAYER met4 ;
        RECT 68.675000 8.900000 68.995000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 9.330000 68.995000 9.650000 ;
      LAYER met4 ;
        RECT 68.675000 9.330000 68.995000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 9.760000 68.995000 10.080000 ;
      LAYER met4 ;
        RECT 68.675000 9.760000 68.995000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 10.190000 69.400000 10.510000 ;
      LAYER met4 ;
        RECT 69.080000 10.190000 69.400000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 10.620000 69.400000 10.940000 ;
      LAYER met4 ;
        RECT 69.080000 10.620000 69.400000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 11.050000 69.400000 11.370000 ;
      LAYER met4 ;
        RECT 69.080000 11.050000 69.400000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 11.480000 69.400000 11.800000 ;
      LAYER met4 ;
        RECT 69.080000 11.480000 69.400000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 11.910000 69.400000 12.230000 ;
      LAYER met4 ;
        RECT 69.080000 11.910000 69.400000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 12.340000 69.400000 12.660000 ;
      LAYER met4 ;
        RECT 69.080000 12.340000 69.400000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 12.770000 69.400000 13.090000 ;
      LAYER met4 ;
        RECT 69.080000 12.770000 69.400000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 13.200000 69.400000 13.520000 ;
      LAYER met4 ;
        RECT 69.080000 13.200000 69.400000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 8.900000 69.400000 9.220000 ;
      LAYER met4 ;
        RECT 69.080000 8.900000 69.400000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 9.330000 69.400000 9.650000 ;
      LAYER met4 ;
        RECT 69.080000 9.330000 69.400000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 9.760000 69.400000 10.080000 ;
      LAYER met4 ;
        RECT 69.080000 9.760000 69.400000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 10.190000 69.805000 10.510000 ;
      LAYER met4 ;
        RECT 69.485000 10.190000 69.805000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 10.620000 69.805000 10.940000 ;
      LAYER met4 ;
        RECT 69.485000 10.620000 69.805000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 11.050000 69.805000 11.370000 ;
      LAYER met4 ;
        RECT 69.485000 11.050000 69.805000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 11.480000 69.805000 11.800000 ;
      LAYER met4 ;
        RECT 69.485000 11.480000 69.805000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 11.910000 69.805000 12.230000 ;
      LAYER met4 ;
        RECT 69.485000 11.910000 69.805000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 12.340000 69.805000 12.660000 ;
      LAYER met4 ;
        RECT 69.485000 12.340000 69.805000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 12.770000 69.805000 13.090000 ;
      LAYER met4 ;
        RECT 69.485000 12.770000 69.805000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 13.200000 69.805000 13.520000 ;
      LAYER met4 ;
        RECT 69.485000 13.200000 69.805000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 8.900000 69.805000 9.220000 ;
      LAYER met4 ;
        RECT 69.485000 8.900000 69.805000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 9.330000 69.805000 9.650000 ;
      LAYER met4 ;
        RECT 69.485000 9.330000 69.805000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 9.760000 69.805000 10.080000 ;
      LAYER met4 ;
        RECT 69.485000 9.760000 69.805000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 10.190000 70.210000 10.510000 ;
      LAYER met4 ;
        RECT 69.890000 10.190000 70.210000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 10.620000 70.210000 10.940000 ;
      LAYER met4 ;
        RECT 69.890000 10.620000 70.210000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 11.050000 70.210000 11.370000 ;
      LAYER met4 ;
        RECT 69.890000 11.050000 70.210000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 11.480000 70.210000 11.800000 ;
      LAYER met4 ;
        RECT 69.890000 11.480000 70.210000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 11.910000 70.210000 12.230000 ;
      LAYER met4 ;
        RECT 69.890000 11.910000 70.210000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 12.340000 70.210000 12.660000 ;
      LAYER met4 ;
        RECT 69.890000 12.340000 70.210000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 12.770000 70.210000 13.090000 ;
      LAYER met4 ;
        RECT 69.890000 12.770000 70.210000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 13.200000 70.210000 13.520000 ;
      LAYER met4 ;
        RECT 69.890000 13.200000 70.210000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 8.900000 70.210000 9.220000 ;
      LAYER met4 ;
        RECT 69.890000 8.900000 70.210000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 9.330000 70.210000 9.650000 ;
      LAYER met4 ;
        RECT 69.890000 9.330000 70.210000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 9.760000 70.210000 10.080000 ;
      LAYER met4 ;
        RECT 69.890000 9.760000 70.210000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 10.190000 7.355000 10.510000 ;
      LAYER met4 ;
        RECT 7.035000 10.190000 7.355000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 10.620000 7.355000 10.940000 ;
      LAYER met4 ;
        RECT 7.035000 10.620000 7.355000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 11.050000 7.355000 11.370000 ;
      LAYER met4 ;
        RECT 7.035000 11.050000 7.355000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 11.480000 7.355000 11.800000 ;
      LAYER met4 ;
        RECT 7.035000 11.480000 7.355000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 11.910000 7.355000 12.230000 ;
      LAYER met4 ;
        RECT 7.035000 11.910000 7.355000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 12.340000 7.355000 12.660000 ;
      LAYER met4 ;
        RECT 7.035000 12.340000 7.355000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 12.770000 7.355000 13.090000 ;
      LAYER met4 ;
        RECT 7.035000 12.770000 7.355000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 13.200000 7.355000 13.520000 ;
      LAYER met4 ;
        RECT 7.035000 13.200000 7.355000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 8.900000 7.355000 9.220000 ;
      LAYER met4 ;
        RECT 7.035000 8.900000 7.355000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 9.330000 7.355000 9.650000 ;
      LAYER met4 ;
        RECT 7.035000 9.330000 7.355000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 9.760000 7.355000 10.080000 ;
      LAYER met4 ;
        RECT 7.035000 9.760000 7.355000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 10.190000 7.760000 10.510000 ;
      LAYER met4 ;
        RECT 7.440000 10.190000 7.760000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 10.620000 7.760000 10.940000 ;
      LAYER met4 ;
        RECT 7.440000 10.620000 7.760000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 11.050000 7.760000 11.370000 ;
      LAYER met4 ;
        RECT 7.440000 11.050000 7.760000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 11.480000 7.760000 11.800000 ;
      LAYER met4 ;
        RECT 7.440000 11.480000 7.760000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 11.910000 7.760000 12.230000 ;
      LAYER met4 ;
        RECT 7.440000 11.910000 7.760000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 12.340000 7.760000 12.660000 ;
      LAYER met4 ;
        RECT 7.440000 12.340000 7.760000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 12.770000 7.760000 13.090000 ;
      LAYER met4 ;
        RECT 7.440000 12.770000 7.760000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 13.200000 7.760000 13.520000 ;
      LAYER met4 ;
        RECT 7.440000 13.200000 7.760000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 8.900000 7.760000 9.220000 ;
      LAYER met4 ;
        RECT 7.440000 8.900000 7.760000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 9.330000 7.760000 9.650000 ;
      LAYER met4 ;
        RECT 7.440000 9.330000 7.760000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 9.760000 7.760000 10.080000 ;
      LAYER met4 ;
        RECT 7.440000 9.760000 7.760000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 10.190000 8.165000 10.510000 ;
      LAYER met4 ;
        RECT 7.845000 10.190000 8.165000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 10.620000 8.165000 10.940000 ;
      LAYER met4 ;
        RECT 7.845000 10.620000 8.165000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 11.050000 8.165000 11.370000 ;
      LAYER met4 ;
        RECT 7.845000 11.050000 8.165000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 11.480000 8.165000 11.800000 ;
      LAYER met4 ;
        RECT 7.845000 11.480000 8.165000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 11.910000 8.165000 12.230000 ;
      LAYER met4 ;
        RECT 7.845000 11.910000 8.165000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 12.340000 8.165000 12.660000 ;
      LAYER met4 ;
        RECT 7.845000 12.340000 8.165000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 12.770000 8.165000 13.090000 ;
      LAYER met4 ;
        RECT 7.845000 12.770000 8.165000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 13.200000 8.165000 13.520000 ;
      LAYER met4 ;
        RECT 7.845000 13.200000 8.165000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 8.900000 8.165000 9.220000 ;
      LAYER met4 ;
        RECT 7.845000 8.900000 8.165000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 9.330000 8.165000 9.650000 ;
      LAYER met4 ;
        RECT 7.845000 9.330000 8.165000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 9.760000 8.165000 10.080000 ;
      LAYER met4 ;
        RECT 7.845000 9.760000 8.165000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 10.190000 70.615000 10.510000 ;
      LAYER met4 ;
        RECT 70.295000 10.190000 70.615000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 10.620000 70.615000 10.940000 ;
      LAYER met4 ;
        RECT 70.295000 10.620000 70.615000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 11.050000 70.615000 11.370000 ;
      LAYER met4 ;
        RECT 70.295000 11.050000 70.615000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 11.480000 70.615000 11.800000 ;
      LAYER met4 ;
        RECT 70.295000 11.480000 70.615000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 11.910000 70.615000 12.230000 ;
      LAYER met4 ;
        RECT 70.295000 11.910000 70.615000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 12.340000 70.615000 12.660000 ;
      LAYER met4 ;
        RECT 70.295000 12.340000 70.615000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 12.770000 70.615000 13.090000 ;
      LAYER met4 ;
        RECT 70.295000 12.770000 70.615000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 13.200000 70.615000 13.520000 ;
      LAYER met4 ;
        RECT 70.295000 13.200000 70.615000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 8.900000 70.615000 9.220000 ;
      LAYER met4 ;
        RECT 70.295000 8.900000 70.615000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 9.330000 70.615000 9.650000 ;
      LAYER met4 ;
        RECT 70.295000 9.330000 70.615000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 9.760000 70.615000 10.080000 ;
      LAYER met4 ;
        RECT 70.295000 9.760000 70.615000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 10.190000 71.020000 10.510000 ;
      LAYER met4 ;
        RECT 70.700000 10.190000 71.020000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 10.620000 71.020000 10.940000 ;
      LAYER met4 ;
        RECT 70.700000 10.620000 71.020000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 11.050000 71.020000 11.370000 ;
      LAYER met4 ;
        RECT 70.700000 11.050000 71.020000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 11.480000 71.020000 11.800000 ;
      LAYER met4 ;
        RECT 70.700000 11.480000 71.020000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 11.910000 71.020000 12.230000 ;
      LAYER met4 ;
        RECT 70.700000 11.910000 71.020000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 12.340000 71.020000 12.660000 ;
      LAYER met4 ;
        RECT 70.700000 12.340000 71.020000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 12.770000 71.020000 13.090000 ;
      LAYER met4 ;
        RECT 70.700000 12.770000 71.020000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 13.200000 71.020000 13.520000 ;
      LAYER met4 ;
        RECT 70.700000 13.200000 71.020000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 8.900000 71.020000 9.220000 ;
      LAYER met4 ;
        RECT 70.700000 8.900000 71.020000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 9.330000 71.020000 9.650000 ;
      LAYER met4 ;
        RECT 70.700000 9.330000 71.020000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 9.760000 71.020000 10.080000 ;
      LAYER met4 ;
        RECT 70.700000 9.760000 71.020000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 10.190000 71.425000 10.510000 ;
      LAYER met4 ;
        RECT 71.105000 10.190000 71.425000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 10.620000 71.425000 10.940000 ;
      LAYER met4 ;
        RECT 71.105000 10.620000 71.425000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 11.050000 71.425000 11.370000 ;
      LAYER met4 ;
        RECT 71.105000 11.050000 71.425000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 11.480000 71.425000 11.800000 ;
      LAYER met4 ;
        RECT 71.105000 11.480000 71.425000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 11.910000 71.425000 12.230000 ;
      LAYER met4 ;
        RECT 71.105000 11.910000 71.425000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 12.340000 71.425000 12.660000 ;
      LAYER met4 ;
        RECT 71.105000 12.340000 71.425000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 12.770000 71.425000 13.090000 ;
      LAYER met4 ;
        RECT 71.105000 12.770000 71.425000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 13.200000 71.425000 13.520000 ;
      LAYER met4 ;
        RECT 71.105000 13.200000 71.425000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 8.900000 71.425000 9.220000 ;
      LAYER met4 ;
        RECT 71.105000 8.900000 71.425000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 9.330000 71.425000 9.650000 ;
      LAYER met4 ;
        RECT 71.105000 9.330000 71.425000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 9.760000 71.425000 10.080000 ;
      LAYER met4 ;
        RECT 71.105000 9.760000 71.425000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 10.190000 71.830000 10.510000 ;
      LAYER met4 ;
        RECT 71.510000 10.190000 71.830000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 10.620000 71.830000 10.940000 ;
      LAYER met4 ;
        RECT 71.510000 10.620000 71.830000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 11.050000 71.830000 11.370000 ;
      LAYER met4 ;
        RECT 71.510000 11.050000 71.830000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 11.480000 71.830000 11.800000 ;
      LAYER met4 ;
        RECT 71.510000 11.480000 71.830000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 11.910000 71.830000 12.230000 ;
      LAYER met4 ;
        RECT 71.510000 11.910000 71.830000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 12.340000 71.830000 12.660000 ;
      LAYER met4 ;
        RECT 71.510000 12.340000 71.830000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 12.770000 71.830000 13.090000 ;
      LAYER met4 ;
        RECT 71.510000 12.770000 71.830000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 13.200000 71.830000 13.520000 ;
      LAYER met4 ;
        RECT 71.510000 13.200000 71.830000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 8.900000 71.830000 9.220000 ;
      LAYER met4 ;
        RECT 71.510000 8.900000 71.830000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 9.330000 71.830000 9.650000 ;
      LAYER met4 ;
        RECT 71.510000 9.330000 71.830000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 9.760000 71.830000 10.080000 ;
      LAYER met4 ;
        RECT 71.510000 9.760000 71.830000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 10.190000 72.235000 10.510000 ;
      LAYER met4 ;
        RECT 71.915000 10.190000 72.235000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 10.620000 72.235000 10.940000 ;
      LAYER met4 ;
        RECT 71.915000 10.620000 72.235000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 11.050000 72.235000 11.370000 ;
      LAYER met4 ;
        RECT 71.915000 11.050000 72.235000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 11.480000 72.235000 11.800000 ;
      LAYER met4 ;
        RECT 71.915000 11.480000 72.235000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 11.910000 72.235000 12.230000 ;
      LAYER met4 ;
        RECT 71.915000 11.910000 72.235000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 12.340000 72.235000 12.660000 ;
      LAYER met4 ;
        RECT 71.915000 12.340000 72.235000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 12.770000 72.235000 13.090000 ;
      LAYER met4 ;
        RECT 71.915000 12.770000 72.235000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 13.200000 72.235000 13.520000 ;
      LAYER met4 ;
        RECT 71.915000 13.200000 72.235000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 8.900000 72.235000 9.220000 ;
      LAYER met4 ;
        RECT 71.915000 8.900000 72.235000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 9.330000 72.235000 9.650000 ;
      LAYER met4 ;
        RECT 71.915000 9.330000 72.235000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 9.760000 72.235000 10.080000 ;
      LAYER met4 ;
        RECT 71.915000 9.760000 72.235000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 10.190000 72.640000 10.510000 ;
      LAYER met4 ;
        RECT 72.320000 10.190000 72.640000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 10.620000 72.640000 10.940000 ;
      LAYER met4 ;
        RECT 72.320000 10.620000 72.640000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 11.050000 72.640000 11.370000 ;
      LAYER met4 ;
        RECT 72.320000 11.050000 72.640000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 11.480000 72.640000 11.800000 ;
      LAYER met4 ;
        RECT 72.320000 11.480000 72.640000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 11.910000 72.640000 12.230000 ;
      LAYER met4 ;
        RECT 72.320000 11.910000 72.640000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 12.340000 72.640000 12.660000 ;
      LAYER met4 ;
        RECT 72.320000 12.340000 72.640000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 12.770000 72.640000 13.090000 ;
      LAYER met4 ;
        RECT 72.320000 12.770000 72.640000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 13.200000 72.640000 13.520000 ;
      LAYER met4 ;
        RECT 72.320000 13.200000 72.640000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 8.900000 72.640000 9.220000 ;
      LAYER met4 ;
        RECT 72.320000 8.900000 72.640000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 9.330000 72.640000 9.650000 ;
      LAYER met4 ;
        RECT 72.320000 9.330000 72.640000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 9.760000 72.640000 10.080000 ;
      LAYER met4 ;
        RECT 72.320000 9.760000 72.640000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 10.190000 73.045000 10.510000 ;
      LAYER met4 ;
        RECT 72.725000 10.190000 73.045000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 10.620000 73.045000 10.940000 ;
      LAYER met4 ;
        RECT 72.725000 10.620000 73.045000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 11.050000 73.045000 11.370000 ;
      LAYER met4 ;
        RECT 72.725000 11.050000 73.045000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 11.480000 73.045000 11.800000 ;
      LAYER met4 ;
        RECT 72.725000 11.480000 73.045000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 11.910000 73.045000 12.230000 ;
      LAYER met4 ;
        RECT 72.725000 11.910000 73.045000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 12.340000 73.045000 12.660000 ;
      LAYER met4 ;
        RECT 72.725000 12.340000 73.045000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 12.770000 73.045000 13.090000 ;
      LAYER met4 ;
        RECT 72.725000 12.770000 73.045000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 13.200000 73.045000 13.520000 ;
      LAYER met4 ;
        RECT 72.725000 13.200000 73.045000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 8.900000 73.045000 9.220000 ;
      LAYER met4 ;
        RECT 72.725000 8.900000 73.045000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 9.330000 73.045000 9.650000 ;
      LAYER met4 ;
        RECT 72.725000 9.330000 73.045000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 9.760000 73.045000 10.080000 ;
      LAYER met4 ;
        RECT 72.725000 9.760000 73.045000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 10.190000 73.450000 10.510000 ;
      LAYER met4 ;
        RECT 73.130000 10.190000 73.450000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 10.620000 73.450000 10.940000 ;
      LAYER met4 ;
        RECT 73.130000 10.620000 73.450000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 11.050000 73.450000 11.370000 ;
      LAYER met4 ;
        RECT 73.130000 11.050000 73.450000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 11.480000 73.450000 11.800000 ;
      LAYER met4 ;
        RECT 73.130000 11.480000 73.450000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 11.910000 73.450000 12.230000 ;
      LAYER met4 ;
        RECT 73.130000 11.910000 73.450000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 12.340000 73.450000 12.660000 ;
      LAYER met4 ;
        RECT 73.130000 12.340000 73.450000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 12.770000 73.450000 13.090000 ;
      LAYER met4 ;
        RECT 73.130000 12.770000 73.450000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 13.200000 73.450000 13.520000 ;
      LAYER met4 ;
        RECT 73.130000 13.200000 73.450000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 8.900000 73.450000 9.220000 ;
      LAYER met4 ;
        RECT 73.130000 8.900000 73.450000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 9.330000 73.450000 9.650000 ;
      LAYER met4 ;
        RECT 73.130000 9.330000 73.450000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 9.760000 73.450000 10.080000 ;
      LAYER met4 ;
        RECT 73.130000 9.760000 73.450000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 10.190000 73.855000 10.510000 ;
      LAYER met4 ;
        RECT 73.535000 10.190000 73.855000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 10.620000 73.855000 10.940000 ;
      LAYER met4 ;
        RECT 73.535000 10.620000 73.855000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 11.050000 73.855000 11.370000 ;
      LAYER met4 ;
        RECT 73.535000 11.050000 73.855000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 11.480000 73.855000 11.800000 ;
      LAYER met4 ;
        RECT 73.535000 11.480000 73.855000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 11.910000 73.855000 12.230000 ;
      LAYER met4 ;
        RECT 73.535000 11.910000 73.855000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 12.340000 73.855000 12.660000 ;
      LAYER met4 ;
        RECT 73.535000 12.340000 73.855000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 12.770000 73.855000 13.090000 ;
      LAYER met4 ;
        RECT 73.535000 12.770000 73.855000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 13.200000 73.855000 13.520000 ;
      LAYER met4 ;
        RECT 73.535000 13.200000 73.855000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 8.900000 73.855000 9.220000 ;
      LAYER met4 ;
        RECT 73.535000 8.900000 73.855000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 9.330000 73.855000 9.650000 ;
      LAYER met4 ;
        RECT 73.535000 9.330000 73.855000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 9.760000 73.855000 10.080000 ;
      LAYER met4 ;
        RECT 73.535000 9.760000 73.855000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 10.190000 74.260000 10.510000 ;
      LAYER met4 ;
        RECT 73.940000 10.190000 74.260000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 10.620000 74.260000 10.940000 ;
      LAYER met4 ;
        RECT 73.940000 10.620000 74.260000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 11.050000 74.260000 11.370000 ;
      LAYER met4 ;
        RECT 73.940000 11.050000 74.260000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 11.480000 74.260000 11.800000 ;
      LAYER met4 ;
        RECT 73.940000 11.480000 74.260000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 11.910000 74.260000 12.230000 ;
      LAYER met4 ;
        RECT 73.940000 11.910000 74.260000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 12.340000 74.260000 12.660000 ;
      LAYER met4 ;
        RECT 73.940000 12.340000 74.260000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 12.770000 74.260000 13.090000 ;
      LAYER met4 ;
        RECT 73.940000 12.770000 74.260000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 13.200000 74.260000 13.520000 ;
      LAYER met4 ;
        RECT 73.940000 13.200000 74.260000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 8.900000 74.260000 9.220000 ;
      LAYER met4 ;
        RECT 73.940000 8.900000 74.260000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 9.330000 74.260000 9.650000 ;
      LAYER met4 ;
        RECT 73.940000 9.330000 74.260000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 9.760000 74.260000 10.080000 ;
      LAYER met4 ;
        RECT 73.940000 9.760000 74.260000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 10.190000 8.570000 10.510000 ;
      LAYER met4 ;
        RECT 8.250000 10.190000 8.570000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 10.620000 8.570000 10.940000 ;
      LAYER met4 ;
        RECT 8.250000 10.620000 8.570000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 11.050000 8.570000 11.370000 ;
      LAYER met4 ;
        RECT 8.250000 11.050000 8.570000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 11.480000 8.570000 11.800000 ;
      LAYER met4 ;
        RECT 8.250000 11.480000 8.570000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 11.910000 8.570000 12.230000 ;
      LAYER met4 ;
        RECT 8.250000 11.910000 8.570000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 12.340000 8.570000 12.660000 ;
      LAYER met4 ;
        RECT 8.250000 12.340000 8.570000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 12.770000 8.570000 13.090000 ;
      LAYER met4 ;
        RECT 8.250000 12.770000 8.570000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 13.200000 8.570000 13.520000 ;
      LAYER met4 ;
        RECT 8.250000 13.200000 8.570000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 8.900000 8.570000 9.220000 ;
      LAYER met4 ;
        RECT 8.250000 8.900000 8.570000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 9.330000 8.570000 9.650000 ;
      LAYER met4 ;
        RECT 8.250000 9.330000 8.570000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 9.760000 8.570000 10.080000 ;
      LAYER met4 ;
        RECT 8.250000 9.760000 8.570000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 10.190000 8.975000 10.510000 ;
      LAYER met4 ;
        RECT 8.655000 10.190000 8.975000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 10.620000 8.975000 10.940000 ;
      LAYER met4 ;
        RECT 8.655000 10.620000 8.975000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 11.050000 8.975000 11.370000 ;
      LAYER met4 ;
        RECT 8.655000 11.050000 8.975000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 11.480000 8.975000 11.800000 ;
      LAYER met4 ;
        RECT 8.655000 11.480000 8.975000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 11.910000 8.975000 12.230000 ;
      LAYER met4 ;
        RECT 8.655000 11.910000 8.975000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 12.340000 8.975000 12.660000 ;
      LAYER met4 ;
        RECT 8.655000 12.340000 8.975000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 12.770000 8.975000 13.090000 ;
      LAYER met4 ;
        RECT 8.655000 12.770000 8.975000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 13.200000 8.975000 13.520000 ;
      LAYER met4 ;
        RECT 8.655000 13.200000 8.975000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 8.900000 8.975000 9.220000 ;
      LAYER met4 ;
        RECT 8.655000 8.900000 8.975000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 9.330000 8.975000 9.650000 ;
      LAYER met4 ;
        RECT 8.655000 9.330000 8.975000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 9.760000 8.975000 10.080000 ;
      LAYER met4 ;
        RECT 8.655000 9.760000 8.975000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 10.190000 9.380000 10.510000 ;
      LAYER met4 ;
        RECT 9.060000 10.190000 9.380000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 10.620000 9.380000 10.940000 ;
      LAYER met4 ;
        RECT 9.060000 10.620000 9.380000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 11.050000 9.380000 11.370000 ;
      LAYER met4 ;
        RECT 9.060000 11.050000 9.380000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 11.480000 9.380000 11.800000 ;
      LAYER met4 ;
        RECT 9.060000 11.480000 9.380000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 11.910000 9.380000 12.230000 ;
      LAYER met4 ;
        RECT 9.060000 11.910000 9.380000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 12.340000 9.380000 12.660000 ;
      LAYER met4 ;
        RECT 9.060000 12.340000 9.380000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 12.770000 9.380000 13.090000 ;
      LAYER met4 ;
        RECT 9.060000 12.770000 9.380000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 13.200000 9.380000 13.520000 ;
      LAYER met4 ;
        RECT 9.060000 13.200000 9.380000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 8.900000 9.380000 9.220000 ;
      LAYER met4 ;
        RECT 9.060000 8.900000 9.380000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 9.330000 9.380000 9.650000 ;
      LAYER met4 ;
        RECT 9.060000 9.330000 9.380000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 9.760000 9.380000 10.080000 ;
      LAYER met4 ;
        RECT 9.060000 9.760000 9.380000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 10.190000 9.785000 10.510000 ;
      LAYER met4 ;
        RECT 9.465000 10.190000 9.785000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 10.620000 9.785000 10.940000 ;
      LAYER met4 ;
        RECT 9.465000 10.620000 9.785000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 11.050000 9.785000 11.370000 ;
      LAYER met4 ;
        RECT 9.465000 11.050000 9.785000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 11.480000 9.785000 11.800000 ;
      LAYER met4 ;
        RECT 9.465000 11.480000 9.785000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 11.910000 9.785000 12.230000 ;
      LAYER met4 ;
        RECT 9.465000 11.910000 9.785000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 12.340000 9.785000 12.660000 ;
      LAYER met4 ;
        RECT 9.465000 12.340000 9.785000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 12.770000 9.785000 13.090000 ;
      LAYER met4 ;
        RECT 9.465000 12.770000 9.785000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 13.200000 9.785000 13.520000 ;
      LAYER met4 ;
        RECT 9.465000 13.200000 9.785000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 8.900000 9.785000 9.220000 ;
      LAYER met4 ;
        RECT 9.465000 8.900000 9.785000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 9.330000 9.785000 9.650000 ;
      LAYER met4 ;
        RECT 9.465000 9.330000 9.785000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 9.760000 9.785000 10.080000 ;
      LAYER met4 ;
        RECT 9.465000 9.760000 9.785000 10.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 10.190000 10.190000 10.510000 ;
      LAYER met4 ;
        RECT 9.870000 10.190000 10.190000 10.510000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 10.620000 10.190000 10.940000 ;
      LAYER met4 ;
        RECT 9.870000 10.620000 10.190000 10.940000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 11.050000 10.190000 11.370000 ;
      LAYER met4 ;
        RECT 9.870000 11.050000 10.190000 11.370000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 11.480000 10.190000 11.800000 ;
      LAYER met4 ;
        RECT 9.870000 11.480000 10.190000 11.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 11.910000 10.190000 12.230000 ;
      LAYER met4 ;
        RECT 9.870000 11.910000 10.190000 12.230000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 12.340000 10.190000 12.660000 ;
      LAYER met4 ;
        RECT 9.870000 12.340000 10.190000 12.660000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 12.770000 10.190000 13.090000 ;
      LAYER met4 ;
        RECT 9.870000 12.770000 10.190000 13.090000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 13.200000 10.190000 13.520000 ;
      LAYER met4 ;
        RECT 9.870000 13.200000 10.190000 13.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 8.900000 10.190000 9.220000 ;
      LAYER met4 ;
        RECT 9.870000 8.900000 10.190000 9.220000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 9.330000 10.190000 9.650000 ;
      LAYER met4 ;
        RECT 9.870000 9.330000 10.190000 9.650000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 9.760000 10.190000 10.080000 ;
      LAYER met4 ;
        RECT 9.870000 9.760000 10.190000 10.080000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 47.735000 75.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met3 ;
      RECT 0.495000 8.890000 74.290000 13.530000 ;
    LAYER met4 ;
      RECT 0.000000  2.035000 75.000000  47.965000 ;
      RECT 0.000000 51.745000 75.000000  52.725000 ;
      RECT 0.000000 56.505000 75.000000 200.000000 ;
    LAYER met5 ;
      RECT 0.000000  2.135000 72.130000   8.985000 ;
      RECT 0.000000  8.985000 75.000000  13.435000 ;
      RECT 0.000000 13.435000 72.435000  19.885000 ;
      RECT 0.000000 19.885000 75.000000  24.335000 ;
      RECT 0.000000 24.335000 72.130000  36.835000 ;
      RECT 0.000000 36.835000 75.000000  40.085000 ;
      RECT 0.000000 40.085000 72.130000  96.585000 ;
      RECT 0.000000 96.585000 75.000000 200.000000 ;
  END
END sky130_fd_io__overlay_vccd_hvc
END LIBRARY
