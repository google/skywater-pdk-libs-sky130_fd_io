/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_IO__TOP_GPIO_OVTV2_PP_SYMBOL_V
`define SKY130_FD_IO__TOP_GPIO_OVTV2_PP_SYMBOL_V

/**
 * top_gpio_ovtv2: General Purpose I/0.
 *
 * Verilog stub (with power pins) for graphical symbol definition
 * generation.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_io__top_gpio_ovtv2 (
           //# {{data|Data Signals}}
           input        SLOW            ,
           output       IN              ,
           input        INP_DIS         ,
           output       IN_H            ,
           input        OUT             ,
           inout        PAD             ,
           inout        PAD_A_ESD_0_H   ,
           inout        PAD_A_ESD_1_H   ,
           inout        PAD_A_NOESD_H   ,

           //# {{control|Control Signals}}
           inout        AMUXBUS_A       ,
           inout        AMUXBUS_B       ,
           input        ANALOG_EN       ,
           input        ANALOG_POL      ,
           input        ANALOG_SEL      ,
           input  [2:0] DM              ,
           input        ENABLE_H        ,
           input        ENABLE_INP_H    ,
           input        ENABLE_VDDA_H   ,
           input        ENABLE_VDDIO    ,
           input        ENABLE_VSWITCH_H,
           input        HLD_H_N         ,
           input        HLD_OVR         ,
           input        HYS_TRIM        ,
           input  [1:0] IB_MODE_SEL     ,
           input        OE_N            ,
           input  [1:0] SLEW_CTL        ,

           //# {{power|Power}}
           input        VTRIP_SEL       ,
           inout        VSWITCH         ,
           inout        VCCD            ,
           inout        VCCHIB          ,
           inout        VDDA            ,
           inout        VDDIO           ,
           inout        VDDIO_Q         ,
           output       TIE_HI_ESD      ,
           input        VINREF          ,
           inout        VSSA            ,
           inout        VSSD            ,
           inout        VSSIO           ,
           inout        VSSIO_Q         ,
           output       TIE_LO_ESD
       );
endmodule

`default_nettype wire
`endif  // SKY130_FD_IO__TOP_GPIO_OVTV2_PP_SYMBOL_V
