# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__top_refgen_new
  CLASS BLOCK ;
  FOREIGN sky130_fd_io__top_refgen_new ;
  ORIGIN  0.620000  0.000000 ;
  SIZE  93.72500 BY  253.7150 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 63.465000 0.000000 63.725000 67.115000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 64.215000 0.000000 64.475000 65.625000 ;
    END
  END AMUXBUS_B
  PIN DFT_REFGEN
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.215000 0.000000 67.475000 236.650000 ;
    END
  END DFT_REFGEN
  PIN ENABLE_H
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.215000 0.000000 70.475000 15.535000 ;
    END
  END ENABLE_H
  PIN ENABLE_VDDA_H
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.965000 0.000000 68.225000 234.180000 ;
    END
  END ENABLE_VDDA_H
  PIN HLD_H_N
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.555000 0.000000 20.815000 14.810000 ;
    END
  END HLD_H_N
  PIN IBUF_SEL
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.250000 0.000000 38.510000 22.530000 ;
    END
  END IBUF_SEL
  PIN REFLEAK_BIAS
    DIRECTION INOUT ;
    PORT
      LAYER met1 ;
        RECT 0.000000 199.485000 7.485000 199.715000 ;
    END
  END REFLEAK_BIAS
  PIN VCCD
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000000 46.015000 31.300000 58.995000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000000 11.670000 55.235000 17.860000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 83.360000 21.960000 84.750000 50.130000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    PORT
      LAYER met1 ;
        RECT 37.420000 205.620000 38.505000 205.805000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 1.835000 25.250000 10.660000 31.440000 ;
    END
  END VDDIO_Q
  PIN VINREF
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 0.080000 28.495000 14.480000 28.755000 ;
    END
  END VINREF
  PIN VINREF_DFT
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 81.590000 0.000000 82.230000 49.025000 ;
    END
  END VINREF_DFT
  PIN VOHREF
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.005000 0.000000 35.265000 4.425000 ;
    END
  END VOHREF
  PIN VOH_SEL[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.965000 0.000000 65.225000 83.625000 ;
    END
  END VOH_SEL[0]
  PIN VOH_SEL[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.715000 0.000000 65.975000 236.010000 ;
    END
  END VOH_SEL[1]
  PIN VOH_SEL[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.465000 0.000000 66.725000 236.330000 ;
    END
  END VOH_SEL[2]
  PIN VOUTREF
    DIRECTION OUTPUT ;
    PORT
      LAYER met1 ;
        RECT 0.000000 200.680000 40.510000 200.940000 ;
    END
  END VOUTREF
  PIN VOUTREF_DFT
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 80.090000 0.000000 80.730000 59.975000 ;
    END
  END VOUTREF_DFT
  PIN VREF_SEL[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.715000 0.000000 68.975000 15.430000 ;
    END
  END VREF_SEL[0]
  PIN VREF_SEL[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.465000 0.000000 69.725000 16.050000 ;
    END
  END VREF_SEL[1]
  PIN VREG_EN
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 60.400000 0.000000 60.660000 16.695000 ;
    END
  END VREG_EN
  PIN VSSA
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 85.430000 36.720000 86.950000 52.700000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 42.275000 32.040000 58.995000 38.625000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    PORT
      LAYER met1 ;
        RECT 37.420000 205.185000 38.505000 205.370000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    PORT
      LAYER met1 ;
        RECT 37.420000 204.755000 38.505000 204.940000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 77.565000 7.300000 78.575000 44.560000 ;
    END
  END VSWITCH
  PIN VTRIP_SEL
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.400000 0.000000 18.660000 22.530000 ;
    END
  END VTRIP_SEL
  OBS
    LAYER li1 ;
      RECT -0.290000 0.130000 93.075000 253.585000 ;
    LAYER met1 ;
      RECT -0.290000   0.070000 93.105000  28.215000 ;
      RECT -0.290000  28.215000 -0.200000  29.035000 ;
      RECT -0.290000  29.035000 93.105000 199.205000 ;
      RECT -0.290000 199.205000 -0.280000 199.995000 ;
      RECT -0.290000 199.995000 93.105000 200.400000 ;
      RECT -0.290000 200.400000 -0.280000 201.220000 ;
      RECT -0.290000 201.220000 93.105000 204.475000 ;
      RECT -0.290000 204.475000 37.140000 206.085000 ;
      RECT -0.290000 206.085000 93.105000 253.645000 ;
      RECT  7.765000 199.205000 93.105000 199.995000 ;
      RECT 14.760000  28.215000 93.105000  29.035000 ;
      RECT 38.785000 204.475000 93.105000 206.085000 ;
      RECT 40.790000 200.400000 93.105000 201.220000 ;
    LAYER met2 ;
      RECT -0.590000   1.825000 18.120000  22.810000 ;
      RECT -0.590000  22.810000 63.185000  67.395000 ;
      RECT -0.590000  67.395000 64.685000  83.905000 ;
      RECT -0.590000  83.905000 65.435000 236.290000 ;
      RECT -0.590000 236.290000 66.185000 236.610000 ;
      RECT -0.590000 236.610000 66.935000 236.930000 ;
      RECT -0.590000 236.930000 89.620000 253.400000 ;
      RECT 18.940000   1.825000 20.275000  15.090000 ;
      RECT 18.940000  15.090000 37.970000  22.810000 ;
      RECT 21.095000   1.825000 34.725000   4.705000 ;
      RECT 21.095000   4.705000 37.970000  15.090000 ;
      RECT 35.545000   1.825000 37.970000   4.705000 ;
      RECT 38.790000   1.825000 60.120000  16.975000 ;
      RECT 38.790000  16.975000 63.185000  22.810000 ;
      RECT 60.940000   1.825000 63.185000  16.975000 ;
      RECT 64.005000  65.905000 64.685000  67.395000 ;
      RECT 67.755000 234.460000 89.620000 236.930000 ;
      RECT 68.505000  15.710000 69.185000  16.330000 ;
      RECT 68.505000  16.330000 77.285000  44.840000 ;
      RECT 68.505000  44.840000 79.810000  60.255000 ;
      RECT 68.505000  60.255000 89.620000 234.460000 ;
      RECT 70.005000  15.815000 77.285000  16.330000 ;
      RECT 70.755000   1.825000 79.810000   7.020000 ;
      RECT 70.755000   7.020000 77.285000  15.815000 ;
      RECT 78.855000   7.020000 79.810000  44.840000 ;
      RECT 81.010000   1.825000 81.310000  49.305000 ;
      RECT 81.010000  49.305000 83.080000  50.410000 ;
      RECT 81.010000  50.410000 85.150000  52.980000 ;
      RECT 81.010000  52.980000 89.620000  60.255000 ;
      RECT 82.510000   1.825000 89.620000  21.680000 ;
      RECT 82.510000  21.680000 83.080000  49.305000 ;
      RECT 85.030000  21.680000 89.620000  36.440000 ;
      RECT 85.030000  36.440000 85.150000  50.410000 ;
      RECT 87.230000  36.440000 89.620000  52.980000 ;
    LAYER met3 ;
      RECT  0.000000  5.830000 89.645000  11.270000 ;
      RECT  0.000000 18.260000 89.645000  24.850000 ;
      RECT  0.000000 24.850000  1.435000  31.840000 ;
      RECT  0.000000 31.840000 41.875000  39.025000 ;
      RECT  0.000000 39.025000 89.645000  45.615000 ;
      RECT  0.000000 59.395000 89.645000 206.260000 ;
      RECT 11.060000 24.850000 89.645000  31.640000 ;
      RECT 11.060000 31.640000 41.875000  31.840000 ;
      RECT 31.700000 45.615000 89.645000  59.395000 ;
      RECT 55.635000 11.270000 89.645000  18.260000 ;
      RECT 59.395000 31.640000 89.645000  39.025000 ;
    LAYER met4 ;
      RECT 64.400000 104.305000 65.245000 109.790000 ;
  END
END sky130_fd_io__top_refgen_new
END LIBRARY
