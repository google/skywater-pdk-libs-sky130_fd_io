# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__overlay_vssa_hvc
  CLASS BLOCK ;
  FOREIGN sky130_fd_io__overlay_vssa_hvc ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  75.00000 BY  200.0000 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 75.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 75.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 8.985000 75.000000 13.435000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 2.135000 75.000000 7.385000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035000 15.035000 75.000000 18.285000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 70.035000 75.000000 94.985000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 64.185000 75.000000 68.435000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.525000 51.655000 0.845000 51.975000 ;
      LAYER met4 ;
        RECT 0.525000 51.655000 0.845000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 52.075000 0.845000 52.395000 ;
      LAYER met4 ;
        RECT 0.525000 52.075000 0.845000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525000 52.495000 0.845000 52.815000 ;
      LAYER met4 ;
        RECT 0.525000 52.495000 0.845000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.560000 47.740000 0.880000 48.060000 ;
      LAYER met4 ;
        RECT 0.560000 47.740000 0.880000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.560000 56.410000 0.880000 56.730000 ;
      LAYER met4 ;
        RECT 0.560000 56.410000 0.880000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 51.655000 1.255000 51.975000 ;
      LAYER met4 ;
        RECT 0.935000 51.655000 1.255000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 52.075000 1.255000 52.395000 ;
      LAYER met4 ;
        RECT 0.935000 52.075000 1.255000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935000 52.495000 1.255000 52.815000 ;
      LAYER met4 ;
        RECT 0.935000 52.495000 1.255000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.965000 47.740000 1.285000 48.060000 ;
      LAYER met4 ;
        RECT 0.965000 47.740000 1.285000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.965000 56.410000 1.285000 56.730000 ;
      LAYER met4 ;
        RECT 0.965000 56.410000 1.285000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000000 36.760000 1.320000 37.080000 ;
      LAYER met4 ;
        RECT 1.000000 36.760000 1.320000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000000 37.200000 1.320000 37.520000 ;
      LAYER met4 ;
        RECT 1.000000 37.200000 1.320000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000000 37.640000 1.320000 37.960000 ;
      LAYER met4 ;
        RECT 1.000000 37.640000 1.320000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000000 38.080000 1.320000 38.400000 ;
      LAYER met4 ;
        RECT 1.000000 38.080000 1.320000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000000 38.520000 1.320000 38.840000 ;
      LAYER met4 ;
        RECT 1.000000 38.520000 1.320000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000000 38.960000 1.320000 39.280000 ;
      LAYER met4 ;
        RECT 1.000000 38.960000 1.320000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000000 39.400000 1.320000 39.720000 ;
      LAYER met4 ;
        RECT 1.000000 39.400000 1.320000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000000 39.840000 1.320000 40.160000 ;
      LAYER met4 ;
        RECT 1.000000 39.840000 1.320000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 51.655000 1.665000 51.975000 ;
      LAYER met4 ;
        RECT 1.345000 51.655000 1.665000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 52.075000 1.665000 52.395000 ;
      LAYER met4 ;
        RECT 1.345000 52.075000 1.665000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345000 52.495000 1.665000 52.815000 ;
      LAYER met4 ;
        RECT 1.345000 52.495000 1.665000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.370000 47.740000 1.690000 48.060000 ;
      LAYER met4 ;
        RECT 1.370000 47.740000 1.690000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.370000 56.410000 1.690000 56.730000 ;
      LAYER met4 ;
        RECT 1.370000 56.410000 1.690000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405000 36.760000 1.725000 37.080000 ;
      LAYER met4 ;
        RECT 1.405000 36.760000 1.725000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405000 37.200000 1.725000 37.520000 ;
      LAYER met4 ;
        RECT 1.405000 37.200000 1.725000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405000 37.640000 1.725000 37.960000 ;
      LAYER met4 ;
        RECT 1.405000 37.640000 1.725000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405000 38.080000 1.725000 38.400000 ;
      LAYER met4 ;
        RECT 1.405000 38.080000 1.725000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405000 38.520000 1.725000 38.840000 ;
      LAYER met4 ;
        RECT 1.405000 38.520000 1.725000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405000 38.960000 1.725000 39.280000 ;
      LAYER met4 ;
        RECT 1.405000 38.960000 1.725000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405000 39.400000 1.725000 39.720000 ;
      LAYER met4 ;
        RECT 1.405000 39.400000 1.725000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405000 39.840000 1.725000 40.160000 ;
      LAYER met4 ;
        RECT 1.405000 39.840000 1.725000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 51.655000 2.075000 51.975000 ;
      LAYER met4 ;
        RECT 1.755000 51.655000 2.075000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 52.075000 2.075000 52.395000 ;
      LAYER met4 ;
        RECT 1.755000 52.075000 2.075000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755000 52.495000 2.075000 52.815000 ;
      LAYER met4 ;
        RECT 1.755000 52.495000 2.075000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.775000 47.740000 2.095000 48.060000 ;
      LAYER met4 ;
        RECT 1.775000 47.740000 2.095000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.775000 56.410000 2.095000 56.730000 ;
      LAYER met4 ;
        RECT 1.775000 56.410000 2.095000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810000 36.760000 2.130000 37.080000 ;
      LAYER met4 ;
        RECT 1.810000 36.760000 2.130000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810000 37.200000 2.130000 37.520000 ;
      LAYER met4 ;
        RECT 1.810000 37.200000 2.130000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810000 37.640000 2.130000 37.960000 ;
      LAYER met4 ;
        RECT 1.810000 37.640000 2.130000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810000 38.080000 2.130000 38.400000 ;
      LAYER met4 ;
        RECT 1.810000 38.080000 2.130000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810000 38.520000 2.130000 38.840000 ;
      LAYER met4 ;
        RECT 1.810000 38.520000 2.130000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810000 38.960000 2.130000 39.280000 ;
      LAYER met4 ;
        RECT 1.810000 38.960000 2.130000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810000 39.400000 2.130000 39.720000 ;
      LAYER met4 ;
        RECT 1.810000 39.400000 2.130000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810000 39.840000 2.130000 40.160000 ;
      LAYER met4 ;
        RECT 1.810000 39.840000 2.130000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 51.655000 10.595000 51.975000 ;
      LAYER met4 ;
        RECT 10.275000 51.655000 10.595000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 52.075000 10.595000 52.395000 ;
      LAYER met4 ;
        RECT 10.275000 52.075000 10.595000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275000 52.495000 10.595000 52.815000 ;
      LAYER met4 ;
        RECT 10.275000 52.495000 10.595000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 47.740000 10.600000 48.060000 ;
      LAYER met4 ;
        RECT 10.280000 47.740000 10.600000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280000 56.410000 10.600000 56.730000 ;
      LAYER met4 ;
        RECT 10.280000 56.410000 10.600000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315000 36.760000 10.635000 37.080000 ;
      LAYER met4 ;
        RECT 10.315000 36.760000 10.635000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315000 37.200000 10.635000 37.520000 ;
      LAYER met4 ;
        RECT 10.315000 37.200000 10.635000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315000 37.640000 10.635000 37.960000 ;
      LAYER met4 ;
        RECT 10.315000 37.640000 10.635000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315000 38.080000 10.635000 38.400000 ;
      LAYER met4 ;
        RECT 10.315000 38.080000 10.635000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315000 38.520000 10.635000 38.840000 ;
      LAYER met4 ;
        RECT 10.315000 38.520000 10.635000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315000 38.960000 10.635000 39.280000 ;
      LAYER met4 ;
        RECT 10.315000 38.960000 10.635000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315000 39.400000 10.635000 39.720000 ;
      LAYER met4 ;
        RECT 10.315000 39.400000 10.635000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315000 39.840000 10.635000 40.160000 ;
      LAYER met4 ;
        RECT 10.315000 39.840000 10.635000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 51.655000 11.000000 51.975000 ;
      LAYER met4 ;
        RECT 10.680000 51.655000 11.000000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 52.075000 11.000000 52.395000 ;
      LAYER met4 ;
        RECT 10.680000 52.075000 11.000000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680000 52.495000 11.000000 52.815000 ;
      LAYER met4 ;
        RECT 10.680000 52.495000 11.000000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 47.740000 11.005000 48.060000 ;
      LAYER met4 ;
        RECT 10.685000 47.740000 11.005000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685000 56.410000 11.005000 56.730000 ;
      LAYER met4 ;
        RECT 10.685000 56.410000 11.005000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720000 36.760000 11.040000 37.080000 ;
      LAYER met4 ;
        RECT 10.720000 36.760000 11.040000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720000 37.200000 11.040000 37.520000 ;
      LAYER met4 ;
        RECT 10.720000 37.200000 11.040000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720000 37.640000 11.040000 37.960000 ;
      LAYER met4 ;
        RECT 10.720000 37.640000 11.040000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720000 38.080000 11.040000 38.400000 ;
      LAYER met4 ;
        RECT 10.720000 38.080000 11.040000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720000 38.520000 11.040000 38.840000 ;
      LAYER met4 ;
        RECT 10.720000 38.520000 11.040000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720000 38.960000 11.040000 39.280000 ;
      LAYER met4 ;
        RECT 10.720000 38.960000 11.040000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720000 39.400000 11.040000 39.720000 ;
      LAYER met4 ;
        RECT 10.720000 39.400000 11.040000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720000 39.840000 11.040000 40.160000 ;
      LAYER met4 ;
        RECT 10.720000 39.840000 11.040000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 51.655000 11.405000 51.975000 ;
      LAYER met4 ;
        RECT 11.085000 51.655000 11.405000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 52.075000 11.405000 52.395000 ;
      LAYER met4 ;
        RECT 11.085000 52.075000 11.405000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085000 52.495000 11.405000 52.815000 ;
      LAYER met4 ;
        RECT 11.085000 52.495000 11.405000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 47.740000 11.410000 48.060000 ;
      LAYER met4 ;
        RECT 11.090000 47.740000 11.410000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090000 56.410000 11.410000 56.730000 ;
      LAYER met4 ;
        RECT 11.090000 56.410000 11.410000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125000 36.760000 11.445000 37.080000 ;
      LAYER met4 ;
        RECT 11.125000 36.760000 11.445000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125000 37.200000 11.445000 37.520000 ;
      LAYER met4 ;
        RECT 11.125000 37.200000 11.445000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125000 37.640000 11.445000 37.960000 ;
      LAYER met4 ;
        RECT 11.125000 37.640000 11.445000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125000 38.080000 11.445000 38.400000 ;
      LAYER met4 ;
        RECT 11.125000 38.080000 11.445000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125000 38.520000 11.445000 38.840000 ;
      LAYER met4 ;
        RECT 11.125000 38.520000 11.445000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125000 38.960000 11.445000 39.280000 ;
      LAYER met4 ;
        RECT 11.125000 38.960000 11.445000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125000 39.400000 11.445000 39.720000 ;
      LAYER met4 ;
        RECT 11.125000 39.400000 11.445000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125000 39.840000 11.445000 40.160000 ;
      LAYER met4 ;
        RECT 11.125000 39.840000 11.445000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 51.655000 11.810000 51.975000 ;
      LAYER met4 ;
        RECT 11.490000 51.655000 11.810000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 52.075000 11.810000 52.395000 ;
      LAYER met4 ;
        RECT 11.490000 52.075000 11.810000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490000 52.495000 11.810000 52.815000 ;
      LAYER met4 ;
        RECT 11.490000 52.495000 11.810000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 47.740000 11.815000 48.060000 ;
      LAYER met4 ;
        RECT 11.495000 47.740000 11.815000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495000 56.410000 11.815000 56.730000 ;
      LAYER met4 ;
        RECT 11.495000 56.410000 11.815000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530000 36.760000 11.850000 37.080000 ;
      LAYER met4 ;
        RECT 11.530000 36.760000 11.850000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530000 37.200000 11.850000 37.520000 ;
      LAYER met4 ;
        RECT 11.530000 37.200000 11.850000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530000 37.640000 11.850000 37.960000 ;
      LAYER met4 ;
        RECT 11.530000 37.640000 11.850000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530000 38.080000 11.850000 38.400000 ;
      LAYER met4 ;
        RECT 11.530000 38.080000 11.850000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530000 38.520000 11.850000 38.840000 ;
      LAYER met4 ;
        RECT 11.530000 38.520000 11.850000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530000 38.960000 11.850000 39.280000 ;
      LAYER met4 ;
        RECT 11.530000 38.960000 11.850000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530000 39.400000 11.850000 39.720000 ;
      LAYER met4 ;
        RECT 11.530000 39.400000 11.850000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530000 39.840000 11.850000 40.160000 ;
      LAYER met4 ;
        RECT 11.530000 39.840000 11.850000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 51.655000 12.215000 51.975000 ;
      LAYER met4 ;
        RECT 11.895000 51.655000 12.215000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 52.075000 12.215000 52.395000 ;
      LAYER met4 ;
        RECT 11.895000 52.075000 12.215000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895000 52.495000 12.215000 52.815000 ;
      LAYER met4 ;
        RECT 11.895000 52.495000 12.215000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 47.740000 12.220000 48.060000 ;
      LAYER met4 ;
        RECT 11.900000 47.740000 12.220000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900000 56.410000 12.220000 56.730000 ;
      LAYER met4 ;
        RECT 11.900000 56.410000 12.220000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935000 36.760000 12.255000 37.080000 ;
      LAYER met4 ;
        RECT 11.935000 36.760000 12.255000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935000 37.200000 12.255000 37.520000 ;
      LAYER met4 ;
        RECT 11.935000 37.200000 12.255000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935000 37.640000 12.255000 37.960000 ;
      LAYER met4 ;
        RECT 11.935000 37.640000 12.255000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935000 38.080000 12.255000 38.400000 ;
      LAYER met4 ;
        RECT 11.935000 38.080000 12.255000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935000 38.520000 12.255000 38.840000 ;
      LAYER met4 ;
        RECT 11.935000 38.520000 12.255000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935000 38.960000 12.255000 39.280000 ;
      LAYER met4 ;
        RECT 11.935000 38.960000 12.255000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935000 39.400000 12.255000 39.720000 ;
      LAYER met4 ;
        RECT 11.935000 39.400000 12.255000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935000 39.840000 12.255000 40.160000 ;
      LAYER met4 ;
        RECT 11.935000 39.840000 12.255000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 51.655000 12.620000 51.975000 ;
      LAYER met4 ;
        RECT 12.300000 51.655000 12.620000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 52.075000 12.620000 52.395000 ;
      LAYER met4 ;
        RECT 12.300000 52.075000 12.620000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300000 52.495000 12.620000 52.815000 ;
      LAYER met4 ;
        RECT 12.300000 52.495000 12.620000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 47.740000 12.625000 48.060000 ;
      LAYER met4 ;
        RECT 12.305000 47.740000 12.625000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305000 56.410000 12.625000 56.730000 ;
      LAYER met4 ;
        RECT 12.305000 56.410000 12.625000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340000 36.760000 12.660000 37.080000 ;
      LAYER met4 ;
        RECT 12.340000 36.760000 12.660000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340000 37.200000 12.660000 37.520000 ;
      LAYER met4 ;
        RECT 12.340000 37.200000 12.660000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340000 37.640000 12.660000 37.960000 ;
      LAYER met4 ;
        RECT 12.340000 37.640000 12.660000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340000 38.080000 12.660000 38.400000 ;
      LAYER met4 ;
        RECT 12.340000 38.080000 12.660000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340000 38.520000 12.660000 38.840000 ;
      LAYER met4 ;
        RECT 12.340000 38.520000 12.660000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340000 38.960000 12.660000 39.280000 ;
      LAYER met4 ;
        RECT 12.340000 38.960000 12.660000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340000 39.400000 12.660000 39.720000 ;
      LAYER met4 ;
        RECT 12.340000 39.400000 12.660000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340000 39.840000 12.660000 40.160000 ;
      LAYER met4 ;
        RECT 12.340000 39.840000 12.660000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 51.655000 13.025000 51.975000 ;
      LAYER met4 ;
        RECT 12.705000 51.655000 13.025000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 52.075000 13.025000 52.395000 ;
      LAYER met4 ;
        RECT 12.705000 52.075000 13.025000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705000 52.495000 13.025000 52.815000 ;
      LAYER met4 ;
        RECT 12.705000 52.495000 13.025000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 47.740000 13.030000 48.060000 ;
      LAYER met4 ;
        RECT 12.710000 47.740000 13.030000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710000 56.410000 13.030000 56.730000 ;
      LAYER met4 ;
        RECT 12.710000 56.410000 13.030000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745000 36.760000 13.065000 37.080000 ;
      LAYER met4 ;
        RECT 12.745000 36.760000 13.065000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745000 37.200000 13.065000 37.520000 ;
      LAYER met4 ;
        RECT 12.745000 37.200000 13.065000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745000 37.640000 13.065000 37.960000 ;
      LAYER met4 ;
        RECT 12.745000 37.640000 13.065000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745000 38.080000 13.065000 38.400000 ;
      LAYER met4 ;
        RECT 12.745000 38.080000 13.065000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745000 38.520000 13.065000 38.840000 ;
      LAYER met4 ;
        RECT 12.745000 38.520000 13.065000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745000 38.960000 13.065000 39.280000 ;
      LAYER met4 ;
        RECT 12.745000 38.960000 13.065000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745000 39.400000 13.065000 39.720000 ;
      LAYER met4 ;
        RECT 12.745000 39.400000 13.065000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745000 39.840000 13.065000 40.160000 ;
      LAYER met4 ;
        RECT 12.745000 39.840000 13.065000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 51.655000 13.430000 51.975000 ;
      LAYER met4 ;
        RECT 13.110000 51.655000 13.430000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 52.075000 13.430000 52.395000 ;
      LAYER met4 ;
        RECT 13.110000 52.075000 13.430000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110000 52.495000 13.430000 52.815000 ;
      LAYER met4 ;
        RECT 13.110000 52.495000 13.430000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 47.740000 13.435000 48.060000 ;
      LAYER met4 ;
        RECT 13.115000 47.740000 13.435000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115000 56.410000 13.435000 56.730000 ;
      LAYER met4 ;
        RECT 13.115000 56.410000 13.435000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150000 36.760000 13.470000 37.080000 ;
      LAYER met4 ;
        RECT 13.150000 36.760000 13.470000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150000 37.200000 13.470000 37.520000 ;
      LAYER met4 ;
        RECT 13.150000 37.200000 13.470000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150000 37.640000 13.470000 37.960000 ;
      LAYER met4 ;
        RECT 13.150000 37.640000 13.470000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150000 38.080000 13.470000 38.400000 ;
      LAYER met4 ;
        RECT 13.150000 38.080000 13.470000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150000 38.520000 13.470000 38.840000 ;
      LAYER met4 ;
        RECT 13.150000 38.520000 13.470000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150000 38.960000 13.470000 39.280000 ;
      LAYER met4 ;
        RECT 13.150000 38.960000 13.470000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150000 39.400000 13.470000 39.720000 ;
      LAYER met4 ;
        RECT 13.150000 39.400000 13.470000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150000 39.840000 13.470000 40.160000 ;
      LAYER met4 ;
        RECT 13.150000 39.840000 13.470000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 51.655000 13.835000 51.975000 ;
      LAYER met4 ;
        RECT 13.515000 51.655000 13.835000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 52.075000 13.835000 52.395000 ;
      LAYER met4 ;
        RECT 13.515000 52.075000 13.835000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515000 52.495000 13.835000 52.815000 ;
      LAYER met4 ;
        RECT 13.515000 52.495000 13.835000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 47.740000 13.840000 48.060000 ;
      LAYER met4 ;
        RECT 13.520000 47.740000 13.840000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520000 56.410000 13.840000 56.730000 ;
      LAYER met4 ;
        RECT 13.520000 56.410000 13.840000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555000 36.760000 13.875000 37.080000 ;
      LAYER met4 ;
        RECT 13.555000 36.760000 13.875000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555000 37.200000 13.875000 37.520000 ;
      LAYER met4 ;
        RECT 13.555000 37.200000 13.875000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555000 37.640000 13.875000 37.960000 ;
      LAYER met4 ;
        RECT 13.555000 37.640000 13.875000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555000 38.080000 13.875000 38.400000 ;
      LAYER met4 ;
        RECT 13.555000 38.080000 13.875000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555000 38.520000 13.875000 38.840000 ;
      LAYER met4 ;
        RECT 13.555000 38.520000 13.875000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555000 38.960000 13.875000 39.280000 ;
      LAYER met4 ;
        RECT 13.555000 38.960000 13.875000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555000 39.400000 13.875000 39.720000 ;
      LAYER met4 ;
        RECT 13.555000 39.400000 13.875000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555000 39.840000 13.875000 40.160000 ;
      LAYER met4 ;
        RECT 13.555000 39.840000 13.875000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 51.655000 14.240000 51.975000 ;
      LAYER met4 ;
        RECT 13.920000 51.655000 14.240000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 52.075000 14.240000 52.395000 ;
      LAYER met4 ;
        RECT 13.920000 52.075000 14.240000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920000 52.495000 14.240000 52.815000 ;
      LAYER met4 ;
        RECT 13.920000 52.495000 14.240000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 47.740000 14.245000 48.060000 ;
      LAYER met4 ;
        RECT 13.925000 47.740000 14.245000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925000 56.410000 14.245000 56.730000 ;
      LAYER met4 ;
        RECT 13.925000 56.410000 14.245000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960000 36.760000 14.280000 37.080000 ;
      LAYER met4 ;
        RECT 13.960000 36.760000 14.280000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960000 37.200000 14.280000 37.520000 ;
      LAYER met4 ;
        RECT 13.960000 37.200000 14.280000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960000 37.640000 14.280000 37.960000 ;
      LAYER met4 ;
        RECT 13.960000 37.640000 14.280000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960000 38.080000 14.280000 38.400000 ;
      LAYER met4 ;
        RECT 13.960000 38.080000 14.280000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960000 38.520000 14.280000 38.840000 ;
      LAYER met4 ;
        RECT 13.960000 38.520000 14.280000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960000 38.960000 14.280000 39.280000 ;
      LAYER met4 ;
        RECT 13.960000 38.960000 14.280000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960000 39.400000 14.280000 39.720000 ;
      LAYER met4 ;
        RECT 13.960000 39.400000 14.280000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960000 39.840000 14.280000 40.160000 ;
      LAYER met4 ;
        RECT 13.960000 39.840000 14.280000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 51.655000 14.645000 51.975000 ;
      LAYER met4 ;
        RECT 14.325000 51.655000 14.645000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 52.075000 14.645000 52.395000 ;
      LAYER met4 ;
        RECT 14.325000 52.075000 14.645000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325000 52.495000 14.645000 52.815000 ;
      LAYER met4 ;
        RECT 14.325000 52.495000 14.645000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 47.740000 14.650000 48.060000 ;
      LAYER met4 ;
        RECT 14.330000 47.740000 14.650000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330000 56.410000 14.650000 56.730000 ;
      LAYER met4 ;
        RECT 14.330000 56.410000 14.650000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365000 36.760000 14.685000 37.080000 ;
      LAYER met4 ;
        RECT 14.365000 36.760000 14.685000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365000 37.200000 14.685000 37.520000 ;
      LAYER met4 ;
        RECT 14.365000 37.200000 14.685000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365000 37.640000 14.685000 37.960000 ;
      LAYER met4 ;
        RECT 14.365000 37.640000 14.685000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365000 38.080000 14.685000 38.400000 ;
      LAYER met4 ;
        RECT 14.365000 38.080000 14.685000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365000 38.520000 14.685000 38.840000 ;
      LAYER met4 ;
        RECT 14.365000 38.520000 14.685000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365000 38.960000 14.685000 39.280000 ;
      LAYER met4 ;
        RECT 14.365000 38.960000 14.685000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365000 39.400000 14.685000 39.720000 ;
      LAYER met4 ;
        RECT 14.365000 39.400000 14.685000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365000 39.840000 14.685000 40.160000 ;
      LAYER met4 ;
        RECT 14.365000 39.840000 14.685000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 51.655000 15.050000 51.975000 ;
      LAYER met4 ;
        RECT 14.730000 51.655000 15.050000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 52.075000 15.050000 52.395000 ;
      LAYER met4 ;
        RECT 14.730000 52.075000 15.050000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730000 52.495000 15.050000 52.815000 ;
      LAYER met4 ;
        RECT 14.730000 52.495000 15.050000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 47.740000 15.055000 48.060000 ;
      LAYER met4 ;
        RECT 14.735000 47.740000 15.055000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735000 56.410000 15.055000 56.730000 ;
      LAYER met4 ;
        RECT 14.735000 56.410000 15.055000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770000 36.760000 15.090000 37.080000 ;
      LAYER met4 ;
        RECT 14.770000 36.760000 15.090000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770000 37.200000 15.090000 37.520000 ;
      LAYER met4 ;
        RECT 14.770000 37.200000 15.090000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770000 37.640000 15.090000 37.960000 ;
      LAYER met4 ;
        RECT 14.770000 37.640000 15.090000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770000 38.080000 15.090000 38.400000 ;
      LAYER met4 ;
        RECT 14.770000 38.080000 15.090000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770000 38.520000 15.090000 38.840000 ;
      LAYER met4 ;
        RECT 14.770000 38.520000 15.090000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770000 38.960000 15.090000 39.280000 ;
      LAYER met4 ;
        RECT 14.770000 38.960000 15.090000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770000 39.400000 15.090000 39.720000 ;
      LAYER met4 ;
        RECT 14.770000 39.400000 15.090000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770000 39.840000 15.090000 40.160000 ;
      LAYER met4 ;
        RECT 14.770000 39.840000 15.090000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 51.655000 15.455000 51.975000 ;
      LAYER met4 ;
        RECT 15.135000 51.655000 15.455000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 52.075000 15.455000 52.395000 ;
      LAYER met4 ;
        RECT 15.135000 52.075000 15.455000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135000 52.495000 15.455000 52.815000 ;
      LAYER met4 ;
        RECT 15.135000 52.495000 15.455000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 47.740000 15.460000 48.060000 ;
      LAYER met4 ;
        RECT 15.140000 47.740000 15.460000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140000 56.410000 15.460000 56.730000 ;
      LAYER met4 ;
        RECT 15.140000 56.410000 15.460000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175000 36.760000 15.495000 37.080000 ;
      LAYER met4 ;
        RECT 15.175000 36.760000 15.495000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175000 37.200000 15.495000 37.520000 ;
      LAYER met4 ;
        RECT 15.175000 37.200000 15.495000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175000 37.640000 15.495000 37.960000 ;
      LAYER met4 ;
        RECT 15.175000 37.640000 15.495000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175000 38.080000 15.495000 38.400000 ;
      LAYER met4 ;
        RECT 15.175000 38.080000 15.495000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175000 38.520000 15.495000 38.840000 ;
      LAYER met4 ;
        RECT 15.175000 38.520000 15.495000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175000 38.960000 15.495000 39.280000 ;
      LAYER met4 ;
        RECT 15.175000 38.960000 15.495000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175000 39.400000 15.495000 39.720000 ;
      LAYER met4 ;
        RECT 15.175000 39.400000 15.495000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175000 39.840000 15.495000 40.160000 ;
      LAYER met4 ;
        RECT 15.175000 39.840000 15.495000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 51.655000 15.860000 51.975000 ;
      LAYER met4 ;
        RECT 15.540000 51.655000 15.860000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 52.075000 15.860000 52.395000 ;
      LAYER met4 ;
        RECT 15.540000 52.075000 15.860000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540000 52.495000 15.860000 52.815000 ;
      LAYER met4 ;
        RECT 15.540000 52.495000 15.860000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 47.740000 15.865000 48.060000 ;
      LAYER met4 ;
        RECT 15.545000 47.740000 15.865000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545000 56.410000 15.865000 56.730000 ;
      LAYER met4 ;
        RECT 15.545000 56.410000 15.865000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580000 36.760000 15.900000 37.080000 ;
      LAYER met4 ;
        RECT 15.580000 36.760000 15.900000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580000 37.200000 15.900000 37.520000 ;
      LAYER met4 ;
        RECT 15.580000 37.200000 15.900000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580000 37.640000 15.900000 37.960000 ;
      LAYER met4 ;
        RECT 15.580000 37.640000 15.900000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580000 38.080000 15.900000 38.400000 ;
      LAYER met4 ;
        RECT 15.580000 38.080000 15.900000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580000 38.520000 15.900000 38.840000 ;
      LAYER met4 ;
        RECT 15.580000 38.520000 15.900000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580000 38.960000 15.900000 39.280000 ;
      LAYER met4 ;
        RECT 15.580000 38.960000 15.900000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580000 39.400000 15.900000 39.720000 ;
      LAYER met4 ;
        RECT 15.580000 39.400000 15.900000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580000 39.840000 15.900000 40.160000 ;
      LAYER met4 ;
        RECT 15.580000 39.840000 15.900000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 51.655000 16.265000 51.975000 ;
      LAYER met4 ;
        RECT 15.945000 51.655000 16.265000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 52.075000 16.265000 52.395000 ;
      LAYER met4 ;
        RECT 15.945000 52.075000 16.265000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945000 52.495000 16.265000 52.815000 ;
      LAYER met4 ;
        RECT 15.945000 52.495000 16.265000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 47.740000 16.270000 48.060000 ;
      LAYER met4 ;
        RECT 15.950000 47.740000 16.270000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950000 56.410000 16.270000 56.730000 ;
      LAYER met4 ;
        RECT 15.950000 56.410000 16.270000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 36.760000 16.305000 37.080000 ;
      LAYER met4 ;
        RECT 15.985000 36.760000 16.305000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 37.200000 16.305000 37.520000 ;
      LAYER met4 ;
        RECT 15.985000 37.200000 16.305000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 37.640000 16.305000 37.960000 ;
      LAYER met4 ;
        RECT 15.985000 37.640000 16.305000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 38.080000 16.305000 38.400000 ;
      LAYER met4 ;
        RECT 15.985000 38.080000 16.305000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 38.520000 16.305000 38.840000 ;
      LAYER met4 ;
        RECT 15.985000 38.520000 16.305000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 38.960000 16.305000 39.280000 ;
      LAYER met4 ;
        RECT 15.985000 38.960000 16.305000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 39.400000 16.305000 39.720000 ;
      LAYER met4 ;
        RECT 15.985000 39.400000 16.305000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985000 39.840000 16.305000 40.160000 ;
      LAYER met4 ;
        RECT 15.985000 39.840000 16.305000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 51.655000 16.670000 51.975000 ;
      LAYER met4 ;
        RECT 16.350000 51.655000 16.670000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 52.075000 16.670000 52.395000 ;
      LAYER met4 ;
        RECT 16.350000 52.075000 16.670000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350000 52.495000 16.670000 52.815000 ;
      LAYER met4 ;
        RECT 16.350000 52.495000 16.670000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 47.740000 16.675000 48.060000 ;
      LAYER met4 ;
        RECT 16.355000 47.740000 16.675000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355000 56.410000 16.675000 56.730000 ;
      LAYER met4 ;
        RECT 16.355000 56.410000 16.675000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390000 36.760000 16.710000 37.080000 ;
      LAYER met4 ;
        RECT 16.390000 36.760000 16.710000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390000 37.200000 16.710000 37.520000 ;
      LAYER met4 ;
        RECT 16.390000 37.200000 16.710000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390000 37.640000 16.710000 37.960000 ;
      LAYER met4 ;
        RECT 16.390000 37.640000 16.710000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390000 38.080000 16.710000 38.400000 ;
      LAYER met4 ;
        RECT 16.390000 38.080000 16.710000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390000 38.520000 16.710000 38.840000 ;
      LAYER met4 ;
        RECT 16.390000 38.520000 16.710000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390000 38.960000 16.710000 39.280000 ;
      LAYER met4 ;
        RECT 16.390000 38.960000 16.710000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390000 39.400000 16.710000 39.720000 ;
      LAYER met4 ;
        RECT 16.390000 39.400000 16.710000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390000 39.840000 16.710000 40.160000 ;
      LAYER met4 ;
        RECT 16.390000 39.840000 16.710000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 51.655000 17.075000 51.975000 ;
      LAYER met4 ;
        RECT 16.755000 51.655000 17.075000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 52.075000 17.075000 52.395000 ;
      LAYER met4 ;
        RECT 16.755000 52.075000 17.075000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755000 52.495000 17.075000 52.815000 ;
      LAYER met4 ;
        RECT 16.755000 52.495000 17.075000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 47.740000 17.080000 48.060000 ;
      LAYER met4 ;
        RECT 16.760000 47.740000 17.080000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760000 56.410000 17.080000 56.730000 ;
      LAYER met4 ;
        RECT 16.760000 56.410000 17.080000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795000 36.760000 17.115000 37.080000 ;
      LAYER met4 ;
        RECT 16.795000 36.760000 17.115000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795000 37.200000 17.115000 37.520000 ;
      LAYER met4 ;
        RECT 16.795000 37.200000 17.115000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795000 37.640000 17.115000 37.960000 ;
      LAYER met4 ;
        RECT 16.795000 37.640000 17.115000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795000 38.080000 17.115000 38.400000 ;
      LAYER met4 ;
        RECT 16.795000 38.080000 17.115000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795000 38.520000 17.115000 38.840000 ;
      LAYER met4 ;
        RECT 16.795000 38.520000 17.115000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795000 38.960000 17.115000 39.280000 ;
      LAYER met4 ;
        RECT 16.795000 38.960000 17.115000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795000 39.400000 17.115000 39.720000 ;
      LAYER met4 ;
        RECT 16.795000 39.400000 17.115000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795000 39.840000 17.115000 40.160000 ;
      LAYER met4 ;
        RECT 16.795000 39.840000 17.115000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 51.655000 17.480000 51.975000 ;
      LAYER met4 ;
        RECT 17.160000 51.655000 17.480000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 52.075000 17.480000 52.395000 ;
      LAYER met4 ;
        RECT 17.160000 52.075000 17.480000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160000 52.495000 17.480000 52.815000 ;
      LAYER met4 ;
        RECT 17.160000 52.495000 17.480000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 47.740000 17.485000 48.060000 ;
      LAYER met4 ;
        RECT 17.165000 47.740000 17.485000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165000 56.410000 17.485000 56.730000 ;
      LAYER met4 ;
        RECT 17.165000 56.410000 17.485000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200000 36.760000 17.520000 37.080000 ;
      LAYER met4 ;
        RECT 17.200000 36.760000 17.520000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200000 37.200000 17.520000 37.520000 ;
      LAYER met4 ;
        RECT 17.200000 37.200000 17.520000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200000 37.640000 17.520000 37.960000 ;
      LAYER met4 ;
        RECT 17.200000 37.640000 17.520000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200000 38.080000 17.520000 38.400000 ;
      LAYER met4 ;
        RECT 17.200000 38.080000 17.520000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200000 38.520000 17.520000 38.840000 ;
      LAYER met4 ;
        RECT 17.200000 38.520000 17.520000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200000 38.960000 17.520000 39.280000 ;
      LAYER met4 ;
        RECT 17.200000 38.960000 17.520000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200000 39.400000 17.520000 39.720000 ;
      LAYER met4 ;
        RECT 17.200000 39.400000 17.520000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200000 39.840000 17.520000 40.160000 ;
      LAYER met4 ;
        RECT 17.200000 39.840000 17.520000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 51.655000 17.885000 51.975000 ;
      LAYER met4 ;
        RECT 17.565000 51.655000 17.885000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 52.075000 17.885000 52.395000 ;
      LAYER met4 ;
        RECT 17.565000 52.075000 17.885000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565000 52.495000 17.885000 52.815000 ;
      LAYER met4 ;
        RECT 17.565000 52.495000 17.885000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 47.740000 17.890000 48.060000 ;
      LAYER met4 ;
        RECT 17.570000 47.740000 17.890000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570000 56.410000 17.890000 56.730000 ;
      LAYER met4 ;
        RECT 17.570000 56.410000 17.890000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605000 36.760000 17.925000 37.080000 ;
      LAYER met4 ;
        RECT 17.605000 36.760000 17.925000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605000 37.200000 17.925000 37.520000 ;
      LAYER met4 ;
        RECT 17.605000 37.200000 17.925000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605000 37.640000 17.925000 37.960000 ;
      LAYER met4 ;
        RECT 17.605000 37.640000 17.925000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605000 38.080000 17.925000 38.400000 ;
      LAYER met4 ;
        RECT 17.605000 38.080000 17.925000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605000 38.520000 17.925000 38.840000 ;
      LAYER met4 ;
        RECT 17.605000 38.520000 17.925000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605000 38.960000 17.925000 39.280000 ;
      LAYER met4 ;
        RECT 17.605000 38.960000 17.925000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605000 39.400000 17.925000 39.720000 ;
      LAYER met4 ;
        RECT 17.605000 39.400000 17.925000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605000 39.840000 17.925000 40.160000 ;
      LAYER met4 ;
        RECT 17.605000 39.840000 17.925000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 51.655000 18.290000 51.975000 ;
      LAYER met4 ;
        RECT 17.970000 51.655000 18.290000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 52.075000 18.290000 52.395000 ;
      LAYER met4 ;
        RECT 17.970000 52.075000 18.290000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970000 52.495000 18.290000 52.815000 ;
      LAYER met4 ;
        RECT 17.970000 52.495000 18.290000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 47.740000 18.295000 48.060000 ;
      LAYER met4 ;
        RECT 17.975000 47.740000 18.295000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975000 56.410000 18.295000 56.730000 ;
      LAYER met4 ;
        RECT 17.975000 56.410000 18.295000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010000 36.760000 18.330000 37.080000 ;
      LAYER met4 ;
        RECT 18.010000 36.760000 18.330000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010000 37.200000 18.330000 37.520000 ;
      LAYER met4 ;
        RECT 18.010000 37.200000 18.330000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010000 37.640000 18.330000 37.960000 ;
      LAYER met4 ;
        RECT 18.010000 37.640000 18.330000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010000 38.080000 18.330000 38.400000 ;
      LAYER met4 ;
        RECT 18.010000 38.080000 18.330000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010000 38.520000 18.330000 38.840000 ;
      LAYER met4 ;
        RECT 18.010000 38.520000 18.330000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010000 38.960000 18.330000 39.280000 ;
      LAYER met4 ;
        RECT 18.010000 38.960000 18.330000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010000 39.400000 18.330000 39.720000 ;
      LAYER met4 ;
        RECT 18.010000 39.400000 18.330000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010000 39.840000 18.330000 40.160000 ;
      LAYER met4 ;
        RECT 18.010000 39.840000 18.330000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 51.655000 18.695000 51.975000 ;
      LAYER met4 ;
        RECT 18.375000 51.655000 18.695000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 52.075000 18.695000 52.395000 ;
      LAYER met4 ;
        RECT 18.375000 52.075000 18.695000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375000 52.495000 18.695000 52.815000 ;
      LAYER met4 ;
        RECT 18.375000 52.495000 18.695000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 47.740000 18.700000 48.060000 ;
      LAYER met4 ;
        RECT 18.380000 47.740000 18.700000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380000 56.410000 18.700000 56.730000 ;
      LAYER met4 ;
        RECT 18.380000 56.410000 18.700000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415000 36.760000 18.735000 37.080000 ;
      LAYER met4 ;
        RECT 18.415000 36.760000 18.735000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415000 37.200000 18.735000 37.520000 ;
      LAYER met4 ;
        RECT 18.415000 37.200000 18.735000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415000 37.640000 18.735000 37.960000 ;
      LAYER met4 ;
        RECT 18.415000 37.640000 18.735000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415000 38.080000 18.735000 38.400000 ;
      LAYER met4 ;
        RECT 18.415000 38.080000 18.735000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415000 38.520000 18.735000 38.840000 ;
      LAYER met4 ;
        RECT 18.415000 38.520000 18.735000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415000 38.960000 18.735000 39.280000 ;
      LAYER met4 ;
        RECT 18.415000 38.960000 18.735000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415000 39.400000 18.735000 39.720000 ;
      LAYER met4 ;
        RECT 18.415000 39.400000 18.735000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415000 39.840000 18.735000 40.160000 ;
      LAYER met4 ;
        RECT 18.415000 39.840000 18.735000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 51.655000 19.100000 51.975000 ;
      LAYER met4 ;
        RECT 18.780000 51.655000 19.100000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 52.075000 19.100000 52.395000 ;
      LAYER met4 ;
        RECT 18.780000 52.075000 19.100000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780000 52.495000 19.100000 52.815000 ;
      LAYER met4 ;
        RECT 18.780000 52.495000 19.100000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 47.740000 19.105000 48.060000 ;
      LAYER met4 ;
        RECT 18.785000 47.740000 19.105000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785000 56.410000 19.105000 56.730000 ;
      LAYER met4 ;
        RECT 18.785000 56.410000 19.105000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820000 36.760000 19.140000 37.080000 ;
      LAYER met4 ;
        RECT 18.820000 36.760000 19.140000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820000 37.200000 19.140000 37.520000 ;
      LAYER met4 ;
        RECT 18.820000 37.200000 19.140000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820000 37.640000 19.140000 37.960000 ;
      LAYER met4 ;
        RECT 18.820000 37.640000 19.140000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820000 38.080000 19.140000 38.400000 ;
      LAYER met4 ;
        RECT 18.820000 38.080000 19.140000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820000 38.520000 19.140000 38.840000 ;
      LAYER met4 ;
        RECT 18.820000 38.520000 19.140000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820000 38.960000 19.140000 39.280000 ;
      LAYER met4 ;
        RECT 18.820000 38.960000 19.140000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820000 39.400000 19.140000 39.720000 ;
      LAYER met4 ;
        RECT 18.820000 39.400000 19.140000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820000 39.840000 19.140000 40.160000 ;
      LAYER met4 ;
        RECT 18.820000 39.840000 19.140000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 51.655000 19.505000 51.975000 ;
      LAYER met4 ;
        RECT 19.185000 51.655000 19.505000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 52.075000 19.505000 52.395000 ;
      LAYER met4 ;
        RECT 19.185000 52.075000 19.505000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185000 52.495000 19.505000 52.815000 ;
      LAYER met4 ;
        RECT 19.185000 52.495000 19.505000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 47.740000 19.510000 48.060000 ;
      LAYER met4 ;
        RECT 19.190000 47.740000 19.510000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190000 56.410000 19.510000 56.730000 ;
      LAYER met4 ;
        RECT 19.190000 56.410000 19.510000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225000 36.760000 19.545000 37.080000 ;
      LAYER met4 ;
        RECT 19.225000 36.760000 19.545000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225000 37.200000 19.545000 37.520000 ;
      LAYER met4 ;
        RECT 19.225000 37.200000 19.545000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225000 37.640000 19.545000 37.960000 ;
      LAYER met4 ;
        RECT 19.225000 37.640000 19.545000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225000 38.080000 19.545000 38.400000 ;
      LAYER met4 ;
        RECT 19.225000 38.080000 19.545000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225000 38.520000 19.545000 38.840000 ;
      LAYER met4 ;
        RECT 19.225000 38.520000 19.545000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225000 38.960000 19.545000 39.280000 ;
      LAYER met4 ;
        RECT 19.225000 38.960000 19.545000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225000 39.400000 19.545000 39.720000 ;
      LAYER met4 ;
        RECT 19.225000 39.400000 19.545000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225000 39.840000 19.545000 40.160000 ;
      LAYER met4 ;
        RECT 19.225000 39.840000 19.545000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 51.655000 19.910000 51.975000 ;
      LAYER met4 ;
        RECT 19.590000 51.655000 19.910000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 52.075000 19.910000 52.395000 ;
      LAYER met4 ;
        RECT 19.590000 52.075000 19.910000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590000 52.495000 19.910000 52.815000 ;
      LAYER met4 ;
        RECT 19.590000 52.495000 19.910000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 47.740000 19.915000 48.060000 ;
      LAYER met4 ;
        RECT 19.595000 47.740000 19.915000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595000 56.410000 19.915000 56.730000 ;
      LAYER met4 ;
        RECT 19.595000 56.410000 19.915000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630000 36.760000 19.950000 37.080000 ;
      LAYER met4 ;
        RECT 19.630000 36.760000 19.950000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630000 37.200000 19.950000 37.520000 ;
      LAYER met4 ;
        RECT 19.630000 37.200000 19.950000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630000 37.640000 19.950000 37.960000 ;
      LAYER met4 ;
        RECT 19.630000 37.640000 19.950000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630000 38.080000 19.950000 38.400000 ;
      LAYER met4 ;
        RECT 19.630000 38.080000 19.950000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630000 38.520000 19.950000 38.840000 ;
      LAYER met4 ;
        RECT 19.630000 38.520000 19.950000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630000 38.960000 19.950000 39.280000 ;
      LAYER met4 ;
        RECT 19.630000 38.960000 19.950000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630000 39.400000 19.950000 39.720000 ;
      LAYER met4 ;
        RECT 19.630000 39.400000 19.950000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630000 39.840000 19.950000 40.160000 ;
      LAYER met4 ;
        RECT 19.630000 39.840000 19.950000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 51.655000 20.315000 51.975000 ;
      LAYER met4 ;
        RECT 19.995000 51.655000 20.315000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 52.075000 20.315000 52.395000 ;
      LAYER met4 ;
        RECT 19.995000 52.075000 20.315000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995000 52.495000 20.315000 52.815000 ;
      LAYER met4 ;
        RECT 19.995000 52.495000 20.315000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 51.655000 2.485000 51.975000 ;
      LAYER met4 ;
        RECT 2.165000 51.655000 2.485000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 52.075000 2.485000 52.395000 ;
      LAYER met4 ;
        RECT 2.165000 52.075000 2.485000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165000 52.495000 2.485000 52.815000 ;
      LAYER met4 ;
        RECT 2.165000 52.495000 2.485000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.180000 47.740000 2.500000 48.060000 ;
      LAYER met4 ;
        RECT 2.180000 47.740000 2.500000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.180000 56.410000 2.500000 56.730000 ;
      LAYER met4 ;
        RECT 2.180000 56.410000 2.500000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 36.760000 2.535000 37.080000 ;
      LAYER met4 ;
        RECT 2.215000 36.760000 2.535000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 37.200000 2.535000 37.520000 ;
      LAYER met4 ;
        RECT 2.215000 37.200000 2.535000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 37.640000 2.535000 37.960000 ;
      LAYER met4 ;
        RECT 2.215000 37.640000 2.535000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 38.080000 2.535000 38.400000 ;
      LAYER met4 ;
        RECT 2.215000 38.080000 2.535000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 38.520000 2.535000 38.840000 ;
      LAYER met4 ;
        RECT 2.215000 38.520000 2.535000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 38.960000 2.535000 39.280000 ;
      LAYER met4 ;
        RECT 2.215000 38.960000 2.535000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 39.400000 2.535000 39.720000 ;
      LAYER met4 ;
        RECT 2.215000 39.400000 2.535000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215000 39.840000 2.535000 40.160000 ;
      LAYER met4 ;
        RECT 2.215000 39.840000 2.535000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 51.655000 2.895000 51.975000 ;
      LAYER met4 ;
        RECT 2.575000 51.655000 2.895000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 52.075000 2.895000 52.395000 ;
      LAYER met4 ;
        RECT 2.575000 52.075000 2.895000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575000 52.495000 2.895000 52.815000 ;
      LAYER met4 ;
        RECT 2.575000 52.495000 2.895000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.585000 47.740000 2.905000 48.060000 ;
      LAYER met4 ;
        RECT 2.585000 47.740000 2.905000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.585000 56.410000 2.905000 56.730000 ;
      LAYER met4 ;
        RECT 2.585000 56.410000 2.905000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620000 36.760000 2.940000 37.080000 ;
      LAYER met4 ;
        RECT 2.620000 36.760000 2.940000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620000 37.200000 2.940000 37.520000 ;
      LAYER met4 ;
        RECT 2.620000 37.200000 2.940000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620000 37.640000 2.940000 37.960000 ;
      LAYER met4 ;
        RECT 2.620000 37.640000 2.940000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620000 38.080000 2.940000 38.400000 ;
      LAYER met4 ;
        RECT 2.620000 38.080000 2.940000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620000 38.520000 2.940000 38.840000 ;
      LAYER met4 ;
        RECT 2.620000 38.520000 2.940000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620000 38.960000 2.940000 39.280000 ;
      LAYER met4 ;
        RECT 2.620000 38.960000 2.940000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620000 39.400000 2.940000 39.720000 ;
      LAYER met4 ;
        RECT 2.620000 39.400000 2.940000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620000 39.840000 2.940000 40.160000 ;
      LAYER met4 ;
        RECT 2.620000 39.840000 2.940000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 51.655000 3.305000 51.975000 ;
      LAYER met4 ;
        RECT 2.985000 51.655000 3.305000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 52.075000 3.305000 52.395000 ;
      LAYER met4 ;
        RECT 2.985000 52.075000 3.305000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985000 52.495000 3.305000 52.815000 ;
      LAYER met4 ;
        RECT 2.985000 52.495000 3.305000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 47.740000 3.310000 48.060000 ;
      LAYER met4 ;
        RECT 2.990000 47.740000 3.310000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990000 56.410000 3.310000 56.730000 ;
      LAYER met4 ;
        RECT 2.990000 56.410000 3.310000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 47.740000 20.320000 48.060000 ;
      LAYER met4 ;
        RECT 20.000000 47.740000 20.320000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000000 56.410000 20.320000 56.730000 ;
      LAYER met4 ;
        RECT 20.000000 56.410000 20.320000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035000 36.760000 20.355000 37.080000 ;
      LAYER met4 ;
        RECT 20.035000 36.760000 20.355000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035000 37.200000 20.355000 37.520000 ;
      LAYER met4 ;
        RECT 20.035000 37.200000 20.355000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035000 37.640000 20.355000 37.960000 ;
      LAYER met4 ;
        RECT 20.035000 37.640000 20.355000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035000 38.080000 20.355000 38.400000 ;
      LAYER met4 ;
        RECT 20.035000 38.080000 20.355000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035000 38.520000 20.355000 38.840000 ;
      LAYER met4 ;
        RECT 20.035000 38.520000 20.355000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035000 38.960000 20.355000 39.280000 ;
      LAYER met4 ;
        RECT 20.035000 38.960000 20.355000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035000 39.400000 20.355000 39.720000 ;
      LAYER met4 ;
        RECT 20.035000 39.400000 20.355000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035000 39.840000 20.355000 40.160000 ;
      LAYER met4 ;
        RECT 20.035000 39.840000 20.355000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 51.655000 20.720000 51.975000 ;
      LAYER met4 ;
        RECT 20.400000 51.655000 20.720000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 52.075000 20.720000 52.395000 ;
      LAYER met4 ;
        RECT 20.400000 52.075000 20.720000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400000 52.495000 20.720000 52.815000 ;
      LAYER met4 ;
        RECT 20.400000 52.495000 20.720000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 47.740000 20.725000 48.060000 ;
      LAYER met4 ;
        RECT 20.405000 47.740000 20.725000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405000 56.410000 20.725000 56.730000 ;
      LAYER met4 ;
        RECT 20.405000 56.410000 20.725000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440000 36.760000 20.760000 37.080000 ;
      LAYER met4 ;
        RECT 20.440000 36.760000 20.760000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440000 37.200000 20.760000 37.520000 ;
      LAYER met4 ;
        RECT 20.440000 37.200000 20.760000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440000 37.640000 20.760000 37.960000 ;
      LAYER met4 ;
        RECT 20.440000 37.640000 20.760000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440000 38.080000 20.760000 38.400000 ;
      LAYER met4 ;
        RECT 20.440000 38.080000 20.760000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440000 38.520000 20.760000 38.840000 ;
      LAYER met4 ;
        RECT 20.440000 38.520000 20.760000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440000 38.960000 20.760000 39.280000 ;
      LAYER met4 ;
        RECT 20.440000 38.960000 20.760000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440000 39.400000 20.760000 39.720000 ;
      LAYER met4 ;
        RECT 20.440000 39.400000 20.760000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440000 39.840000 20.760000 40.160000 ;
      LAYER met4 ;
        RECT 20.440000 39.840000 20.760000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 51.655000 21.125000 51.975000 ;
      LAYER met4 ;
        RECT 20.805000 51.655000 21.125000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 52.075000 21.125000 52.395000 ;
      LAYER met4 ;
        RECT 20.805000 52.075000 21.125000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805000 52.495000 21.125000 52.815000 ;
      LAYER met4 ;
        RECT 20.805000 52.495000 21.125000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 47.740000 21.130000 48.060000 ;
      LAYER met4 ;
        RECT 20.810000 47.740000 21.130000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810000 56.410000 21.130000 56.730000 ;
      LAYER met4 ;
        RECT 20.810000 56.410000 21.130000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845000 36.760000 21.165000 37.080000 ;
      LAYER met4 ;
        RECT 20.845000 36.760000 21.165000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845000 37.200000 21.165000 37.520000 ;
      LAYER met4 ;
        RECT 20.845000 37.200000 21.165000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845000 37.640000 21.165000 37.960000 ;
      LAYER met4 ;
        RECT 20.845000 37.640000 21.165000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845000 38.080000 21.165000 38.400000 ;
      LAYER met4 ;
        RECT 20.845000 38.080000 21.165000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845000 38.520000 21.165000 38.840000 ;
      LAYER met4 ;
        RECT 20.845000 38.520000 21.165000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845000 38.960000 21.165000 39.280000 ;
      LAYER met4 ;
        RECT 20.845000 38.960000 21.165000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845000 39.400000 21.165000 39.720000 ;
      LAYER met4 ;
        RECT 20.845000 39.400000 21.165000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845000 39.840000 21.165000 40.160000 ;
      LAYER met4 ;
        RECT 20.845000 39.840000 21.165000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 51.655000 21.530000 51.975000 ;
      LAYER met4 ;
        RECT 21.210000 51.655000 21.530000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 52.075000 21.530000 52.395000 ;
      LAYER met4 ;
        RECT 21.210000 52.075000 21.530000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210000 52.495000 21.530000 52.815000 ;
      LAYER met4 ;
        RECT 21.210000 52.495000 21.530000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 47.740000 21.535000 48.060000 ;
      LAYER met4 ;
        RECT 21.215000 47.740000 21.535000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215000 56.410000 21.535000 56.730000 ;
      LAYER met4 ;
        RECT 21.215000 56.410000 21.535000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245000 36.760000 21.565000 37.080000 ;
      LAYER met4 ;
        RECT 21.245000 36.760000 21.565000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245000 37.200000 21.565000 37.520000 ;
      LAYER met4 ;
        RECT 21.245000 37.200000 21.565000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245000 37.640000 21.565000 37.960000 ;
      LAYER met4 ;
        RECT 21.245000 37.640000 21.565000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245000 38.080000 21.565000 38.400000 ;
      LAYER met4 ;
        RECT 21.245000 38.080000 21.565000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245000 38.520000 21.565000 38.840000 ;
      LAYER met4 ;
        RECT 21.245000 38.520000 21.565000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245000 38.960000 21.565000 39.280000 ;
      LAYER met4 ;
        RECT 21.245000 38.960000 21.565000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245000 39.400000 21.565000 39.720000 ;
      LAYER met4 ;
        RECT 21.245000 39.400000 21.565000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245000 39.840000 21.565000 40.160000 ;
      LAYER met4 ;
        RECT 21.245000 39.840000 21.565000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 51.655000 21.935000 51.975000 ;
      LAYER met4 ;
        RECT 21.615000 51.655000 21.935000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 52.075000 21.935000 52.395000 ;
      LAYER met4 ;
        RECT 21.615000 52.075000 21.935000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615000 52.495000 21.935000 52.815000 ;
      LAYER met4 ;
        RECT 21.615000 52.495000 21.935000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 47.740000 21.940000 48.060000 ;
      LAYER met4 ;
        RECT 21.620000 47.740000 21.940000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620000 56.410000 21.940000 56.730000 ;
      LAYER met4 ;
        RECT 21.620000 56.410000 21.940000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645000 36.760000 21.965000 37.080000 ;
      LAYER met4 ;
        RECT 21.645000 36.760000 21.965000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645000 37.200000 21.965000 37.520000 ;
      LAYER met4 ;
        RECT 21.645000 37.200000 21.965000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645000 37.640000 21.965000 37.960000 ;
      LAYER met4 ;
        RECT 21.645000 37.640000 21.965000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645000 38.080000 21.965000 38.400000 ;
      LAYER met4 ;
        RECT 21.645000 38.080000 21.965000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645000 38.520000 21.965000 38.840000 ;
      LAYER met4 ;
        RECT 21.645000 38.520000 21.965000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645000 38.960000 21.965000 39.280000 ;
      LAYER met4 ;
        RECT 21.645000 38.960000 21.965000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645000 39.400000 21.965000 39.720000 ;
      LAYER met4 ;
        RECT 21.645000 39.400000 21.965000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645000 39.840000 21.965000 40.160000 ;
      LAYER met4 ;
        RECT 21.645000 39.840000 21.965000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 51.655000 22.340000 51.975000 ;
      LAYER met4 ;
        RECT 22.020000 51.655000 22.340000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 52.075000 22.340000 52.395000 ;
      LAYER met4 ;
        RECT 22.020000 52.075000 22.340000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020000 52.495000 22.340000 52.815000 ;
      LAYER met4 ;
        RECT 22.020000 52.495000 22.340000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 47.740000 22.345000 48.060000 ;
      LAYER met4 ;
        RECT 22.025000 47.740000 22.345000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025000 56.410000 22.345000 56.730000 ;
      LAYER met4 ;
        RECT 22.025000 56.410000 22.345000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045000 36.760000 22.365000 37.080000 ;
      LAYER met4 ;
        RECT 22.045000 36.760000 22.365000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045000 37.200000 22.365000 37.520000 ;
      LAYER met4 ;
        RECT 22.045000 37.200000 22.365000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045000 37.640000 22.365000 37.960000 ;
      LAYER met4 ;
        RECT 22.045000 37.640000 22.365000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045000 38.080000 22.365000 38.400000 ;
      LAYER met4 ;
        RECT 22.045000 38.080000 22.365000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045000 38.520000 22.365000 38.840000 ;
      LAYER met4 ;
        RECT 22.045000 38.520000 22.365000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045000 38.960000 22.365000 39.280000 ;
      LAYER met4 ;
        RECT 22.045000 38.960000 22.365000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045000 39.400000 22.365000 39.720000 ;
      LAYER met4 ;
        RECT 22.045000 39.400000 22.365000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045000 39.840000 22.365000 40.160000 ;
      LAYER met4 ;
        RECT 22.045000 39.840000 22.365000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 51.655000 22.745000 51.975000 ;
      LAYER met4 ;
        RECT 22.425000 51.655000 22.745000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 52.075000 22.745000 52.395000 ;
      LAYER met4 ;
        RECT 22.425000 52.075000 22.745000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425000 52.495000 22.745000 52.815000 ;
      LAYER met4 ;
        RECT 22.425000 52.495000 22.745000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 47.740000 22.750000 48.060000 ;
      LAYER met4 ;
        RECT 22.430000 47.740000 22.750000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430000 56.410000 22.750000 56.730000 ;
      LAYER met4 ;
        RECT 22.430000 56.410000 22.750000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445000 36.760000 22.765000 37.080000 ;
      LAYER met4 ;
        RECT 22.445000 36.760000 22.765000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445000 37.200000 22.765000 37.520000 ;
      LAYER met4 ;
        RECT 22.445000 37.200000 22.765000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445000 37.640000 22.765000 37.960000 ;
      LAYER met4 ;
        RECT 22.445000 37.640000 22.765000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445000 38.080000 22.765000 38.400000 ;
      LAYER met4 ;
        RECT 22.445000 38.080000 22.765000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445000 38.520000 22.765000 38.840000 ;
      LAYER met4 ;
        RECT 22.445000 38.520000 22.765000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445000 38.960000 22.765000 39.280000 ;
      LAYER met4 ;
        RECT 22.445000 38.960000 22.765000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445000 39.400000 22.765000 39.720000 ;
      LAYER met4 ;
        RECT 22.445000 39.400000 22.765000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445000 39.840000 22.765000 40.160000 ;
      LAYER met4 ;
        RECT 22.445000 39.840000 22.765000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 51.655000 23.150000 51.975000 ;
      LAYER met4 ;
        RECT 22.830000 51.655000 23.150000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 52.075000 23.150000 52.395000 ;
      LAYER met4 ;
        RECT 22.830000 52.075000 23.150000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830000 52.495000 23.150000 52.815000 ;
      LAYER met4 ;
        RECT 22.830000 52.495000 23.150000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 47.740000 23.155000 48.060000 ;
      LAYER met4 ;
        RECT 22.835000 47.740000 23.155000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835000 56.410000 23.155000 56.730000 ;
      LAYER met4 ;
        RECT 22.835000 56.410000 23.155000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845000 36.760000 23.165000 37.080000 ;
      LAYER met4 ;
        RECT 22.845000 36.760000 23.165000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845000 37.200000 23.165000 37.520000 ;
      LAYER met4 ;
        RECT 22.845000 37.200000 23.165000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845000 37.640000 23.165000 37.960000 ;
      LAYER met4 ;
        RECT 22.845000 37.640000 23.165000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845000 38.080000 23.165000 38.400000 ;
      LAYER met4 ;
        RECT 22.845000 38.080000 23.165000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845000 38.520000 23.165000 38.840000 ;
      LAYER met4 ;
        RECT 22.845000 38.520000 23.165000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845000 38.960000 23.165000 39.280000 ;
      LAYER met4 ;
        RECT 22.845000 38.960000 23.165000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845000 39.400000 23.165000 39.720000 ;
      LAYER met4 ;
        RECT 22.845000 39.400000 23.165000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845000 39.840000 23.165000 40.160000 ;
      LAYER met4 ;
        RECT 22.845000 39.840000 23.165000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 51.655000 23.555000 51.975000 ;
      LAYER met4 ;
        RECT 23.235000 51.655000 23.555000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 52.075000 23.555000 52.395000 ;
      LAYER met4 ;
        RECT 23.235000 52.075000 23.555000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235000 52.495000 23.555000 52.815000 ;
      LAYER met4 ;
        RECT 23.235000 52.495000 23.555000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 47.740000 23.560000 48.060000 ;
      LAYER met4 ;
        RECT 23.240000 47.740000 23.560000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240000 56.410000 23.560000 56.730000 ;
      LAYER met4 ;
        RECT 23.240000 56.410000 23.560000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245000 36.760000 23.565000 37.080000 ;
      LAYER met4 ;
        RECT 23.245000 36.760000 23.565000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245000 37.200000 23.565000 37.520000 ;
      LAYER met4 ;
        RECT 23.245000 37.200000 23.565000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245000 37.640000 23.565000 37.960000 ;
      LAYER met4 ;
        RECT 23.245000 37.640000 23.565000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245000 38.080000 23.565000 38.400000 ;
      LAYER met4 ;
        RECT 23.245000 38.080000 23.565000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245000 38.520000 23.565000 38.840000 ;
      LAYER met4 ;
        RECT 23.245000 38.520000 23.565000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245000 38.960000 23.565000 39.280000 ;
      LAYER met4 ;
        RECT 23.245000 38.960000 23.565000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245000 39.400000 23.565000 39.720000 ;
      LAYER met4 ;
        RECT 23.245000 39.400000 23.565000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245000 39.840000 23.565000 40.160000 ;
      LAYER met4 ;
        RECT 23.245000 39.840000 23.565000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 51.655000 23.960000 51.975000 ;
      LAYER met4 ;
        RECT 23.640000 51.655000 23.960000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 52.075000 23.960000 52.395000 ;
      LAYER met4 ;
        RECT 23.640000 52.075000 23.960000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640000 52.495000 23.960000 52.815000 ;
      LAYER met4 ;
        RECT 23.640000 52.495000 23.960000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 36.760000 23.965000 37.080000 ;
      LAYER met4 ;
        RECT 23.645000 36.760000 23.965000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 37.200000 23.965000 37.520000 ;
      LAYER met4 ;
        RECT 23.645000 37.200000 23.965000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 37.640000 23.965000 37.960000 ;
      LAYER met4 ;
        RECT 23.645000 37.640000 23.965000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 38.080000 23.965000 38.400000 ;
      LAYER met4 ;
        RECT 23.645000 38.080000 23.965000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 38.520000 23.965000 38.840000 ;
      LAYER met4 ;
        RECT 23.645000 38.520000 23.965000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 38.960000 23.965000 39.280000 ;
      LAYER met4 ;
        RECT 23.645000 38.960000 23.965000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 39.400000 23.965000 39.720000 ;
      LAYER met4 ;
        RECT 23.645000 39.400000 23.965000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 39.840000 23.965000 40.160000 ;
      LAYER met4 ;
        RECT 23.645000 39.840000 23.965000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 47.740000 23.965000 48.060000 ;
      LAYER met4 ;
        RECT 23.645000 47.740000 23.965000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645000 56.410000 23.965000 56.730000 ;
      LAYER met4 ;
        RECT 23.645000 56.410000 23.965000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 36.760000 24.365000 37.080000 ;
      LAYER met4 ;
        RECT 24.045000 36.760000 24.365000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 37.200000 24.365000 37.520000 ;
      LAYER met4 ;
        RECT 24.045000 37.200000 24.365000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 37.640000 24.365000 37.960000 ;
      LAYER met4 ;
        RECT 24.045000 37.640000 24.365000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 38.080000 24.365000 38.400000 ;
      LAYER met4 ;
        RECT 24.045000 38.080000 24.365000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 38.520000 24.365000 38.840000 ;
      LAYER met4 ;
        RECT 24.045000 38.520000 24.365000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 38.960000 24.365000 39.280000 ;
      LAYER met4 ;
        RECT 24.045000 38.960000 24.365000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 39.400000 24.365000 39.720000 ;
      LAYER met4 ;
        RECT 24.045000 39.400000 24.365000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 39.840000 24.365000 40.160000 ;
      LAYER met4 ;
        RECT 24.045000 39.840000 24.365000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 47.740000 24.365000 48.060000 ;
      LAYER met4 ;
        RECT 24.045000 47.740000 24.365000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 51.655000 24.365000 51.975000 ;
      LAYER met4 ;
        RECT 24.045000 51.655000 24.365000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 52.075000 24.365000 52.395000 ;
      LAYER met4 ;
        RECT 24.045000 52.075000 24.365000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 52.495000 24.365000 52.815000 ;
      LAYER met4 ;
        RECT 24.045000 52.495000 24.365000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045000 56.410000 24.365000 56.730000 ;
      LAYER met4 ;
        RECT 24.045000 56.410000 24.365000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 36.760000 3.345000 37.080000 ;
      LAYER met4 ;
        RECT 3.025000 36.760000 3.345000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 37.200000 3.345000 37.520000 ;
      LAYER met4 ;
        RECT 3.025000 37.200000 3.345000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 37.640000 3.345000 37.960000 ;
      LAYER met4 ;
        RECT 3.025000 37.640000 3.345000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 38.080000 3.345000 38.400000 ;
      LAYER met4 ;
        RECT 3.025000 38.080000 3.345000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 38.520000 3.345000 38.840000 ;
      LAYER met4 ;
        RECT 3.025000 38.520000 3.345000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 38.960000 3.345000 39.280000 ;
      LAYER met4 ;
        RECT 3.025000 38.960000 3.345000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 39.400000 3.345000 39.720000 ;
      LAYER met4 ;
        RECT 3.025000 39.400000 3.345000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025000 39.840000 3.345000 40.160000 ;
      LAYER met4 ;
        RECT 3.025000 39.840000 3.345000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 51.655000 3.710000 51.975000 ;
      LAYER met4 ;
        RECT 3.390000 51.655000 3.710000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 52.075000 3.710000 52.395000 ;
      LAYER met4 ;
        RECT 3.390000 52.075000 3.710000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390000 52.495000 3.710000 52.815000 ;
      LAYER met4 ;
        RECT 3.390000 52.495000 3.710000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 47.740000 3.715000 48.060000 ;
      LAYER met4 ;
        RECT 3.395000 47.740000 3.715000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395000 56.410000 3.715000 56.730000 ;
      LAYER met4 ;
        RECT 3.395000 56.410000 3.715000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430000 36.760000 3.750000 37.080000 ;
      LAYER met4 ;
        RECT 3.430000 36.760000 3.750000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430000 37.200000 3.750000 37.520000 ;
      LAYER met4 ;
        RECT 3.430000 37.200000 3.750000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430000 37.640000 3.750000 37.960000 ;
      LAYER met4 ;
        RECT 3.430000 37.640000 3.750000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430000 38.080000 3.750000 38.400000 ;
      LAYER met4 ;
        RECT 3.430000 38.080000 3.750000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430000 38.520000 3.750000 38.840000 ;
      LAYER met4 ;
        RECT 3.430000 38.520000 3.750000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430000 38.960000 3.750000 39.280000 ;
      LAYER met4 ;
        RECT 3.430000 38.960000 3.750000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430000 39.400000 3.750000 39.720000 ;
      LAYER met4 ;
        RECT 3.430000 39.400000 3.750000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430000 39.840000 3.750000 40.160000 ;
      LAYER met4 ;
        RECT 3.430000 39.840000 3.750000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 51.655000 4.115000 51.975000 ;
      LAYER met4 ;
        RECT 3.795000 51.655000 4.115000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 52.075000 4.115000 52.395000 ;
      LAYER met4 ;
        RECT 3.795000 52.075000 4.115000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795000 52.495000 4.115000 52.815000 ;
      LAYER met4 ;
        RECT 3.795000 52.495000 4.115000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 47.740000 4.120000 48.060000 ;
      LAYER met4 ;
        RECT 3.800000 47.740000 4.120000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800000 56.410000 4.120000 56.730000 ;
      LAYER met4 ;
        RECT 3.800000 56.410000 4.120000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835000 36.760000 4.155000 37.080000 ;
      LAYER met4 ;
        RECT 3.835000 36.760000 4.155000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835000 37.200000 4.155000 37.520000 ;
      LAYER met4 ;
        RECT 3.835000 37.200000 4.155000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835000 37.640000 4.155000 37.960000 ;
      LAYER met4 ;
        RECT 3.835000 37.640000 4.155000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835000 38.080000 4.155000 38.400000 ;
      LAYER met4 ;
        RECT 3.835000 38.080000 4.155000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835000 38.520000 4.155000 38.840000 ;
      LAYER met4 ;
        RECT 3.835000 38.520000 4.155000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835000 38.960000 4.155000 39.280000 ;
      LAYER met4 ;
        RECT 3.835000 38.960000 4.155000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835000 39.400000 4.155000 39.720000 ;
      LAYER met4 ;
        RECT 3.835000 39.400000 4.155000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835000 39.840000 4.155000 40.160000 ;
      LAYER met4 ;
        RECT 3.835000 39.840000 4.155000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 51.655000 4.520000 51.975000 ;
      LAYER met4 ;
        RECT 4.200000 51.655000 4.520000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 52.075000 4.520000 52.395000 ;
      LAYER met4 ;
        RECT 4.200000 52.075000 4.520000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200000 52.495000 4.520000 52.815000 ;
      LAYER met4 ;
        RECT 4.200000 52.495000 4.520000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 47.740000 4.525000 48.060000 ;
      LAYER met4 ;
        RECT 4.205000 47.740000 4.525000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205000 56.410000 4.525000 56.730000 ;
      LAYER met4 ;
        RECT 4.205000 56.410000 4.525000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240000 36.760000 4.560000 37.080000 ;
      LAYER met4 ;
        RECT 4.240000 36.760000 4.560000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240000 37.200000 4.560000 37.520000 ;
      LAYER met4 ;
        RECT 4.240000 37.200000 4.560000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240000 37.640000 4.560000 37.960000 ;
      LAYER met4 ;
        RECT 4.240000 37.640000 4.560000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240000 38.080000 4.560000 38.400000 ;
      LAYER met4 ;
        RECT 4.240000 38.080000 4.560000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240000 38.520000 4.560000 38.840000 ;
      LAYER met4 ;
        RECT 4.240000 38.520000 4.560000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240000 38.960000 4.560000 39.280000 ;
      LAYER met4 ;
        RECT 4.240000 38.960000 4.560000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240000 39.400000 4.560000 39.720000 ;
      LAYER met4 ;
        RECT 4.240000 39.400000 4.560000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240000 39.840000 4.560000 40.160000 ;
      LAYER met4 ;
        RECT 4.240000 39.840000 4.560000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 51.655000 4.925000 51.975000 ;
      LAYER met4 ;
        RECT 4.605000 51.655000 4.925000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 52.075000 4.925000 52.395000 ;
      LAYER met4 ;
        RECT 4.605000 52.075000 4.925000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605000 52.495000 4.925000 52.815000 ;
      LAYER met4 ;
        RECT 4.605000 52.495000 4.925000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 47.740000 4.930000 48.060000 ;
      LAYER met4 ;
        RECT 4.610000 47.740000 4.930000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610000 56.410000 4.930000 56.730000 ;
      LAYER met4 ;
        RECT 4.610000 56.410000 4.930000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645000 36.760000 4.965000 37.080000 ;
      LAYER met4 ;
        RECT 4.645000 36.760000 4.965000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645000 37.200000 4.965000 37.520000 ;
      LAYER met4 ;
        RECT 4.645000 37.200000 4.965000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645000 37.640000 4.965000 37.960000 ;
      LAYER met4 ;
        RECT 4.645000 37.640000 4.965000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645000 38.080000 4.965000 38.400000 ;
      LAYER met4 ;
        RECT 4.645000 38.080000 4.965000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645000 38.520000 4.965000 38.840000 ;
      LAYER met4 ;
        RECT 4.645000 38.520000 4.965000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645000 38.960000 4.965000 39.280000 ;
      LAYER met4 ;
        RECT 4.645000 38.960000 4.965000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645000 39.400000 4.965000 39.720000 ;
      LAYER met4 ;
        RECT 4.645000 39.400000 4.965000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645000 39.840000 4.965000 40.160000 ;
      LAYER met4 ;
        RECT 4.645000 39.840000 4.965000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 51.655000 5.330000 51.975000 ;
      LAYER met4 ;
        RECT 5.010000 51.655000 5.330000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 52.075000 5.330000 52.395000 ;
      LAYER met4 ;
        RECT 5.010000 52.075000 5.330000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010000 52.495000 5.330000 52.815000 ;
      LAYER met4 ;
        RECT 5.010000 52.495000 5.330000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 47.740000 5.335000 48.060000 ;
      LAYER met4 ;
        RECT 5.015000 47.740000 5.335000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015000 56.410000 5.335000 56.730000 ;
      LAYER met4 ;
        RECT 5.015000 56.410000 5.335000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050000 36.760000 5.370000 37.080000 ;
      LAYER met4 ;
        RECT 5.050000 36.760000 5.370000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050000 37.200000 5.370000 37.520000 ;
      LAYER met4 ;
        RECT 5.050000 37.200000 5.370000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050000 37.640000 5.370000 37.960000 ;
      LAYER met4 ;
        RECT 5.050000 37.640000 5.370000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050000 38.080000 5.370000 38.400000 ;
      LAYER met4 ;
        RECT 5.050000 38.080000 5.370000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050000 38.520000 5.370000 38.840000 ;
      LAYER met4 ;
        RECT 5.050000 38.520000 5.370000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050000 38.960000 5.370000 39.280000 ;
      LAYER met4 ;
        RECT 5.050000 38.960000 5.370000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050000 39.400000 5.370000 39.720000 ;
      LAYER met4 ;
        RECT 5.050000 39.400000 5.370000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050000 39.840000 5.370000 40.160000 ;
      LAYER met4 ;
        RECT 5.050000 39.840000 5.370000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 51.655000 5.735000 51.975000 ;
      LAYER met4 ;
        RECT 5.415000 51.655000 5.735000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 52.075000 5.735000 52.395000 ;
      LAYER met4 ;
        RECT 5.415000 52.075000 5.735000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415000 52.495000 5.735000 52.815000 ;
      LAYER met4 ;
        RECT 5.415000 52.495000 5.735000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 47.740000 5.740000 48.060000 ;
      LAYER met4 ;
        RECT 5.420000 47.740000 5.740000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420000 56.410000 5.740000 56.730000 ;
      LAYER met4 ;
        RECT 5.420000 56.410000 5.740000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455000 36.760000 5.775000 37.080000 ;
      LAYER met4 ;
        RECT 5.455000 36.760000 5.775000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455000 37.200000 5.775000 37.520000 ;
      LAYER met4 ;
        RECT 5.455000 37.200000 5.775000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455000 37.640000 5.775000 37.960000 ;
      LAYER met4 ;
        RECT 5.455000 37.640000 5.775000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455000 38.080000 5.775000 38.400000 ;
      LAYER met4 ;
        RECT 5.455000 38.080000 5.775000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455000 38.520000 5.775000 38.840000 ;
      LAYER met4 ;
        RECT 5.455000 38.520000 5.775000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455000 38.960000 5.775000 39.280000 ;
      LAYER met4 ;
        RECT 5.455000 38.960000 5.775000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455000 39.400000 5.775000 39.720000 ;
      LAYER met4 ;
        RECT 5.455000 39.400000 5.775000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455000 39.840000 5.775000 40.160000 ;
      LAYER met4 ;
        RECT 5.455000 39.840000 5.775000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 51.655000 6.140000 51.975000 ;
      LAYER met4 ;
        RECT 5.820000 51.655000 6.140000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 52.075000 6.140000 52.395000 ;
      LAYER met4 ;
        RECT 5.820000 52.075000 6.140000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820000 52.495000 6.140000 52.815000 ;
      LAYER met4 ;
        RECT 5.820000 52.495000 6.140000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 47.740000 6.145000 48.060000 ;
      LAYER met4 ;
        RECT 5.825000 47.740000 6.145000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825000 56.410000 6.145000 56.730000 ;
      LAYER met4 ;
        RECT 5.825000 56.410000 6.145000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860000 36.760000 6.180000 37.080000 ;
      LAYER met4 ;
        RECT 5.860000 36.760000 6.180000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860000 37.200000 6.180000 37.520000 ;
      LAYER met4 ;
        RECT 5.860000 37.200000 6.180000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860000 37.640000 6.180000 37.960000 ;
      LAYER met4 ;
        RECT 5.860000 37.640000 6.180000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860000 38.080000 6.180000 38.400000 ;
      LAYER met4 ;
        RECT 5.860000 38.080000 6.180000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860000 38.520000 6.180000 38.840000 ;
      LAYER met4 ;
        RECT 5.860000 38.520000 6.180000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860000 38.960000 6.180000 39.280000 ;
      LAYER met4 ;
        RECT 5.860000 38.960000 6.180000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860000 39.400000 6.180000 39.720000 ;
      LAYER met4 ;
        RECT 5.860000 39.400000 6.180000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860000 39.840000 6.180000 40.160000 ;
      LAYER met4 ;
        RECT 5.860000 39.840000 6.180000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 36.760000 50.740000 37.080000 ;
      LAYER met4 ;
        RECT 50.420000 36.760000 50.740000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 37.200000 50.740000 37.520000 ;
      LAYER met4 ;
        RECT 50.420000 37.200000 50.740000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 37.640000 50.740000 37.960000 ;
      LAYER met4 ;
        RECT 50.420000 37.640000 50.740000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 38.080000 50.740000 38.400000 ;
      LAYER met4 ;
        RECT 50.420000 38.080000 50.740000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 38.520000 50.740000 38.840000 ;
      LAYER met4 ;
        RECT 50.420000 38.520000 50.740000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 38.960000 50.740000 39.280000 ;
      LAYER met4 ;
        RECT 50.420000 38.960000 50.740000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 39.400000 50.740000 39.720000 ;
      LAYER met4 ;
        RECT 50.420000 39.400000 50.740000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 39.840000 50.740000 40.160000 ;
      LAYER met4 ;
        RECT 50.420000 39.840000 50.740000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 47.740000 50.740000 48.060000 ;
      LAYER met4 ;
        RECT 50.420000 47.740000 50.740000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 51.655000 50.740000 51.975000 ;
      LAYER met4 ;
        RECT 50.420000 51.655000 50.740000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 52.075000 50.740000 52.395000 ;
      LAYER met4 ;
        RECT 50.420000 52.075000 50.740000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 52.495000 50.740000 52.815000 ;
      LAYER met4 ;
        RECT 50.420000 52.495000 50.740000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420000 56.410000 50.740000 56.730000 ;
      LAYER met4 ;
        RECT 50.420000 56.410000 50.740000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.825000 47.740000 51.145000 48.060000 ;
      LAYER met4 ;
        RECT 50.825000 47.740000 51.145000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.825000 56.410000 51.145000 56.730000 ;
      LAYER met4 ;
        RECT 50.825000 56.410000 51.145000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 36.760000 51.150000 37.080000 ;
      LAYER met4 ;
        RECT 50.830000 36.760000 51.150000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 37.200000 51.150000 37.520000 ;
      LAYER met4 ;
        RECT 50.830000 37.200000 51.150000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 37.640000 51.150000 37.960000 ;
      LAYER met4 ;
        RECT 50.830000 37.640000 51.150000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 38.080000 51.150000 38.400000 ;
      LAYER met4 ;
        RECT 50.830000 38.080000 51.150000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 38.520000 51.150000 38.840000 ;
      LAYER met4 ;
        RECT 50.830000 38.520000 51.150000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 38.960000 51.150000 39.280000 ;
      LAYER met4 ;
        RECT 50.830000 38.960000 51.150000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 39.400000 51.150000 39.720000 ;
      LAYER met4 ;
        RECT 50.830000 39.400000 51.150000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 39.840000 51.150000 40.160000 ;
      LAYER met4 ;
        RECT 50.830000 39.840000 51.150000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 51.655000 51.150000 51.975000 ;
      LAYER met4 ;
        RECT 50.830000 51.655000 51.150000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 52.075000 51.150000 52.395000 ;
      LAYER met4 ;
        RECT 50.830000 52.075000 51.150000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830000 52.495000 51.150000 52.815000 ;
      LAYER met4 ;
        RECT 50.830000 52.495000 51.150000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.230000 47.740000 51.550000 48.060000 ;
      LAYER met4 ;
        RECT 51.230000 47.740000 51.550000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.230000 56.410000 51.550000 56.730000 ;
      LAYER met4 ;
        RECT 51.230000 56.410000 51.550000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 36.760000 51.560000 37.080000 ;
      LAYER met4 ;
        RECT 51.240000 36.760000 51.560000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 37.200000 51.560000 37.520000 ;
      LAYER met4 ;
        RECT 51.240000 37.200000 51.560000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 37.640000 51.560000 37.960000 ;
      LAYER met4 ;
        RECT 51.240000 37.640000 51.560000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 38.080000 51.560000 38.400000 ;
      LAYER met4 ;
        RECT 51.240000 38.080000 51.560000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 38.520000 51.560000 38.840000 ;
      LAYER met4 ;
        RECT 51.240000 38.520000 51.560000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 38.960000 51.560000 39.280000 ;
      LAYER met4 ;
        RECT 51.240000 38.960000 51.560000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 39.400000 51.560000 39.720000 ;
      LAYER met4 ;
        RECT 51.240000 39.400000 51.560000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 39.840000 51.560000 40.160000 ;
      LAYER met4 ;
        RECT 51.240000 39.840000 51.560000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 51.655000 51.560000 51.975000 ;
      LAYER met4 ;
        RECT 51.240000 51.655000 51.560000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 52.075000 51.560000 52.395000 ;
      LAYER met4 ;
        RECT 51.240000 52.075000 51.560000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240000 52.495000 51.560000 52.815000 ;
      LAYER met4 ;
        RECT 51.240000 52.495000 51.560000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.635000 47.740000 51.955000 48.060000 ;
      LAYER met4 ;
        RECT 51.635000 47.740000 51.955000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.635000 56.410000 51.955000 56.730000 ;
      LAYER met4 ;
        RECT 51.635000 56.410000 51.955000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 36.760000 51.970000 37.080000 ;
      LAYER met4 ;
        RECT 51.650000 36.760000 51.970000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 37.200000 51.970000 37.520000 ;
      LAYER met4 ;
        RECT 51.650000 37.200000 51.970000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 37.640000 51.970000 37.960000 ;
      LAYER met4 ;
        RECT 51.650000 37.640000 51.970000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 38.080000 51.970000 38.400000 ;
      LAYER met4 ;
        RECT 51.650000 38.080000 51.970000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 38.520000 51.970000 38.840000 ;
      LAYER met4 ;
        RECT 51.650000 38.520000 51.970000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 38.960000 51.970000 39.280000 ;
      LAYER met4 ;
        RECT 51.650000 38.960000 51.970000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 39.400000 51.970000 39.720000 ;
      LAYER met4 ;
        RECT 51.650000 39.400000 51.970000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 39.840000 51.970000 40.160000 ;
      LAYER met4 ;
        RECT 51.650000 39.840000 51.970000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 51.655000 51.970000 51.975000 ;
      LAYER met4 ;
        RECT 51.650000 51.655000 51.970000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 52.075000 51.970000 52.395000 ;
      LAYER met4 ;
        RECT 51.650000 52.075000 51.970000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650000 52.495000 51.970000 52.815000 ;
      LAYER met4 ;
        RECT 51.650000 52.495000 51.970000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.040000 47.740000 52.360000 48.060000 ;
      LAYER met4 ;
        RECT 52.040000 47.740000 52.360000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.040000 56.410000 52.360000 56.730000 ;
      LAYER met4 ;
        RECT 52.040000 56.410000 52.360000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 36.760000 52.380000 37.080000 ;
      LAYER met4 ;
        RECT 52.060000 36.760000 52.380000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 37.200000 52.380000 37.520000 ;
      LAYER met4 ;
        RECT 52.060000 37.200000 52.380000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 37.640000 52.380000 37.960000 ;
      LAYER met4 ;
        RECT 52.060000 37.640000 52.380000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 38.080000 52.380000 38.400000 ;
      LAYER met4 ;
        RECT 52.060000 38.080000 52.380000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 38.520000 52.380000 38.840000 ;
      LAYER met4 ;
        RECT 52.060000 38.520000 52.380000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 38.960000 52.380000 39.280000 ;
      LAYER met4 ;
        RECT 52.060000 38.960000 52.380000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 39.400000 52.380000 39.720000 ;
      LAYER met4 ;
        RECT 52.060000 39.400000 52.380000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 39.840000 52.380000 40.160000 ;
      LAYER met4 ;
        RECT 52.060000 39.840000 52.380000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 51.655000 52.380000 51.975000 ;
      LAYER met4 ;
        RECT 52.060000 51.655000 52.380000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 52.075000 52.380000 52.395000 ;
      LAYER met4 ;
        RECT 52.060000 52.075000 52.380000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060000 52.495000 52.380000 52.815000 ;
      LAYER met4 ;
        RECT 52.060000 52.495000 52.380000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.445000 47.740000 52.765000 48.060000 ;
      LAYER met4 ;
        RECT 52.445000 47.740000 52.765000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.445000 56.410000 52.765000 56.730000 ;
      LAYER met4 ;
        RECT 52.445000 56.410000 52.765000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 36.760000 52.790000 37.080000 ;
      LAYER met4 ;
        RECT 52.470000 36.760000 52.790000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 37.200000 52.790000 37.520000 ;
      LAYER met4 ;
        RECT 52.470000 37.200000 52.790000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 37.640000 52.790000 37.960000 ;
      LAYER met4 ;
        RECT 52.470000 37.640000 52.790000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 38.080000 52.790000 38.400000 ;
      LAYER met4 ;
        RECT 52.470000 38.080000 52.790000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 38.520000 52.790000 38.840000 ;
      LAYER met4 ;
        RECT 52.470000 38.520000 52.790000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 38.960000 52.790000 39.280000 ;
      LAYER met4 ;
        RECT 52.470000 38.960000 52.790000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 39.400000 52.790000 39.720000 ;
      LAYER met4 ;
        RECT 52.470000 39.400000 52.790000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 39.840000 52.790000 40.160000 ;
      LAYER met4 ;
        RECT 52.470000 39.840000 52.790000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 51.655000 52.790000 51.975000 ;
      LAYER met4 ;
        RECT 52.470000 51.655000 52.790000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 52.075000 52.790000 52.395000 ;
      LAYER met4 ;
        RECT 52.470000 52.075000 52.790000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470000 52.495000 52.790000 52.815000 ;
      LAYER met4 ;
        RECT 52.470000 52.495000 52.790000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.850000 47.740000 53.170000 48.060000 ;
      LAYER met4 ;
        RECT 52.850000 47.740000 53.170000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.850000 56.410000 53.170000 56.730000 ;
      LAYER met4 ;
        RECT 52.850000 56.410000 53.170000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 36.760000 53.200000 37.080000 ;
      LAYER met4 ;
        RECT 52.880000 36.760000 53.200000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 37.200000 53.200000 37.520000 ;
      LAYER met4 ;
        RECT 52.880000 37.200000 53.200000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 37.640000 53.200000 37.960000 ;
      LAYER met4 ;
        RECT 52.880000 37.640000 53.200000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 38.080000 53.200000 38.400000 ;
      LAYER met4 ;
        RECT 52.880000 38.080000 53.200000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 38.520000 53.200000 38.840000 ;
      LAYER met4 ;
        RECT 52.880000 38.520000 53.200000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 38.960000 53.200000 39.280000 ;
      LAYER met4 ;
        RECT 52.880000 38.960000 53.200000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 39.400000 53.200000 39.720000 ;
      LAYER met4 ;
        RECT 52.880000 39.400000 53.200000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 39.840000 53.200000 40.160000 ;
      LAYER met4 ;
        RECT 52.880000 39.840000 53.200000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 51.655000 53.200000 51.975000 ;
      LAYER met4 ;
        RECT 52.880000 51.655000 53.200000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 52.075000 53.200000 52.395000 ;
      LAYER met4 ;
        RECT 52.880000 52.075000 53.200000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880000 52.495000 53.200000 52.815000 ;
      LAYER met4 ;
        RECT 52.880000 52.495000 53.200000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.255000 47.740000 53.575000 48.060000 ;
      LAYER met4 ;
        RECT 53.255000 47.740000 53.575000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.255000 56.410000 53.575000 56.730000 ;
      LAYER met4 ;
        RECT 53.255000 56.410000 53.575000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 36.760000 53.605000 37.080000 ;
      LAYER met4 ;
        RECT 53.285000 36.760000 53.605000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 37.200000 53.605000 37.520000 ;
      LAYER met4 ;
        RECT 53.285000 37.200000 53.605000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 37.640000 53.605000 37.960000 ;
      LAYER met4 ;
        RECT 53.285000 37.640000 53.605000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 38.080000 53.605000 38.400000 ;
      LAYER met4 ;
        RECT 53.285000 38.080000 53.605000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 38.520000 53.605000 38.840000 ;
      LAYER met4 ;
        RECT 53.285000 38.520000 53.605000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 38.960000 53.605000 39.280000 ;
      LAYER met4 ;
        RECT 53.285000 38.960000 53.605000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 39.400000 53.605000 39.720000 ;
      LAYER met4 ;
        RECT 53.285000 39.400000 53.605000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 39.840000 53.605000 40.160000 ;
      LAYER met4 ;
        RECT 53.285000 39.840000 53.605000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 51.655000 53.605000 51.975000 ;
      LAYER met4 ;
        RECT 53.285000 51.655000 53.605000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 52.075000 53.605000 52.395000 ;
      LAYER met4 ;
        RECT 53.285000 52.075000 53.605000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285000 52.495000 53.605000 52.815000 ;
      LAYER met4 ;
        RECT 53.285000 52.495000 53.605000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.660000 47.740000 53.980000 48.060000 ;
      LAYER met4 ;
        RECT 53.660000 47.740000 53.980000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.660000 56.410000 53.980000 56.730000 ;
      LAYER met4 ;
        RECT 53.660000 56.410000 53.980000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 36.760000 54.010000 37.080000 ;
      LAYER met4 ;
        RECT 53.690000 36.760000 54.010000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 37.200000 54.010000 37.520000 ;
      LAYER met4 ;
        RECT 53.690000 37.200000 54.010000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 37.640000 54.010000 37.960000 ;
      LAYER met4 ;
        RECT 53.690000 37.640000 54.010000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 38.080000 54.010000 38.400000 ;
      LAYER met4 ;
        RECT 53.690000 38.080000 54.010000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 38.520000 54.010000 38.840000 ;
      LAYER met4 ;
        RECT 53.690000 38.520000 54.010000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 38.960000 54.010000 39.280000 ;
      LAYER met4 ;
        RECT 53.690000 38.960000 54.010000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 39.400000 54.010000 39.720000 ;
      LAYER met4 ;
        RECT 53.690000 39.400000 54.010000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 39.840000 54.010000 40.160000 ;
      LAYER met4 ;
        RECT 53.690000 39.840000 54.010000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 51.655000 54.010000 51.975000 ;
      LAYER met4 ;
        RECT 53.690000 51.655000 54.010000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 52.075000 54.010000 52.395000 ;
      LAYER met4 ;
        RECT 53.690000 52.075000 54.010000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690000 52.495000 54.010000 52.815000 ;
      LAYER met4 ;
        RECT 53.690000 52.495000 54.010000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 47.740000 54.385000 48.060000 ;
      LAYER met4 ;
        RECT 54.065000 47.740000 54.385000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.065000 56.410000 54.385000 56.730000 ;
      LAYER met4 ;
        RECT 54.065000 56.410000 54.385000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 36.760000 54.415000 37.080000 ;
      LAYER met4 ;
        RECT 54.095000 36.760000 54.415000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 37.200000 54.415000 37.520000 ;
      LAYER met4 ;
        RECT 54.095000 37.200000 54.415000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 37.640000 54.415000 37.960000 ;
      LAYER met4 ;
        RECT 54.095000 37.640000 54.415000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 38.080000 54.415000 38.400000 ;
      LAYER met4 ;
        RECT 54.095000 38.080000 54.415000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 38.520000 54.415000 38.840000 ;
      LAYER met4 ;
        RECT 54.095000 38.520000 54.415000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 38.960000 54.415000 39.280000 ;
      LAYER met4 ;
        RECT 54.095000 38.960000 54.415000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 39.400000 54.415000 39.720000 ;
      LAYER met4 ;
        RECT 54.095000 39.400000 54.415000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 39.840000 54.415000 40.160000 ;
      LAYER met4 ;
        RECT 54.095000 39.840000 54.415000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 51.655000 54.415000 51.975000 ;
      LAYER met4 ;
        RECT 54.095000 51.655000 54.415000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 52.075000 54.415000 52.395000 ;
      LAYER met4 ;
        RECT 54.095000 52.075000 54.415000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095000 52.495000 54.415000 52.815000 ;
      LAYER met4 ;
        RECT 54.095000 52.495000 54.415000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.470000 47.740000 54.790000 48.060000 ;
      LAYER met4 ;
        RECT 54.470000 47.740000 54.790000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.470000 56.410000 54.790000 56.730000 ;
      LAYER met4 ;
        RECT 54.470000 56.410000 54.790000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 36.760000 54.820000 37.080000 ;
      LAYER met4 ;
        RECT 54.500000 36.760000 54.820000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 37.200000 54.820000 37.520000 ;
      LAYER met4 ;
        RECT 54.500000 37.200000 54.820000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 37.640000 54.820000 37.960000 ;
      LAYER met4 ;
        RECT 54.500000 37.640000 54.820000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 38.080000 54.820000 38.400000 ;
      LAYER met4 ;
        RECT 54.500000 38.080000 54.820000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 38.520000 54.820000 38.840000 ;
      LAYER met4 ;
        RECT 54.500000 38.520000 54.820000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 38.960000 54.820000 39.280000 ;
      LAYER met4 ;
        RECT 54.500000 38.960000 54.820000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 39.400000 54.820000 39.720000 ;
      LAYER met4 ;
        RECT 54.500000 39.400000 54.820000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 39.840000 54.820000 40.160000 ;
      LAYER met4 ;
        RECT 54.500000 39.840000 54.820000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 51.655000 54.820000 51.975000 ;
      LAYER met4 ;
        RECT 54.500000 51.655000 54.820000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 52.075000 54.820000 52.395000 ;
      LAYER met4 ;
        RECT 54.500000 52.075000 54.820000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500000 52.495000 54.820000 52.815000 ;
      LAYER met4 ;
        RECT 54.500000 52.495000 54.820000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.875000 47.740000 55.195000 48.060000 ;
      LAYER met4 ;
        RECT 54.875000 47.740000 55.195000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.875000 56.410000 55.195000 56.730000 ;
      LAYER met4 ;
        RECT 54.875000 56.410000 55.195000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 36.760000 55.225000 37.080000 ;
      LAYER met4 ;
        RECT 54.905000 36.760000 55.225000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 37.200000 55.225000 37.520000 ;
      LAYER met4 ;
        RECT 54.905000 37.200000 55.225000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 37.640000 55.225000 37.960000 ;
      LAYER met4 ;
        RECT 54.905000 37.640000 55.225000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 38.080000 55.225000 38.400000 ;
      LAYER met4 ;
        RECT 54.905000 38.080000 55.225000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 38.520000 55.225000 38.840000 ;
      LAYER met4 ;
        RECT 54.905000 38.520000 55.225000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 38.960000 55.225000 39.280000 ;
      LAYER met4 ;
        RECT 54.905000 38.960000 55.225000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 39.400000 55.225000 39.720000 ;
      LAYER met4 ;
        RECT 54.905000 39.400000 55.225000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 39.840000 55.225000 40.160000 ;
      LAYER met4 ;
        RECT 54.905000 39.840000 55.225000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 51.655000 55.225000 51.975000 ;
      LAYER met4 ;
        RECT 54.905000 51.655000 55.225000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 52.075000 55.225000 52.395000 ;
      LAYER met4 ;
        RECT 54.905000 52.075000 55.225000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905000 52.495000 55.225000 52.815000 ;
      LAYER met4 ;
        RECT 54.905000 52.495000 55.225000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.280000 47.740000 55.600000 48.060000 ;
      LAYER met4 ;
        RECT 55.280000 47.740000 55.600000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.280000 56.410000 55.600000 56.730000 ;
      LAYER met4 ;
        RECT 55.280000 56.410000 55.600000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 36.760000 55.630000 37.080000 ;
      LAYER met4 ;
        RECT 55.310000 36.760000 55.630000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 37.200000 55.630000 37.520000 ;
      LAYER met4 ;
        RECT 55.310000 37.200000 55.630000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 37.640000 55.630000 37.960000 ;
      LAYER met4 ;
        RECT 55.310000 37.640000 55.630000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 38.080000 55.630000 38.400000 ;
      LAYER met4 ;
        RECT 55.310000 38.080000 55.630000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 38.520000 55.630000 38.840000 ;
      LAYER met4 ;
        RECT 55.310000 38.520000 55.630000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 38.960000 55.630000 39.280000 ;
      LAYER met4 ;
        RECT 55.310000 38.960000 55.630000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 39.400000 55.630000 39.720000 ;
      LAYER met4 ;
        RECT 55.310000 39.400000 55.630000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 39.840000 55.630000 40.160000 ;
      LAYER met4 ;
        RECT 55.310000 39.840000 55.630000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 51.655000 55.630000 51.975000 ;
      LAYER met4 ;
        RECT 55.310000 51.655000 55.630000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 52.075000 55.630000 52.395000 ;
      LAYER met4 ;
        RECT 55.310000 52.075000 55.630000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310000 52.495000 55.630000 52.815000 ;
      LAYER met4 ;
        RECT 55.310000 52.495000 55.630000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.685000 47.740000 56.005000 48.060000 ;
      LAYER met4 ;
        RECT 55.685000 47.740000 56.005000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.685000 56.410000 56.005000 56.730000 ;
      LAYER met4 ;
        RECT 55.685000 56.410000 56.005000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 36.760000 56.035000 37.080000 ;
      LAYER met4 ;
        RECT 55.715000 36.760000 56.035000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 37.200000 56.035000 37.520000 ;
      LAYER met4 ;
        RECT 55.715000 37.200000 56.035000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 37.640000 56.035000 37.960000 ;
      LAYER met4 ;
        RECT 55.715000 37.640000 56.035000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 38.080000 56.035000 38.400000 ;
      LAYER met4 ;
        RECT 55.715000 38.080000 56.035000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 38.520000 56.035000 38.840000 ;
      LAYER met4 ;
        RECT 55.715000 38.520000 56.035000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 38.960000 56.035000 39.280000 ;
      LAYER met4 ;
        RECT 55.715000 38.960000 56.035000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 39.400000 56.035000 39.720000 ;
      LAYER met4 ;
        RECT 55.715000 39.400000 56.035000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 39.840000 56.035000 40.160000 ;
      LAYER met4 ;
        RECT 55.715000 39.840000 56.035000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 51.655000 56.035000 51.975000 ;
      LAYER met4 ;
        RECT 55.715000 51.655000 56.035000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 52.075000 56.035000 52.395000 ;
      LAYER met4 ;
        RECT 55.715000 52.075000 56.035000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715000 52.495000 56.035000 52.815000 ;
      LAYER met4 ;
        RECT 55.715000 52.495000 56.035000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.090000 47.740000 56.410000 48.060000 ;
      LAYER met4 ;
        RECT 56.090000 47.740000 56.410000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.090000 56.410000 56.410000 56.730000 ;
      LAYER met4 ;
        RECT 56.090000 56.410000 56.410000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 36.760000 56.440000 37.080000 ;
      LAYER met4 ;
        RECT 56.120000 36.760000 56.440000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 37.200000 56.440000 37.520000 ;
      LAYER met4 ;
        RECT 56.120000 37.200000 56.440000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 37.640000 56.440000 37.960000 ;
      LAYER met4 ;
        RECT 56.120000 37.640000 56.440000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 38.080000 56.440000 38.400000 ;
      LAYER met4 ;
        RECT 56.120000 38.080000 56.440000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 38.520000 56.440000 38.840000 ;
      LAYER met4 ;
        RECT 56.120000 38.520000 56.440000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 38.960000 56.440000 39.280000 ;
      LAYER met4 ;
        RECT 56.120000 38.960000 56.440000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 39.400000 56.440000 39.720000 ;
      LAYER met4 ;
        RECT 56.120000 39.400000 56.440000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 39.840000 56.440000 40.160000 ;
      LAYER met4 ;
        RECT 56.120000 39.840000 56.440000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 51.655000 56.440000 51.975000 ;
      LAYER met4 ;
        RECT 56.120000 51.655000 56.440000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 52.075000 56.440000 52.395000 ;
      LAYER met4 ;
        RECT 56.120000 52.075000 56.440000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120000 52.495000 56.440000 52.815000 ;
      LAYER met4 ;
        RECT 56.120000 52.495000 56.440000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.495000 47.740000 56.815000 48.060000 ;
      LAYER met4 ;
        RECT 56.495000 47.740000 56.815000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.495000 56.410000 56.815000 56.730000 ;
      LAYER met4 ;
        RECT 56.495000 56.410000 56.815000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 36.760000 56.845000 37.080000 ;
      LAYER met4 ;
        RECT 56.525000 36.760000 56.845000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 37.200000 56.845000 37.520000 ;
      LAYER met4 ;
        RECT 56.525000 37.200000 56.845000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 37.640000 56.845000 37.960000 ;
      LAYER met4 ;
        RECT 56.525000 37.640000 56.845000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 38.080000 56.845000 38.400000 ;
      LAYER met4 ;
        RECT 56.525000 38.080000 56.845000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 38.520000 56.845000 38.840000 ;
      LAYER met4 ;
        RECT 56.525000 38.520000 56.845000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 38.960000 56.845000 39.280000 ;
      LAYER met4 ;
        RECT 56.525000 38.960000 56.845000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 39.400000 56.845000 39.720000 ;
      LAYER met4 ;
        RECT 56.525000 39.400000 56.845000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 39.840000 56.845000 40.160000 ;
      LAYER met4 ;
        RECT 56.525000 39.840000 56.845000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 51.655000 56.845000 51.975000 ;
      LAYER met4 ;
        RECT 56.525000 51.655000 56.845000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 52.075000 56.845000 52.395000 ;
      LAYER met4 ;
        RECT 56.525000 52.075000 56.845000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525000 52.495000 56.845000 52.815000 ;
      LAYER met4 ;
        RECT 56.525000 52.495000 56.845000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.900000 47.740000 57.220000 48.060000 ;
      LAYER met4 ;
        RECT 56.900000 47.740000 57.220000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.900000 56.410000 57.220000 56.730000 ;
      LAYER met4 ;
        RECT 56.900000 56.410000 57.220000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 36.760000 57.250000 37.080000 ;
      LAYER met4 ;
        RECT 56.930000 36.760000 57.250000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 37.200000 57.250000 37.520000 ;
      LAYER met4 ;
        RECT 56.930000 37.200000 57.250000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 37.640000 57.250000 37.960000 ;
      LAYER met4 ;
        RECT 56.930000 37.640000 57.250000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 38.080000 57.250000 38.400000 ;
      LAYER met4 ;
        RECT 56.930000 38.080000 57.250000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 38.520000 57.250000 38.840000 ;
      LAYER met4 ;
        RECT 56.930000 38.520000 57.250000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 38.960000 57.250000 39.280000 ;
      LAYER met4 ;
        RECT 56.930000 38.960000 57.250000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 39.400000 57.250000 39.720000 ;
      LAYER met4 ;
        RECT 56.930000 39.400000 57.250000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 39.840000 57.250000 40.160000 ;
      LAYER met4 ;
        RECT 56.930000 39.840000 57.250000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 51.655000 57.250000 51.975000 ;
      LAYER met4 ;
        RECT 56.930000 51.655000 57.250000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 52.075000 57.250000 52.395000 ;
      LAYER met4 ;
        RECT 56.930000 52.075000 57.250000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930000 52.495000 57.250000 52.815000 ;
      LAYER met4 ;
        RECT 56.930000 52.495000 57.250000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.305000 47.740000 57.625000 48.060000 ;
      LAYER met4 ;
        RECT 57.305000 47.740000 57.625000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.305000 56.410000 57.625000 56.730000 ;
      LAYER met4 ;
        RECT 57.305000 56.410000 57.625000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 36.760000 57.655000 37.080000 ;
      LAYER met4 ;
        RECT 57.335000 36.760000 57.655000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 37.200000 57.655000 37.520000 ;
      LAYER met4 ;
        RECT 57.335000 37.200000 57.655000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 37.640000 57.655000 37.960000 ;
      LAYER met4 ;
        RECT 57.335000 37.640000 57.655000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 38.080000 57.655000 38.400000 ;
      LAYER met4 ;
        RECT 57.335000 38.080000 57.655000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 38.520000 57.655000 38.840000 ;
      LAYER met4 ;
        RECT 57.335000 38.520000 57.655000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 38.960000 57.655000 39.280000 ;
      LAYER met4 ;
        RECT 57.335000 38.960000 57.655000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 39.400000 57.655000 39.720000 ;
      LAYER met4 ;
        RECT 57.335000 39.400000 57.655000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 39.840000 57.655000 40.160000 ;
      LAYER met4 ;
        RECT 57.335000 39.840000 57.655000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 51.655000 57.655000 51.975000 ;
      LAYER met4 ;
        RECT 57.335000 51.655000 57.655000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 52.075000 57.655000 52.395000 ;
      LAYER met4 ;
        RECT 57.335000 52.075000 57.655000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335000 52.495000 57.655000 52.815000 ;
      LAYER met4 ;
        RECT 57.335000 52.495000 57.655000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.710000 47.740000 58.030000 48.060000 ;
      LAYER met4 ;
        RECT 57.710000 47.740000 58.030000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.710000 56.410000 58.030000 56.730000 ;
      LAYER met4 ;
        RECT 57.710000 56.410000 58.030000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 36.760000 58.060000 37.080000 ;
      LAYER met4 ;
        RECT 57.740000 36.760000 58.060000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 37.200000 58.060000 37.520000 ;
      LAYER met4 ;
        RECT 57.740000 37.200000 58.060000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 37.640000 58.060000 37.960000 ;
      LAYER met4 ;
        RECT 57.740000 37.640000 58.060000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 38.080000 58.060000 38.400000 ;
      LAYER met4 ;
        RECT 57.740000 38.080000 58.060000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 38.520000 58.060000 38.840000 ;
      LAYER met4 ;
        RECT 57.740000 38.520000 58.060000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 38.960000 58.060000 39.280000 ;
      LAYER met4 ;
        RECT 57.740000 38.960000 58.060000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 39.400000 58.060000 39.720000 ;
      LAYER met4 ;
        RECT 57.740000 39.400000 58.060000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 39.840000 58.060000 40.160000 ;
      LAYER met4 ;
        RECT 57.740000 39.840000 58.060000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 51.655000 58.060000 51.975000 ;
      LAYER met4 ;
        RECT 57.740000 51.655000 58.060000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 52.075000 58.060000 52.395000 ;
      LAYER met4 ;
        RECT 57.740000 52.075000 58.060000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740000 52.495000 58.060000 52.815000 ;
      LAYER met4 ;
        RECT 57.740000 52.495000 58.060000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.115000 47.740000 58.435000 48.060000 ;
      LAYER met4 ;
        RECT 58.115000 47.740000 58.435000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.115000 56.410000 58.435000 56.730000 ;
      LAYER met4 ;
        RECT 58.115000 56.410000 58.435000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 36.760000 58.465000 37.080000 ;
      LAYER met4 ;
        RECT 58.145000 36.760000 58.465000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 37.200000 58.465000 37.520000 ;
      LAYER met4 ;
        RECT 58.145000 37.200000 58.465000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 37.640000 58.465000 37.960000 ;
      LAYER met4 ;
        RECT 58.145000 37.640000 58.465000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 38.080000 58.465000 38.400000 ;
      LAYER met4 ;
        RECT 58.145000 38.080000 58.465000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 38.520000 58.465000 38.840000 ;
      LAYER met4 ;
        RECT 58.145000 38.520000 58.465000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 38.960000 58.465000 39.280000 ;
      LAYER met4 ;
        RECT 58.145000 38.960000 58.465000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 39.400000 58.465000 39.720000 ;
      LAYER met4 ;
        RECT 58.145000 39.400000 58.465000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 39.840000 58.465000 40.160000 ;
      LAYER met4 ;
        RECT 58.145000 39.840000 58.465000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 51.655000 58.465000 51.975000 ;
      LAYER met4 ;
        RECT 58.145000 51.655000 58.465000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 52.075000 58.465000 52.395000 ;
      LAYER met4 ;
        RECT 58.145000 52.075000 58.465000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145000 52.495000 58.465000 52.815000 ;
      LAYER met4 ;
        RECT 58.145000 52.495000 58.465000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.520000 47.740000 58.840000 48.060000 ;
      LAYER met4 ;
        RECT 58.520000 47.740000 58.840000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.520000 56.410000 58.840000 56.730000 ;
      LAYER met4 ;
        RECT 58.520000 56.410000 58.840000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 36.760000 58.870000 37.080000 ;
      LAYER met4 ;
        RECT 58.550000 36.760000 58.870000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 37.200000 58.870000 37.520000 ;
      LAYER met4 ;
        RECT 58.550000 37.200000 58.870000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 37.640000 58.870000 37.960000 ;
      LAYER met4 ;
        RECT 58.550000 37.640000 58.870000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 38.080000 58.870000 38.400000 ;
      LAYER met4 ;
        RECT 58.550000 38.080000 58.870000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 38.520000 58.870000 38.840000 ;
      LAYER met4 ;
        RECT 58.550000 38.520000 58.870000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 38.960000 58.870000 39.280000 ;
      LAYER met4 ;
        RECT 58.550000 38.960000 58.870000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 39.400000 58.870000 39.720000 ;
      LAYER met4 ;
        RECT 58.550000 39.400000 58.870000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 39.840000 58.870000 40.160000 ;
      LAYER met4 ;
        RECT 58.550000 39.840000 58.870000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 51.655000 58.870000 51.975000 ;
      LAYER met4 ;
        RECT 58.550000 51.655000 58.870000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 52.075000 58.870000 52.395000 ;
      LAYER met4 ;
        RECT 58.550000 52.075000 58.870000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550000 52.495000 58.870000 52.815000 ;
      LAYER met4 ;
        RECT 58.550000 52.495000 58.870000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.925000 47.740000 59.245000 48.060000 ;
      LAYER met4 ;
        RECT 58.925000 47.740000 59.245000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.925000 56.410000 59.245000 56.730000 ;
      LAYER met4 ;
        RECT 58.925000 56.410000 59.245000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 36.760000 59.275000 37.080000 ;
      LAYER met4 ;
        RECT 58.955000 36.760000 59.275000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 37.200000 59.275000 37.520000 ;
      LAYER met4 ;
        RECT 58.955000 37.200000 59.275000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 37.640000 59.275000 37.960000 ;
      LAYER met4 ;
        RECT 58.955000 37.640000 59.275000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 38.080000 59.275000 38.400000 ;
      LAYER met4 ;
        RECT 58.955000 38.080000 59.275000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 38.520000 59.275000 38.840000 ;
      LAYER met4 ;
        RECT 58.955000 38.520000 59.275000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 38.960000 59.275000 39.280000 ;
      LAYER met4 ;
        RECT 58.955000 38.960000 59.275000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 39.400000 59.275000 39.720000 ;
      LAYER met4 ;
        RECT 58.955000 39.400000 59.275000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 39.840000 59.275000 40.160000 ;
      LAYER met4 ;
        RECT 58.955000 39.840000 59.275000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 51.655000 59.275000 51.975000 ;
      LAYER met4 ;
        RECT 58.955000 51.655000 59.275000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 52.075000 59.275000 52.395000 ;
      LAYER met4 ;
        RECT 58.955000 52.075000 59.275000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955000 52.495000 59.275000 52.815000 ;
      LAYER met4 ;
        RECT 58.955000 52.495000 59.275000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.330000 47.740000 59.650000 48.060000 ;
      LAYER met4 ;
        RECT 59.330000 47.740000 59.650000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.330000 56.410000 59.650000 56.730000 ;
      LAYER met4 ;
        RECT 59.330000 56.410000 59.650000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 36.760000 59.680000 37.080000 ;
      LAYER met4 ;
        RECT 59.360000 36.760000 59.680000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 37.200000 59.680000 37.520000 ;
      LAYER met4 ;
        RECT 59.360000 37.200000 59.680000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 37.640000 59.680000 37.960000 ;
      LAYER met4 ;
        RECT 59.360000 37.640000 59.680000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 38.080000 59.680000 38.400000 ;
      LAYER met4 ;
        RECT 59.360000 38.080000 59.680000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 38.520000 59.680000 38.840000 ;
      LAYER met4 ;
        RECT 59.360000 38.520000 59.680000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 38.960000 59.680000 39.280000 ;
      LAYER met4 ;
        RECT 59.360000 38.960000 59.680000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 39.400000 59.680000 39.720000 ;
      LAYER met4 ;
        RECT 59.360000 39.400000 59.680000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 39.840000 59.680000 40.160000 ;
      LAYER met4 ;
        RECT 59.360000 39.840000 59.680000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 51.655000 59.680000 51.975000 ;
      LAYER met4 ;
        RECT 59.360000 51.655000 59.680000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 52.075000 59.680000 52.395000 ;
      LAYER met4 ;
        RECT 59.360000 52.075000 59.680000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360000 52.495000 59.680000 52.815000 ;
      LAYER met4 ;
        RECT 59.360000 52.495000 59.680000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.735000 47.740000 60.055000 48.060000 ;
      LAYER met4 ;
        RECT 59.735000 47.740000 60.055000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.735000 56.410000 60.055000 56.730000 ;
      LAYER met4 ;
        RECT 59.735000 56.410000 60.055000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 36.760000 60.085000 37.080000 ;
      LAYER met4 ;
        RECT 59.765000 36.760000 60.085000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 37.200000 60.085000 37.520000 ;
      LAYER met4 ;
        RECT 59.765000 37.200000 60.085000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 37.640000 60.085000 37.960000 ;
      LAYER met4 ;
        RECT 59.765000 37.640000 60.085000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 38.080000 60.085000 38.400000 ;
      LAYER met4 ;
        RECT 59.765000 38.080000 60.085000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 38.520000 60.085000 38.840000 ;
      LAYER met4 ;
        RECT 59.765000 38.520000 60.085000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 38.960000 60.085000 39.280000 ;
      LAYER met4 ;
        RECT 59.765000 38.960000 60.085000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 39.400000 60.085000 39.720000 ;
      LAYER met4 ;
        RECT 59.765000 39.400000 60.085000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 39.840000 60.085000 40.160000 ;
      LAYER met4 ;
        RECT 59.765000 39.840000 60.085000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 51.655000 60.085000 51.975000 ;
      LAYER met4 ;
        RECT 59.765000 51.655000 60.085000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 52.075000 60.085000 52.395000 ;
      LAYER met4 ;
        RECT 59.765000 52.075000 60.085000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765000 52.495000 60.085000 52.815000 ;
      LAYER met4 ;
        RECT 59.765000 52.495000 60.085000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 51.655000 6.545000 51.975000 ;
      LAYER met4 ;
        RECT 6.225000 51.655000 6.545000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 52.075000 6.545000 52.395000 ;
      LAYER met4 ;
        RECT 6.225000 52.075000 6.545000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225000 52.495000 6.545000 52.815000 ;
      LAYER met4 ;
        RECT 6.225000 52.495000 6.545000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 47.740000 6.550000 48.060000 ;
      LAYER met4 ;
        RECT 6.230000 47.740000 6.550000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230000 56.410000 6.550000 56.730000 ;
      LAYER met4 ;
        RECT 6.230000 56.410000 6.550000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265000 36.760000 6.585000 37.080000 ;
      LAYER met4 ;
        RECT 6.265000 36.760000 6.585000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265000 37.200000 6.585000 37.520000 ;
      LAYER met4 ;
        RECT 6.265000 37.200000 6.585000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265000 37.640000 6.585000 37.960000 ;
      LAYER met4 ;
        RECT 6.265000 37.640000 6.585000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265000 38.080000 6.585000 38.400000 ;
      LAYER met4 ;
        RECT 6.265000 38.080000 6.585000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265000 38.520000 6.585000 38.840000 ;
      LAYER met4 ;
        RECT 6.265000 38.520000 6.585000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265000 38.960000 6.585000 39.280000 ;
      LAYER met4 ;
        RECT 6.265000 38.960000 6.585000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265000 39.400000 6.585000 39.720000 ;
      LAYER met4 ;
        RECT 6.265000 39.400000 6.585000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265000 39.840000 6.585000 40.160000 ;
      LAYER met4 ;
        RECT 6.265000 39.840000 6.585000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 51.655000 6.950000 51.975000 ;
      LAYER met4 ;
        RECT 6.630000 51.655000 6.950000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 52.075000 6.950000 52.395000 ;
      LAYER met4 ;
        RECT 6.630000 52.075000 6.950000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630000 52.495000 6.950000 52.815000 ;
      LAYER met4 ;
        RECT 6.630000 52.495000 6.950000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 47.740000 6.955000 48.060000 ;
      LAYER met4 ;
        RECT 6.635000 47.740000 6.955000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635000 56.410000 6.955000 56.730000 ;
      LAYER met4 ;
        RECT 6.635000 56.410000 6.955000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670000 36.760000 6.990000 37.080000 ;
      LAYER met4 ;
        RECT 6.670000 36.760000 6.990000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670000 37.200000 6.990000 37.520000 ;
      LAYER met4 ;
        RECT 6.670000 37.200000 6.990000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670000 37.640000 6.990000 37.960000 ;
      LAYER met4 ;
        RECT 6.670000 37.640000 6.990000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670000 38.080000 6.990000 38.400000 ;
      LAYER met4 ;
        RECT 6.670000 38.080000 6.990000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670000 38.520000 6.990000 38.840000 ;
      LAYER met4 ;
        RECT 6.670000 38.520000 6.990000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670000 38.960000 6.990000 39.280000 ;
      LAYER met4 ;
        RECT 6.670000 38.960000 6.990000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670000 39.400000 6.990000 39.720000 ;
      LAYER met4 ;
        RECT 6.670000 39.400000 6.990000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670000 39.840000 6.990000 40.160000 ;
      LAYER met4 ;
        RECT 6.670000 39.840000 6.990000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.140000 47.740000 60.460000 48.060000 ;
      LAYER met4 ;
        RECT 60.140000 47.740000 60.460000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.140000 56.410000 60.460000 56.730000 ;
      LAYER met4 ;
        RECT 60.140000 56.410000 60.460000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 36.760000 60.490000 37.080000 ;
      LAYER met4 ;
        RECT 60.170000 36.760000 60.490000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 37.200000 60.490000 37.520000 ;
      LAYER met4 ;
        RECT 60.170000 37.200000 60.490000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 37.640000 60.490000 37.960000 ;
      LAYER met4 ;
        RECT 60.170000 37.640000 60.490000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 38.080000 60.490000 38.400000 ;
      LAYER met4 ;
        RECT 60.170000 38.080000 60.490000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 38.520000 60.490000 38.840000 ;
      LAYER met4 ;
        RECT 60.170000 38.520000 60.490000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 38.960000 60.490000 39.280000 ;
      LAYER met4 ;
        RECT 60.170000 38.960000 60.490000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 39.400000 60.490000 39.720000 ;
      LAYER met4 ;
        RECT 60.170000 39.400000 60.490000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 39.840000 60.490000 40.160000 ;
      LAYER met4 ;
        RECT 60.170000 39.840000 60.490000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 51.655000 60.490000 51.975000 ;
      LAYER met4 ;
        RECT 60.170000 51.655000 60.490000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 52.075000 60.490000 52.395000 ;
      LAYER met4 ;
        RECT 60.170000 52.075000 60.490000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170000 52.495000 60.490000 52.815000 ;
      LAYER met4 ;
        RECT 60.170000 52.495000 60.490000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.545000 47.740000 60.865000 48.060000 ;
      LAYER met4 ;
        RECT 60.545000 47.740000 60.865000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.545000 56.410000 60.865000 56.730000 ;
      LAYER met4 ;
        RECT 60.545000 56.410000 60.865000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 36.760000 60.895000 37.080000 ;
      LAYER met4 ;
        RECT 60.575000 36.760000 60.895000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 37.200000 60.895000 37.520000 ;
      LAYER met4 ;
        RECT 60.575000 37.200000 60.895000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 37.640000 60.895000 37.960000 ;
      LAYER met4 ;
        RECT 60.575000 37.640000 60.895000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 38.080000 60.895000 38.400000 ;
      LAYER met4 ;
        RECT 60.575000 38.080000 60.895000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 38.520000 60.895000 38.840000 ;
      LAYER met4 ;
        RECT 60.575000 38.520000 60.895000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 38.960000 60.895000 39.280000 ;
      LAYER met4 ;
        RECT 60.575000 38.960000 60.895000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 39.400000 60.895000 39.720000 ;
      LAYER met4 ;
        RECT 60.575000 39.400000 60.895000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 39.840000 60.895000 40.160000 ;
      LAYER met4 ;
        RECT 60.575000 39.840000 60.895000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 51.655000 60.895000 51.975000 ;
      LAYER met4 ;
        RECT 60.575000 51.655000 60.895000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 52.075000 60.895000 52.395000 ;
      LAYER met4 ;
        RECT 60.575000 52.075000 60.895000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575000 52.495000 60.895000 52.815000 ;
      LAYER met4 ;
        RECT 60.575000 52.495000 60.895000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 47.740000 61.270000 48.060000 ;
      LAYER met4 ;
        RECT 60.950000 47.740000 61.270000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.950000 56.410000 61.270000 56.730000 ;
      LAYER met4 ;
        RECT 60.950000 56.410000 61.270000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 36.760000 61.300000 37.080000 ;
      LAYER met4 ;
        RECT 60.980000 36.760000 61.300000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 37.200000 61.300000 37.520000 ;
      LAYER met4 ;
        RECT 60.980000 37.200000 61.300000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 37.640000 61.300000 37.960000 ;
      LAYER met4 ;
        RECT 60.980000 37.640000 61.300000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 38.080000 61.300000 38.400000 ;
      LAYER met4 ;
        RECT 60.980000 38.080000 61.300000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 38.520000 61.300000 38.840000 ;
      LAYER met4 ;
        RECT 60.980000 38.520000 61.300000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 38.960000 61.300000 39.280000 ;
      LAYER met4 ;
        RECT 60.980000 38.960000 61.300000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 39.400000 61.300000 39.720000 ;
      LAYER met4 ;
        RECT 60.980000 39.400000 61.300000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 39.840000 61.300000 40.160000 ;
      LAYER met4 ;
        RECT 60.980000 39.840000 61.300000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 51.655000 61.300000 51.975000 ;
      LAYER met4 ;
        RECT 60.980000 51.655000 61.300000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 52.075000 61.300000 52.395000 ;
      LAYER met4 ;
        RECT 60.980000 52.075000 61.300000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980000 52.495000 61.300000 52.815000 ;
      LAYER met4 ;
        RECT 60.980000 52.495000 61.300000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.355000 47.740000 61.675000 48.060000 ;
      LAYER met4 ;
        RECT 61.355000 47.740000 61.675000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.355000 56.410000 61.675000 56.730000 ;
      LAYER met4 ;
        RECT 61.355000 56.410000 61.675000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 36.760000 61.705000 37.080000 ;
      LAYER met4 ;
        RECT 61.385000 36.760000 61.705000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 37.200000 61.705000 37.520000 ;
      LAYER met4 ;
        RECT 61.385000 37.200000 61.705000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 37.640000 61.705000 37.960000 ;
      LAYER met4 ;
        RECT 61.385000 37.640000 61.705000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 38.080000 61.705000 38.400000 ;
      LAYER met4 ;
        RECT 61.385000 38.080000 61.705000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 38.520000 61.705000 38.840000 ;
      LAYER met4 ;
        RECT 61.385000 38.520000 61.705000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 38.960000 61.705000 39.280000 ;
      LAYER met4 ;
        RECT 61.385000 38.960000 61.705000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 39.400000 61.705000 39.720000 ;
      LAYER met4 ;
        RECT 61.385000 39.400000 61.705000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 39.840000 61.705000 40.160000 ;
      LAYER met4 ;
        RECT 61.385000 39.840000 61.705000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 51.655000 61.705000 51.975000 ;
      LAYER met4 ;
        RECT 61.385000 51.655000 61.705000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 52.075000 61.705000 52.395000 ;
      LAYER met4 ;
        RECT 61.385000 52.075000 61.705000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385000 52.495000 61.705000 52.815000 ;
      LAYER met4 ;
        RECT 61.385000 52.495000 61.705000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.760000 47.740000 62.080000 48.060000 ;
      LAYER met4 ;
        RECT 61.760000 47.740000 62.080000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.760000 56.410000 62.080000 56.730000 ;
      LAYER met4 ;
        RECT 61.760000 56.410000 62.080000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 36.760000 62.110000 37.080000 ;
      LAYER met4 ;
        RECT 61.790000 36.760000 62.110000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 37.200000 62.110000 37.520000 ;
      LAYER met4 ;
        RECT 61.790000 37.200000 62.110000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 37.640000 62.110000 37.960000 ;
      LAYER met4 ;
        RECT 61.790000 37.640000 62.110000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 38.080000 62.110000 38.400000 ;
      LAYER met4 ;
        RECT 61.790000 38.080000 62.110000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 38.520000 62.110000 38.840000 ;
      LAYER met4 ;
        RECT 61.790000 38.520000 62.110000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 38.960000 62.110000 39.280000 ;
      LAYER met4 ;
        RECT 61.790000 38.960000 62.110000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 39.400000 62.110000 39.720000 ;
      LAYER met4 ;
        RECT 61.790000 39.400000 62.110000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 39.840000 62.110000 40.160000 ;
      LAYER met4 ;
        RECT 61.790000 39.840000 62.110000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 51.655000 62.110000 51.975000 ;
      LAYER met4 ;
        RECT 61.790000 51.655000 62.110000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 52.075000 62.110000 52.395000 ;
      LAYER met4 ;
        RECT 61.790000 52.075000 62.110000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790000 52.495000 62.110000 52.815000 ;
      LAYER met4 ;
        RECT 61.790000 52.495000 62.110000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.165000 47.740000 62.485000 48.060000 ;
      LAYER met4 ;
        RECT 62.165000 47.740000 62.485000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.165000 56.410000 62.485000 56.730000 ;
      LAYER met4 ;
        RECT 62.165000 56.410000 62.485000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 36.760000 62.515000 37.080000 ;
      LAYER met4 ;
        RECT 62.195000 36.760000 62.515000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 37.200000 62.515000 37.520000 ;
      LAYER met4 ;
        RECT 62.195000 37.200000 62.515000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 37.640000 62.515000 37.960000 ;
      LAYER met4 ;
        RECT 62.195000 37.640000 62.515000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 38.080000 62.515000 38.400000 ;
      LAYER met4 ;
        RECT 62.195000 38.080000 62.515000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 38.520000 62.515000 38.840000 ;
      LAYER met4 ;
        RECT 62.195000 38.520000 62.515000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 38.960000 62.515000 39.280000 ;
      LAYER met4 ;
        RECT 62.195000 38.960000 62.515000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 39.400000 62.515000 39.720000 ;
      LAYER met4 ;
        RECT 62.195000 39.400000 62.515000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 39.840000 62.515000 40.160000 ;
      LAYER met4 ;
        RECT 62.195000 39.840000 62.515000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 51.655000 62.515000 51.975000 ;
      LAYER met4 ;
        RECT 62.195000 51.655000 62.515000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 52.075000 62.515000 52.395000 ;
      LAYER met4 ;
        RECT 62.195000 52.075000 62.515000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195000 52.495000 62.515000 52.815000 ;
      LAYER met4 ;
        RECT 62.195000 52.495000 62.515000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.570000 47.740000 62.890000 48.060000 ;
      LAYER met4 ;
        RECT 62.570000 47.740000 62.890000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.570000 56.410000 62.890000 56.730000 ;
      LAYER met4 ;
        RECT 62.570000 56.410000 62.890000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 36.760000 62.920000 37.080000 ;
      LAYER met4 ;
        RECT 62.600000 36.760000 62.920000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 37.200000 62.920000 37.520000 ;
      LAYER met4 ;
        RECT 62.600000 37.200000 62.920000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 37.640000 62.920000 37.960000 ;
      LAYER met4 ;
        RECT 62.600000 37.640000 62.920000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 38.080000 62.920000 38.400000 ;
      LAYER met4 ;
        RECT 62.600000 38.080000 62.920000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 38.520000 62.920000 38.840000 ;
      LAYER met4 ;
        RECT 62.600000 38.520000 62.920000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 38.960000 62.920000 39.280000 ;
      LAYER met4 ;
        RECT 62.600000 38.960000 62.920000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 39.400000 62.920000 39.720000 ;
      LAYER met4 ;
        RECT 62.600000 39.400000 62.920000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 39.840000 62.920000 40.160000 ;
      LAYER met4 ;
        RECT 62.600000 39.840000 62.920000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 51.655000 62.920000 51.975000 ;
      LAYER met4 ;
        RECT 62.600000 51.655000 62.920000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 52.075000 62.920000 52.395000 ;
      LAYER met4 ;
        RECT 62.600000 52.075000 62.920000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600000 52.495000 62.920000 52.815000 ;
      LAYER met4 ;
        RECT 62.600000 52.495000 62.920000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.975000 47.740000 63.295000 48.060000 ;
      LAYER met4 ;
        RECT 62.975000 47.740000 63.295000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.975000 56.410000 63.295000 56.730000 ;
      LAYER met4 ;
        RECT 62.975000 56.410000 63.295000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 36.760000 63.325000 37.080000 ;
      LAYER met4 ;
        RECT 63.005000 36.760000 63.325000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 37.200000 63.325000 37.520000 ;
      LAYER met4 ;
        RECT 63.005000 37.200000 63.325000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 37.640000 63.325000 37.960000 ;
      LAYER met4 ;
        RECT 63.005000 37.640000 63.325000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 38.080000 63.325000 38.400000 ;
      LAYER met4 ;
        RECT 63.005000 38.080000 63.325000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 38.520000 63.325000 38.840000 ;
      LAYER met4 ;
        RECT 63.005000 38.520000 63.325000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 38.960000 63.325000 39.280000 ;
      LAYER met4 ;
        RECT 63.005000 38.960000 63.325000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 39.400000 63.325000 39.720000 ;
      LAYER met4 ;
        RECT 63.005000 39.400000 63.325000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 39.840000 63.325000 40.160000 ;
      LAYER met4 ;
        RECT 63.005000 39.840000 63.325000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 51.655000 63.325000 51.975000 ;
      LAYER met4 ;
        RECT 63.005000 51.655000 63.325000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 52.075000 63.325000 52.395000 ;
      LAYER met4 ;
        RECT 63.005000 52.075000 63.325000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005000 52.495000 63.325000 52.815000 ;
      LAYER met4 ;
        RECT 63.005000 52.495000 63.325000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.380000 47.740000 63.700000 48.060000 ;
      LAYER met4 ;
        RECT 63.380000 47.740000 63.700000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.380000 56.410000 63.700000 56.730000 ;
      LAYER met4 ;
        RECT 63.380000 56.410000 63.700000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 36.760000 63.730000 37.080000 ;
      LAYER met4 ;
        RECT 63.410000 36.760000 63.730000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 37.200000 63.730000 37.520000 ;
      LAYER met4 ;
        RECT 63.410000 37.200000 63.730000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 37.640000 63.730000 37.960000 ;
      LAYER met4 ;
        RECT 63.410000 37.640000 63.730000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 38.080000 63.730000 38.400000 ;
      LAYER met4 ;
        RECT 63.410000 38.080000 63.730000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 38.520000 63.730000 38.840000 ;
      LAYER met4 ;
        RECT 63.410000 38.520000 63.730000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 38.960000 63.730000 39.280000 ;
      LAYER met4 ;
        RECT 63.410000 38.960000 63.730000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 39.400000 63.730000 39.720000 ;
      LAYER met4 ;
        RECT 63.410000 39.400000 63.730000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 39.840000 63.730000 40.160000 ;
      LAYER met4 ;
        RECT 63.410000 39.840000 63.730000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 51.655000 63.730000 51.975000 ;
      LAYER met4 ;
        RECT 63.410000 51.655000 63.730000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 52.075000 63.730000 52.395000 ;
      LAYER met4 ;
        RECT 63.410000 52.075000 63.730000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410000 52.495000 63.730000 52.815000 ;
      LAYER met4 ;
        RECT 63.410000 52.495000 63.730000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.785000 47.740000 64.105000 48.060000 ;
      LAYER met4 ;
        RECT 63.785000 47.740000 64.105000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.785000 56.410000 64.105000 56.730000 ;
      LAYER met4 ;
        RECT 63.785000 56.410000 64.105000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 36.760000 64.135000 37.080000 ;
      LAYER met4 ;
        RECT 63.815000 36.760000 64.135000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 37.200000 64.135000 37.520000 ;
      LAYER met4 ;
        RECT 63.815000 37.200000 64.135000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 37.640000 64.135000 37.960000 ;
      LAYER met4 ;
        RECT 63.815000 37.640000 64.135000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 38.080000 64.135000 38.400000 ;
      LAYER met4 ;
        RECT 63.815000 38.080000 64.135000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 38.520000 64.135000 38.840000 ;
      LAYER met4 ;
        RECT 63.815000 38.520000 64.135000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 38.960000 64.135000 39.280000 ;
      LAYER met4 ;
        RECT 63.815000 38.960000 64.135000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 39.400000 64.135000 39.720000 ;
      LAYER met4 ;
        RECT 63.815000 39.400000 64.135000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 39.840000 64.135000 40.160000 ;
      LAYER met4 ;
        RECT 63.815000 39.840000 64.135000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 51.655000 64.135000 51.975000 ;
      LAYER met4 ;
        RECT 63.815000 51.655000 64.135000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 52.075000 64.135000 52.395000 ;
      LAYER met4 ;
        RECT 63.815000 52.075000 64.135000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815000 52.495000 64.135000 52.815000 ;
      LAYER met4 ;
        RECT 63.815000 52.495000 64.135000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190000 47.740000 64.510000 48.060000 ;
      LAYER met4 ;
        RECT 64.190000 47.740000 64.510000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190000 56.410000 64.510000 56.730000 ;
      LAYER met4 ;
        RECT 64.190000 56.410000 64.510000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 36.760000 64.540000 37.080000 ;
      LAYER met4 ;
        RECT 64.220000 36.760000 64.540000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 37.200000 64.540000 37.520000 ;
      LAYER met4 ;
        RECT 64.220000 37.200000 64.540000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 37.640000 64.540000 37.960000 ;
      LAYER met4 ;
        RECT 64.220000 37.640000 64.540000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 38.080000 64.540000 38.400000 ;
      LAYER met4 ;
        RECT 64.220000 38.080000 64.540000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 38.520000 64.540000 38.840000 ;
      LAYER met4 ;
        RECT 64.220000 38.520000 64.540000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 38.960000 64.540000 39.280000 ;
      LAYER met4 ;
        RECT 64.220000 38.960000 64.540000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 39.400000 64.540000 39.720000 ;
      LAYER met4 ;
        RECT 64.220000 39.400000 64.540000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 39.840000 64.540000 40.160000 ;
      LAYER met4 ;
        RECT 64.220000 39.840000 64.540000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 51.655000 64.540000 51.975000 ;
      LAYER met4 ;
        RECT 64.220000 51.655000 64.540000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 52.075000 64.540000 52.395000 ;
      LAYER met4 ;
        RECT 64.220000 52.075000 64.540000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220000 52.495000 64.540000 52.815000 ;
      LAYER met4 ;
        RECT 64.220000 52.495000 64.540000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.595000 47.740000 64.915000 48.060000 ;
      LAYER met4 ;
        RECT 64.595000 47.740000 64.915000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.595000 56.410000 64.915000 56.730000 ;
      LAYER met4 ;
        RECT 64.595000 56.410000 64.915000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 36.760000 64.945000 37.080000 ;
      LAYER met4 ;
        RECT 64.625000 36.760000 64.945000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 37.200000 64.945000 37.520000 ;
      LAYER met4 ;
        RECT 64.625000 37.200000 64.945000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 37.640000 64.945000 37.960000 ;
      LAYER met4 ;
        RECT 64.625000 37.640000 64.945000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 38.080000 64.945000 38.400000 ;
      LAYER met4 ;
        RECT 64.625000 38.080000 64.945000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 38.520000 64.945000 38.840000 ;
      LAYER met4 ;
        RECT 64.625000 38.520000 64.945000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 38.960000 64.945000 39.280000 ;
      LAYER met4 ;
        RECT 64.625000 38.960000 64.945000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 39.400000 64.945000 39.720000 ;
      LAYER met4 ;
        RECT 64.625000 39.400000 64.945000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 39.840000 64.945000 40.160000 ;
      LAYER met4 ;
        RECT 64.625000 39.840000 64.945000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 51.655000 64.945000 51.975000 ;
      LAYER met4 ;
        RECT 64.625000 51.655000 64.945000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 52.075000 64.945000 52.395000 ;
      LAYER met4 ;
        RECT 64.625000 52.075000 64.945000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625000 52.495000 64.945000 52.815000 ;
      LAYER met4 ;
        RECT 64.625000 52.495000 64.945000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.000000 47.740000 65.320000 48.060000 ;
      LAYER met4 ;
        RECT 65.000000 47.740000 65.320000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.000000 56.410000 65.320000 56.730000 ;
      LAYER met4 ;
        RECT 65.000000 56.410000 65.320000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 36.760000 65.350000 37.080000 ;
      LAYER met4 ;
        RECT 65.030000 36.760000 65.350000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 37.200000 65.350000 37.520000 ;
      LAYER met4 ;
        RECT 65.030000 37.200000 65.350000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 37.640000 65.350000 37.960000 ;
      LAYER met4 ;
        RECT 65.030000 37.640000 65.350000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 38.080000 65.350000 38.400000 ;
      LAYER met4 ;
        RECT 65.030000 38.080000 65.350000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 38.520000 65.350000 38.840000 ;
      LAYER met4 ;
        RECT 65.030000 38.520000 65.350000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 38.960000 65.350000 39.280000 ;
      LAYER met4 ;
        RECT 65.030000 38.960000 65.350000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 39.400000 65.350000 39.720000 ;
      LAYER met4 ;
        RECT 65.030000 39.400000 65.350000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 39.840000 65.350000 40.160000 ;
      LAYER met4 ;
        RECT 65.030000 39.840000 65.350000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 51.655000 65.350000 51.975000 ;
      LAYER met4 ;
        RECT 65.030000 51.655000 65.350000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 52.075000 65.350000 52.395000 ;
      LAYER met4 ;
        RECT 65.030000 52.075000 65.350000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030000 52.495000 65.350000 52.815000 ;
      LAYER met4 ;
        RECT 65.030000 52.495000 65.350000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.405000 47.740000 65.725000 48.060000 ;
      LAYER met4 ;
        RECT 65.405000 47.740000 65.725000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.405000 56.410000 65.725000 56.730000 ;
      LAYER met4 ;
        RECT 65.405000 56.410000 65.725000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 36.760000 65.755000 37.080000 ;
      LAYER met4 ;
        RECT 65.435000 36.760000 65.755000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 37.200000 65.755000 37.520000 ;
      LAYER met4 ;
        RECT 65.435000 37.200000 65.755000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 37.640000 65.755000 37.960000 ;
      LAYER met4 ;
        RECT 65.435000 37.640000 65.755000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 38.080000 65.755000 38.400000 ;
      LAYER met4 ;
        RECT 65.435000 38.080000 65.755000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 38.520000 65.755000 38.840000 ;
      LAYER met4 ;
        RECT 65.435000 38.520000 65.755000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 38.960000 65.755000 39.280000 ;
      LAYER met4 ;
        RECT 65.435000 38.960000 65.755000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 39.400000 65.755000 39.720000 ;
      LAYER met4 ;
        RECT 65.435000 39.400000 65.755000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 39.840000 65.755000 40.160000 ;
      LAYER met4 ;
        RECT 65.435000 39.840000 65.755000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 51.655000 65.755000 51.975000 ;
      LAYER met4 ;
        RECT 65.435000 51.655000 65.755000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 52.075000 65.755000 52.395000 ;
      LAYER met4 ;
        RECT 65.435000 52.075000 65.755000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435000 52.495000 65.755000 52.815000 ;
      LAYER met4 ;
        RECT 65.435000 52.495000 65.755000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810000 47.740000 66.130000 48.060000 ;
      LAYER met4 ;
        RECT 65.810000 47.740000 66.130000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810000 56.410000 66.130000 56.730000 ;
      LAYER met4 ;
        RECT 65.810000 56.410000 66.130000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 36.760000 66.160000 37.080000 ;
      LAYER met4 ;
        RECT 65.840000 36.760000 66.160000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 37.200000 66.160000 37.520000 ;
      LAYER met4 ;
        RECT 65.840000 37.200000 66.160000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 37.640000 66.160000 37.960000 ;
      LAYER met4 ;
        RECT 65.840000 37.640000 66.160000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 38.080000 66.160000 38.400000 ;
      LAYER met4 ;
        RECT 65.840000 38.080000 66.160000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 38.520000 66.160000 38.840000 ;
      LAYER met4 ;
        RECT 65.840000 38.520000 66.160000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 38.960000 66.160000 39.280000 ;
      LAYER met4 ;
        RECT 65.840000 38.960000 66.160000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 39.400000 66.160000 39.720000 ;
      LAYER met4 ;
        RECT 65.840000 39.400000 66.160000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 39.840000 66.160000 40.160000 ;
      LAYER met4 ;
        RECT 65.840000 39.840000 66.160000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 51.655000 66.160000 51.975000 ;
      LAYER met4 ;
        RECT 65.840000 51.655000 66.160000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 52.075000 66.160000 52.395000 ;
      LAYER met4 ;
        RECT 65.840000 52.075000 66.160000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840000 52.495000 66.160000 52.815000 ;
      LAYER met4 ;
        RECT 65.840000 52.495000 66.160000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.215000 47.740000 66.535000 48.060000 ;
      LAYER met4 ;
        RECT 66.215000 47.740000 66.535000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.215000 56.410000 66.535000 56.730000 ;
      LAYER met4 ;
        RECT 66.215000 56.410000 66.535000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 36.760000 66.565000 37.080000 ;
      LAYER met4 ;
        RECT 66.245000 36.760000 66.565000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 37.200000 66.565000 37.520000 ;
      LAYER met4 ;
        RECT 66.245000 37.200000 66.565000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 37.640000 66.565000 37.960000 ;
      LAYER met4 ;
        RECT 66.245000 37.640000 66.565000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 38.080000 66.565000 38.400000 ;
      LAYER met4 ;
        RECT 66.245000 38.080000 66.565000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 38.520000 66.565000 38.840000 ;
      LAYER met4 ;
        RECT 66.245000 38.520000 66.565000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 38.960000 66.565000 39.280000 ;
      LAYER met4 ;
        RECT 66.245000 38.960000 66.565000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 39.400000 66.565000 39.720000 ;
      LAYER met4 ;
        RECT 66.245000 39.400000 66.565000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 39.840000 66.565000 40.160000 ;
      LAYER met4 ;
        RECT 66.245000 39.840000 66.565000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 51.655000 66.565000 51.975000 ;
      LAYER met4 ;
        RECT 66.245000 51.655000 66.565000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 52.075000 66.565000 52.395000 ;
      LAYER met4 ;
        RECT 66.245000 52.075000 66.565000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245000 52.495000 66.565000 52.815000 ;
      LAYER met4 ;
        RECT 66.245000 52.495000 66.565000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.620000 47.740000 66.940000 48.060000 ;
      LAYER met4 ;
        RECT 66.620000 47.740000 66.940000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.620000 56.410000 66.940000 56.730000 ;
      LAYER met4 ;
        RECT 66.620000 56.410000 66.940000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 36.760000 66.970000 37.080000 ;
      LAYER met4 ;
        RECT 66.650000 36.760000 66.970000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 37.200000 66.970000 37.520000 ;
      LAYER met4 ;
        RECT 66.650000 37.200000 66.970000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 37.640000 66.970000 37.960000 ;
      LAYER met4 ;
        RECT 66.650000 37.640000 66.970000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 38.080000 66.970000 38.400000 ;
      LAYER met4 ;
        RECT 66.650000 38.080000 66.970000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 38.520000 66.970000 38.840000 ;
      LAYER met4 ;
        RECT 66.650000 38.520000 66.970000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 38.960000 66.970000 39.280000 ;
      LAYER met4 ;
        RECT 66.650000 38.960000 66.970000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 39.400000 66.970000 39.720000 ;
      LAYER met4 ;
        RECT 66.650000 39.400000 66.970000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 39.840000 66.970000 40.160000 ;
      LAYER met4 ;
        RECT 66.650000 39.840000 66.970000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 51.655000 66.970000 51.975000 ;
      LAYER met4 ;
        RECT 66.650000 51.655000 66.970000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 52.075000 66.970000 52.395000 ;
      LAYER met4 ;
        RECT 66.650000 52.075000 66.970000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650000 52.495000 66.970000 52.815000 ;
      LAYER met4 ;
        RECT 66.650000 52.495000 66.970000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.025000 47.740000 67.345000 48.060000 ;
      LAYER met4 ;
        RECT 67.025000 47.740000 67.345000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.025000 56.410000 67.345000 56.730000 ;
      LAYER met4 ;
        RECT 67.025000 56.410000 67.345000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 36.760000 67.375000 37.080000 ;
      LAYER met4 ;
        RECT 67.055000 36.760000 67.375000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 37.200000 67.375000 37.520000 ;
      LAYER met4 ;
        RECT 67.055000 37.200000 67.375000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 37.640000 67.375000 37.960000 ;
      LAYER met4 ;
        RECT 67.055000 37.640000 67.375000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 38.080000 67.375000 38.400000 ;
      LAYER met4 ;
        RECT 67.055000 38.080000 67.375000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 38.520000 67.375000 38.840000 ;
      LAYER met4 ;
        RECT 67.055000 38.520000 67.375000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 38.960000 67.375000 39.280000 ;
      LAYER met4 ;
        RECT 67.055000 38.960000 67.375000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 39.400000 67.375000 39.720000 ;
      LAYER met4 ;
        RECT 67.055000 39.400000 67.375000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 39.840000 67.375000 40.160000 ;
      LAYER met4 ;
        RECT 67.055000 39.840000 67.375000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 51.655000 67.375000 51.975000 ;
      LAYER met4 ;
        RECT 67.055000 51.655000 67.375000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 52.075000 67.375000 52.395000 ;
      LAYER met4 ;
        RECT 67.055000 52.075000 67.375000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055000 52.495000 67.375000 52.815000 ;
      LAYER met4 ;
        RECT 67.055000 52.495000 67.375000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.430000 47.740000 67.750000 48.060000 ;
      LAYER met4 ;
        RECT 67.430000 47.740000 67.750000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.430000 56.410000 67.750000 56.730000 ;
      LAYER met4 ;
        RECT 67.430000 56.410000 67.750000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 36.760000 67.780000 37.080000 ;
      LAYER met4 ;
        RECT 67.460000 36.760000 67.780000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 37.200000 67.780000 37.520000 ;
      LAYER met4 ;
        RECT 67.460000 37.200000 67.780000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 37.640000 67.780000 37.960000 ;
      LAYER met4 ;
        RECT 67.460000 37.640000 67.780000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 38.080000 67.780000 38.400000 ;
      LAYER met4 ;
        RECT 67.460000 38.080000 67.780000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 38.520000 67.780000 38.840000 ;
      LAYER met4 ;
        RECT 67.460000 38.520000 67.780000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 38.960000 67.780000 39.280000 ;
      LAYER met4 ;
        RECT 67.460000 38.960000 67.780000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 39.400000 67.780000 39.720000 ;
      LAYER met4 ;
        RECT 67.460000 39.400000 67.780000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 39.840000 67.780000 40.160000 ;
      LAYER met4 ;
        RECT 67.460000 39.840000 67.780000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 51.655000 67.780000 51.975000 ;
      LAYER met4 ;
        RECT 67.460000 51.655000 67.780000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 52.075000 67.780000 52.395000 ;
      LAYER met4 ;
        RECT 67.460000 52.075000 67.780000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460000 52.495000 67.780000 52.815000 ;
      LAYER met4 ;
        RECT 67.460000 52.495000 67.780000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.835000 47.740000 68.155000 48.060000 ;
      LAYER met4 ;
        RECT 67.835000 47.740000 68.155000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.835000 56.410000 68.155000 56.730000 ;
      LAYER met4 ;
        RECT 67.835000 56.410000 68.155000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 36.760000 68.185000 37.080000 ;
      LAYER met4 ;
        RECT 67.865000 36.760000 68.185000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 37.200000 68.185000 37.520000 ;
      LAYER met4 ;
        RECT 67.865000 37.200000 68.185000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 37.640000 68.185000 37.960000 ;
      LAYER met4 ;
        RECT 67.865000 37.640000 68.185000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 38.080000 68.185000 38.400000 ;
      LAYER met4 ;
        RECT 67.865000 38.080000 68.185000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 38.520000 68.185000 38.840000 ;
      LAYER met4 ;
        RECT 67.865000 38.520000 68.185000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 38.960000 68.185000 39.280000 ;
      LAYER met4 ;
        RECT 67.865000 38.960000 68.185000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 39.400000 68.185000 39.720000 ;
      LAYER met4 ;
        RECT 67.865000 39.400000 68.185000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 39.840000 68.185000 40.160000 ;
      LAYER met4 ;
        RECT 67.865000 39.840000 68.185000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 51.655000 68.185000 51.975000 ;
      LAYER met4 ;
        RECT 67.865000 51.655000 68.185000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 52.075000 68.185000 52.395000 ;
      LAYER met4 ;
        RECT 67.865000 52.075000 68.185000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865000 52.495000 68.185000 52.815000 ;
      LAYER met4 ;
        RECT 67.865000 52.495000 68.185000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.240000 47.740000 68.560000 48.060000 ;
      LAYER met4 ;
        RECT 68.240000 47.740000 68.560000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.240000 56.410000 68.560000 56.730000 ;
      LAYER met4 ;
        RECT 68.240000 56.410000 68.560000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 36.760000 68.590000 37.080000 ;
      LAYER met4 ;
        RECT 68.270000 36.760000 68.590000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 37.200000 68.590000 37.520000 ;
      LAYER met4 ;
        RECT 68.270000 37.200000 68.590000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 37.640000 68.590000 37.960000 ;
      LAYER met4 ;
        RECT 68.270000 37.640000 68.590000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 38.080000 68.590000 38.400000 ;
      LAYER met4 ;
        RECT 68.270000 38.080000 68.590000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 38.520000 68.590000 38.840000 ;
      LAYER met4 ;
        RECT 68.270000 38.520000 68.590000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 38.960000 68.590000 39.280000 ;
      LAYER met4 ;
        RECT 68.270000 38.960000 68.590000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 39.400000 68.590000 39.720000 ;
      LAYER met4 ;
        RECT 68.270000 39.400000 68.590000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 39.840000 68.590000 40.160000 ;
      LAYER met4 ;
        RECT 68.270000 39.840000 68.590000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 51.655000 68.590000 51.975000 ;
      LAYER met4 ;
        RECT 68.270000 51.655000 68.590000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 52.075000 68.590000 52.395000 ;
      LAYER met4 ;
        RECT 68.270000 52.075000 68.590000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270000 52.495000 68.590000 52.815000 ;
      LAYER met4 ;
        RECT 68.270000 52.495000 68.590000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.645000 47.740000 68.965000 48.060000 ;
      LAYER met4 ;
        RECT 68.645000 47.740000 68.965000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.645000 56.410000 68.965000 56.730000 ;
      LAYER met4 ;
        RECT 68.645000 56.410000 68.965000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 36.760000 68.995000 37.080000 ;
      LAYER met4 ;
        RECT 68.675000 36.760000 68.995000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 37.200000 68.995000 37.520000 ;
      LAYER met4 ;
        RECT 68.675000 37.200000 68.995000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 37.640000 68.995000 37.960000 ;
      LAYER met4 ;
        RECT 68.675000 37.640000 68.995000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 38.080000 68.995000 38.400000 ;
      LAYER met4 ;
        RECT 68.675000 38.080000 68.995000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 38.520000 68.995000 38.840000 ;
      LAYER met4 ;
        RECT 68.675000 38.520000 68.995000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 38.960000 68.995000 39.280000 ;
      LAYER met4 ;
        RECT 68.675000 38.960000 68.995000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 39.400000 68.995000 39.720000 ;
      LAYER met4 ;
        RECT 68.675000 39.400000 68.995000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 39.840000 68.995000 40.160000 ;
      LAYER met4 ;
        RECT 68.675000 39.840000 68.995000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 51.655000 68.995000 51.975000 ;
      LAYER met4 ;
        RECT 68.675000 51.655000 68.995000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 52.075000 68.995000 52.395000 ;
      LAYER met4 ;
        RECT 68.675000 52.075000 68.995000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675000 52.495000 68.995000 52.815000 ;
      LAYER met4 ;
        RECT 68.675000 52.495000 68.995000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 47.740000 69.370000 48.060000 ;
      LAYER met4 ;
        RECT 69.050000 47.740000 69.370000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.050000 56.410000 69.370000 56.730000 ;
      LAYER met4 ;
        RECT 69.050000 56.410000 69.370000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 36.760000 69.400000 37.080000 ;
      LAYER met4 ;
        RECT 69.080000 36.760000 69.400000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 37.200000 69.400000 37.520000 ;
      LAYER met4 ;
        RECT 69.080000 37.200000 69.400000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 37.640000 69.400000 37.960000 ;
      LAYER met4 ;
        RECT 69.080000 37.640000 69.400000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 38.080000 69.400000 38.400000 ;
      LAYER met4 ;
        RECT 69.080000 38.080000 69.400000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 38.520000 69.400000 38.840000 ;
      LAYER met4 ;
        RECT 69.080000 38.520000 69.400000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 38.960000 69.400000 39.280000 ;
      LAYER met4 ;
        RECT 69.080000 38.960000 69.400000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 39.400000 69.400000 39.720000 ;
      LAYER met4 ;
        RECT 69.080000 39.400000 69.400000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 39.840000 69.400000 40.160000 ;
      LAYER met4 ;
        RECT 69.080000 39.840000 69.400000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 51.655000 69.400000 51.975000 ;
      LAYER met4 ;
        RECT 69.080000 51.655000 69.400000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 52.075000 69.400000 52.395000 ;
      LAYER met4 ;
        RECT 69.080000 52.075000 69.400000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080000 52.495000 69.400000 52.815000 ;
      LAYER met4 ;
        RECT 69.080000 52.495000 69.400000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.455000 47.740000 69.775000 48.060000 ;
      LAYER met4 ;
        RECT 69.455000 47.740000 69.775000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.455000 56.410000 69.775000 56.730000 ;
      LAYER met4 ;
        RECT 69.455000 56.410000 69.775000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 36.760000 69.805000 37.080000 ;
      LAYER met4 ;
        RECT 69.485000 36.760000 69.805000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 37.200000 69.805000 37.520000 ;
      LAYER met4 ;
        RECT 69.485000 37.200000 69.805000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 37.640000 69.805000 37.960000 ;
      LAYER met4 ;
        RECT 69.485000 37.640000 69.805000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 38.080000 69.805000 38.400000 ;
      LAYER met4 ;
        RECT 69.485000 38.080000 69.805000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 38.520000 69.805000 38.840000 ;
      LAYER met4 ;
        RECT 69.485000 38.520000 69.805000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 38.960000 69.805000 39.280000 ;
      LAYER met4 ;
        RECT 69.485000 38.960000 69.805000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 39.400000 69.805000 39.720000 ;
      LAYER met4 ;
        RECT 69.485000 39.400000 69.805000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 39.840000 69.805000 40.160000 ;
      LAYER met4 ;
        RECT 69.485000 39.840000 69.805000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 51.655000 69.805000 51.975000 ;
      LAYER met4 ;
        RECT 69.485000 51.655000 69.805000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 52.075000 69.805000 52.395000 ;
      LAYER met4 ;
        RECT 69.485000 52.075000 69.805000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485000 52.495000 69.805000 52.815000 ;
      LAYER met4 ;
        RECT 69.485000 52.495000 69.805000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.860000 47.740000 70.180000 48.060000 ;
      LAYER met4 ;
        RECT 69.860000 47.740000 70.180000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.860000 56.410000 70.180000 56.730000 ;
      LAYER met4 ;
        RECT 69.860000 56.410000 70.180000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 36.760000 70.210000 37.080000 ;
      LAYER met4 ;
        RECT 69.890000 36.760000 70.210000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 37.200000 70.210000 37.520000 ;
      LAYER met4 ;
        RECT 69.890000 37.200000 70.210000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 37.640000 70.210000 37.960000 ;
      LAYER met4 ;
        RECT 69.890000 37.640000 70.210000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 38.080000 70.210000 38.400000 ;
      LAYER met4 ;
        RECT 69.890000 38.080000 70.210000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 38.520000 70.210000 38.840000 ;
      LAYER met4 ;
        RECT 69.890000 38.520000 70.210000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 38.960000 70.210000 39.280000 ;
      LAYER met4 ;
        RECT 69.890000 38.960000 70.210000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 39.400000 70.210000 39.720000 ;
      LAYER met4 ;
        RECT 69.890000 39.400000 70.210000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 39.840000 70.210000 40.160000 ;
      LAYER met4 ;
        RECT 69.890000 39.840000 70.210000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 51.655000 70.210000 51.975000 ;
      LAYER met4 ;
        RECT 69.890000 51.655000 70.210000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 52.075000 70.210000 52.395000 ;
      LAYER met4 ;
        RECT 69.890000 52.075000 70.210000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890000 52.495000 70.210000 52.815000 ;
      LAYER met4 ;
        RECT 69.890000 52.495000 70.210000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 51.655000 7.355000 51.975000 ;
      LAYER met4 ;
        RECT 7.035000 51.655000 7.355000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 52.075000 7.355000 52.395000 ;
      LAYER met4 ;
        RECT 7.035000 52.075000 7.355000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035000 52.495000 7.355000 52.815000 ;
      LAYER met4 ;
        RECT 7.035000 52.495000 7.355000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 47.740000 7.360000 48.060000 ;
      LAYER met4 ;
        RECT 7.040000 47.740000 7.360000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040000 56.410000 7.360000 56.730000 ;
      LAYER met4 ;
        RECT 7.040000 56.410000 7.360000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075000 36.760000 7.395000 37.080000 ;
      LAYER met4 ;
        RECT 7.075000 36.760000 7.395000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075000 37.200000 7.395000 37.520000 ;
      LAYER met4 ;
        RECT 7.075000 37.200000 7.395000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075000 37.640000 7.395000 37.960000 ;
      LAYER met4 ;
        RECT 7.075000 37.640000 7.395000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075000 38.080000 7.395000 38.400000 ;
      LAYER met4 ;
        RECT 7.075000 38.080000 7.395000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075000 38.520000 7.395000 38.840000 ;
      LAYER met4 ;
        RECT 7.075000 38.520000 7.395000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075000 38.960000 7.395000 39.280000 ;
      LAYER met4 ;
        RECT 7.075000 38.960000 7.395000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075000 39.400000 7.395000 39.720000 ;
      LAYER met4 ;
        RECT 7.075000 39.400000 7.395000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075000 39.840000 7.395000 40.160000 ;
      LAYER met4 ;
        RECT 7.075000 39.840000 7.395000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 51.655000 7.760000 51.975000 ;
      LAYER met4 ;
        RECT 7.440000 51.655000 7.760000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 52.075000 7.760000 52.395000 ;
      LAYER met4 ;
        RECT 7.440000 52.075000 7.760000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440000 52.495000 7.760000 52.815000 ;
      LAYER met4 ;
        RECT 7.440000 52.495000 7.760000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 47.740000 7.765000 48.060000 ;
      LAYER met4 ;
        RECT 7.445000 47.740000 7.765000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445000 56.410000 7.765000 56.730000 ;
      LAYER met4 ;
        RECT 7.445000 56.410000 7.765000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480000 36.760000 7.800000 37.080000 ;
      LAYER met4 ;
        RECT 7.480000 36.760000 7.800000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480000 37.200000 7.800000 37.520000 ;
      LAYER met4 ;
        RECT 7.480000 37.200000 7.800000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480000 37.640000 7.800000 37.960000 ;
      LAYER met4 ;
        RECT 7.480000 37.640000 7.800000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480000 38.080000 7.800000 38.400000 ;
      LAYER met4 ;
        RECT 7.480000 38.080000 7.800000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480000 38.520000 7.800000 38.840000 ;
      LAYER met4 ;
        RECT 7.480000 38.520000 7.800000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480000 38.960000 7.800000 39.280000 ;
      LAYER met4 ;
        RECT 7.480000 38.960000 7.800000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480000 39.400000 7.800000 39.720000 ;
      LAYER met4 ;
        RECT 7.480000 39.400000 7.800000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480000 39.840000 7.800000 40.160000 ;
      LAYER met4 ;
        RECT 7.480000 39.840000 7.800000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 51.655000 8.165000 51.975000 ;
      LAYER met4 ;
        RECT 7.845000 51.655000 8.165000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 52.075000 8.165000 52.395000 ;
      LAYER met4 ;
        RECT 7.845000 52.075000 8.165000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845000 52.495000 8.165000 52.815000 ;
      LAYER met4 ;
        RECT 7.845000 52.495000 8.165000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 47.740000 8.170000 48.060000 ;
      LAYER met4 ;
        RECT 7.850000 47.740000 8.170000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850000 56.410000 8.170000 56.730000 ;
      LAYER met4 ;
        RECT 7.850000 56.410000 8.170000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 36.760000 8.205000 37.080000 ;
      LAYER met4 ;
        RECT 7.885000 36.760000 8.205000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 37.200000 8.205000 37.520000 ;
      LAYER met4 ;
        RECT 7.885000 37.200000 8.205000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 37.640000 8.205000 37.960000 ;
      LAYER met4 ;
        RECT 7.885000 37.640000 8.205000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 38.080000 8.205000 38.400000 ;
      LAYER met4 ;
        RECT 7.885000 38.080000 8.205000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 38.520000 8.205000 38.840000 ;
      LAYER met4 ;
        RECT 7.885000 38.520000 8.205000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 38.960000 8.205000 39.280000 ;
      LAYER met4 ;
        RECT 7.885000 38.960000 8.205000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 39.400000 8.205000 39.720000 ;
      LAYER met4 ;
        RECT 7.885000 39.400000 8.205000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885000 39.840000 8.205000 40.160000 ;
      LAYER met4 ;
        RECT 7.885000 39.840000 8.205000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.265000 47.740000 70.585000 48.060000 ;
      LAYER met4 ;
        RECT 70.265000 47.740000 70.585000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.265000 56.410000 70.585000 56.730000 ;
      LAYER met4 ;
        RECT 70.265000 56.410000 70.585000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 36.760000 70.615000 37.080000 ;
      LAYER met4 ;
        RECT 70.295000 36.760000 70.615000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 37.200000 70.615000 37.520000 ;
      LAYER met4 ;
        RECT 70.295000 37.200000 70.615000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 37.640000 70.615000 37.960000 ;
      LAYER met4 ;
        RECT 70.295000 37.640000 70.615000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 38.080000 70.615000 38.400000 ;
      LAYER met4 ;
        RECT 70.295000 38.080000 70.615000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 38.520000 70.615000 38.840000 ;
      LAYER met4 ;
        RECT 70.295000 38.520000 70.615000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 38.960000 70.615000 39.280000 ;
      LAYER met4 ;
        RECT 70.295000 38.960000 70.615000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 39.400000 70.615000 39.720000 ;
      LAYER met4 ;
        RECT 70.295000 39.400000 70.615000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 39.840000 70.615000 40.160000 ;
      LAYER met4 ;
        RECT 70.295000 39.840000 70.615000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 51.655000 70.615000 51.975000 ;
      LAYER met4 ;
        RECT 70.295000 51.655000 70.615000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 52.075000 70.615000 52.395000 ;
      LAYER met4 ;
        RECT 70.295000 52.075000 70.615000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295000 52.495000 70.615000 52.815000 ;
      LAYER met4 ;
        RECT 70.295000 52.495000 70.615000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.670000 47.740000 70.990000 48.060000 ;
      LAYER met4 ;
        RECT 70.670000 47.740000 70.990000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.670000 56.410000 70.990000 56.730000 ;
      LAYER met4 ;
        RECT 70.670000 56.410000 70.990000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 36.760000 71.020000 37.080000 ;
      LAYER met4 ;
        RECT 70.700000 36.760000 71.020000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 37.200000 71.020000 37.520000 ;
      LAYER met4 ;
        RECT 70.700000 37.200000 71.020000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 37.640000 71.020000 37.960000 ;
      LAYER met4 ;
        RECT 70.700000 37.640000 71.020000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 38.080000 71.020000 38.400000 ;
      LAYER met4 ;
        RECT 70.700000 38.080000 71.020000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 38.520000 71.020000 38.840000 ;
      LAYER met4 ;
        RECT 70.700000 38.520000 71.020000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 38.960000 71.020000 39.280000 ;
      LAYER met4 ;
        RECT 70.700000 38.960000 71.020000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 39.400000 71.020000 39.720000 ;
      LAYER met4 ;
        RECT 70.700000 39.400000 71.020000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 39.840000 71.020000 40.160000 ;
      LAYER met4 ;
        RECT 70.700000 39.840000 71.020000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 51.655000 71.020000 51.975000 ;
      LAYER met4 ;
        RECT 70.700000 51.655000 71.020000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 52.075000 71.020000 52.395000 ;
      LAYER met4 ;
        RECT 70.700000 52.075000 71.020000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700000 52.495000 71.020000 52.815000 ;
      LAYER met4 ;
        RECT 70.700000 52.495000 71.020000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.075000 47.740000 71.395000 48.060000 ;
      LAYER met4 ;
        RECT 71.075000 47.740000 71.395000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.075000 56.410000 71.395000 56.730000 ;
      LAYER met4 ;
        RECT 71.075000 56.410000 71.395000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 36.760000 71.425000 37.080000 ;
      LAYER met4 ;
        RECT 71.105000 36.760000 71.425000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 37.200000 71.425000 37.520000 ;
      LAYER met4 ;
        RECT 71.105000 37.200000 71.425000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 37.640000 71.425000 37.960000 ;
      LAYER met4 ;
        RECT 71.105000 37.640000 71.425000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 38.080000 71.425000 38.400000 ;
      LAYER met4 ;
        RECT 71.105000 38.080000 71.425000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 38.520000 71.425000 38.840000 ;
      LAYER met4 ;
        RECT 71.105000 38.520000 71.425000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 38.960000 71.425000 39.280000 ;
      LAYER met4 ;
        RECT 71.105000 38.960000 71.425000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 39.400000 71.425000 39.720000 ;
      LAYER met4 ;
        RECT 71.105000 39.400000 71.425000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 39.840000 71.425000 40.160000 ;
      LAYER met4 ;
        RECT 71.105000 39.840000 71.425000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 51.655000 71.425000 51.975000 ;
      LAYER met4 ;
        RECT 71.105000 51.655000 71.425000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 52.075000 71.425000 52.395000 ;
      LAYER met4 ;
        RECT 71.105000 52.075000 71.425000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105000 52.495000 71.425000 52.815000 ;
      LAYER met4 ;
        RECT 71.105000 52.495000 71.425000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.480000 47.740000 71.800000 48.060000 ;
      LAYER met4 ;
        RECT 71.480000 47.740000 71.800000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.480000 56.410000 71.800000 56.730000 ;
      LAYER met4 ;
        RECT 71.480000 56.410000 71.800000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 36.760000 71.830000 37.080000 ;
      LAYER met4 ;
        RECT 71.510000 36.760000 71.830000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 37.200000 71.830000 37.520000 ;
      LAYER met4 ;
        RECT 71.510000 37.200000 71.830000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 37.640000 71.830000 37.960000 ;
      LAYER met4 ;
        RECT 71.510000 37.640000 71.830000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 38.080000 71.830000 38.400000 ;
      LAYER met4 ;
        RECT 71.510000 38.080000 71.830000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 38.520000 71.830000 38.840000 ;
      LAYER met4 ;
        RECT 71.510000 38.520000 71.830000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 38.960000 71.830000 39.280000 ;
      LAYER met4 ;
        RECT 71.510000 38.960000 71.830000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 39.400000 71.830000 39.720000 ;
      LAYER met4 ;
        RECT 71.510000 39.400000 71.830000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 39.840000 71.830000 40.160000 ;
      LAYER met4 ;
        RECT 71.510000 39.840000 71.830000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 51.655000 71.830000 51.975000 ;
      LAYER met4 ;
        RECT 71.510000 51.655000 71.830000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 52.075000 71.830000 52.395000 ;
      LAYER met4 ;
        RECT 71.510000 52.075000 71.830000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510000 52.495000 71.830000 52.815000 ;
      LAYER met4 ;
        RECT 71.510000 52.495000 71.830000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.890000 47.740000 72.210000 48.060000 ;
      LAYER met4 ;
        RECT 71.890000 47.740000 72.210000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.890000 56.410000 72.210000 56.730000 ;
      LAYER met4 ;
        RECT 71.890000 56.410000 72.210000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 36.760000 72.235000 37.080000 ;
      LAYER met4 ;
        RECT 71.915000 36.760000 72.235000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 37.200000 72.235000 37.520000 ;
      LAYER met4 ;
        RECT 71.915000 37.200000 72.235000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 37.640000 72.235000 37.960000 ;
      LAYER met4 ;
        RECT 71.915000 37.640000 72.235000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 38.080000 72.235000 38.400000 ;
      LAYER met4 ;
        RECT 71.915000 38.080000 72.235000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 38.520000 72.235000 38.840000 ;
      LAYER met4 ;
        RECT 71.915000 38.520000 72.235000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 38.960000 72.235000 39.280000 ;
      LAYER met4 ;
        RECT 71.915000 38.960000 72.235000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 39.400000 72.235000 39.720000 ;
      LAYER met4 ;
        RECT 71.915000 39.400000 72.235000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 39.840000 72.235000 40.160000 ;
      LAYER met4 ;
        RECT 71.915000 39.840000 72.235000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 51.655000 72.235000 51.975000 ;
      LAYER met4 ;
        RECT 71.915000 51.655000 72.235000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 52.075000 72.235000 52.395000 ;
      LAYER met4 ;
        RECT 71.915000 52.075000 72.235000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915000 52.495000 72.235000 52.815000 ;
      LAYER met4 ;
        RECT 71.915000 52.495000 72.235000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.300000 47.740000 72.620000 48.060000 ;
      LAYER met4 ;
        RECT 72.300000 47.740000 72.620000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.300000 56.410000 72.620000 56.730000 ;
      LAYER met4 ;
        RECT 72.300000 56.410000 72.620000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 36.760000 72.640000 37.080000 ;
      LAYER met4 ;
        RECT 72.320000 36.760000 72.640000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 37.200000 72.640000 37.520000 ;
      LAYER met4 ;
        RECT 72.320000 37.200000 72.640000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 37.640000 72.640000 37.960000 ;
      LAYER met4 ;
        RECT 72.320000 37.640000 72.640000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 38.080000 72.640000 38.400000 ;
      LAYER met4 ;
        RECT 72.320000 38.080000 72.640000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 38.520000 72.640000 38.840000 ;
      LAYER met4 ;
        RECT 72.320000 38.520000 72.640000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 38.960000 72.640000 39.280000 ;
      LAYER met4 ;
        RECT 72.320000 38.960000 72.640000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 39.400000 72.640000 39.720000 ;
      LAYER met4 ;
        RECT 72.320000 39.400000 72.640000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 39.840000 72.640000 40.160000 ;
      LAYER met4 ;
        RECT 72.320000 39.840000 72.640000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 51.655000 72.640000 51.975000 ;
      LAYER met4 ;
        RECT 72.320000 51.655000 72.640000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 52.075000 72.640000 52.395000 ;
      LAYER met4 ;
        RECT 72.320000 52.075000 72.640000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320000 52.495000 72.640000 52.815000 ;
      LAYER met4 ;
        RECT 72.320000 52.495000 72.640000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.710000 47.740000 73.030000 48.060000 ;
      LAYER met4 ;
        RECT 72.710000 47.740000 73.030000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.710000 56.410000 73.030000 56.730000 ;
      LAYER met4 ;
        RECT 72.710000 56.410000 73.030000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 36.760000 73.045000 37.080000 ;
      LAYER met4 ;
        RECT 72.725000 36.760000 73.045000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 37.200000 73.045000 37.520000 ;
      LAYER met4 ;
        RECT 72.725000 37.200000 73.045000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 37.640000 73.045000 37.960000 ;
      LAYER met4 ;
        RECT 72.725000 37.640000 73.045000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 38.080000 73.045000 38.400000 ;
      LAYER met4 ;
        RECT 72.725000 38.080000 73.045000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 38.520000 73.045000 38.840000 ;
      LAYER met4 ;
        RECT 72.725000 38.520000 73.045000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 38.960000 73.045000 39.280000 ;
      LAYER met4 ;
        RECT 72.725000 38.960000 73.045000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 39.400000 73.045000 39.720000 ;
      LAYER met4 ;
        RECT 72.725000 39.400000 73.045000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 39.840000 73.045000 40.160000 ;
      LAYER met4 ;
        RECT 72.725000 39.840000 73.045000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 51.655000 73.045000 51.975000 ;
      LAYER met4 ;
        RECT 72.725000 51.655000 73.045000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 52.075000 73.045000 52.395000 ;
      LAYER met4 ;
        RECT 72.725000 52.075000 73.045000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725000 52.495000 73.045000 52.815000 ;
      LAYER met4 ;
        RECT 72.725000 52.495000 73.045000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.120000 47.740000 73.440000 48.060000 ;
      LAYER met4 ;
        RECT 73.120000 47.740000 73.440000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.120000 56.410000 73.440000 56.730000 ;
      LAYER met4 ;
        RECT 73.120000 56.410000 73.440000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 36.760000 73.450000 37.080000 ;
      LAYER met4 ;
        RECT 73.130000 36.760000 73.450000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 37.200000 73.450000 37.520000 ;
      LAYER met4 ;
        RECT 73.130000 37.200000 73.450000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 37.640000 73.450000 37.960000 ;
      LAYER met4 ;
        RECT 73.130000 37.640000 73.450000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 38.080000 73.450000 38.400000 ;
      LAYER met4 ;
        RECT 73.130000 38.080000 73.450000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 38.520000 73.450000 38.840000 ;
      LAYER met4 ;
        RECT 73.130000 38.520000 73.450000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 38.960000 73.450000 39.280000 ;
      LAYER met4 ;
        RECT 73.130000 38.960000 73.450000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 39.400000 73.450000 39.720000 ;
      LAYER met4 ;
        RECT 73.130000 39.400000 73.450000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 39.840000 73.450000 40.160000 ;
      LAYER met4 ;
        RECT 73.130000 39.840000 73.450000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 51.655000 73.450000 51.975000 ;
      LAYER met4 ;
        RECT 73.130000 51.655000 73.450000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 52.075000 73.450000 52.395000 ;
      LAYER met4 ;
        RECT 73.130000 52.075000 73.450000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130000 52.495000 73.450000 52.815000 ;
      LAYER met4 ;
        RECT 73.130000 52.495000 73.450000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530000 47.740000 73.850000 48.060000 ;
      LAYER met4 ;
        RECT 73.530000 47.740000 73.850000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530000 56.410000 73.850000 56.730000 ;
      LAYER met4 ;
        RECT 73.530000 56.410000 73.850000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 36.760000 73.855000 37.080000 ;
      LAYER met4 ;
        RECT 73.535000 36.760000 73.855000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 37.200000 73.855000 37.520000 ;
      LAYER met4 ;
        RECT 73.535000 37.200000 73.855000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 37.640000 73.855000 37.960000 ;
      LAYER met4 ;
        RECT 73.535000 37.640000 73.855000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 38.080000 73.855000 38.400000 ;
      LAYER met4 ;
        RECT 73.535000 38.080000 73.855000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 38.520000 73.855000 38.840000 ;
      LAYER met4 ;
        RECT 73.535000 38.520000 73.855000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 38.960000 73.855000 39.280000 ;
      LAYER met4 ;
        RECT 73.535000 38.960000 73.855000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 39.400000 73.855000 39.720000 ;
      LAYER met4 ;
        RECT 73.535000 39.400000 73.855000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 39.840000 73.855000 40.160000 ;
      LAYER met4 ;
        RECT 73.535000 39.840000 73.855000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 51.655000 73.855000 51.975000 ;
      LAYER met4 ;
        RECT 73.535000 51.655000 73.855000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 52.075000 73.855000 52.395000 ;
      LAYER met4 ;
        RECT 73.535000 52.075000 73.855000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535000 52.495000 73.855000 52.815000 ;
      LAYER met4 ;
        RECT 73.535000 52.495000 73.855000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 36.760000 74.260000 37.080000 ;
      LAYER met4 ;
        RECT 73.940000 36.760000 74.260000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 37.200000 74.260000 37.520000 ;
      LAYER met4 ;
        RECT 73.940000 37.200000 74.260000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 37.640000 74.260000 37.960000 ;
      LAYER met4 ;
        RECT 73.940000 37.640000 74.260000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 38.080000 74.260000 38.400000 ;
      LAYER met4 ;
        RECT 73.940000 38.080000 74.260000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 38.520000 74.260000 38.840000 ;
      LAYER met4 ;
        RECT 73.940000 38.520000 74.260000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 38.960000 74.260000 39.280000 ;
      LAYER met4 ;
        RECT 73.940000 38.960000 74.260000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 39.400000 74.260000 39.720000 ;
      LAYER met4 ;
        RECT 73.940000 39.400000 74.260000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 39.840000 74.260000 40.160000 ;
      LAYER met4 ;
        RECT 73.940000 39.840000 74.260000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 47.740000 74.260000 48.060000 ;
      LAYER met4 ;
        RECT 73.940000 47.740000 74.260000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 51.655000 74.260000 51.975000 ;
      LAYER met4 ;
        RECT 73.940000 51.655000 74.260000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 52.075000 74.260000 52.395000 ;
      LAYER met4 ;
        RECT 73.940000 52.075000 74.260000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 52.495000 74.260000 52.815000 ;
      LAYER met4 ;
        RECT 73.940000 52.495000 74.260000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940000 56.410000 74.260000 56.730000 ;
      LAYER met4 ;
        RECT 73.940000 56.410000 74.260000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 51.655000 8.570000 51.975000 ;
      LAYER met4 ;
        RECT 8.250000 51.655000 8.570000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 52.075000 8.570000 52.395000 ;
      LAYER met4 ;
        RECT 8.250000 52.075000 8.570000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250000 52.495000 8.570000 52.815000 ;
      LAYER met4 ;
        RECT 8.250000 52.495000 8.570000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 47.740000 8.575000 48.060000 ;
      LAYER met4 ;
        RECT 8.255000 47.740000 8.575000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255000 56.410000 8.575000 56.730000 ;
      LAYER met4 ;
        RECT 8.255000 56.410000 8.575000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290000 36.760000 8.610000 37.080000 ;
      LAYER met4 ;
        RECT 8.290000 36.760000 8.610000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290000 37.200000 8.610000 37.520000 ;
      LAYER met4 ;
        RECT 8.290000 37.200000 8.610000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290000 37.640000 8.610000 37.960000 ;
      LAYER met4 ;
        RECT 8.290000 37.640000 8.610000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290000 38.080000 8.610000 38.400000 ;
      LAYER met4 ;
        RECT 8.290000 38.080000 8.610000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290000 38.520000 8.610000 38.840000 ;
      LAYER met4 ;
        RECT 8.290000 38.520000 8.610000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290000 38.960000 8.610000 39.280000 ;
      LAYER met4 ;
        RECT 8.290000 38.960000 8.610000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290000 39.400000 8.610000 39.720000 ;
      LAYER met4 ;
        RECT 8.290000 39.400000 8.610000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290000 39.840000 8.610000 40.160000 ;
      LAYER met4 ;
        RECT 8.290000 39.840000 8.610000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 51.655000 8.975000 51.975000 ;
      LAYER met4 ;
        RECT 8.655000 51.655000 8.975000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 52.075000 8.975000 52.395000 ;
      LAYER met4 ;
        RECT 8.655000 52.075000 8.975000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655000 52.495000 8.975000 52.815000 ;
      LAYER met4 ;
        RECT 8.655000 52.495000 8.975000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 47.740000 8.980000 48.060000 ;
      LAYER met4 ;
        RECT 8.660000 47.740000 8.980000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660000 56.410000 8.980000 56.730000 ;
      LAYER met4 ;
        RECT 8.660000 56.410000 8.980000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695000 36.760000 9.015000 37.080000 ;
      LAYER met4 ;
        RECT 8.695000 36.760000 9.015000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695000 37.200000 9.015000 37.520000 ;
      LAYER met4 ;
        RECT 8.695000 37.200000 9.015000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695000 37.640000 9.015000 37.960000 ;
      LAYER met4 ;
        RECT 8.695000 37.640000 9.015000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695000 38.080000 9.015000 38.400000 ;
      LAYER met4 ;
        RECT 8.695000 38.080000 9.015000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695000 38.520000 9.015000 38.840000 ;
      LAYER met4 ;
        RECT 8.695000 38.520000 9.015000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695000 38.960000 9.015000 39.280000 ;
      LAYER met4 ;
        RECT 8.695000 38.960000 9.015000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695000 39.400000 9.015000 39.720000 ;
      LAYER met4 ;
        RECT 8.695000 39.400000 9.015000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695000 39.840000 9.015000 40.160000 ;
      LAYER met4 ;
        RECT 8.695000 39.840000 9.015000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 51.655000 9.380000 51.975000 ;
      LAYER met4 ;
        RECT 9.060000 51.655000 9.380000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 52.075000 9.380000 52.395000 ;
      LAYER met4 ;
        RECT 9.060000 52.075000 9.380000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060000 52.495000 9.380000 52.815000 ;
      LAYER met4 ;
        RECT 9.060000 52.495000 9.380000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 47.740000 9.385000 48.060000 ;
      LAYER met4 ;
        RECT 9.065000 47.740000 9.385000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065000 56.410000 9.385000 56.730000 ;
      LAYER met4 ;
        RECT 9.065000 56.410000 9.385000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100000 36.760000 9.420000 37.080000 ;
      LAYER met4 ;
        RECT 9.100000 36.760000 9.420000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100000 37.200000 9.420000 37.520000 ;
      LAYER met4 ;
        RECT 9.100000 37.200000 9.420000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100000 37.640000 9.420000 37.960000 ;
      LAYER met4 ;
        RECT 9.100000 37.640000 9.420000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100000 38.080000 9.420000 38.400000 ;
      LAYER met4 ;
        RECT 9.100000 38.080000 9.420000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100000 38.520000 9.420000 38.840000 ;
      LAYER met4 ;
        RECT 9.100000 38.520000 9.420000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100000 38.960000 9.420000 39.280000 ;
      LAYER met4 ;
        RECT 9.100000 38.960000 9.420000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100000 39.400000 9.420000 39.720000 ;
      LAYER met4 ;
        RECT 9.100000 39.400000 9.420000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100000 39.840000 9.420000 40.160000 ;
      LAYER met4 ;
        RECT 9.100000 39.840000 9.420000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 51.655000 9.785000 51.975000 ;
      LAYER met4 ;
        RECT 9.465000 51.655000 9.785000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 52.075000 9.785000 52.395000 ;
      LAYER met4 ;
        RECT 9.465000 52.075000 9.785000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465000 52.495000 9.785000 52.815000 ;
      LAYER met4 ;
        RECT 9.465000 52.495000 9.785000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 47.740000 9.790000 48.060000 ;
      LAYER met4 ;
        RECT 9.470000 47.740000 9.790000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470000 56.410000 9.790000 56.730000 ;
      LAYER met4 ;
        RECT 9.470000 56.410000 9.790000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505000 36.760000 9.825000 37.080000 ;
      LAYER met4 ;
        RECT 9.505000 36.760000 9.825000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505000 37.200000 9.825000 37.520000 ;
      LAYER met4 ;
        RECT 9.505000 37.200000 9.825000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505000 37.640000 9.825000 37.960000 ;
      LAYER met4 ;
        RECT 9.505000 37.640000 9.825000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505000 38.080000 9.825000 38.400000 ;
      LAYER met4 ;
        RECT 9.505000 38.080000 9.825000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505000 38.520000 9.825000 38.840000 ;
      LAYER met4 ;
        RECT 9.505000 38.520000 9.825000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505000 38.960000 9.825000 39.280000 ;
      LAYER met4 ;
        RECT 9.505000 38.960000 9.825000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505000 39.400000 9.825000 39.720000 ;
      LAYER met4 ;
        RECT 9.505000 39.400000 9.825000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505000 39.840000 9.825000 40.160000 ;
      LAYER met4 ;
        RECT 9.505000 39.840000 9.825000 40.160000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 51.655000 10.190000 51.975000 ;
      LAYER met4 ;
        RECT 9.870000 51.655000 10.190000 51.975000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 52.075000 10.190000 52.395000 ;
      LAYER met4 ;
        RECT 9.870000 52.075000 10.190000 52.395000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870000 52.495000 10.190000 52.815000 ;
      LAYER met4 ;
        RECT 9.870000 52.495000 10.190000 52.815000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 47.740000 10.195000 48.060000 ;
      LAYER met4 ;
        RECT 9.875000 47.740000 10.195000 48.060000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875000 56.410000 10.195000 56.730000 ;
      LAYER met4 ;
        RECT 9.875000 56.410000 10.195000 56.730000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910000 36.760000 10.230000 37.080000 ;
      LAYER met4 ;
        RECT 9.910000 36.760000 10.230000 37.080000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910000 37.200000 10.230000 37.520000 ;
      LAYER met4 ;
        RECT 9.910000 37.200000 10.230000 37.520000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910000 37.640000 10.230000 37.960000 ;
      LAYER met4 ;
        RECT 9.910000 37.640000 10.230000 37.960000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910000 38.080000 10.230000 38.400000 ;
      LAYER met4 ;
        RECT 9.910000 38.080000 10.230000 38.400000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910000 38.520000 10.230000 38.840000 ;
      LAYER met4 ;
        RECT 9.910000 38.520000 10.230000 38.840000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910000 38.960000 10.230000 39.280000 ;
      LAYER met4 ;
        RECT 9.910000 38.960000 10.230000 39.280000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910000 39.400000 10.230000 39.720000 ;
      LAYER met4 ;
        RECT 9.910000 39.400000 10.230000 39.720000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910000 39.840000 10.230000 40.160000 ;
      LAYER met4 ;
        RECT 9.910000 39.840000 10.230000 40.160000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 41.685000 75.000000 46.135000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 25.935000 75.000000 30.385000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730000 58.335000 75.000000 62.585000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730000 31.985000 75.000000 35.235000 ;
    END
  END VSWITCH
  OBS
    LAYER met3 ;
      RECT 0.495000 36.740000 74.290000 56.730000 ;
    LAYER met4 ;
      RECT 0.000000  2.035000 75.000000  47.965000 ;
      RECT 0.000000 51.745000 75.000000  52.725000 ;
      RECT 0.000000 56.505000 75.000000 200.000000 ;
    LAYER met5 ;
      RECT 0.000000  2.135000 72.130000  15.035000 ;
      RECT 0.000000 15.035000 72.435000  19.885000 ;
      RECT 0.000000 19.885000 75.000000  24.335000 ;
      RECT 0.000000 24.335000 72.130000  36.835000 ;
      RECT 0.000000 36.835000 75.000000  40.085000 ;
      RECT 0.000000 40.085000 72.130000  47.735000 ;
      RECT 0.000000 47.735000 75.000000  56.735000 ;
      RECT 0.000000 56.735000 72.130000  96.585000 ;
      RECT 0.000000 96.585000 75.000000 200.000000 ;
  END
END sky130_fd_io__overlay_vssa_hvc
END LIBRARY
