/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_IO__TOP_POWER_HVC_WPADV2_PP_BLACKBOX_V
`define SKY130_FD_IO__TOP_POWER_HVC_WPADV2_PP_BLACKBOX_V

/**
 * top_power_hvc_wpadv2: A power pad with an ESD high-voltage clamp.
 *
 * Verilog stub definition (black box with power pins).
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_io__top_power_hvc_wpadv2 (
           P_PAD      ,
           AMUXBUS_A  ,
           AMUXBUS_B  ,
           OGC_HVC    ,
           DRN_HVC    ,
           SRC_BDY_HVC,
           P_CORE     ,
           VDDIO      ,
           VDDIO_Q    ,
           VDDA       ,
           VCCD       ,
           VSWITCH    ,
           VCCHIB     ,
           VSSA       ,
           VSSD       ,
           VSSIO_Q    ,
           VSSIO
       );

inout P_PAD      ;
inout AMUXBUS_A  ;
inout AMUXBUS_B  ;
inout OGC_HVC    ;
inout DRN_HVC    ;
inout SRC_BDY_HVC;
inout P_CORE     ;
inout VDDIO      ;
inout VDDIO_Q    ;
inout VDDA       ;
inout VCCD       ;
inout VSWITCH    ;
inout VCCHIB     ;
inout VSSA       ;
inout VSSD       ;
inout VSSIO_Q    ;
inout VSSIO      ;
endmodule

`default_nettype wire
`endif  // SKY130_FD_IO__TOP_POWER_HVC_WPADV2_PP_BLACKBOX_V
